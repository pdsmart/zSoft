-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b87fa",
             1 => x"f80d0b0b",
             2 => x"0b93e904",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"cd040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b93b0",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b83be",
           162 => x"bc738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93b50400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0bac",
           171 => x"cc2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0bab",
           179 => x"ab2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"96040b0b",
           269 => x"0b8ca604",
           270 => x"0b0b0b8c",
           271 => x"b6040b0b",
           272 => x"0b8cc604",
           273 => x"0b0b0b8c",
           274 => x"d6040b0b",
           275 => x"0b8ce604",
           276 => x"0b0b0b8c",
           277 => x"f6040b0b",
           278 => x"0b8d8604",
           279 => x"0b0b0b8d",
           280 => x"96040b0b",
           281 => x"0b8da604",
           282 => x"0b0b0b8d",
           283 => x"b6040b0b",
           284 => x"0b8dc604",
           285 => x"0b0b0b8d",
           286 => x"d7040b0b",
           287 => x"0b8de804",
           288 => x"0b0b0b8d",
           289 => x"f9040b0b",
           290 => x"0b8e8a04",
           291 => x"0b0b0b8e",
           292 => x"9b040b0b",
           293 => x"0b8eac04",
           294 => x"0b0b0b8e",
           295 => x"bd040b0b",
           296 => x"0b8ece04",
           297 => x"0b0b0b8e",
           298 => x"df040b0b",
           299 => x"0b8ef004",
           300 => x"0b0b0b8f",
           301 => x"81040b0b",
           302 => x"0b8f9204",
           303 => x"0b0b0b8f",
           304 => x"a3040b0b",
           305 => x"0b8fb404",
           306 => x"0b0b0b8f",
           307 => x"c5040b0b",
           308 => x"0b8fd604",
           309 => x"0b0b0b8f",
           310 => x"e7040b0b",
           311 => x"0b8ff804",
           312 => x"0b0b0b90",
           313 => x"89040b0b",
           314 => x"0b909a04",
           315 => x"0b0b0b90",
           316 => x"ab040b0b",
           317 => x"0b90bc04",
           318 => x"0b0b0b90",
           319 => x"cd040b0b",
           320 => x"0b90de04",
           321 => x"0b0b0b90",
           322 => x"ef040b0b",
           323 => x"0b918004",
           324 => x"0b0b0b91",
           325 => x"91040b0b",
           326 => x"0b91a204",
           327 => x"0b0b0b91",
           328 => x"b3040b0b",
           329 => x"0b91c404",
           330 => x"0b0b0b91",
           331 => x"d5040b0b",
           332 => x"0b91e604",
           333 => x"0b0b0b91",
           334 => x"f7040b0b",
           335 => x"0b928804",
           336 => x"0b0b0b92",
           337 => x"99040b0b",
           338 => x"0b92aa04",
           339 => x"0b0b0b92",
           340 => x"bb040b0b",
           341 => x"0b92cb04",
           342 => x"0b0b0b92",
           343 => x"dc040b0b",
           344 => x"0b92ed04",
           345 => x"0b0b0b92",
           346 => x"fe04ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0484ba98",
           386 => x"0c80d5f6",
           387 => x"2d84ba98",
           388 => x"0880c080",
           389 => x"900484ba",
           390 => x"980ca2ee",
           391 => x"2d84ba98",
           392 => x"0880c080",
           393 => x"900484ba",
           394 => x"980ca0f3",
           395 => x"2d84ba98",
           396 => x"0880c080",
           397 => x"900484ba",
           398 => x"980ca0e0",
           399 => x"2d84ba98",
           400 => x"0880c080",
           401 => x"900484ba",
           402 => x"980c94a3",
           403 => x"2d84ba98",
           404 => x"0880c080",
           405 => x"900484ba",
           406 => x"980ca1f6",
           407 => x"2d84ba98",
           408 => x"0880c080",
           409 => x"900484ba",
           410 => x"980caf86",
           411 => x"2d84ba98",
           412 => x"0880c080",
           413 => x"900484ba",
           414 => x"980cad82",
           415 => x"2d84ba98",
           416 => x"0880c080",
           417 => x"900484ba",
           418 => x"980c9488",
           419 => x"2d84ba98",
           420 => x"0880c080",
           421 => x"900484ba",
           422 => x"980c95a8",
           423 => x"2d84ba98",
           424 => x"0880c080",
           425 => x"900484ba",
           426 => x"980c95d1",
           427 => x"2d84ba98",
           428 => x"0880c080",
           429 => x"900484ba",
           430 => x"980cb18a",
           431 => x"2d84ba98",
           432 => x"0880c080",
           433 => x"900484ba",
           434 => x"980c80d4",
           435 => x"db2d84ba",
           436 => x"980880c0",
           437 => x"80900484",
           438 => x"ba980c80",
           439 => x"d5c02d84",
           440 => x"ba980880",
           441 => x"c0809004",
           442 => x"84ba980c",
           443 => x"80d2972d",
           444 => x"84ba9808",
           445 => x"80c08090",
           446 => x"0484ba98",
           447 => x"0c80d3ca",
           448 => x"2d84ba98",
           449 => x"0880c080",
           450 => x"900484ba",
           451 => x"980c82c9",
           452 => x"f72d84ba",
           453 => x"980880c0",
           454 => x"80900484",
           455 => x"ba980c82",
           456 => x"e3c92d84",
           457 => x"ba980880",
           458 => x"c0809004",
           459 => x"84ba980c",
           460 => x"82d2e72d",
           461 => x"84ba9808",
           462 => x"80c08090",
           463 => x"0484ba98",
           464 => x"0c82d889",
           465 => x"2d84ba98",
           466 => x"0880c080",
           467 => x"900484ba",
           468 => x"980c82ed",
           469 => x"e62d84ba",
           470 => x"980880c0",
           471 => x"80900484",
           472 => x"ba980c82",
           473 => x"faee2d84",
           474 => x"ba980880",
           475 => x"c0809004",
           476 => x"84ba980c",
           477 => x"82dfd02d",
           478 => x"84ba9808",
           479 => x"80c08090",
           480 => x"0484ba98",
           481 => x"0c82f287",
           482 => x"2d84ba98",
           483 => x"0880c080",
           484 => x"900484ba",
           485 => x"980c82f3",
           486 => x"d42d84ba",
           487 => x"980880c0",
           488 => x"80900484",
           489 => x"ba980c82",
           490 => x"f4a92d84",
           491 => x"ba980880",
           492 => x"c0809004",
           493 => x"84ba980c",
           494 => x"8384eb2d",
           495 => x"84ba9808",
           496 => x"80c08090",
           497 => x"0484ba98",
           498 => x"0c82ffb0",
           499 => x"2d84ba98",
           500 => x"0880c080",
           501 => x"900484ba",
           502 => x"980c838b",
           503 => x"cf2d84ba",
           504 => x"980880c0",
           505 => x"80900484",
           506 => x"ba980c82",
           507 => x"f6862d84",
           508 => x"ba980880",
           509 => x"c0809004",
           510 => x"84ba980c",
           511 => x"8394c62d",
           512 => x"84ba9808",
           513 => x"80c08090",
           514 => x"0484ba98",
           515 => x"0c8395d1",
           516 => x"2d84ba98",
           517 => x"0880c080",
           518 => x"900484ba",
           519 => x"980c82e6",
           520 => x"992d84ba",
           521 => x"980880c0",
           522 => x"80900484",
           523 => x"ba980c82",
           524 => x"e4b02d84",
           525 => x"ba980880",
           526 => x"c0809004",
           527 => x"84ba980c",
           528 => x"82e7d72d",
           529 => x"84ba9808",
           530 => x"80c08090",
           531 => x"0484ba98",
           532 => x"0c82f6f0",
           533 => x"2d84ba98",
           534 => x"0880c080",
           535 => x"900484ba",
           536 => x"980c8396",
           537 => x"e32d84ba",
           538 => x"980880c0",
           539 => x"80900484",
           540 => x"ba980c83",
           541 => x"9ac02d84",
           542 => x"ba980880",
           543 => x"c0809004",
           544 => x"84ba980c",
           545 => x"83a1b22d",
           546 => x"84ba9808",
           547 => x"80c08090",
           548 => x"0484ba98",
           549 => x"0c82c7c8",
           550 => x"2d84ba98",
           551 => x"0880c080",
           552 => x"900484ba",
           553 => x"980c83a4",
           554 => x"db2d84ba",
           555 => x"980880c0",
           556 => x"80900484",
           557 => x"ba980c83",
           558 => x"b9dc2d84",
           559 => x"ba980880",
           560 => x"c0809004",
           561 => x"84ba980c",
           562 => x"83b88e2d",
           563 => x"84ba9808",
           564 => x"80c08090",
           565 => x"0484ba98",
           566 => x"0c81f4ac",
           567 => x"2d84ba98",
           568 => x"0880c080",
           569 => x"900484ba",
           570 => x"980c81f5",
           571 => x"ab2d84ba",
           572 => x"980880c0",
           573 => x"80900484",
           574 => x"ba980c81",
           575 => x"f6aa2d84",
           576 => x"ba980880",
           577 => x"c0809004",
           578 => x"84ba980c",
           579 => x"80d0992d",
           580 => x"84ba9808",
           581 => x"80c08090",
           582 => x"0484ba98",
           583 => x"0c80d1e9",
           584 => x"2d84ba98",
           585 => x"0880c080",
           586 => x"900484ba",
           587 => x"980c80d7",
           588 => x"942d84ba",
           589 => x"980880c0",
           590 => x"80900484",
           591 => x"ba980cb1",
           592 => x"9a2d84ba",
           593 => x"980880c0",
           594 => x"80900484",
           595 => x"ba980c81",
           596 => x"dbca2d84",
           597 => x"ba980880",
           598 => x"c0809004",
           599 => x"84ba980c",
           600 => x"81dd852d",
           601 => x"84ba9808",
           602 => x"80c08090",
           603 => x"0484ba98",
           604 => x"0c81f286",
           605 => x"2d84ba98",
           606 => x"0880c080",
           607 => x"900484ba",
           608 => x"980c81d5",
           609 => x"da2d84ba",
           610 => x"980880c0",
           611 => x"8090043c",
           612 => x"04101010",
           613 => x"10101010",
           614 => x"10101010",
           615 => x"10101010",
           616 => x"10101010",
           617 => x"10101010",
           618 => x"10101010",
           619 => x"10101010",
           620 => x"53510400",
           621 => x"007381ff",
           622 => x"06738306",
           623 => x"09810583",
           624 => x"05101010",
           625 => x"2b0772fc",
           626 => x"060c5151",
           627 => x"04727280",
           628 => x"728106ff",
           629 => x"05097206",
           630 => x"05711052",
           631 => x"720a100a",
           632 => x"5372ed38",
           633 => x"51515351",
           634 => x"0484ba8c",
           635 => x"7084d5f8",
           636 => x"278e3880",
           637 => x"71708405",
           638 => x"530c0b0b",
           639 => x"0b93ec04",
           640 => x"8c815180",
           641 => x"cec40400",
           642 => x"fc3d0d87",
           643 => x"3d707084",
           644 => x"05520856",
           645 => x"53745284",
           646 => x"d5f00851",
           647 => x"81c53f86",
           648 => x"3d0d04fa",
           649 => x"3d0d787a",
           650 => x"7c851133",
           651 => x"81328106",
           652 => x"80732507",
           653 => x"56585557",
           654 => x"80527272",
           655 => x"2e098106",
           656 => x"80d338ff",
           657 => x"1477748a",
           658 => x"32703070",
           659 => x"72079f2a",
           660 => x"51555556",
           661 => x"54807425",
           662 => x"b7387180",
           663 => x"2eb23875",
           664 => x"518efa3f",
           665 => x"84ba8c08",
           666 => x"5384ba8c",
           667 => x"08ff2eae",
           668 => x"3884ba8c",
           669 => x"08757081",
           670 => x"055734ff",
           671 => x"14738a32",
           672 => x"70307072",
           673 => x"079f2a51",
           674 => x"54545473",
           675 => x"8024cb38",
           676 => x"80753476",
           677 => x"527184ba",
           678 => x"8c0c883d",
           679 => x"0d04800b",
           680 => x"84ba8c0c",
           681 => x"883d0d04",
           682 => x"f53d0d7d",
           683 => x"54860284",
           684 => x"05990534",
           685 => x"7356fe0a",
           686 => x"588e3d88",
           687 => x"05537e52",
           688 => x"8d3de405",
           689 => x"519d3f73",
           690 => x"19548074",
           691 => x"348d3d0d",
           692 => x"04fd3d0d",
           693 => x"863d8805",
           694 => x"53765275",
           695 => x"51853f85",
           696 => x"3d0d04f1",
           697 => x"3d0d6163",
           698 => x"65425d5d",
           699 => x"80708c1f",
           700 => x"0c851e33",
           701 => x"70812a81",
           702 => x"32810655",
           703 => x"555bff54",
           704 => x"727b2e09",
           705 => x"810680d2",
           706 => x"387b3357",
           707 => x"767b2e80",
           708 => x"c538811c",
           709 => x"7b810654",
           710 => x"5c72802e",
           711 => x"818138d0",
           712 => x"175f7e89",
           713 => x"2681a338",
           714 => x"76b03270",
           715 => x"30708025",
           716 => x"51545578",
           717 => x"ae387280",
           718 => x"2ea9387a",
           719 => x"832a7081",
           720 => x"32810640",
           721 => x"547e802e",
           722 => x"9e387a82",
           723 => x"80075b7b",
           724 => x"335776ff",
           725 => x"bd388c1d",
           726 => x"08547384",
           727 => x"ba8c0c91",
           728 => x"3d0d047a",
           729 => x"832a5478",
           730 => x"10101079",
           731 => x"10057098",
           732 => x"2b70982c",
           733 => x"19708180",
           734 => x"0a298b0a",
           735 => x"0570982c",
           736 => x"525a5b56",
           737 => x"5f807924",
           738 => x"81863873",
           739 => x"81065372",
           740 => x"ffbd3878",
           741 => x"7c335858",
           742 => x"76fef738",
           743 => x"ffb83976",
           744 => x"a52e0981",
           745 => x"06933881",
           746 => x"73745a5a",
           747 => x"5b8a7c33",
           748 => x"585a76fe",
           749 => x"dd38ff9e",
           750 => x"397c5276",
           751 => x"518baf3f",
           752 => x"7b335776",
           753 => x"fecc38ff",
           754 => x"8d397a83",
           755 => x"2a708106",
           756 => x"5455788a",
           757 => x"38817074",
           758 => x"0640547e",
           759 => x"9538e017",
           760 => x"537280d8",
           761 => x"26973872",
           762 => x"101083ca",
           763 => x"cc055473",
           764 => x"080473e0",
           765 => x"18545980",
           766 => x"d87327eb",
           767 => x"387c5276",
           768 => x"518aeb3f",
           769 => x"807c3358",
           770 => x"5b76fe86",
           771 => x"38fec739",
           772 => x"80ff59fe",
           773 => x"f639885a",
           774 => x"7f608405",
           775 => x"71087d83",
           776 => x"ffcf065e",
           777 => x"58415484",
           778 => x"ba9c5e79",
           779 => x"52755193",
           780 => x"9a3f84ba",
           781 => x"8c0881ff",
           782 => x"0684ba8c",
           783 => x"0818df05",
           784 => x"56537289",
           785 => x"26883884",
           786 => x"ba8c08b0",
           787 => x"0555747e",
           788 => x"70810540",
           789 => x"34795275",
           790 => x"5190ca3f",
           791 => x"84ba8c08",
           792 => x"5684ba8c",
           793 => x"08c5387d",
           794 => x"84ba9c31",
           795 => x"982b7bb2",
           796 => x"0640567e",
           797 => x"802e8f38",
           798 => x"77848080",
           799 => x"29fc8080",
           800 => x"0570902c",
           801 => x"59557a86",
           802 => x"2a708106",
           803 => x"555f7380",
           804 => x"2e9e3877",
           805 => x"84808029",
           806 => x"f8808005",
           807 => x"5379902e",
           808 => x"8b387784",
           809 => x"808029fc",
           810 => x"80800553",
           811 => x"72902c58",
           812 => x"7a832a70",
           813 => x"81065455",
           814 => x"72802e9e",
           815 => x"3875982c",
           816 => x"7081ff06",
           817 => x"54547873",
           818 => x"2486cc38",
           819 => x"7a83fff7",
           820 => x"0670832a",
           821 => x"71862a41",
           822 => x"565b7481",
           823 => x"06547380",
           824 => x"2e85f038",
           825 => x"77793190",
           826 => x"2b70902c",
           827 => x"7c838006",
           828 => x"56595373",
           829 => x"802e8596",
           830 => x"387a812a",
           831 => x"81065473",
           832 => x"85eb387a",
           833 => x"842a8106",
           834 => x"54738698",
           835 => x"387a852a",
           836 => x"81065473",
           837 => x"8697387e",
           838 => x"81065473",
           839 => x"858f387a",
           840 => x"882a8106",
           841 => x"5f7e802e",
           842 => x"b2387778",
           843 => x"84808029",
           844 => x"fc808005",
           845 => x"70902c5a",
           846 => x"40548074",
           847 => x"259d387c",
           848 => x"52b05188",
           849 => x"a93f7778",
           850 => x"84808029",
           851 => x"fc808005",
           852 => x"70902c5a",
           853 => x"40547380",
           854 => x"24e53874",
           855 => x"81065372",
           856 => x"802eb238",
           857 => x"78798180",
           858 => x"0a2981ff",
           859 => x"0a057098",
           860 => x"2c5b5555",
           861 => x"8075259d",
           862 => x"387c52b0",
           863 => x"5187ef3f",
           864 => x"78798180",
           865 => x"0a2981ff",
           866 => x"0a057098",
           867 => x"2c5b5555",
           868 => x"748024e5",
           869 => x"387a872a",
           870 => x"7081065c",
           871 => x"557a802e",
           872 => x"81b93876",
           873 => x"80e32e84",
           874 => x"d8387680",
           875 => x"f32e81ca",
           876 => x"387680d3",
           877 => x"2e81e238",
           878 => x"7d84ba9c",
           879 => x"2e96387c",
           880 => x"52ff1e70",
           881 => x"33525e87",
           882 => x"a53f7d84",
           883 => x"ba9c2e09",
           884 => x"8106ec38",
           885 => x"7481065b",
           886 => x"7a802efc",
           887 => x"a7387778",
           888 => x"84808029",
           889 => x"fc808005",
           890 => x"70902c5a",
           891 => x"40558075",
           892 => x"25fc9138",
           893 => x"7c52a051",
           894 => x"86f43fe2",
           895 => x"397a9007",
           896 => x"5b7aa007",
           897 => x"7c33585b",
           898 => x"76fa8738",
           899 => x"fac8397a",
           900 => x"80c0075b",
           901 => x"80f85790",
           902 => x"60618405",
           903 => x"71087e83",
           904 => x"ffcf065f",
           905 => x"5942555a",
           906 => x"fbfd397f",
           907 => x"60840577",
           908 => x"fe800a06",
           909 => x"83133370",
           910 => x"982b7207",
           911 => x"7c848080",
           912 => x"29fc8080",
           913 => x"0570902c",
           914 => x"5e525a56",
           915 => x"57415f7a",
           916 => x"872a7081",
           917 => x"065c557a",
           918 => x"fec93877",
           919 => x"78848080",
           920 => x"29fc8080",
           921 => x"0570902c",
           922 => x"5a545f80",
           923 => x"7f25feb3",
           924 => x"387c52a0",
           925 => x"5185f73f",
           926 => x"e239ff1a",
           927 => x"7083ffff",
           928 => x"065b5779",
           929 => x"83ffff2e",
           930 => x"feca387c",
           931 => x"52757081",
           932 => x"05573351",
           933 => x"85d83fe2",
           934 => x"39ff1a70",
           935 => x"83ffff06",
           936 => x"5b547983",
           937 => x"ffff2efe",
           938 => x"ab387c52",
           939 => x"75708105",
           940 => x"57335185",
           941 => x"b93fe239",
           942 => x"75fc0a06",
           943 => x"81fc0a07",
           944 => x"78848080",
           945 => x"29fc8080",
           946 => x"0570902c",
           947 => x"5a585680",
           948 => x"e37b872a",
           949 => x"7081065d",
           950 => x"56577afd",
           951 => x"c638fefb",
           952 => x"397f6084",
           953 => x"05710870",
           954 => x"53404156",
           955 => x"807e2482",
           956 => x"df387a83",
           957 => x"ffbf065b",
           958 => x"84ba9c5e",
           959 => x"faad397a",
           960 => x"84077c33",
           961 => x"585b76f8",
           962 => x"8938f8ca",
           963 => x"397a8807",
           964 => x"5b807c33",
           965 => x"585976f7",
           966 => x"f938f8ba",
           967 => x"397f6084",
           968 => x"05710877",
           969 => x"81065658",
           970 => x"415f7282",
           971 => x"8a387551",
           972 => x"87f63f84",
           973 => x"ba8c0883",
           974 => x"ffff0678",
           975 => x"7131902b",
           976 => x"545a7290",
           977 => x"2c58fe87",
           978 => x"397a80c0",
           979 => x"077c3358",
           980 => x"5b76f7be",
           981 => x"38f7ff39",
           982 => x"7f608405",
           983 => x"71087781",
           984 => x"065d5841",
           985 => x"547981cf",
           986 => x"38755187",
           987 => x"bb3f84ba",
           988 => x"8c0883ff",
           989 => x"ff067871",
           990 => x"31902b54",
           991 => x"5ac4397a",
           992 => x"8180077c",
           993 => x"33585b76",
           994 => x"f78838f7",
           995 => x"c9397778",
           996 => x"84808029",
           997 => x"fc808005",
           998 => x"70902c5a",
           999 => x"54548074",
          1000 => x"25fad638",
          1001 => x"7c52a051",
          1002 => x"83c43fe2",
          1003 => x"397c52b0",
          1004 => x"5183bb3f",
          1005 => x"79902e09",
          1006 => x"8106fae3",
          1007 => x"387c5276",
          1008 => x"5183ab3f",
          1009 => x"7a882a81",
          1010 => x"065f7e80",
          1011 => x"2efb8c38",
          1012 => x"fad83975",
          1013 => x"982c7871",
          1014 => x"31902b70",
          1015 => x"902c7d83",
          1016 => x"8006575a",
          1017 => x"515373fa",
          1018 => x"9038ffa2",
          1019 => x"397c52ad",
          1020 => x"5182fb3f",
          1021 => x"7e810654",
          1022 => x"73802efa",
          1023 => x"a238ffad",
          1024 => x"397c5275",
          1025 => x"982a5182",
          1026 => x"e53f7481",
          1027 => x"065b7a80",
          1028 => x"2ef7f138",
          1029 => x"fbc83978",
          1030 => x"7431982b",
          1031 => x"70982c5a",
          1032 => x"53f9b739",
          1033 => x"7c52ab51",
          1034 => x"82c43fc8",
          1035 => x"397c52a0",
          1036 => x"5182bb3f",
          1037 => x"ffbe3978",
          1038 => x"52755188",
          1039 => x"8b3f84ba",
          1040 => x"8c0883ff",
          1041 => x"ff067871",
          1042 => x"31902b54",
          1043 => x"5afdf339",
          1044 => x"7a82077e",
          1045 => x"307183ff",
          1046 => x"bf065257",
          1047 => x"5bfd9939",
          1048 => x"fe3d0d84",
          1049 => x"d5ec0853",
          1050 => x"75527451",
          1051 => x"f3b53f84",
          1052 => x"3d0d04fa",
          1053 => x"3d0d7855",
          1054 => x"800b84d5",
          1055 => x"f0088511",
          1056 => x"3370812a",
          1057 => x"81327081",
          1058 => x"06515658",
          1059 => x"5557ff56",
          1060 => x"72772e09",
          1061 => x"810680d5",
          1062 => x"38747081",
          1063 => x"05563353",
          1064 => x"72772eb0",
          1065 => x"3884d5f0",
          1066 => x"08527251",
          1067 => x"90140853",
          1068 => x"722d84ba",
          1069 => x"8c08802e",
          1070 => x"8338ff57",
          1071 => x"74708105",
          1072 => x"56335372",
          1073 => x"802e8838",
          1074 => x"84d5f008",
          1075 => x"54d73984",
          1076 => x"d5f00854",
          1077 => x"84d5f008",
          1078 => x"528a5190",
          1079 => x"14085574",
          1080 => x"2d84ba8c",
          1081 => x"08802e83",
          1082 => x"38ff5776",
          1083 => x"567584ba",
          1084 => x"8c0c883d",
          1085 => x"0d04fa3d",
          1086 => x"0d787a56",
          1087 => x"54800b85",
          1088 => x"16337081",
          1089 => x"2a813270",
          1090 => x"81065155",
          1091 => x"5757ff56",
          1092 => x"72772e09",
          1093 => x"81069238",
          1094 => x"73708105",
          1095 => x"55335372",
          1096 => x"772e0981",
          1097 => x"06983876",
          1098 => x"567584ba",
          1099 => x"8c0c883d",
          1100 => x"0d047370",
          1101 => x"81055533",
          1102 => x"5372802e",
          1103 => x"ea387452",
          1104 => x"72519015",
          1105 => x"0853722d",
          1106 => x"84ba8c08",
          1107 => x"802ee338",
          1108 => x"ff747081",
          1109 => x"05563354",
          1110 => x"5772e338",
          1111 => x"ca39ff3d",
          1112 => x"0d84d5f0",
          1113 => x"08527351",
          1114 => x"853f833d",
          1115 => x"0d04fa3d",
          1116 => x"0d787a85",
          1117 => x"11337081",
          1118 => x"2a813281",
          1119 => x"06565656",
          1120 => x"57ff5672",
          1121 => x"ae387382",
          1122 => x"2a810654",
          1123 => x"73802eac",
          1124 => x"388c1508",
          1125 => x"53728816",
          1126 => x"08259138",
          1127 => x"74085676",
          1128 => x"76347408",
          1129 => x"8105750c",
          1130 => x"8c150853",
          1131 => x"81138c16",
          1132 => x"0c765675",
          1133 => x"84ba8c0c",
          1134 => x"883d0d04",
          1135 => x"74527681",
          1136 => x"ff065190",
          1137 => x"15085473",
          1138 => x"2dff5684",
          1139 => x"ba8c08e3",
          1140 => x"388c1508",
          1141 => x"81058c16",
          1142 => x"0c7656d7",
          1143 => x"39fb3d0d",
          1144 => x"77851133",
          1145 => x"7081ff06",
          1146 => x"70813281",
          1147 => x"06555556",
          1148 => x"56ff5471",
          1149 => x"b3387286",
          1150 => x"2a810652",
          1151 => x"71b33872",
          1152 => x"822a8106",
          1153 => x"5271802e",
          1154 => x"80c33875",
          1155 => x"08703353",
          1156 => x"5371802e",
          1157 => x"80f03881",
          1158 => x"13760c8c",
          1159 => x"16088105",
          1160 => x"8c170c71",
          1161 => x"81ff0654",
          1162 => x"7384ba8c",
          1163 => x"0c873d0d",
          1164 => x"0474ffbf",
          1165 => x"06537285",
          1166 => x"17348c16",
          1167 => x"0881058c",
          1168 => x"170c8416",
          1169 => x"3384ba8c",
          1170 => x"0c873d0d",
          1171 => x"04755194",
          1172 => x"16085574",
          1173 => x"2d84ba8c",
          1174 => x"085284ba",
          1175 => x"8c088025",
          1176 => x"ffb93885",
          1177 => x"16337090",
          1178 => x"07545284",
          1179 => x"ba8c08ff",
          1180 => x"2e853871",
          1181 => x"a0075372",
          1182 => x"851734ff",
          1183 => x"547384ba",
          1184 => x"8c0c873d",
          1185 => x"0d0474a0",
          1186 => x"07537285",
          1187 => x"1734ff54",
          1188 => x"ec39fd3d",
          1189 => x"0d757771",
          1190 => x"54545471",
          1191 => x"70810553",
          1192 => x"335170f7",
          1193 => x"38ff1252",
          1194 => x"72708105",
          1195 => x"54335170",
          1196 => x"72708105",
          1197 => x"543470f0",
          1198 => x"387384ba",
          1199 => x"8c0c853d",
          1200 => x"0d04fc3d",
          1201 => x"0d767971",
          1202 => x"7a555552",
          1203 => x"5470802e",
          1204 => x"9d387372",
          1205 => x"27a13870",
          1206 => x"802e9338",
          1207 => x"71708105",
          1208 => x"53337370",
          1209 => x"81055534",
          1210 => x"ff115170",
          1211 => x"ef387384",
          1212 => x"ba8c0c86",
          1213 => x"3d0d0470",
          1214 => x"12557375",
          1215 => x"27d93870",
          1216 => x"14755353",
          1217 => x"ff13ff13",
          1218 => x"53537133",
          1219 => x"7334ff11",
          1220 => x"5170802e",
          1221 => x"d938ff13",
          1222 => x"ff135353",
          1223 => x"71337334",
          1224 => x"ff115170",
          1225 => x"df38c739",
          1226 => x"fe3d0d74",
          1227 => x"70535371",
          1228 => x"70810553",
          1229 => x"335170f7",
          1230 => x"38ff1270",
          1231 => x"743184ba",
          1232 => x"8c0c5184",
          1233 => x"3d0d04fd",
          1234 => x"3d0d7577",
          1235 => x"71545454",
          1236 => x"72708105",
          1237 => x"54335170",
          1238 => x"72708105",
          1239 => x"543470f0",
          1240 => x"387384ba",
          1241 => x"8c0c853d",
          1242 => x"0d04fd3d",
          1243 => x"0d757871",
          1244 => x"79555552",
          1245 => x"5470802e",
          1246 => x"93387170",
          1247 => x"81055333",
          1248 => x"73708105",
          1249 => x"5534ff11",
          1250 => x"5170ef38",
          1251 => x"7384ba8c",
          1252 => x"0c853d0d",
          1253 => x"04fc3d0d",
          1254 => x"76787a55",
          1255 => x"56547280",
          1256 => x"2ea13873",
          1257 => x"33757081",
          1258 => x"05573352",
          1259 => x"5271712e",
          1260 => x"0981069a",
          1261 => x"38811454",
          1262 => x"71802eb7",
          1263 => x"38ff1353",
          1264 => x"72e13880",
          1265 => x"517084ba",
          1266 => x"8c0c863d",
          1267 => x"0d047280",
          1268 => x"2ef13873",
          1269 => x"3353ff51",
          1270 => x"72802ee9",
          1271 => x"38ff1533",
          1272 => x"52815171",
          1273 => x"802ede38",
          1274 => x"72723184",
          1275 => x"ba8c0c86",
          1276 => x"3d0d0471",
          1277 => x"84ba8c0c",
          1278 => x"863d0d04",
          1279 => x"fb3d0d77",
          1280 => x"79537052",
          1281 => x"5680c13f",
          1282 => x"84ba8c08",
          1283 => x"84ba8c08",
          1284 => x"81055255",
          1285 => x"81b3b33f",
          1286 => x"84ba8c08",
          1287 => x"5484ba8c",
          1288 => x"08802e9b",
          1289 => x"3884ba8c",
          1290 => x"08155480",
          1291 => x"74347453",
          1292 => x"755284ba",
          1293 => x"8c0851fe",
          1294 => x"b13f84ba",
          1295 => x"8c085473",
          1296 => x"84ba8c0c",
          1297 => x"873d0d04",
          1298 => x"fd3d0d75",
          1299 => x"77717154",
          1300 => x"55535471",
          1301 => x"802e9f38",
          1302 => x"72708105",
          1303 => x"54335170",
          1304 => x"802e8c38",
          1305 => x"ff125271",
          1306 => x"ff2e0981",
          1307 => x"06ea38ff",
          1308 => x"13707531",
          1309 => x"52527084",
          1310 => x"ba8c0c85",
          1311 => x"3d0d04fd",
          1312 => x"3d0d7577",
          1313 => x"79725553",
          1314 => x"54547080",
          1315 => x"2e8e3872",
          1316 => x"72708105",
          1317 => x"5434ff11",
          1318 => x"5170f438",
          1319 => x"7384ba8c",
          1320 => x"0c853d0d",
          1321 => x"04fa3d0d",
          1322 => x"787a5854",
          1323 => x"a0527680",
          1324 => x"2e8b3876",
          1325 => x"5180f53f",
          1326 => x"84ba8c08",
          1327 => x"52e01253",
          1328 => x"73802e8d",
          1329 => x"38735180",
          1330 => x"e33f7184",
          1331 => x"ba8c0831",
          1332 => x"53805272",
          1333 => x"9f2680cb",
          1334 => x"38735272",
          1335 => x"9f2e80c3",
          1336 => x"38811374",
          1337 => x"712aa072",
          1338 => x"3176712b",
          1339 => x"57545455",
          1340 => x"80567476",
          1341 => x"2ea83872",
          1342 => x"10749f2a",
          1343 => x"07741077",
          1344 => x"07787231",
          1345 => x"ff119f2c",
          1346 => x"7081067b",
          1347 => x"72067571",
          1348 => x"31ff1c5c",
          1349 => x"56525255",
          1350 => x"58555374",
          1351 => x"da387310",
          1352 => x"76075271",
          1353 => x"84ba8c0c",
          1354 => x"883d0d04",
          1355 => x"fc3d0d76",
          1356 => x"70fc8080",
          1357 => x"06703070",
          1358 => x"72078025",
          1359 => x"70842b90",
          1360 => x"71317571",
          1361 => x"2a7083fe",
          1362 => x"80067030",
          1363 => x"70802583",
          1364 => x"2b887131",
          1365 => x"74712a70",
          1366 => x"81f00670",
          1367 => x"30708025",
          1368 => x"822b8471",
          1369 => x"3174712a",
          1370 => x"5553751b",
          1371 => x"05738c06",
          1372 => x"70307080",
          1373 => x"25108271",
          1374 => x"3177712a",
          1375 => x"70812a81",
          1376 => x"32708106",
          1377 => x"70308274",
          1378 => x"31067519",
          1379 => x"0584ba8c",
          1380 => x"0c515254",
          1381 => x"55515456",
          1382 => x"5a535555",
          1383 => x"55515656",
          1384 => x"56565158",
          1385 => x"56545286",
          1386 => x"3d0d04fd",
          1387 => x"3d0d7577",
          1388 => x"70547153",
          1389 => x"54548194",
          1390 => x"3f84ba8c",
          1391 => x"08732974",
          1392 => x"713184ba",
          1393 => x"8c0c5385",
          1394 => x"3d0d04fa",
          1395 => x"3d0d787a",
          1396 => x"5854a053",
          1397 => x"76802e8b",
          1398 => x"387651fe",
          1399 => x"cf3f84ba",
          1400 => x"8c0853e0",
          1401 => x"13527380",
          1402 => x"2e8d3873",
          1403 => x"51febd3f",
          1404 => x"7284ba8c",
          1405 => x"08315273",
          1406 => x"53719f26",
          1407 => x"80c53880",
          1408 => x"53719f2e",
          1409 => x"be388112",
          1410 => x"74712aa0",
          1411 => x"72317671",
          1412 => x"2b575454",
          1413 => x"55805674",
          1414 => x"762ea838",
          1415 => x"7210749f",
          1416 => x"2a077410",
          1417 => x"77077872",
          1418 => x"31ff119f",
          1419 => x"2c708106",
          1420 => x"7b720675",
          1421 => x"7131ff1c",
          1422 => x"5c565252",
          1423 => x"55585553",
          1424 => x"74da3872",
          1425 => x"84ba8c0c",
          1426 => x"883d0d04",
          1427 => x"fa3d0d78",
          1428 => x"9f2c7a9f",
          1429 => x"2c7a9f2c",
          1430 => x"7b327c9f",
          1431 => x"2c7d3273",
          1432 => x"73327174",
          1433 => x"31577275",
          1434 => x"31565956",
          1435 => x"595556fc",
          1436 => x"b43f84ba",
          1437 => x"8c087532",
          1438 => x"753184ba",
          1439 => x"8c0c883d",
          1440 => x"0d04f73d",
          1441 => x"0d7b7d5b",
          1442 => x"5780707b",
          1443 => x"0c770870",
          1444 => x"33565659",
          1445 => x"73a02e09",
          1446 => x"81068f38",
          1447 => x"81157078",
          1448 => x"0c703355",
          1449 => x"5573a02e",
          1450 => x"f33873ad",
          1451 => x"2e80f538",
          1452 => x"73b02e81",
          1453 => x"8338d014",
          1454 => x"58805677",
          1455 => x"892680db",
          1456 => x"388a5880",
          1457 => x"56a07427",
          1458 => x"80c43880",
          1459 => x"e0742789",
          1460 => x"38e01470",
          1461 => x"81ff0655",
          1462 => x"53d01470",
          1463 => x"81ff0651",
          1464 => x"53907327",
          1465 => x"8f38f913",
          1466 => x"7081ff06",
          1467 => x"54548973",
          1468 => x"27818938",
          1469 => x"72782781",
          1470 => x"83387776",
          1471 => x"29138116",
          1472 => x"70790c70",
          1473 => x"33565656",
          1474 => x"73a026ff",
          1475 => x"be387880",
          1476 => x"2e843875",
          1477 => x"3056757a",
          1478 => x"0c815675",
          1479 => x"84ba8c0c",
          1480 => x"8b3d0d04",
          1481 => x"81701670",
          1482 => x"790c7033",
          1483 => x"56565973",
          1484 => x"b02e0981",
          1485 => x"06feff38",
          1486 => x"81157078",
          1487 => x"0c703355",
          1488 => x"557380e2",
          1489 => x"2ea63890",
          1490 => x"587380f8",
          1491 => x"2ea03881",
          1492 => x"56a07427",
          1493 => x"c638d014",
          1494 => x"53805688",
          1495 => x"58897327",
          1496 => x"fee13875",
          1497 => x"84ba8c0c",
          1498 => x"8b3d0d04",
          1499 => x"82588115",
          1500 => x"70780c70",
          1501 => x"33555580",
          1502 => x"56feca39",
          1503 => x"800b84ba",
          1504 => x"8c0c8b3d",
          1505 => x"0d04f73d",
          1506 => x"0d7b7d5b",
          1507 => x"5780707b",
          1508 => x"0c770870",
          1509 => x"33565659",
          1510 => x"73a02e09",
          1511 => x"81068f38",
          1512 => x"81157078",
          1513 => x"0c703355",
          1514 => x"5573a02e",
          1515 => x"f33873ad",
          1516 => x"2e80f538",
          1517 => x"73b02e81",
          1518 => x"8338d014",
          1519 => x"58805677",
          1520 => x"892680db",
          1521 => x"388a5880",
          1522 => x"56a07427",
          1523 => x"80c43880",
          1524 => x"e0742789",
          1525 => x"38e01470",
          1526 => x"81ff0655",
          1527 => x"53d01470",
          1528 => x"81ff0651",
          1529 => x"53907327",
          1530 => x"8f38f913",
          1531 => x"7081ff06",
          1532 => x"54548973",
          1533 => x"27818938",
          1534 => x"72782781",
          1535 => x"83387776",
          1536 => x"29138116",
          1537 => x"70790c70",
          1538 => x"33565656",
          1539 => x"73a026ff",
          1540 => x"be387880",
          1541 => x"2e843875",
          1542 => x"3056757a",
          1543 => x"0c815675",
          1544 => x"84ba8c0c",
          1545 => x"8b3d0d04",
          1546 => x"81701670",
          1547 => x"790c7033",
          1548 => x"56565973",
          1549 => x"b02e0981",
          1550 => x"06feff38",
          1551 => x"81157078",
          1552 => x"0c703355",
          1553 => x"557380e2",
          1554 => x"2ea63890",
          1555 => x"587380f8",
          1556 => x"2ea03881",
          1557 => x"56a07427",
          1558 => x"c638d014",
          1559 => x"53805688",
          1560 => x"58897327",
          1561 => x"fee13875",
          1562 => x"84ba8c0c",
          1563 => x"8b3d0d04",
          1564 => x"82588115",
          1565 => x"70780c70",
          1566 => x"33555580",
          1567 => x"56feca39",
          1568 => x"800b84ba",
          1569 => x"8c0c8b3d",
          1570 => x"0d0480d6",
          1571 => x"dc3f84ba",
          1572 => x"8c0881ff",
          1573 => x"0684ba8c",
          1574 => x"0c04ff3d",
          1575 => x"0d735271",
          1576 => x"93268c38",
          1577 => x"71101083",
          1578 => x"becc0552",
          1579 => x"71080483",
          1580 => x"cee451ef",
          1581 => x"be3f833d",
          1582 => x"0d0483ce",
          1583 => x"f451efb3",
          1584 => x"3f833d0d",
          1585 => x"0483cf8c",
          1586 => x"51efa83f",
          1587 => x"833d0d04",
          1588 => x"83cfa451",
          1589 => x"ef9d3f83",
          1590 => x"3d0d0483",
          1591 => x"cfbc51ef",
          1592 => x"923f833d",
          1593 => x"0d0483cf",
          1594 => x"cc51ef87",
          1595 => x"3f833d0d",
          1596 => x"0483cfec",
          1597 => x"51eefc3f",
          1598 => x"833d0d04",
          1599 => x"83cffc51",
          1600 => x"eef13f83",
          1601 => x"3d0d0483",
          1602 => x"d0a451ee",
          1603 => x"e63f833d",
          1604 => x"0d0483d0",
          1605 => x"b851eedb",
          1606 => x"3f833d0d",
          1607 => x"0483d0d4",
          1608 => x"51eed03f",
          1609 => x"833d0d04",
          1610 => x"83d0ec51",
          1611 => x"eec53f83",
          1612 => x"3d0d0483",
          1613 => x"d18451ee",
          1614 => x"ba3f833d",
          1615 => x"0d0483d1",
          1616 => x"9c51eeaf",
          1617 => x"3f833d0d",
          1618 => x"0483d1ac",
          1619 => x"51eea43f",
          1620 => x"833d0d04",
          1621 => x"83d1c051",
          1622 => x"ee993f83",
          1623 => x"3d0d0483",
          1624 => x"d1d051ee",
          1625 => x"8e3f833d",
          1626 => x"0d0483d1",
          1627 => x"e051ee83",
          1628 => x"3f833d0d",
          1629 => x"0483d1f0",
          1630 => x"51edf83f",
          1631 => x"833d0d04",
          1632 => x"83d28051",
          1633 => x"eded3f83",
          1634 => x"3d0d0483",
          1635 => x"d28c51ed",
          1636 => x"e23f833d",
          1637 => x"0d04ec3d",
          1638 => x"0d660284",
          1639 => x"0580e305",
          1640 => x"335b5880",
          1641 => x"68793070",
          1642 => x"7b077325",
          1643 => x"51575759",
          1644 => x"78577587",
          1645 => x"ff268338",
          1646 => x"81577477",
          1647 => x"077081ff",
          1648 => x"06515593",
          1649 => x"577480e2",
          1650 => x"38815377",
          1651 => x"528c3d70",
          1652 => x"52588296",
          1653 => x"a23f84ba",
          1654 => x"8c085784",
          1655 => x"ba8c0880",
          1656 => x"2e80d038",
          1657 => x"775182af",
          1658 => x"e03f7630",
          1659 => x"70780780",
          1660 => x"257b3070",
          1661 => x"9f2a7206",
          1662 => x"53575758",
          1663 => x"77802eaa",
          1664 => x"3887c098",
          1665 => x"88085574",
          1666 => x"87e72680",
          1667 => x"e0387452",
          1668 => x"7887e829",
          1669 => x"51f58e3f",
          1670 => x"84ba8c08",
          1671 => x"5483d2bc",
          1672 => x"53785283",
          1673 => x"d29851df",
          1674 => x"df3f7684",
          1675 => x"ba8c0c96",
          1676 => x"3d0d0484",
          1677 => x"ba8c0887",
          1678 => x"c098880c",
          1679 => x"84ba8c08",
          1680 => x"59963dd4",
          1681 => x"05548480",
          1682 => x"53755277",
          1683 => x"51829e97",
          1684 => x"3f84ba8c",
          1685 => x"085784ba",
          1686 => x"8c08ff88",
          1687 => x"387a5574",
          1688 => x"802eff80",
          1689 => x"38741975",
          1690 => x"175759d5",
          1691 => x"3987e852",
          1692 => x"7451f4b1",
          1693 => x"3f84ba8c",
          1694 => x"08527851",
          1695 => x"f4a73f84",
          1696 => x"ba8c0854",
          1697 => x"83d2bc53",
          1698 => x"785283d2",
          1699 => x"9851def8",
          1700 => x"3fff9739",
          1701 => x"f83d0d7c",
          1702 => x"028405b7",
          1703 => x"05335859",
          1704 => x"ff588053",
          1705 => x"7b527a51",
          1706 => x"fdec3f84",
          1707 => x"ba8c088b",
          1708 => x"3876802e",
          1709 => x"91387681",
          1710 => x"2e8a3877",
          1711 => x"84ba8c0c",
          1712 => x"8a3d0d04",
          1713 => x"780484d5",
          1714 => x"ec566155",
          1715 => x"605484ba",
          1716 => x"8c537f52",
          1717 => x"7e51782d",
          1718 => x"84ba8c08",
          1719 => x"84ba8c0c",
          1720 => x"8a3d0d04",
          1721 => x"f33d0d7f",
          1722 => x"6163028c",
          1723 => x"0580cf05",
          1724 => x"33737315",
          1725 => x"68415f5c",
          1726 => x"5c5f5d5e",
          1727 => x"78802e83",
          1728 => x"82387a52",
          1729 => x"83d2c451",
          1730 => x"ddfe3f83",
          1731 => x"d2cc51dd",
          1732 => x"f73f8054",
          1733 => x"737927b2",
          1734 => x"387c902e",
          1735 => x"81ed387c",
          1736 => x"a02e82a8",
          1737 => x"38731853",
          1738 => x"727a2781",
          1739 => x"a7387233",
          1740 => x"5283d2d0",
          1741 => x"51ddd13f",
          1742 => x"811484d5",
          1743 => x"f0085354",
          1744 => x"a051ecaa",
          1745 => x"3f787426",
          1746 => x"dc3883d2",
          1747 => x"d851ddb8",
          1748 => x"3f805675",
          1749 => x"792780c0",
          1750 => x"38751870",
          1751 => x"33555380",
          1752 => x"55727a27",
          1753 => x"83388155",
          1754 => x"80539f74",
          1755 => x"27833881",
          1756 => x"53747306",
          1757 => x"7081ff06",
          1758 => x"56577480",
          1759 => x"2e883880",
          1760 => x"fe742781",
          1761 => x"ee3884d5",
          1762 => x"f00852a0",
          1763 => x"51ebdf3f",
          1764 => x"81165678",
          1765 => x"7626c238",
          1766 => x"83d2dc51",
          1767 => x"e9d53f78",
          1768 => x"18791c5c",
          1769 => x"5880519d",
          1770 => x"b23f84ba",
          1771 => x"8c08982b",
          1772 => x"70982c58",
          1773 => x"5476a02e",
          1774 => x"81ee3876",
          1775 => x"9b2e82c3",
          1776 => x"387b1e57",
          1777 => x"767826fe",
          1778 => x"b938ff0b",
          1779 => x"84ba8c0c",
          1780 => x"8f3d0d04",
          1781 => x"83d2e051",
          1782 => x"dcae3f81",
          1783 => x"1484d5f0",
          1784 => x"085354a0",
          1785 => x"51eb873f",
          1786 => x"787426fe",
          1787 => x"b838feda",
          1788 => x"3983d2f0",
          1789 => x"51dc913f",
          1790 => x"821484d5",
          1791 => x"f0085354",
          1792 => x"a051eaea",
          1793 => x"3f737927",
          1794 => x"fec03873",
          1795 => x"1853727a",
          1796 => x"27df3872",
          1797 => x"225283d2",
          1798 => x"e451dbec",
          1799 => x"3f821484",
          1800 => x"d5f00853",
          1801 => x"54a051ea",
          1802 => x"c53f7874",
          1803 => x"26dd38fe",
          1804 => x"993983d2",
          1805 => x"ec51dbd0",
          1806 => x"3f841484",
          1807 => x"d5f00853",
          1808 => x"54a051ea",
          1809 => x"a93f7379",
          1810 => x"27fdff38",
          1811 => x"73185372",
          1812 => x"7a27df38",
          1813 => x"72085283",
          1814 => x"d2c451db",
          1815 => x"ab3f8414",
          1816 => x"84d5f008",
          1817 => x"5354a051",
          1818 => x"ea843f78",
          1819 => x"7426dd38",
          1820 => x"fdd83984",
          1821 => x"d5f00852",
          1822 => x"7351e9f2",
          1823 => x"3f811656",
          1824 => x"fe913980",
          1825 => x"cee33f84",
          1826 => x"ba8c0881",
          1827 => x"ff065388",
          1828 => x"5972a82e",
          1829 => x"fcec38a0",
          1830 => x"597280d0",
          1831 => x"2e098106",
          1832 => x"fce03890",
          1833 => x"59fcdb39",
          1834 => x"80519baf",
          1835 => x"3f84ba8c",
          1836 => x"08982b70",
          1837 => x"982c70a0",
          1838 => x"32703072",
          1839 => x"9b327030",
          1840 => x"70720773",
          1841 => x"75070651",
          1842 => x"55585957",
          1843 => x"58537280",
          1844 => x"25fde838",
          1845 => x"80519b83",
          1846 => x"3f84ba8c",
          1847 => x"08982b70",
          1848 => x"982c70a0",
          1849 => x"32703072",
          1850 => x"9b327030",
          1851 => x"70720773",
          1852 => x"75070651",
          1853 => x"55585957",
          1854 => x"58538073",
          1855 => x"24ffa938",
          1856 => x"fdb93980",
          1857 => x"0b84ba8c",
          1858 => x"0c8f3d0d",
          1859 => x"04fe3d0d",
          1860 => x"87c09680",
          1861 => x"0853aad1",
          1862 => x"3f81519c",
          1863 => x"f73f83d3",
          1864 => x"b4519d88",
          1865 => x"3f80519c",
          1866 => x"eb3f7281",
          1867 => x"2a708106",
          1868 => x"51527182",
          1869 => x"b7387282",
          1870 => x"2a708106",
          1871 => x"51527182",
          1872 => x"89387283",
          1873 => x"2a708106",
          1874 => x"51527181",
          1875 => x"db387284",
          1876 => x"2a708106",
          1877 => x"51527181",
          1878 => x"ad387285",
          1879 => x"2a708106",
          1880 => x"51527180",
          1881 => x"ff387286",
          1882 => x"2a708106",
          1883 => x"51527180",
          1884 => x"d2387287",
          1885 => x"2a708106",
          1886 => x"515271a9",
          1887 => x"3872882a",
          1888 => x"81065372",
          1889 => x"8838a9e9",
          1890 => x"3f843d0d",
          1891 => x"0481519c",
          1892 => x"833f83d3",
          1893 => x"cc519c94",
          1894 => x"3f80519b",
          1895 => x"f73fa9d1",
          1896 => x"3f843d0d",
          1897 => x"0481519b",
          1898 => x"eb3f83d3",
          1899 => x"e0519bfc",
          1900 => x"3f80519b",
          1901 => x"df3f7288",
          1902 => x"2a810653",
          1903 => x"72802ec6",
          1904 => x"38cb3981",
          1905 => x"519bcd3f",
          1906 => x"83d3f451",
          1907 => x"9bde3f80",
          1908 => x"519bc13f",
          1909 => x"72872a70",
          1910 => x"81065152",
          1911 => x"71802eff",
          1912 => x"9c38c239",
          1913 => x"81519bac",
          1914 => x"3f83d488",
          1915 => x"519bbd3f",
          1916 => x"80519ba0",
          1917 => x"3f72862a",
          1918 => x"70810651",
          1919 => x"5271802e",
          1920 => x"fef038ff",
          1921 => x"be398151",
          1922 => x"9b8a3f83",
          1923 => x"d49c519b",
          1924 => x"9b3f8051",
          1925 => x"9afe3f72",
          1926 => x"852a7081",
          1927 => x"06515271",
          1928 => x"802efec2",
          1929 => x"38ffbd39",
          1930 => x"81519ae8",
          1931 => x"3f83d4b0",
          1932 => x"519af93f",
          1933 => x"80519adc",
          1934 => x"3f72842a",
          1935 => x"70810651",
          1936 => x"5271802e",
          1937 => x"fe9438ff",
          1938 => x"bd398151",
          1939 => x"9ac63f83",
          1940 => x"d4c4519a",
          1941 => x"d73f8051",
          1942 => x"9aba3f72",
          1943 => x"832a7081",
          1944 => x"06515271",
          1945 => x"802efde6",
          1946 => x"38ffbd39",
          1947 => x"81519aa4",
          1948 => x"3f83d4d4",
          1949 => x"519ab53f",
          1950 => x"80519a98",
          1951 => x"3f72822a",
          1952 => x"70810651",
          1953 => x"5271802e",
          1954 => x"fdb838ff",
          1955 => x"bd39ca3d",
          1956 => x"0d807041",
          1957 => x"41ff6184",
          1958 => x"d1980c42",
          1959 => x"81526051",
          1960 => x"81b6d53f",
          1961 => x"84ba8c08",
          1962 => x"81ff069b",
          1963 => x"3d405978",
          1964 => x"612e84b1",
          1965 => x"3883d5a8",
          1966 => x"51e3b83f",
          1967 => x"983d4383",
          1968 => x"d5e051d6",
          1969 => x"c33f7e48",
          1970 => x"80f85380",
          1971 => x"527e51eb",
          1972 => x"ae3f0b0b",
          1973 => x"83ef8033",
          1974 => x"7081ff06",
          1975 => x"5b597980",
          1976 => x"2e82f138",
          1977 => x"79812e83",
          1978 => x"88387881",
          1979 => x"ff065e7d",
          1980 => x"822e83c1",
          1981 => x"3867705a",
          1982 => x"5a79802e",
          1983 => x"83dc3879",
          1984 => x"335c7ba0",
          1985 => x"2e098106",
          1986 => x"8c38811a",
          1987 => x"70335d5a",
          1988 => x"7ba02ef6",
          1989 => x"38805c7b",
          1990 => x"9b26be38",
          1991 => x"7b902983",
          1992 => x"ef840570",
          1993 => x"08525be7",
          1994 => x"ff3f84ba",
          1995 => x"8c0884ba",
          1996 => x"8c08547a",
          1997 => x"537b0852",
          1998 => x"5de8da3f",
          1999 => x"84ba8c08",
          2000 => x"8b38841b",
          2001 => x"335e7d81",
          2002 => x"2e838038",
          2003 => x"811c7081",
          2004 => x"ff065d5b",
          2005 => x"9b7c27c4",
          2006 => x"389a3d33",
          2007 => x"5c7b802e",
          2008 => x"fedd3880",
          2009 => x"f8527e51",
          2010 => x"e9923f84",
          2011 => x"ba8c085e",
          2012 => x"84ba8c08",
          2013 => x"802e8dd3",
          2014 => x"3884ba8c",
          2015 => x"0848b83d",
          2016 => x"ff800551",
          2017 => x"91933f84",
          2018 => x"ba8c0860",
          2019 => x"62065c5c",
          2020 => x"7a802e81",
          2021 => x"843884ba",
          2022 => x"8c0851e7",
          2023 => x"8b3f84ba",
          2024 => x"8c088f26",
          2025 => x"80f33881",
          2026 => x"0ba53d5e",
          2027 => x"5b7a822e",
          2028 => x"8d8f387a",
          2029 => x"82248cec",
          2030 => x"387a812e",
          2031 => x"82ee387b",
          2032 => x"54805383",
          2033 => x"d5e4527c",
          2034 => x"51d5dd3f",
          2035 => x"83f2c858",
          2036 => x"84babc57",
          2037 => x"7d566755",
          2038 => x"80549080",
          2039 => x"0a539080",
          2040 => x"0a527c51",
          2041 => x"f5ae3f84",
          2042 => x"ba8c0884",
          2043 => x"ba8c0809",
          2044 => x"70307072",
          2045 => x"07802551",
          2046 => x"5b5b4280",
          2047 => x"5a7a8326",
          2048 => x"8338815a",
          2049 => x"787a0659",
          2050 => x"78802e8d",
          2051 => x"38811b70",
          2052 => x"81ff065c",
          2053 => x"5a7aff95",
          2054 => x"387f8132",
          2055 => x"61813207",
          2056 => x"5d7c81f8",
          2057 => x"3861ff2e",
          2058 => x"81f2387d",
          2059 => x"518195aa",
          2060 => x"3f83d5e0",
          2061 => x"51d3d13f",
          2062 => x"7e4880f8",
          2063 => x"5380527e",
          2064 => x"51e8bc3f",
          2065 => x"0b0b83ef",
          2066 => x"80337081",
          2067 => x"ff065b59",
          2068 => x"79fd9138",
          2069 => x"815383d5",
          2070 => x"8c5284d1",
          2071 => x"9c518289",
          2072 => x"963f84ba",
          2073 => x"8c0880c5",
          2074 => x"38810b0b",
          2075 => x"0b83ef80",
          2076 => x"3484d19c",
          2077 => x"5380f852",
          2078 => x"7e5182f7",
          2079 => x"913f84ba",
          2080 => x"8c08802e",
          2081 => x"a03884ba",
          2082 => x"8c0851df",
          2083 => x"e63f0b0b",
          2084 => x"83ef8033",
          2085 => x"7081ff06",
          2086 => x"5f597d82",
          2087 => x"2e098106",
          2088 => x"fcd33891",
          2089 => x"3984d19c",
          2090 => x"5182a29d",
          2091 => x"3f820b0b",
          2092 => x"0b83ef80",
          2093 => x"3483d59c",
          2094 => x"5380f852",
          2095 => x"7e51a7ce",
          2096 => x"3f67705a",
          2097 => x"5a79fcb7",
          2098 => x"3890397c",
          2099 => x"1a630c85",
          2100 => x"1b335978",
          2101 => x"818926fd",
          2102 => x"80387810",
          2103 => x"1083bf9c",
          2104 => x"055a7908",
          2105 => x"0483d5ec",
          2106 => x"51df883f",
          2107 => x"9a3d5f83",
          2108 => x"5383d680",
          2109 => x"527e51e4",
          2110 => x"f13f6053",
          2111 => x"7e5284bb",
          2112 => x"b8518285",
          2113 => x"c33f84ba",
          2114 => x"8c08612e",
          2115 => x"098106fb",
          2116 => x"a4388170",
          2117 => x"9a3d4541",
          2118 => x"41fba439",
          2119 => x"83d68451",
          2120 => x"ded13f7d",
          2121 => x"518193b2",
          2122 => x"3ffe8639",
          2123 => x"83d69456",
          2124 => x"7b5583d6",
          2125 => x"98548053",
          2126 => x"83d69c52",
          2127 => x"7c51d2e8",
          2128 => x"3ffd8939",
          2129 => x"818ce33f",
          2130 => x"faf5399a",
          2131 => x"dd3ffaef",
          2132 => x"39815283",
          2133 => x"51bf943f",
          2134 => x"fae53981",
          2135 => x"8e953ffa",
          2136 => x"de3983d6",
          2137 => x"ac51de8b",
          2138 => x"3f805978",
          2139 => x"0483d6c0",
          2140 => x"51de803f",
          2141 => x"d0f33ffa",
          2142 => x"c639b83d",
          2143 => x"ff841153",
          2144 => x"ff800551",
          2145 => x"ec803f84",
          2146 => x"ba8c0880",
          2147 => x"2efab038",
          2148 => x"685283d6",
          2149 => x"dc51d0f0",
          2150 => x"3f685a79",
          2151 => x"2d84ba8c",
          2152 => x"08802efa",
          2153 => x"9a3884ba",
          2154 => x"8c085283",
          2155 => x"d6f851d0",
          2156 => x"d73ffa8b",
          2157 => x"39b83dff",
          2158 => x"841153ff",
          2159 => x"800551eb",
          2160 => x"c53f84ba",
          2161 => x"8c08802e",
          2162 => x"f9f53868",
          2163 => x"5283d794",
          2164 => x"51d0b53f",
          2165 => x"68597804",
          2166 => x"b83dfef4",
          2167 => x"1153ff80",
          2168 => x"0551e99e",
          2169 => x"3f84ba8c",
          2170 => x"08802ef9",
          2171 => x"d238b83d",
          2172 => x"fef01153",
          2173 => x"ff800551",
          2174 => x"e9883f84",
          2175 => x"ba8c0886",
          2176 => x"d0386459",
          2177 => x"78085378",
          2178 => x"5283d7b0",
          2179 => x"51cff93f",
          2180 => x"84d5ec08",
          2181 => x"5380f852",
          2182 => x"7e51d087",
          2183 => x"3f7e487e",
          2184 => x"335978ae",
          2185 => x"2ef99838",
          2186 => x"789f2687",
          2187 => x"d3386484",
          2188 => x"05704659",
          2189 => x"cf39b83d",
          2190 => x"fef41153",
          2191 => x"ff800551",
          2192 => x"e8c03f84",
          2193 => x"ba8c0880",
          2194 => x"2ef8f438",
          2195 => x"b83dfef0",
          2196 => x"1153ff80",
          2197 => x"0551e8aa",
          2198 => x"3f84ba8c",
          2199 => x"0886b038",
          2200 => x"64597822",
          2201 => x"53785283",
          2202 => x"d7c051cf",
          2203 => x"9b3f84d5",
          2204 => x"ec085380",
          2205 => x"f8527e51",
          2206 => x"cfa93f7e",
          2207 => x"487e3359",
          2208 => x"78ae2ef8",
          2209 => x"ba38789f",
          2210 => x"2687ca38",
          2211 => x"64820570",
          2212 => x"4659cf39",
          2213 => x"b83dff84",
          2214 => x"1153ff80",
          2215 => x"0551e9e6",
          2216 => x"3f84ba8c",
          2217 => x"08802ef8",
          2218 => x"9638b83d",
          2219 => x"fefc1153",
          2220 => x"ff800551",
          2221 => x"e9d03f84",
          2222 => x"ba8c0880",
          2223 => x"2ef88038",
          2224 => x"b83dfef8",
          2225 => x"1153ff80",
          2226 => x"0551e9ba",
          2227 => x"3f84ba8c",
          2228 => x"08802ef7",
          2229 => x"ea3883d7",
          2230 => x"cc51ceac",
          2231 => x"3f68675d",
          2232 => x"59787c27",
          2233 => x"838d3865",
          2234 => x"70337a33",
          2235 => x"5f5c5a7a",
          2236 => x"7d2e9538",
          2237 => x"7a557954",
          2238 => x"78335378",
          2239 => x"5283d7dc",
          2240 => x"51ce853f",
          2241 => x"66665b5c",
          2242 => x"8119811b",
          2243 => x"4759d239",
          2244 => x"b83dff84",
          2245 => x"1153ff80",
          2246 => x"0551e8ea",
          2247 => x"3f84ba8c",
          2248 => x"08802ef7",
          2249 => x"9a38b83d",
          2250 => x"fefc1153",
          2251 => x"ff800551",
          2252 => x"e8d43f84",
          2253 => x"ba8c0880",
          2254 => x"2ef78438",
          2255 => x"b83dfef8",
          2256 => x"1153ff80",
          2257 => x"0551e8be",
          2258 => x"3f84ba8c",
          2259 => x"08802ef6",
          2260 => x"ee3883d7",
          2261 => x"f851cdb0",
          2262 => x"3f685a79",
          2263 => x"67278293",
          2264 => x"38655c79",
          2265 => x"7081055b",
          2266 => x"337c3465",
          2267 => x"810546eb",
          2268 => x"39b83dff",
          2269 => x"841153ff",
          2270 => x"800551e8",
          2271 => x"893f84ba",
          2272 => x"8c08802e",
          2273 => x"f6b938b8",
          2274 => x"3dfefc11",
          2275 => x"53ff8005",
          2276 => x"51e7f33f",
          2277 => x"84ba8c08",
          2278 => x"b1386870",
          2279 => x"33545283",
          2280 => x"d88451cc",
          2281 => x"e33f84d5",
          2282 => x"ec085380",
          2283 => x"f8527e51",
          2284 => x"ccf13f7e",
          2285 => x"487e3359",
          2286 => x"78ae2ef6",
          2287 => x"8238789f",
          2288 => x"26849738",
          2289 => x"68810549",
          2290 => x"d1396859",
          2291 => x"0280db05",
          2292 => x"33793468",
          2293 => x"810549b8",
          2294 => x"3dfefc11",
          2295 => x"53ff8005",
          2296 => x"51e7a33f",
          2297 => x"84ba8c08",
          2298 => x"802ef5d3",
          2299 => x"38685902",
          2300 => x"80db0533",
          2301 => x"79346881",
          2302 => x"0549b83d",
          2303 => x"fefc1153",
          2304 => x"ff800551",
          2305 => x"e7803f84",
          2306 => x"ba8c08ff",
          2307 => x"bd38f5af",
          2308 => x"39b83dff",
          2309 => x"841153ff",
          2310 => x"800551e6",
          2311 => x"e93f84ba",
          2312 => x"8c08802e",
          2313 => x"f59938b8",
          2314 => x"3dfefc11",
          2315 => x"53ff8005",
          2316 => x"51e6d33f",
          2317 => x"84ba8c08",
          2318 => x"802ef583",
          2319 => x"38b83dfe",
          2320 => x"f81153ff",
          2321 => x"800551e6",
          2322 => x"bd3f84ba",
          2323 => x"8c088638",
          2324 => x"84ba8c08",
          2325 => x"4683d890",
          2326 => x"51cbad3f",
          2327 => x"68675b59",
          2328 => x"787a278f",
          2329 => x"38655b7a",
          2330 => x"79708405",
          2331 => x"5b0c7979",
          2332 => x"26f5388a",
          2333 => x"51d9e73f",
          2334 => x"f4c539b8",
          2335 => x"3dff8005",
          2336 => x"5187963f",
          2337 => x"84ba8c08",
          2338 => x"b93dff80",
          2339 => x"05525988",
          2340 => x"d83f8153",
          2341 => x"84ba8c08",
          2342 => x"527851e9",
          2343 => x"f93f84ba",
          2344 => x"8c08802e",
          2345 => x"f4993884",
          2346 => x"ba8c0851",
          2347 => x"e7ec3ff4",
          2348 => x"8e39b83d",
          2349 => x"ff841153",
          2350 => x"ff800551",
          2351 => x"e5c83f84",
          2352 => x"ba8c0891",
          2353 => x"3883f390",
          2354 => x"335a7980",
          2355 => x"2e83c038",
          2356 => x"83f2c808",
          2357 => x"49b83dfe",
          2358 => x"fc1153ff",
          2359 => x"800551e5",
          2360 => x"a53f84ba",
          2361 => x"8c089138",
          2362 => x"83f39033",
          2363 => x"5a79802e",
          2364 => x"838a3883",
          2365 => x"f2cc0847",
          2366 => x"b83dfef8",
          2367 => x"1153ff80",
          2368 => x"0551e582",
          2369 => x"3f84ba8c",
          2370 => x"08802ea5",
          2371 => x"3880665c",
          2372 => x"5c7a882e",
          2373 => x"8338815c",
          2374 => x"7a903270",
          2375 => x"30707207",
          2376 => x"9f2a7e06",
          2377 => x"5c5f5d79",
          2378 => x"802e8838",
          2379 => x"7aa02e83",
          2380 => x"38884683",
          2381 => x"d8a051d6",
          2382 => x"ba3f8055",
          2383 => x"68546553",
          2384 => x"66526851",
          2385 => x"eb9e3f83",
          2386 => x"d8ac51d6",
          2387 => x"a63ff2ef",
          2388 => x"39646471",
          2389 => x"0c596484",
          2390 => x"0545b83d",
          2391 => x"fef01153",
          2392 => x"ff800551",
          2393 => x"e29c3f84",
          2394 => x"ba8c0880",
          2395 => x"2ef2d038",
          2396 => x"6464710c",
          2397 => x"59648405",
          2398 => x"45b83dfe",
          2399 => x"f01153ff",
          2400 => x"800551e1",
          2401 => x"fd3f84ba",
          2402 => x"8c08c638",
          2403 => x"f2b13964",
          2404 => x"5e0280ce",
          2405 => x"05227e70",
          2406 => x"82054023",
          2407 => x"7d45b83d",
          2408 => x"fef01153",
          2409 => x"ff800551",
          2410 => x"e1d83f84",
          2411 => x"ba8c0880",
          2412 => x"2ef28c38",
          2413 => x"645e0280",
          2414 => x"ce05227e",
          2415 => x"70820540",
          2416 => x"237d45b8",
          2417 => x"3dfef011",
          2418 => x"53ff8005",
          2419 => x"51e1b33f",
          2420 => x"84ba8c08",
          2421 => x"ffb938f1",
          2422 => x"e639b83d",
          2423 => x"fefc1153",
          2424 => x"ff800551",
          2425 => x"e3a03f84",
          2426 => x"ba8c0880",
          2427 => x"2e81dc38",
          2428 => x"685c0280",
          2429 => x"db05337c",
          2430 => x"34688105",
          2431 => x"49fb9b39",
          2432 => x"b83dfef0",
          2433 => x"1153ff80",
          2434 => x"0551e0f6",
          2435 => x"3f84ba8c",
          2436 => x"08802e81",
          2437 => x"98386464",
          2438 => x"710c5d64",
          2439 => x"84057046",
          2440 => x"59f7e139",
          2441 => x"7a832e09",
          2442 => x"8106f393",
          2443 => x"387b5583",
          2444 => x"d6985480",
          2445 => x"5383d8b8",
          2446 => x"527c51c8",
          2447 => x"eb3ff38c",
          2448 => x"397b527c",
          2449 => x"51da803f",
          2450 => x"f3823983",
          2451 => x"d8c451d4",
          2452 => x"a23ff0eb",
          2453 => x"39b83dfe",
          2454 => x"f01153ff",
          2455 => x"800551e0",
          2456 => x"a13f84ba",
          2457 => x"8c08802e",
          2458 => x"b8386459",
          2459 => x"0280ce05",
          2460 => x"22797082",
          2461 => x"055b2378",
          2462 => x"45f7e739",
          2463 => x"83f39133",
          2464 => x"5c7b802e",
          2465 => x"80cf3883",
          2466 => x"f2d40847",
          2467 => x"fcea3983",
          2468 => x"f391335c",
          2469 => x"7b802ea1",
          2470 => x"3883f2d0",
          2471 => x"0849fcb5",
          2472 => x"3983d8f0",
          2473 => x"51d3cc3f",
          2474 => x"6459f7b6",
          2475 => x"3983d8f0",
          2476 => x"51d3c03f",
          2477 => x"6459f6cc",
          2478 => x"3983f392",
          2479 => x"33597880",
          2480 => x"2ea53883",
          2481 => x"f2d80849",
          2482 => x"fc8b3983",
          2483 => x"d8f051d3",
          2484 => x"a23ff9c6",
          2485 => x"3983f392",
          2486 => x"33597880",
          2487 => x"2e9b3883",
          2488 => x"f2dc0847",
          2489 => x"fc923983",
          2490 => x"f393335e",
          2491 => x"7d802e9b",
          2492 => x"3883f2e0",
          2493 => x"0849fbdd",
          2494 => x"3983f393",
          2495 => x"335e7d80",
          2496 => x"2e9b3883",
          2497 => x"f2e40847",
          2498 => x"fbee3983",
          2499 => x"f38e335d",
          2500 => x"7c802e9b",
          2501 => x"3883f2e8",
          2502 => x"0849fbb9",
          2503 => x"3983f38e",
          2504 => x"335d7c80",
          2505 => x"2e943883",
          2506 => x"f2ec0847",
          2507 => x"fbca3983",
          2508 => x"f2f808fc",
          2509 => x"800549fb",
          2510 => x"9c3983f2",
          2511 => x"f8088805",
          2512 => x"47fbb539",
          2513 => x"f33d0d80",
          2514 => x"0b84babc",
          2515 => x"3487c094",
          2516 => x"8c700856",
          2517 => x"57878480",
          2518 => x"527451da",
          2519 => x"c83f84ba",
          2520 => x"8c08902b",
          2521 => x"77085755",
          2522 => x"87848052",
          2523 => x"7551dab5",
          2524 => x"3f7484ba",
          2525 => x"8c080777",
          2526 => x"0c87c094",
          2527 => x"9c700856",
          2528 => x"57878480",
          2529 => x"527451da",
          2530 => x"9c3f84ba",
          2531 => x"8c08902b",
          2532 => x"77085755",
          2533 => x"87848052",
          2534 => x"7551da89",
          2535 => x"3f7484ba",
          2536 => x"8c080777",
          2537 => x"0c8c8083",
          2538 => x"0b87c094",
          2539 => x"840c8c80",
          2540 => x"830b87c0",
          2541 => x"94940c81",
          2542 => x"bcec5c81",
          2543 => x"c7eb5d83",
          2544 => x"028405a1",
          2545 => x"0534805e",
          2546 => x"84d5ec0b",
          2547 => x"893d7088",
          2548 => x"130c7072",
          2549 => x"0c84d5f0",
          2550 => x"0c56b6f5",
          2551 => x"3f89833f",
          2552 => x"95873fba",
          2553 => x"8d5194fc",
          2554 => x"3f83d2f8",
          2555 => x"5283d2fc",
          2556 => x"51c4953f",
          2557 => x"83f2fc70",
          2558 => x"22525594",
          2559 => x"873f83d3",
          2560 => x"845483d3",
          2561 => x"90538115",
          2562 => x"335283d3",
          2563 => x"9851c3f8",
          2564 => x"3f8d973f",
          2565 => x"ecf83f80",
          2566 => x"04fb3d0d",
          2567 => x"77700856",
          2568 => x"56807552",
          2569 => x"5374732e",
          2570 => x"81833874",
          2571 => x"337081ff",
          2572 => x"06525270",
          2573 => x"a02e0981",
          2574 => x"06913881",
          2575 => x"15703370",
          2576 => x"81ff0653",
          2577 => x"535570a0",
          2578 => x"2ef13871",
          2579 => x"81ff0654",
          2580 => x"73a22e81",
          2581 => x"82387452",
          2582 => x"72812e80",
          2583 => x"e7388072",
          2584 => x"337081ff",
          2585 => x"06535454",
          2586 => x"70a02e83",
          2587 => x"38815470",
          2588 => x"802e8b38",
          2589 => x"73802e86",
          2590 => x"38811252",
          2591 => x"e1398073",
          2592 => x"81ff0652",
          2593 => x"5470a02e",
          2594 => x"09810683",
          2595 => x"38815470",
          2596 => x"a2327030",
          2597 => x"70802576",
          2598 => x"07525253",
          2599 => x"72802e88",
          2600 => x"38807270",
          2601 => x"81055434",
          2602 => x"71760c74",
          2603 => x"517084ba",
          2604 => x"8c0c873d",
          2605 => x"0d047080",
          2606 => x"2ec43873",
          2607 => x"802effbe",
          2608 => x"38811252",
          2609 => x"80723370",
          2610 => x"81ff0653",
          2611 => x"545470a2",
          2612 => x"2ee43881",
          2613 => x"54e03981",
          2614 => x"15558175",
          2615 => x"53537281",
          2616 => x"2e098106",
          2617 => x"fef838dc",
          2618 => x"39fc3d0d",
          2619 => x"76537208",
          2620 => x"8b38800b",
          2621 => x"84ba8c0c",
          2622 => x"863d0d04",
          2623 => x"863dfc05",
          2624 => x"527251da",
          2625 => x"fd3f84ba",
          2626 => x"8c08802e",
          2627 => x"e5387484",
          2628 => x"ba8c0c86",
          2629 => x"3d0d04fc",
          2630 => x"3d0d7682",
          2631 => x"1133ff05",
          2632 => x"52538152",
          2633 => x"708b2681",
          2634 => x"98388313",
          2635 => x"33ff0554",
          2636 => x"8252739e",
          2637 => x"26818a38",
          2638 => x"84133351",
          2639 => x"83527097",
          2640 => x"2680fe38",
          2641 => x"85133354",
          2642 => x"845273bb",
          2643 => x"2680f238",
          2644 => x"86133355",
          2645 => x"855274bb",
          2646 => x"2680e638",
          2647 => x"88132255",
          2648 => x"86527487",
          2649 => x"e72680d9",
          2650 => x"388a1322",
          2651 => x"54875273",
          2652 => x"87e72680",
          2653 => x"cc38810b",
          2654 => x"87c0989c",
          2655 => x"0c722287",
          2656 => x"c098bc0c",
          2657 => x"82133387",
          2658 => x"c098b80c",
          2659 => x"83133387",
          2660 => x"c098b40c",
          2661 => x"84133387",
          2662 => x"c098b00c",
          2663 => x"85133387",
          2664 => x"c098ac0c",
          2665 => x"86133387",
          2666 => x"c098a80c",
          2667 => x"7487c098",
          2668 => x"a40c7387",
          2669 => x"c098a00c",
          2670 => x"800b87c0",
          2671 => x"989c0c80",
          2672 => x"527184ba",
          2673 => x"8c0c863d",
          2674 => x"0d04f33d",
          2675 => x"0d7f5b87",
          2676 => x"c0989c5d",
          2677 => x"817d0c87",
          2678 => x"c098bc08",
          2679 => x"5e7d7b23",
          2680 => x"87c098b8",
          2681 => x"085c7b82",
          2682 => x"1c3487c0",
          2683 => x"98b4085a",
          2684 => x"79831c34",
          2685 => x"87c098b0",
          2686 => x"085c7b84",
          2687 => x"1c3487c0",
          2688 => x"98ac085a",
          2689 => x"79851c34",
          2690 => x"87c098a8",
          2691 => x"085c7b86",
          2692 => x"1c3487c0",
          2693 => x"98a4085c",
          2694 => x"7b881c23",
          2695 => x"87c098a0",
          2696 => x"085a798a",
          2697 => x"1c23807d",
          2698 => x"0c7983ff",
          2699 => x"ff06597b",
          2700 => x"83ffff06",
          2701 => x"58861b33",
          2702 => x"57851b33",
          2703 => x"56841b33",
          2704 => x"55831b33",
          2705 => x"54821b33",
          2706 => x"537d83ff",
          2707 => x"ff065283",
          2708 => x"d8f451ff",
          2709 => x"bfb23f8f",
          2710 => x"3d0d04fe",
          2711 => x"3d0d0293",
          2712 => x"05335372",
          2713 => x"812ea838",
          2714 => x"725180e8",
          2715 => x"b13f84ba",
          2716 => x"8c08982b",
          2717 => x"70982c51",
          2718 => x"5271ff2e",
          2719 => x"09810686",
          2720 => x"3872832e",
          2721 => x"e3387184",
          2722 => x"ba8c0c84",
          2723 => x"3d0d0472",
          2724 => x"5180e88a",
          2725 => x"3f84ba8c",
          2726 => x"08982b70",
          2727 => x"982c5152",
          2728 => x"71ff2e09",
          2729 => x"8106df38",
          2730 => x"725180e7",
          2731 => x"f13f84ba",
          2732 => x"8c08982b",
          2733 => x"70982c51",
          2734 => x"5271ff2e",
          2735 => x"d238c739",
          2736 => x"fd3d0d80",
          2737 => x"70545271",
          2738 => x"882b5481",
          2739 => x"5180e7ce",
          2740 => x"3f84ba8c",
          2741 => x"08982b70",
          2742 => x"982c5152",
          2743 => x"71ff2eeb",
          2744 => x"38737207",
          2745 => x"81145452",
          2746 => x"837325db",
          2747 => x"387184ba",
          2748 => x"8c0c853d",
          2749 => x"0d04fc3d",
          2750 => x"0d029b05",
          2751 => x"3383f2c4",
          2752 => x"337081ff",
          2753 => x"06535555",
          2754 => x"70802e80",
          2755 => x"f43887c0",
          2756 => x"94940870",
          2757 => x"962a7081",
          2758 => x"06535452",
          2759 => x"70802e8c",
          2760 => x"3871912a",
          2761 => x"70810651",
          2762 => x"5170e338",
          2763 => x"72813281",
          2764 => x"06537280",
          2765 => x"2e8a3871",
          2766 => x"932a8106",
          2767 => x"5271cf38",
          2768 => x"7381ff06",
          2769 => x"5187c094",
          2770 => x"80527080",
          2771 => x"2e863887",
          2772 => x"c0949052",
          2773 => x"74720c74",
          2774 => x"84ba8c0c",
          2775 => x"863d0d04",
          2776 => x"71912a70",
          2777 => x"81065151",
          2778 => x"70973872",
          2779 => x"81328106",
          2780 => x"5372802e",
          2781 => x"cb387193",
          2782 => x"2a810652",
          2783 => x"71802ec0",
          2784 => x"3887c094",
          2785 => x"84087096",
          2786 => x"2a708106",
          2787 => x"53545270",
          2788 => x"cf38d839",
          2789 => x"ff3d0d02",
          2790 => x"8f053370",
          2791 => x"30709f2a",
          2792 => x"51525270",
          2793 => x"83f2c434",
          2794 => x"833d0d04",
          2795 => x"fa3d0d78",
          2796 => x"55807533",
          2797 => x"70565257",
          2798 => x"70772e80",
          2799 => x"e7388115",
          2800 => x"83f2c433",
          2801 => x"7081ff06",
          2802 => x"54575571",
          2803 => x"802e80ff",
          2804 => x"3887c094",
          2805 => x"94087096",
          2806 => x"2a708106",
          2807 => x"53545270",
          2808 => x"802e8c38",
          2809 => x"71912a70",
          2810 => x"81065151",
          2811 => x"70e33872",
          2812 => x"81328106",
          2813 => x"5372802e",
          2814 => x"8a387193",
          2815 => x"2a810652",
          2816 => x"71cf3875",
          2817 => x"81ff0651",
          2818 => x"87c09480",
          2819 => x"5270802e",
          2820 => x"863887c0",
          2821 => x"94905273",
          2822 => x"720c8117",
          2823 => x"75335557",
          2824 => x"73ff9b38",
          2825 => x"7684ba8c",
          2826 => x"0c883d0d",
          2827 => x"0471912a",
          2828 => x"70810651",
          2829 => x"51709838",
          2830 => x"72813281",
          2831 => x"06537280",
          2832 => x"2ec13871",
          2833 => x"932a8106",
          2834 => x"5271802e",
          2835 => x"ffb53887",
          2836 => x"c0948408",
          2837 => x"70962a70",
          2838 => x"81065354",
          2839 => x"5270ce38",
          2840 => x"d739ff3d",
          2841 => x"0d87c09e",
          2842 => x"8008709c",
          2843 => x"2a8a0652",
          2844 => x"5270802e",
          2845 => x"84ab3887",
          2846 => x"c09ea408",
          2847 => x"83f2c80c",
          2848 => x"87c09ea8",
          2849 => x"0883f2cc",
          2850 => x"0c87c09e",
          2851 => x"940883f2",
          2852 => x"d00c87c0",
          2853 => x"9e980883",
          2854 => x"f2d40c87",
          2855 => x"c09e9c08",
          2856 => x"83f2d80c",
          2857 => x"87c09ea0",
          2858 => x"0883f2dc",
          2859 => x"0c87c09e",
          2860 => x"ac0883f2",
          2861 => x"e00c87c0",
          2862 => x"9eb00883",
          2863 => x"f2e40c87",
          2864 => x"c09eb408",
          2865 => x"83f2e80c",
          2866 => x"87c09eb8",
          2867 => x"0883f2ec",
          2868 => x"0c87c09e",
          2869 => x"bc0883f2",
          2870 => x"f00c87c0",
          2871 => x"9ec00883",
          2872 => x"f2f40c87",
          2873 => x"c09ec408",
          2874 => x"83f2f80c",
          2875 => x"87c09e80",
          2876 => x"08527183",
          2877 => x"f2fc2387",
          2878 => x"c09e8408",
          2879 => x"83f3800c",
          2880 => x"87c09e88",
          2881 => x"0883f384",
          2882 => x"0c87c09e",
          2883 => x"8c0883f3",
          2884 => x"880c810b",
          2885 => x"83f38c34",
          2886 => x"800b87c0",
          2887 => x"9e900870",
          2888 => x"84800a06",
          2889 => x"51525270",
          2890 => x"82fb3871",
          2891 => x"83f38d34",
          2892 => x"800b87c0",
          2893 => x"9e900870",
          2894 => x"88800a06",
          2895 => x"51525270",
          2896 => x"802e8338",
          2897 => x"81527183",
          2898 => x"f38e3480",
          2899 => x"0b87c09e",
          2900 => x"90087090",
          2901 => x"800a0651",
          2902 => x"52527080",
          2903 => x"2e833881",
          2904 => x"527183f3",
          2905 => x"8f34800b",
          2906 => x"87c09e90",
          2907 => x"08708880",
          2908 => x"80065152",
          2909 => x"5270802e",
          2910 => x"83388152",
          2911 => x"7183f390",
          2912 => x"34800b87",
          2913 => x"c09e9008",
          2914 => x"70a08080",
          2915 => x"06515252",
          2916 => x"70802e83",
          2917 => x"38815271",
          2918 => x"83f39134",
          2919 => x"800b87c0",
          2920 => x"9e900870",
          2921 => x"90808006",
          2922 => x"51525270",
          2923 => x"802e8338",
          2924 => x"81527183",
          2925 => x"f3923480",
          2926 => x"0b87c09e",
          2927 => x"90087084",
          2928 => x"80800651",
          2929 => x"52527080",
          2930 => x"2e833881",
          2931 => x"527183f3",
          2932 => x"9334800b",
          2933 => x"87c09e90",
          2934 => x"08708280",
          2935 => x"80065152",
          2936 => x"5270802e",
          2937 => x"83388152",
          2938 => x"7183f394",
          2939 => x"34800b87",
          2940 => x"c09e9008",
          2941 => x"70818080",
          2942 => x"06515252",
          2943 => x"70802e83",
          2944 => x"38815271",
          2945 => x"83f39534",
          2946 => x"800b87c0",
          2947 => x"9e900870",
          2948 => x"80c08006",
          2949 => x"51525270",
          2950 => x"802e8338",
          2951 => x"81527183",
          2952 => x"f3963480",
          2953 => x"0b87c09e",
          2954 => x"900870a0",
          2955 => x"80065152",
          2956 => x"5270802e",
          2957 => x"83388152",
          2958 => x"7183f397",
          2959 => x"3487c09e",
          2960 => x"90089880",
          2961 => x"06708a2a",
          2962 => x"53517183",
          2963 => x"f3983480",
          2964 => x"0b87c09e",
          2965 => x"90087084",
          2966 => x"80065152",
          2967 => x"5270802e",
          2968 => x"83388152",
          2969 => x"7183f399",
          2970 => x"3487c09e",
          2971 => x"900883f0",
          2972 => x"0670842a",
          2973 => x"53517183",
          2974 => x"f39a3480",
          2975 => x"0b87c09e",
          2976 => x"90087088",
          2977 => x"06515252",
          2978 => x"70802e83",
          2979 => x"38815271",
          2980 => x"83f39b34",
          2981 => x"87c09e90",
          2982 => x"08870651",
          2983 => x"7083f39c",
          2984 => x"34833d0d",
          2985 => x"048152fd",
          2986 => x"8239fb3d",
          2987 => x"0d83d98c",
          2988 => x"51ffb6d4",
          2989 => x"3f83f38c",
          2990 => x"33547386",
          2991 => x"aa3883d9",
          2992 => x"a051c3af",
          2993 => x"3f83f38e",
          2994 => x"33557485",
          2995 => x"fa3883f3",
          2996 => x"93335473",
          2997 => x"85d13883",
          2998 => x"f3903356",
          2999 => x"7585a838",
          3000 => x"83f39133",
          3001 => x"557484ff",
          3002 => x"3883f392",
          3003 => x"33547384",
          3004 => x"d63883f3",
          3005 => x"97335675",
          3006 => x"84b33883",
          3007 => x"f39b3354",
          3008 => x"73849038",
          3009 => x"83f39933",
          3010 => x"557483ed",
          3011 => x"3883f38d",
          3012 => x"33567583",
          3013 => x"cf3883f3",
          3014 => x"8f335473",
          3015 => x"83b13883",
          3016 => x"f3943355",
          3017 => x"74839338",
          3018 => x"83f39533",
          3019 => x"567582f4",
          3020 => x"3883f396",
          3021 => x"33547381",
          3022 => x"ec3883d9",
          3023 => x"b851c2b3",
          3024 => x"3f83f2f0",
          3025 => x"085283d9",
          3026 => x"c451ffb5",
          3027 => x"bb3f83f2",
          3028 => x"f4085283",
          3029 => x"d9ec51ff",
          3030 => x"b5ae3f83",
          3031 => x"f2f80852",
          3032 => x"83da9451",
          3033 => x"ffb5a13f",
          3034 => x"83dabc51",
          3035 => x"c2853f83",
          3036 => x"f2fc2252",
          3037 => x"83dac451",
          3038 => x"ffb58d3f",
          3039 => x"83f38008",
          3040 => x"56bd84c0",
          3041 => x"527551ca",
          3042 => x"9c3f84ba",
          3043 => x"8c08bd84",
          3044 => x"c0297671",
          3045 => x"31545484",
          3046 => x"ba8c0852",
          3047 => x"83daec51",
          3048 => x"ffb4e53f",
          3049 => x"83f39333",
          3050 => x"557480c3",
          3051 => x"3883f38e",
          3052 => x"3355748a",
          3053 => x"388a51c3",
          3054 => x"a53f873d",
          3055 => x"0d0483f3",
          3056 => x"880856bd",
          3057 => x"84c05275",
          3058 => x"51c9da3f",
          3059 => x"84ba8c08",
          3060 => x"bd84c029",
          3061 => x"76713154",
          3062 => x"5484ba8c",
          3063 => x"085283db",
          3064 => x"9851ffb4",
          3065 => x"a33f8a51",
          3066 => x"c2f43f87",
          3067 => x"3d0d0483",
          3068 => x"f3840856",
          3069 => x"bd84c052",
          3070 => x"7551c9a9",
          3071 => x"3f84ba8c",
          3072 => x"08bd84c0",
          3073 => x"29767131",
          3074 => x"545484ba",
          3075 => x"8c085283",
          3076 => x"dbc451ff",
          3077 => x"b3f23f83",
          3078 => x"f38e3355",
          3079 => x"74802eff",
          3080 => x"9438ff9a",
          3081 => x"3983dbf0",
          3082 => x"51c0c83f",
          3083 => x"83d9b851",
          3084 => x"c0c13f83",
          3085 => x"f2f00852",
          3086 => x"83d9c451",
          3087 => x"ffb3c93f",
          3088 => x"83f2f408",
          3089 => x"5283d9ec",
          3090 => x"51ffb3bc",
          3091 => x"3f83f2f8",
          3092 => x"085283da",
          3093 => x"9451ffb3",
          3094 => x"af3f83da",
          3095 => x"bc51c093",
          3096 => x"3f83f2fc",
          3097 => x"225283da",
          3098 => x"c451ffb3",
          3099 => x"9b3f83f3",
          3100 => x"800856bd",
          3101 => x"84c05275",
          3102 => x"51c8aa3f",
          3103 => x"84ba8c08",
          3104 => x"bd84c029",
          3105 => x"76713154",
          3106 => x"5484ba8c",
          3107 => x"085283da",
          3108 => x"ec51ffb2",
          3109 => x"f33f83f3",
          3110 => x"93335574",
          3111 => x"802efe8d",
          3112 => x"38fecc39",
          3113 => x"83dbf851",
          3114 => x"ffbfc83f",
          3115 => x"83f39633",
          3116 => x"5473802e",
          3117 => x"fd8438fe",
          3118 => x"ec3983dc",
          3119 => x"8051ffbf",
          3120 => x"b23f83f3",
          3121 => x"95335675",
          3122 => x"802efce5",
          3123 => x"38d63983",
          3124 => x"dc8c51ff",
          3125 => x"bf9d3f83",
          3126 => x"f3943355",
          3127 => x"74802efc",
          3128 => x"c738d739",
          3129 => x"83dc9851",
          3130 => x"ffbf883f",
          3131 => x"83f38f33",
          3132 => x"5473802e",
          3133 => x"fca938d7",
          3134 => x"3983f39a",
          3135 => x"335283dc",
          3136 => x"ac51ffb2",
          3137 => x"833f83f3",
          3138 => x"8d335675",
          3139 => x"802efc86",
          3140 => x"38d23983",
          3141 => x"f39c3352",
          3142 => x"83dccc51",
          3143 => x"ffb1e93f",
          3144 => x"83f39933",
          3145 => x"5574802e",
          3146 => x"fbe338cd",
          3147 => x"3983f398",
          3148 => x"335283dc",
          3149 => x"ec51ffb1",
          3150 => x"cf3f83f3",
          3151 => x"9b335473",
          3152 => x"802efbc0",
          3153 => x"38cd3983",
          3154 => x"f2d80883",
          3155 => x"f2dc0811",
          3156 => x"545283dd",
          3157 => x"8c51ffb1",
          3158 => x"af3f83f3",
          3159 => x"97335675",
          3160 => x"802efb97",
          3161 => x"38c73983",
          3162 => x"f2d00883",
          3163 => x"f2d40811",
          3164 => x"545283dd",
          3165 => x"a851ffb1",
          3166 => x"8f3f83f3",
          3167 => x"92335473",
          3168 => x"802efaee",
          3169 => x"38c13983",
          3170 => x"f2c80883",
          3171 => x"f2cc0811",
          3172 => x"545283dd",
          3173 => x"c451ffb0",
          3174 => x"ef3f83f3",
          3175 => x"91335574",
          3176 => x"802efac5",
          3177 => x"38c13983",
          3178 => x"f2e00883",
          3179 => x"f2e40811",
          3180 => x"545283dd",
          3181 => x"e051ffb0",
          3182 => x"cf3f83f3",
          3183 => x"90335675",
          3184 => x"802efa9c",
          3185 => x"38c13983",
          3186 => x"f2e80883",
          3187 => x"f2ec0811",
          3188 => x"545283dd",
          3189 => x"fc51ffb0",
          3190 => x"af3f83f3",
          3191 => x"93335473",
          3192 => x"802ef9f3",
          3193 => x"38c13983",
          3194 => x"de9851ff",
          3195 => x"b09a3f83",
          3196 => x"d9a051ff",
          3197 => x"bcfd3f83",
          3198 => x"f38e3355",
          3199 => x"74802ef9",
          3200 => x"cd38c439",
          3201 => x"ff3d0d02",
          3202 => x"8e053352",
          3203 => x"7185268c",
          3204 => x"38711010",
          3205 => x"83c3c405",
          3206 => x"52710804",
          3207 => x"83deac51",
          3208 => x"ffafe53f",
          3209 => x"833d0d04",
          3210 => x"83deb451",
          3211 => x"ffafd93f",
          3212 => x"833d0d04",
          3213 => x"83debc51",
          3214 => x"ffafcd3f",
          3215 => x"833d0d04",
          3216 => x"83dec451",
          3217 => x"ffafc13f",
          3218 => x"833d0d04",
          3219 => x"83decc51",
          3220 => x"ffafb53f",
          3221 => x"833d0d04",
          3222 => x"83ded451",
          3223 => x"ffafa93f",
          3224 => x"833d0d04",
          3225 => x"7188800c",
          3226 => x"04800b87",
          3227 => x"c096840c",
          3228 => x"0483f3a0",
          3229 => x"0887c096",
          3230 => x"840c04d9",
          3231 => x"3d0daa3d",
          3232 => x"08ad3d08",
          3233 => x"5a5a8170",
          3234 => x"57588052",
          3235 => x"83f3f808",
          3236 => x"518288d2",
          3237 => x"3f84ba8c",
          3238 => x"0880ed38",
          3239 => x"8b3d57ff",
          3240 => x"0b83f3f8",
          3241 => x"08545580",
          3242 => x"f8527651",
          3243 => x"82d2df3f",
          3244 => x"84ba8c08",
          3245 => x"802ea438",
          3246 => x"7651c0ec",
          3247 => x"3f84ba8c",
          3248 => x"08811757",
          3249 => x"55800b84",
          3250 => x"ba8c0825",
          3251 => x"8e3884ba",
          3252 => x"8c08ff05",
          3253 => x"70185555",
          3254 => x"80743474",
          3255 => x"09703070",
          3256 => x"72079f2a",
          3257 => x"51555578",
          3258 => x"762e8538",
          3259 => x"73ffb038",
          3260 => x"83f3f808",
          3261 => x"8c110853",
          3262 => x"518287ea",
          3263 => x"3f84ba8c",
          3264 => x"088f3878",
          3265 => x"762e9a38",
          3266 => x"7784ba8c",
          3267 => x"0ca93d0d",
          3268 => x"0483e284",
          3269 => x"51ffadf0",
          3270 => x"3f78762e",
          3271 => x"098106e8",
          3272 => x"38765279",
          3273 => x"51c0a03f",
          3274 => x"7951ffbf",
          3275 => x"fb3fab3d",
          3276 => x"085684ba",
          3277 => x"8c087634",
          3278 => x"765283e2",
          3279 => x"b051ffad",
          3280 => x"c73f800b",
          3281 => x"84ba8c0c",
          3282 => x"a93d0d04",
          3283 => x"d83d0dab",
          3284 => x"3d08ad3d",
          3285 => x"0871725d",
          3286 => x"72335757",
          3287 => x"5a5773a0",
          3288 => x"2e819138",
          3289 => x"800b8d3d",
          3290 => x"59567510",
          3291 => x"101083f4",
          3292 => x"80057008",
          3293 => x"5254ffbf",
          3294 => x"af3f84ba",
          3295 => x"8c085379",
          3296 => x"52730851",
          3297 => x"c08f3f84",
          3298 => x"ba8c0890",
          3299 => x"38841433",
          3300 => x"5473812e",
          3301 => x"81883873",
          3302 => x"822e9938",
          3303 => x"81167081",
          3304 => x"ff065754",
          3305 => x"827627c2",
          3306 => x"38805473",
          3307 => x"84ba8c0c",
          3308 => x"aa3d0d04",
          3309 => x"811a5aaa",
          3310 => x"3dff8411",
          3311 => x"53ff8005",
          3312 => x"51c7c33f",
          3313 => x"84ba8c08",
          3314 => x"802ed138",
          3315 => x"ff1b5378",
          3316 => x"527651fd",
          3317 => x"a63f84ba",
          3318 => x"8c0881ff",
          3319 => x"06547380",
          3320 => x"2ec93881",
          3321 => x"167081ff",
          3322 => x"06575482",
          3323 => x"7627fefa",
          3324 => x"38ffb639",
          3325 => x"78337705",
          3326 => x"56767627",
          3327 => x"fee63881",
          3328 => x"15705b70",
          3329 => x"33555573",
          3330 => x"a02e0981",
          3331 => x"06fed538",
          3332 => x"757526eb",
          3333 => x"38800b8d",
          3334 => x"3d5956fe",
          3335 => x"cd397384",
          3336 => x"ba8c0853",
          3337 => x"83f3f808",
          3338 => x"52568285",
          3339 => x"b93f84ba",
          3340 => x"8c0880d0",
          3341 => x"3883f3f8",
          3342 => x"085380f8",
          3343 => x"52775182",
          3344 => x"cfcc3f84",
          3345 => x"ba8c0880",
          3346 => x"2eba3877",
          3347 => x"51ffbdd8",
          3348 => x"3f84ba8c",
          3349 => x"0855800b",
          3350 => x"84ba8c08",
          3351 => x"259d3884",
          3352 => x"ba8c08ff",
          3353 => x"05701958",
          3354 => x"55807734",
          3355 => x"77537552",
          3356 => x"811683e1",
          3357 => x"f85256ff",
          3358 => x"ab8e3f74",
          3359 => x"ff2e0981",
          3360 => x"06ffb238",
          3361 => x"810b84ba",
          3362 => x"8c0caa3d",
          3363 => x"0d04ce3d",
          3364 => x"0db53d08",
          3365 => x"b73d08b9",
          3366 => x"3d085a41",
          3367 => x"5c800bb4",
          3368 => x"3d3483f3",
          3369 => x"fc3383f3",
          3370 => x"f808565d",
          3371 => x"749e3874",
          3372 => x"83f3f433",
          3373 => x"56567480",
          3374 => x"2e82cb38",
          3375 => x"77802e91",
          3376 => x"8d388170",
          3377 => x"77065a57",
          3378 => x"7890a038",
          3379 => x"77802e90",
          3380 => x"fd38933d",
          3381 => x"b43d5f5f",
          3382 => x"8051eaff",
          3383 => x"3f84ba8c",
          3384 => x"08982b70",
          3385 => x"982c5b56",
          3386 => x"79ff2eec",
          3387 => x"387981ff",
          3388 => x"0684d1c8",
          3389 => x"3370982b",
          3390 => x"70982c84",
          3391 => x"d1c43370",
          3392 => x"982b7097",
          3393 => x"2c71982c",
          3394 => x"05701010",
          3395 => x"83ded805",
          3396 => x"70081570",
          3397 => x"3352535c",
          3398 => x"5d46525b",
          3399 => x"585c5981",
          3400 => x"5774792e",
          3401 => x"80cd3878",
          3402 => x"75278187",
          3403 => x"38758180",
          3404 => x"0a2981ff",
          3405 => x"0a057098",
          3406 => x"2c575580",
          3407 => x"762481cb",
          3408 => x"38751016",
          3409 => x"70822b56",
          3410 => x"57800b83",
          3411 => x"dedc1633",
          3412 => x"42577761",
          3413 => x"25913883",
          3414 => x"ded81508",
          3415 => x"18703356",
          3416 => x"4178752e",
          3417 => x"81953876",
          3418 => x"802ec238",
          3419 => x"7584d1c4",
          3420 => x"34815776",
          3421 => x"802e8199",
          3422 => x"38811b70",
          3423 => x"982b7098",
          3424 => x"2c84d1c4",
          3425 => x"3370982b",
          3426 => x"70972c71",
          3427 => x"982c0570",
          3428 => x"822b83de",
          3429 => x"dc11335f",
          3430 => x"535f5d58",
          3431 => x"5d57577a",
          3432 => x"782e8190",
          3433 => x"387684d1",
          3434 => x"c834feac",
          3435 => x"39815776",
          3436 => x"ffba3875",
          3437 => x"81800a29",
          3438 => x"81800a05",
          3439 => x"70982c70",
          3440 => x"81ff0659",
          3441 => x"57417695",
          3442 => x"2680c038",
          3443 => x"75101670",
          3444 => x"822b5155",
          3445 => x"800b83de",
          3446 => x"dc163342",
          3447 => x"57776125",
          3448 => x"ce3883de",
          3449 => x"d8150818",
          3450 => x"70334255",
          3451 => x"78612eff",
          3452 => x"bc387680",
          3453 => x"2effbc38",
          3454 => x"fef23981",
          3455 => x"5776802e",
          3456 => x"feab38fe",
          3457 => x"e7398156",
          3458 => x"fdb23980",
          3459 => x"5776fee9",
          3460 => x"387684d1",
          3461 => x"c8347684",
          3462 => x"d1c43479",
          3463 => x"7e34767f",
          3464 => x"0c625574",
          3465 => x"9526fdb0",
          3466 => x"38741010",
          3467 => x"83c3dc05",
          3468 => x"57760804",
          3469 => x"83dee015",
          3470 => x"087f0c80",
          3471 => x"0b84d1c8",
          3472 => x"34800b84",
          3473 => x"d1c434d9",
          3474 => x"3984d1d0",
          3475 => x"33567580",
          3476 => x"2efd8538",
          3477 => x"84d5f008",
          3478 => x"528851ff",
          3479 => x"b6903f84",
          3480 => x"d1d033ff",
          3481 => x"05577684",
          3482 => x"d1d034fc",
          3483 => x"eb3984d1",
          3484 => x"d0337081",
          3485 => x"ff0684d1",
          3486 => x"cc335b57",
          3487 => x"55757927",
          3488 => x"fcd63884",
          3489 => x"d5f00852",
          3490 => x"81155877",
          3491 => x"84d1d034",
          3492 => x"7b167033",
          3493 => x"5255ffb5",
          3494 => x"d53ffcbc",
          3495 => x"397c932e",
          3496 => x"8bda387c",
          3497 => x"101083f3",
          3498 => x"a8057008",
          3499 => x"5759758f",
          3500 => x"83387584",
          3501 => x"d1cc3475",
          3502 => x"7c3484d1",
          3503 => x"cc3384d1",
          3504 => x"d0335656",
          3505 => x"74802eb6",
          3506 => x"3884d5f0",
          3507 => x"08528851",
          3508 => x"ffb59b3f",
          3509 => x"84d5f008",
          3510 => x"52a051ff",
          3511 => x"b5903f84",
          3512 => x"d5f00852",
          3513 => x"8851ffb5",
          3514 => x"853f84d1",
          3515 => x"d033ff05",
          3516 => x"5b7a84d1",
          3517 => x"d0347a81",
          3518 => x"ff065574",
          3519 => x"cc387b51",
          3520 => x"ffa6853f",
          3521 => x"7584d1d0",
          3522 => x"34fbcd39",
          3523 => x"7c8a3883",
          3524 => x"f3f00856",
          3525 => x"758d9e38",
          3526 => x"7c101083",
          3527 => x"f3a405fc",
          3528 => x"11085755",
          3529 => x"758ef938",
          3530 => x"74085675",
          3531 => x"802efba8",
          3532 => x"387551ff",
          3533 => x"b7f23f84",
          3534 => x"ba8c0884",
          3535 => x"d1cc3484",
          3536 => x"ba8c0881",
          3537 => x"ff068105",
          3538 => x"5375527b",
          3539 => x"51ffb89a",
          3540 => x"3f84d1cc",
          3541 => x"3384d1d0",
          3542 => x"33565674",
          3543 => x"802eff9e",
          3544 => x"3884d5f0",
          3545 => x"08528851",
          3546 => x"ffb4833f",
          3547 => x"84d5f008",
          3548 => x"52a051ff",
          3549 => x"b3f83f84",
          3550 => x"d5f00852",
          3551 => x"8851ffb3",
          3552 => x"ed3f84d1",
          3553 => x"d033ff05",
          3554 => x"557484d1",
          3555 => x"d0347481",
          3556 => x"ff0655c7",
          3557 => x"3984d1d0",
          3558 => x"337081ff",
          3559 => x"0684d1cc",
          3560 => x"335b5755",
          3561 => x"757927fa",
          3562 => x"af3884d5",
          3563 => x"f0085281",
          3564 => x"15577684",
          3565 => x"d1d0347b",
          3566 => x"16703352",
          3567 => x"55ffb3ae",
          3568 => x"3f84d1d0",
          3569 => x"337081ff",
          3570 => x"0684d1cc",
          3571 => x"335a5755",
          3572 => x"757827fa",
          3573 => x"833884d5",
          3574 => x"f0085281",
          3575 => x"15577684",
          3576 => x"d1d0347b",
          3577 => x"16703352",
          3578 => x"55ffb382",
          3579 => x"3f84d1d0",
          3580 => x"337081ff",
          3581 => x"0684d1cc",
          3582 => x"335a5755",
          3583 => x"777626ff",
          3584 => x"a938f9d4",
          3585 => x"3984d1d0",
          3586 => x"3384d1cc",
          3587 => x"33565674",
          3588 => x"762ef9c4",
          3589 => x"38ff155b",
          3590 => x"7a84d1cc",
          3591 => x"3475982b",
          3592 => x"70982c7c",
          3593 => x"81ff0643",
          3594 => x"575a6076",
          3595 => x"2480ef38",
          3596 => x"84d5f008",
          3597 => x"52a051ff",
          3598 => x"b2b43f84",
          3599 => x"d1d03370",
          3600 => x"982b7098",
          3601 => x"2c84d1cc",
          3602 => x"335a5757",
          3603 => x"41747724",
          3604 => x"f9863884",
          3605 => x"d5f00852",
          3606 => x"8851ffb2",
          3607 => x"913f7481",
          3608 => x"800a2981",
          3609 => x"800a0570",
          3610 => x"982c84d1",
          3611 => x"cc335d56",
          3612 => x"5a747b24",
          3613 => x"f8e23884",
          3614 => x"d5f00852",
          3615 => x"8851ffb1",
          3616 => x"ed3f7481",
          3617 => x"800a2981",
          3618 => x"800a0570",
          3619 => x"982c84d1",
          3620 => x"cc335d56",
          3621 => x"5a7a7525",
          3622 => x"ffb938f8",
          3623 => x"bb397b16",
          3624 => x"58811833",
          3625 => x"783484d5",
          3626 => x"f0085277",
          3627 => x"3351ffb1",
          3628 => x"bd3f7581",
          3629 => x"800a2981",
          3630 => x"800a0570",
          3631 => x"982c84d1",
          3632 => x"cc335b57",
          3633 => x"55757925",
          3634 => x"fee6387b",
          3635 => x"16588118",
          3636 => x"33783484",
          3637 => x"d5f00852",
          3638 => x"773351ff",
          3639 => x"b1903f75",
          3640 => x"81800a29",
          3641 => x"81800a05",
          3642 => x"70982c84",
          3643 => x"d1cc335b",
          3644 => x"57557876",
          3645 => x"24ffa738",
          3646 => x"feb63984",
          3647 => x"d1d03355",
          3648 => x"74802ef7",
          3649 => x"d33884d5",
          3650 => x"f0085288",
          3651 => x"51ffb0de",
          3652 => x"3f84d1d0",
          3653 => x"33ff0557",
          3654 => x"7684d1d0",
          3655 => x"347681ff",
          3656 => x"0655dd39",
          3657 => x"84d1cc33",
          3658 => x"7c055f80",
          3659 => x"7f3484d5",
          3660 => x"f008528a",
          3661 => x"51ffb0b6",
          3662 => x"3f84d1cc",
          3663 => x"527b51f4",
          3664 => x"8b3f84ba",
          3665 => x"8c0881ff",
          3666 => x"06587789",
          3667 => x"cf3884d1",
          3668 => x"cc335776",
          3669 => x"802e80d8",
          3670 => x"3883f3fc",
          3671 => x"33701010",
          3672 => x"83f3a405",
          3673 => x"7008575e",
          3674 => x"56748ba0",
          3675 => x"3875822b",
          3676 => x"87fc0683",
          3677 => x"f3a40581",
          3678 => x"18705357",
          3679 => x"5b80e8ca",
          3680 => x"3f84ba8c",
          3681 => x"087b0c83",
          3682 => x"f3fc3370",
          3683 => x"101083f3",
          3684 => x"a4057008",
          3685 => x"57414174",
          3686 => x"8bad3883",
          3687 => x"f3f80856",
          3688 => x"75802e8c",
          3689 => x"3883f3f4",
          3690 => x"33587780",
          3691 => x"2e8bbc38",
          3692 => x"800b84d1",
          3693 => x"d034800b",
          3694 => x"84d1cc34",
          3695 => x"7b84ba8c",
          3696 => x"0cb43d0d",
          3697 => x"0484d1d0",
          3698 => x"33557480",
          3699 => x"2eb63884",
          3700 => x"d5f00852",
          3701 => x"8851ffaf",
          3702 => x"953f84d5",
          3703 => x"f00852a0",
          3704 => x"51ffaf8a",
          3705 => x"3f84d5f0",
          3706 => x"08528851",
          3707 => x"ffaeff3f",
          3708 => x"84d1d033",
          3709 => x"ff055675",
          3710 => x"84d1d034",
          3711 => x"7581ff06",
          3712 => x"5574cc38",
          3713 => x"83d2b851",
          3714 => x"ff9ffd3f",
          3715 => x"800b84d1",
          3716 => x"d034800b",
          3717 => x"84d1cc34",
          3718 => x"f5be3983",
          3719 => x"7c34800b",
          3720 => x"811d3484",
          3721 => x"d1d03355",
          3722 => x"74802eb6",
          3723 => x"3884d5f0",
          3724 => x"08528851",
          3725 => x"ffaeb73f",
          3726 => x"84d5f008",
          3727 => x"52a051ff",
          3728 => x"aeac3f84",
          3729 => x"d5f00852",
          3730 => x"8851ffae",
          3731 => x"a13f84d1",
          3732 => x"d033ff05",
          3733 => x"5d7c84d1",
          3734 => x"d0347c81",
          3735 => x"ff065574",
          3736 => x"cc3883d2",
          3737 => x"b851ff9f",
          3738 => x"9f3f800b",
          3739 => x"84d1d034",
          3740 => x"800b84d1",
          3741 => x"cc347b84",
          3742 => x"ba8c0cb4",
          3743 => x"3d0d0484",
          3744 => x"d1d03370",
          3745 => x"81ff065c",
          3746 => x"567a802e",
          3747 => x"f4ca3884",
          3748 => x"d1cc33ff",
          3749 => x"05597884",
          3750 => x"d1cc34ff",
          3751 => x"16587784",
          3752 => x"d1d03484",
          3753 => x"d5f00852",
          3754 => x"8851ffad",
          3755 => x"c13f84d1",
          3756 => x"d0337098",
          3757 => x"2b70982c",
          3758 => x"84d1cc33",
          3759 => x"5a525b56",
          3760 => x"76762480",
          3761 => x"ef3884d5",
          3762 => x"f00852a0",
          3763 => x"51ffad9e",
          3764 => x"3f84d1d0",
          3765 => x"3370982b",
          3766 => x"70982c84",
          3767 => x"d1cc335d",
          3768 => x"57595674",
          3769 => x"7a24f3f0",
          3770 => x"3884d5f0",
          3771 => x"08528851",
          3772 => x"ffacfb3f",
          3773 => x"7481800a",
          3774 => x"2981800a",
          3775 => x"0570982c",
          3776 => x"84d1cc33",
          3777 => x"5b515574",
          3778 => x"7924f3cc",
          3779 => x"3884d5f0",
          3780 => x"08528851",
          3781 => x"ffacd73f",
          3782 => x"7481800a",
          3783 => x"2981800a",
          3784 => x"0570982c",
          3785 => x"84d1cc33",
          3786 => x"5b515578",
          3787 => x"7525ffb9",
          3788 => x"38f3a539",
          3789 => x"7b165781",
          3790 => x"17337734",
          3791 => x"84d5f008",
          3792 => x"52763351",
          3793 => x"ffaca73f",
          3794 => x"7581800a",
          3795 => x"2981800a",
          3796 => x"0570982c",
          3797 => x"84d1cc33",
          3798 => x"43575b75",
          3799 => x"6125fee6",
          3800 => x"387b1657",
          3801 => x"81173377",
          3802 => x"3484d5f0",
          3803 => x"08527633",
          3804 => x"51ffabfa",
          3805 => x"3f758180",
          3806 => x"0a298180",
          3807 => x"0a057098",
          3808 => x"2c84d1cc",
          3809 => x"3343575b",
          3810 => x"607624ff",
          3811 => x"a738feb6",
          3812 => x"3984d1d0",
          3813 => x"337081ff",
          3814 => x"06585876",
          3815 => x"602ef2b8",
          3816 => x"3884d1cc",
          3817 => x"33557675",
          3818 => x"27ae3874",
          3819 => x"982b7098",
          3820 => x"2c574176",
          3821 => x"7624a138",
          3822 => x"7b165b7a",
          3823 => x"33811c34",
          3824 => x"7581800a",
          3825 => x"2981ff0a",
          3826 => x"0570982c",
          3827 => x"84d1d033",
          3828 => x"52575875",
          3829 => x"7825e138",
          3830 => x"81185574",
          3831 => x"84d1d034",
          3832 => x"7781ff06",
          3833 => x"7c055ab3",
          3834 => x"3d337a34",
          3835 => x"84d1cc33",
          3836 => x"57766025",
          3837 => x"8b388117",
          3838 => x"567584d1",
          3839 => x"cc347557",
          3840 => x"84d1d033",
          3841 => x"7081800a",
          3842 => x"2981ff0a",
          3843 => x"0570982c",
          3844 => x"7981ff06",
          3845 => x"44585c58",
          3846 => x"60762481",
          3847 => x"ef387798",
          3848 => x"2b70982c",
          3849 => x"7881ff06",
          3850 => x"5c575975",
          3851 => x"7a25f1a8",
          3852 => x"3884d5f0",
          3853 => x"08528851",
          3854 => x"ffaab33f",
          3855 => x"7581800a",
          3856 => x"2981800a",
          3857 => x"0570982c",
          3858 => x"84d1cc33",
          3859 => x"57574175",
          3860 => x"7525f184",
          3861 => x"3884d5f0",
          3862 => x"08528851",
          3863 => x"ffaa8f3f",
          3864 => x"7581800a",
          3865 => x"2981800a",
          3866 => x"0570982c",
          3867 => x"84d1cc33",
          3868 => x"57574174",
          3869 => x"7624ffb9",
          3870 => x"38f0dd39",
          3871 => x"83f3a408",
          3872 => x"5675802e",
          3873 => x"f49d3875",
          3874 => x"51ffad9c",
          3875 => x"3f84ba8c",
          3876 => x"0884d1cc",
          3877 => x"3484ba8c",
          3878 => x"0881ff06",
          3879 => x"81055375",
          3880 => x"527b51ff",
          3881 => x"adc43f84",
          3882 => x"d1cc3384",
          3883 => x"d1d03356",
          3884 => x"5674802e",
          3885 => x"f4c83884",
          3886 => x"d5f00852",
          3887 => x"8851ffa9",
          3888 => x"ad3f84d5",
          3889 => x"f00852a0",
          3890 => x"51ffa9a2",
          3891 => x"3f84d5f0",
          3892 => x"08528851",
          3893 => x"ffa9973f",
          3894 => x"84d1d033",
          3895 => x"ff055b7a",
          3896 => x"84d1d034",
          3897 => x"7a81ff06",
          3898 => x"55c739a8",
          3899 => x"5180e1da",
          3900 => x"3f84ba8c",
          3901 => x"0883f3f8",
          3902 => x"0c84ba8c",
          3903 => x"0885a538",
          3904 => x"7683f3f4",
          3905 => x"3477efca",
          3906 => x"3880c339",
          3907 => x"84d5f008",
          3908 => x"527b1670",
          3909 => x"335258ff",
          3910 => x"a8d43f75",
          3911 => x"81800a29",
          3912 => x"81800a05",
          3913 => x"70982c84",
          3914 => x"d1cc3352",
          3915 => x"57577676",
          3916 => x"24da3884",
          3917 => x"d1d03370",
          3918 => x"982b7098",
          3919 => x"2c7981ff",
          3920 => x"065d585a",
          3921 => x"58757a25",
          3922 => x"ef8e38fd",
          3923 => x"e43983f3",
          3924 => x"f808802e",
          3925 => x"eefc3883",
          3926 => x"f3a45793",
          3927 => x"56760855",
          3928 => x"74bb38ff",
          3929 => x"16841858",
          3930 => x"56758025",
          3931 => x"f038800b",
          3932 => x"83f3fc34",
          3933 => x"83f3f808",
          3934 => x"5574802e",
          3935 => x"eed43874",
          3936 => x"5181e8c5",
          3937 => x"3f83f3f8",
          3938 => x"085180da",
          3939 => x"cd3f800b",
          3940 => x"83f3f80c",
          3941 => x"933db43d",
          3942 => x"5f5feebc",
          3943 => x"39745180",
          3944 => x"dab83f80",
          3945 => x"770cff16",
          3946 => x"84185856",
          3947 => x"758025ff",
          3948 => x"ac38ffba",
          3949 => x"397551ff",
          3950 => x"aaee3f84",
          3951 => x"ba8c0884",
          3952 => x"d1cc3484",
          3953 => x"ba8c0881",
          3954 => x"ff068105",
          3955 => x"5375527b",
          3956 => x"51ffab96",
          3957 => x"3f930b84",
          3958 => x"d1cc3384",
          3959 => x"d1d03357",
          3960 => x"575d7480",
          3961 => x"2ef29738",
          3962 => x"84d5f008",
          3963 => x"528851ff",
          3964 => x"a6fc3f84",
          3965 => x"d5f00852",
          3966 => x"a051ffa6",
          3967 => x"f13f84d5",
          3968 => x"f0085288",
          3969 => x"51ffa6e6",
          3970 => x"3f84d1d0",
          3971 => x"33ff055a",
          3972 => x"7984d1d0",
          3973 => x"347981ff",
          3974 => x"0655c739",
          3975 => x"807c3480",
          3976 => x"0b84d1d0",
          3977 => x"34800b84",
          3978 => x"d1cc347b",
          3979 => x"84ba8c0c",
          3980 => x"b43d0d04",
          3981 => x"7551ffa9",
          3982 => x"ef3f84ba",
          3983 => x"8c0884d1",
          3984 => x"cc3484ba",
          3985 => x"8c0881ff",
          3986 => x"06810553",
          3987 => x"75527b51",
          3988 => x"ffaa973f",
          3989 => x"811d7081",
          3990 => x"ff0684d1",
          3991 => x"cc3384d1",
          3992 => x"d0335852",
          3993 => x"5e567480",
          3994 => x"2ef19338",
          3995 => x"84d5f008",
          3996 => x"528851ff",
          3997 => x"a5f83f84",
          3998 => x"d5f00852",
          3999 => x"a051ffa5",
          4000 => x"ed3f84d5",
          4001 => x"f0085288",
          4002 => x"51ffa5e2",
          4003 => x"3f84d1d0",
          4004 => x"33ff0557",
          4005 => x"7684d1d0",
          4006 => x"347681ff",
          4007 => x"0655c739",
          4008 => x"7551ffa9",
          4009 => x"833f84ba",
          4010 => x"8c0884d1",
          4011 => x"cc3484ba",
          4012 => x"8c0881ff",
          4013 => x"06810553",
          4014 => x"75527b51",
          4015 => x"ffa9ab3f",
          4016 => x"ff1d7081",
          4017 => x"ff0684d1",
          4018 => x"cc3384d1",
          4019 => x"d0335858",
          4020 => x"5e587480",
          4021 => x"2ef0a738",
          4022 => x"84d5f008",
          4023 => x"528851ff",
          4024 => x"a58c3f84",
          4025 => x"d5f00852",
          4026 => x"a051ffa5",
          4027 => x"813f84d5",
          4028 => x"f0085288",
          4029 => x"51ffa4f6",
          4030 => x"3f84d1d0",
          4031 => x"33ff0541",
          4032 => x"6084d1d0",
          4033 => x"346081ff",
          4034 => x"0655c739",
          4035 => x"745180d7",
          4036 => x"c93f83f3",
          4037 => x"fc337082",
          4038 => x"2b87fc06",
          4039 => x"83f3a405",
          4040 => x"81197054",
          4041 => x"525c5680",
          4042 => x"dda03f84",
          4043 => x"ba8c087b",
          4044 => x"0c83f3fc",
          4045 => x"33701010",
          4046 => x"83f3a405",
          4047 => x"70085741",
          4048 => x"4174802e",
          4049 => x"f4d53875",
          4050 => x"537b5274",
          4051 => x"51ffa89a",
          4052 => x"3f83f3fc",
          4053 => x"33810570",
          4054 => x"81ff065a",
          4055 => x"56937927",
          4056 => x"82f23877",
          4057 => x"83f3fc34",
          4058 => x"f4b139b4",
          4059 => x"3dfef805",
          4060 => x"5476537b",
          4061 => x"52755181",
          4062 => x"d98f3f83",
          4063 => x"f3f80852",
          4064 => x"8a5182ba",
          4065 => x"d73f83f3",
          4066 => x"f8085181",
          4067 => x"e0c23f80",
          4068 => x"0b84d1d0",
          4069 => x"34800b84",
          4070 => x"d1cc347b",
          4071 => x"84ba8c0c",
          4072 => x"b43d0d04",
          4073 => x"93537752",
          4074 => x"84ba8c08",
          4075 => x"5181cac7",
          4076 => x"3f84ba8c",
          4077 => x"0882a538",
          4078 => x"84ba8c08",
          4079 => x"963d5c5d",
          4080 => x"83f3f808",
          4081 => x"5380f852",
          4082 => x"7a5182b8",
          4083 => x"c13f84ba",
          4084 => x"8c085a84",
          4085 => x"ba8c087b",
          4086 => x"2e098106",
          4087 => x"e9ee3884",
          4088 => x"ba8c0851",
          4089 => x"ffa6c13f",
          4090 => x"84ba8c08",
          4091 => x"56800b84",
          4092 => x"ba8c0825",
          4093 => x"80e33884",
          4094 => x"ba8c08ff",
          4095 => x"05701b58",
          4096 => x"56807734",
          4097 => x"7581ff06",
          4098 => x"83f3fc33",
          4099 => x"70101083",
          4100 => x"f3a40570",
          4101 => x"08584058",
          4102 => x"597480f2",
          4103 => x"3876822b",
          4104 => x"87fc0683",
          4105 => x"f3a40581",
          4106 => x"1a705358",
          4107 => x"5580db9a",
          4108 => x"3f84ba8c",
          4109 => x"08750c83",
          4110 => x"f3fc3370",
          4111 => x"101083f3",
          4112 => x"a4057008",
          4113 => x"57404174",
          4114 => x"a038811d",
          4115 => x"7081ff06",
          4116 => x"5e57937d",
          4117 => x"27833880",
          4118 => x"5d75ff2e",
          4119 => x"098106fe",
          4120 => x"df3877e8",
          4121 => x"ed38f9e6",
          4122 => x"39765379",
          4123 => x"527451ff",
          4124 => x"a5f83f83",
          4125 => x"f3fc3381",
          4126 => x"057081ff",
          4127 => x"065b5793",
          4128 => x"7a2780c8",
          4129 => x"38800b83",
          4130 => x"f3fc34ff",
          4131 => x"bd397451",
          4132 => x"80d4c73f",
          4133 => x"83f3fc33",
          4134 => x"70822b87",
          4135 => x"fc0683f3",
          4136 => x"a405811b",
          4137 => x"70545256",
          4138 => x"5780da9e",
          4139 => x"3f84ba8c",
          4140 => x"08750c83",
          4141 => x"f3fc3370",
          4142 => x"101083f3",
          4143 => x"a4057008",
          4144 => x"57404174",
          4145 => x"802eff82",
          4146 => x"38ff9e39",
          4147 => x"7683f3fc",
          4148 => x"34fef739",
          4149 => x"7583f3fc",
          4150 => x"34f1c039",
          4151 => x"83e1b851",
          4152 => x"ff9f903f",
          4153 => x"77e7eb38",
          4154 => x"f8e439f2",
          4155 => x"3d0d0280",
          4156 => x"c3053302",
          4157 => x"840580c7",
          4158 => x"05335b53",
          4159 => x"72832681",
          4160 => x"8d387281",
          4161 => x"2e818b38",
          4162 => x"81732583",
          4163 => x"9e387282",
          4164 => x"2e82a838",
          4165 => x"87a3a080",
          4166 => x"5987a3b0",
          4167 => x"80705e57",
          4168 => x"80569fa0",
          4169 => x"5879762e",
          4170 => x"90387583",
          4171 => x"f9bc3475",
          4172 => x"83f9bd34",
          4173 => x"7583f9ba",
          4174 => x"2383f9b8",
          4175 => x"3370982b",
          4176 => x"71902b07",
          4177 => x"71882b07",
          4178 => x"71077a7f",
          4179 => x"5656565b",
          4180 => x"78772794",
          4181 => x"38807470",
          4182 => x"8405560c",
          4183 => x"74737084",
          4184 => x"05550c76",
          4185 => x"7426ee38",
          4186 => x"757827a2",
          4187 => x"3883f9b8",
          4188 => x"338498de",
          4189 => x"17797831",
          4190 => x"555555a0",
          4191 => x"0be0e015",
          4192 => x"34747470",
          4193 => x"81055634",
          4194 => x"ff135372",
          4195 => x"ee38903d",
          4196 => x"0d0487a3",
          4197 => x"a0800b83",
          4198 => x"f9bc3370",
          4199 => x"10101183",
          4200 => x"f9bd3371",
          4201 => x"90291174",
          4202 => x"055b4158",
          4203 => x"405987a3",
          4204 => x"b0800b84",
          4205 => x"b8803370",
          4206 => x"81ff0684",
          4207 => x"b7ff3370",
          4208 => x"81ff0683",
          4209 => x"f9ba2270",
          4210 => x"83ffff06",
          4211 => x"7075295d",
          4212 => x"595d585e",
          4213 => x"575b5d73",
          4214 => x"73268738",
          4215 => x"72743175",
          4216 => x"29567981",
          4217 => x"ff067e81",
          4218 => x"ff067c81",
          4219 => x"ff067a83",
          4220 => x"ffff0662",
          4221 => x"81ff0670",
          4222 => x"7529145d",
          4223 => x"4257575b",
          4224 => x"5c747426",
          4225 => x"8f3883f9",
          4226 => x"bc337476",
          4227 => x"3105707d",
          4228 => x"291b595f",
          4229 => x"7683065c",
          4230 => x"7b802efe",
          4231 => x"9c38787d",
          4232 => x"55537277",
          4233 => x"26fec138",
          4234 => x"80737081",
          4235 => x"05553483",
          4236 => x"f9b83374",
          4237 => x"70810556",
          4238 => x"34e83987",
          4239 => x"a3a08059",
          4240 => x"87a3b080",
          4241 => x"7084b880",
          4242 => x"337081ff",
          4243 => x"0684b7ff",
          4244 => x"337081ff",
          4245 => x"0683f9ba",
          4246 => x"22707429",
          4247 => x"5d5b5d57",
          4248 => x"5e565e57",
          4249 => x"74782781",
          4250 => x"df387381",
          4251 => x"ff067381",
          4252 => x"ff067171",
          4253 => x"29185a54",
          4254 => x"5479802e",
          4255 => x"fdbb3880",
          4256 => x"0b83f9bc",
          4257 => x"34800b83",
          4258 => x"f9bd3483",
          4259 => x"f9b83370",
          4260 => x"982b7190",
          4261 => x"2b077188",
          4262 => x"2b077107",
          4263 => x"7a7f5656",
          4264 => x"565b7679",
          4265 => x"26fdae38",
          4266 => x"fdbe3972",
          4267 => x"fce63883",
          4268 => x"f9bc3370",
          4269 => x"81ff0670",
          4270 => x"10101183",
          4271 => x"f9bd3371",
          4272 => x"90291187",
          4273 => x"a3a08011",
          4274 => x"5e575b56",
          4275 => x"565f87a3",
          4276 => x"b0807014",
          4277 => x"84b88033",
          4278 => x"7081ff06",
          4279 => x"84b7ff33",
          4280 => x"7081ff06",
          4281 => x"83f9ba22",
          4282 => x"7083ffff",
          4283 => x"067c7529",
          4284 => x"60055e5a",
          4285 => x"415f585f",
          4286 => x"405e5779",
          4287 => x"73268b38",
          4288 => x"727a3115",
          4289 => x"707d2919",
          4290 => x"57537d81",
          4291 => x"ff067481",
          4292 => x"ff067171",
          4293 => x"297d83ff",
          4294 => x"ff066281",
          4295 => x"ff067075",
          4296 => x"29585f5b",
          4297 => x"5c5d557b",
          4298 => x"78268538",
          4299 => x"77752953",
          4300 => x"79733116",
          4301 => x"7983065b",
          4302 => x"5879fde2",
          4303 => x"38768306",
          4304 => x"5c7bfdda",
          4305 => x"38fbf239",
          4306 => x"7478317b",
          4307 => x"2956fe9a",
          4308 => x"39fb3d0d",
          4309 => x"86ee809c",
          4310 => x"5480f474",
          4311 => x"34ffb074",
          4312 => x"3486ee80",
          4313 => x"98538073",
          4314 => x"34807334",
          4315 => x"86ee8094",
          4316 => x"568a7634",
          4317 => x"807634ff",
          4318 => x"80743486",
          4319 => x"ee808c55",
          4320 => x"ff8a7534",
          4321 => x"87753485",
          4322 => x"75348175",
          4323 => x"34815283",
          4324 => x"51fad83f",
          4325 => x"879087e0",
          4326 => x"70085454",
          4327 => x"81f85687",
          4328 => x"8c81f873",
          4329 => x"77068407",
          4330 => x"54557275",
          4331 => x"34730870",
          4332 => x"80ff0680",
          4333 => x"c0075153",
          4334 => x"72753487",
          4335 => x"9087cc08",
          4336 => x"70770681",
          4337 => x"07515372",
          4338 => x"878c81f3",
          4339 => x"34730881",
          4340 => x"f7068807",
          4341 => x"53727534",
          4342 => x"80d00b84",
          4343 => x"b8803480",
          4344 => x"0b84ba8c",
          4345 => x"0c873d0d",
          4346 => x"0484b880",
          4347 => x"3384ba8c",
          4348 => x"0c04f73d",
          4349 => x"0d02af05",
          4350 => x"33028405",
          4351 => x"b3053384",
          4352 => x"b7ff335b",
          4353 => x"59568153",
          4354 => x"75792682",
          4355 => x"da3884b8",
          4356 => x"803383f9",
          4357 => x"bd3383f9",
          4358 => x"bc337271",
          4359 => x"291287a3",
          4360 => x"a0801183",
          4361 => x"f9ba225f",
          4362 => x"51575971",
          4363 => x"7c290570",
          4364 => x"83ffff06",
          4365 => x"83f89233",
          4366 => x"53575853",
          4367 => x"72812e83",
          4368 => x"c43883f9",
          4369 => x"ba227605",
          4370 => x"557483f9",
          4371 => x"ba2383f9",
          4372 => x"bc337605",
          4373 => x"7081ff06",
          4374 => x"7a81ff06",
          4375 => x"555b5572",
          4376 => x"7a26828c",
          4377 => x"38ff1953",
          4378 => x"7283f9bc",
          4379 => x"3483f9ba",
          4380 => x"227083ff",
          4381 => x"ff0684b7",
          4382 => x"fe335c55",
          4383 => x"57797426",
          4384 => x"82893884",
          4385 => x"b8803376",
          4386 => x"71295458",
          4387 => x"8054729f",
          4388 => x"9f26ac38",
          4389 => x"8498de70",
          4390 => x"145455e0",
          4391 => x"e01333e0",
          4392 => x"e0163472",
          4393 => x"70810554",
          4394 => x"33757081",
          4395 => x"05573481",
          4396 => x"145484b7",
          4397 => x"fd7327e3",
          4398 => x"38739f9f",
          4399 => x"26a13883",
          4400 => x"f9b83384",
          4401 => x"98de1554",
          4402 => x"55a00be0",
          4403 => x"e0143474",
          4404 => x"73708105",
          4405 => x"55348114",
          4406 => x"549f9f74",
          4407 => x"27eb3884",
          4408 => x"b7fe33ff",
          4409 => x"05567583",
          4410 => x"f9ba2375",
          4411 => x"577881ff",
          4412 => x"067783ff",
          4413 => x"ff065454",
          4414 => x"73732681",
          4415 => x"fd387274",
          4416 => x"31810584",
          4417 => x"b8803371",
          4418 => x"71295855",
          4419 => x"57755587",
          4420 => x"a3a08058",
          4421 => x"87a3b080",
          4422 => x"7981ff06",
          4423 => x"7581ff06",
          4424 => x"71712919",
          4425 => x"5c5c5457",
          4426 => x"757927b9",
          4427 => x"388498de",
          4428 => x"1654e0e0",
          4429 => x"14335384",
          4430 => x"b8881333",
          4431 => x"78708105",
          4432 => x"5a347370",
          4433 => x"81055533",
          4434 => x"77708105",
          4435 => x"59348115",
          4436 => x"84b88033",
          4437 => x"84b7ff33",
          4438 => x"71712919",
          4439 => x"565c5a55",
          4440 => x"727526ce",
          4441 => x"38805372",
          4442 => x"84ba8c0c",
          4443 => x"8b3d0d04",
          4444 => x"7483f9bc",
          4445 => x"3483f9ba",
          4446 => x"227083ff",
          4447 => x"ff0684b7",
          4448 => x"fe335c55",
          4449 => x"57737a27",
          4450 => x"fdf93877",
          4451 => x"802efedd",
          4452 => x"387881ff",
          4453 => x"06ff0583",
          4454 => x"f9bc3356",
          4455 => x"5372752e",
          4456 => x"098106fe",
          4457 => x"c8387376",
          4458 => x"31810584",
          4459 => x"b8803371",
          4460 => x"71297872",
          4461 => x"29115652",
          4462 => x"59547373",
          4463 => x"27feae38",
          4464 => x"83f9b833",
          4465 => x"8498de15",
          4466 => x"74763155",
          4467 => x"5656a00b",
          4468 => x"e0e01634",
          4469 => x"75757081",
          4470 => x"055734ff",
          4471 => x"13537280",
          4472 => x"2efe8a38",
          4473 => x"a00be0e0",
          4474 => x"16347575",
          4475 => x"70810557",
          4476 => x"34ff1353",
          4477 => x"72d838fd",
          4478 => x"f439800b",
          4479 => x"84b88033",
          4480 => x"5556fe89",
          4481 => x"3983f9be",
          4482 => x"15335984",
          4483 => x"b8881933",
          4484 => x"743484b7",
          4485 => x"ff3359fc",
          4486 => x"a939fc3d",
          4487 => x"0d760284",
          4488 => x"059f0533",
          4489 => x"53517086",
          4490 => x"269b3870",
          4491 => x"101083c4",
          4492 => x"b4055170",
          4493 => x"080484b8",
          4494 => x"80335171",
          4495 => x"71278638",
          4496 => x"7183f9bd",
          4497 => x"34800b84",
          4498 => x"ba8c0c86",
          4499 => x"3d0d0480",
          4500 => x"0b83f9bd",
          4501 => x"3483f9bc",
          4502 => x"337081ff",
          4503 => x"06545272",
          4504 => x"802ee238",
          4505 => x"ff125170",
          4506 => x"83f9bc34",
          4507 => x"800b84ba",
          4508 => x"8c0c863d",
          4509 => x"0d0483f9",
          4510 => x"bc337073",
          4511 => x"31700970",
          4512 => x"9f2c7206",
          4513 => x"54555354",
          4514 => x"7083f9bc",
          4515 => x"34de3983",
          4516 => x"f9bc3372",
          4517 => x"0584b7ff",
          4518 => x"33ff1155",
          4519 => x"56517075",
          4520 => x"25833870",
          4521 => x"537283f9",
          4522 => x"bc34800b",
          4523 => x"84ba8c0c",
          4524 => x"863d0d04",
          4525 => x"83f9bd33",
          4526 => x"70733170",
          4527 => x"09709f2c",
          4528 => x"72065456",
          4529 => x"53557083",
          4530 => x"f9bd3480",
          4531 => x"0b84ba8c",
          4532 => x"0c863d0d",
          4533 => x"0483f9bd",
          4534 => x"33720584",
          4535 => x"b88033ff",
          4536 => x"11555551",
          4537 => x"70742583",
          4538 => x"38705372",
          4539 => x"83f9bd34",
          4540 => x"800b84ba",
          4541 => x"8c0c863d",
          4542 => x"0d04800b",
          4543 => x"83f9bd34",
          4544 => x"83f9bc33",
          4545 => x"84b7ff33",
          4546 => x"ff055652",
          4547 => x"717525fe",
          4548 => x"b4388112",
          4549 => x"517083f9",
          4550 => x"bc34fed0",
          4551 => x"39ff3d0d",
          4552 => x"028f0533",
          4553 => x"5170b126",
          4554 => x"b3387010",
          4555 => x"1083c4d0",
          4556 => x"05517008",
          4557 => x"0483f9b8",
          4558 => x"337080f0",
          4559 => x"0671842b",
          4560 => x"80f00670",
          4561 => x"72842a07",
          4562 => x"51525351",
          4563 => x"7180f02e",
          4564 => x"0981069c",
          4565 => x"3880f20b",
          4566 => x"83f9b834",
          4567 => x"800b84ba",
          4568 => x"8c0c833d",
          4569 => x"0d0483f9",
          4570 => x"b833819f",
          4571 => x"06900751",
          4572 => x"7083f9b8",
          4573 => x"34800b84",
          4574 => x"ba8c0c83",
          4575 => x"3d0d0483",
          4576 => x"f9b83380",
          4577 => x"f0075170",
          4578 => x"83f9b834",
          4579 => x"e83983f9",
          4580 => x"b83381fe",
          4581 => x"06860751",
          4582 => x"7083f9b8",
          4583 => x"34d73980",
          4584 => x"f10b83f9",
          4585 => x"b834800b",
          4586 => x"84ba8c0c",
          4587 => x"833d0d04",
          4588 => x"83f9b833",
          4589 => x"81fc0684",
          4590 => x"07517083",
          4591 => x"f9b834ff",
          4592 => x"b43983f9",
          4593 => x"b8338707",
          4594 => x"517083f9",
          4595 => x"b834ffa5",
          4596 => x"3983f9b8",
          4597 => x"3381fd06",
          4598 => x"85075170",
          4599 => x"83f9b834",
          4600 => x"ff933983",
          4601 => x"f9b83381",
          4602 => x"fb068307",
          4603 => x"517083f9",
          4604 => x"b834ff81",
          4605 => x"3983f9b8",
          4606 => x"3381f906",
          4607 => x"81075170",
          4608 => x"83f9b834",
          4609 => x"feef3983",
          4610 => x"f9b83381",
          4611 => x"f8065170",
          4612 => x"83f9b834",
          4613 => x"fedf3983",
          4614 => x"f9b83381",
          4615 => x"df0680d0",
          4616 => x"07517083",
          4617 => x"f9b834fe",
          4618 => x"cc3983f9",
          4619 => x"b83381bf",
          4620 => x"06b00751",
          4621 => x"7083f9b8",
          4622 => x"34feba39",
          4623 => x"83f9b833",
          4624 => x"81ef0680",
          4625 => x"e0075170",
          4626 => x"83f9b834",
          4627 => x"fea73983",
          4628 => x"f9b83381",
          4629 => x"cf0680c0",
          4630 => x"07517083",
          4631 => x"f9b834fe",
          4632 => x"943983f9",
          4633 => x"b83381af",
          4634 => x"06a00751",
          4635 => x"7083f9b8",
          4636 => x"34fe8239",
          4637 => x"83f9b833",
          4638 => x"818f0651",
          4639 => x"7083f9b8",
          4640 => x"34fdf239",
          4641 => x"83f9b833",
          4642 => x"81fa0682",
          4643 => x"07517083",
          4644 => x"f9b834fd",
          4645 => x"e039f33d",
          4646 => x"0d02bf05",
          4647 => x"33028405",
          4648 => x"80c30533",
          4649 => x"83f9bc33",
          4650 => x"83f9bb33",
          4651 => x"83f9bd33",
          4652 => x"84b88233",
          4653 => x"43415f5d",
          4654 => x"5b597882",
          4655 => x"2e82a138",
          4656 => x"788224a5",
          4657 => x"3878812e",
          4658 => x"8182387d",
          4659 => x"84b88234",
          4660 => x"800b84b8",
          4661 => x"84347a83",
          4662 => x"f9bc347b",
          4663 => x"83f9ba23",
          4664 => x"7c83f9bd",
          4665 => x"348f3d0d",
          4666 => x"0478832e",
          4667 => x"098106db",
          4668 => x"38800b84",
          4669 => x"b8823481",
          4670 => x"0b84b884",
          4671 => x"34820b83",
          4672 => x"f9bc34a8",
          4673 => x"0b83f9bd",
          4674 => x"34820b83",
          4675 => x"f9ba2379",
          4676 => x"5884b880",
          4677 => x"335784b7",
          4678 => x"ff335684",
          4679 => x"b7fe3355",
          4680 => x"7b547c53",
          4681 => x"7a5283e3",
          4682 => x"c451ff81",
          4683 => x"db3f7d84",
          4684 => x"b8823480",
          4685 => x"0b84b884",
          4686 => x"347a83f9",
          4687 => x"bc347b83",
          4688 => x"f9ba237c",
          4689 => x"83f9bd34",
          4690 => x"8f3d0d04",
          4691 => x"800b84b8",
          4692 => x"8234810b",
          4693 => x"84b88434",
          4694 => x"800b83f9",
          4695 => x"bc34a80b",
          4696 => x"83f9bd34",
          4697 => x"800b83f9",
          4698 => x"ba2384b9",
          4699 => x"8f335884",
          4700 => x"b98e3357",
          4701 => x"84b98d33",
          4702 => x"5679557b",
          4703 => x"547c537a",
          4704 => x"5283e3e0",
          4705 => x"51ff8180",
          4706 => x"3f800b84",
          4707 => x"b98d335a",
          4708 => x"5a797927",
          4709 => x"a5387910",
          4710 => x"84b9e005",
          4711 => x"70225359",
          4712 => x"83e3f851",
          4713 => x"ff80e13f",
          4714 => x"811a7081",
          4715 => x"ff0684b9",
          4716 => x"8d33525b",
          4717 => x"59787a26",
          4718 => x"dd3883d2",
          4719 => x"ec51ff80",
          4720 => x"c73f7d84",
          4721 => x"b8823480",
          4722 => x"0b84b884",
          4723 => x"347a83f9",
          4724 => x"bc347b83",
          4725 => x"f9ba237c",
          4726 => x"83f9bd34",
          4727 => x"8f3d0d04",
          4728 => x"800b84b8",
          4729 => x"8234810b",
          4730 => x"84b88434",
          4731 => x"810b83f9",
          4732 => x"bc34a80b",
          4733 => x"83f9bd34",
          4734 => x"810b83f9",
          4735 => x"ba2383f7",
          4736 => x"f051ff92",
          4737 => x"a33f84ba",
          4738 => x"8c085283",
          4739 => x"e3fc51fe",
          4740 => x"fff63f80",
          4741 => x"5983f7f0",
          4742 => x"51ff928c",
          4743 => x"3f7884ba",
          4744 => x"8c0827fd",
          4745 => x"a63883f7",
          4746 => x"f0193352",
          4747 => x"83e48451",
          4748 => x"feffd53f",
          4749 => x"81197081",
          4750 => x"ff065a5a",
          4751 => x"d839f93d",
          4752 => x"0d7a0284",
          4753 => x"05a70533",
          4754 => x"84b88033",
          4755 => x"83f9bd33",
          4756 => x"83f9bc33",
          4757 => x"72712912",
          4758 => x"87a3a080",
          4759 => x"1183f9ba",
          4760 => x"22535159",
          4761 => x"5c717c29",
          4762 => x"057083ff",
          4763 => x"ff0683f8",
          4764 => x"92335259",
          4765 => x"51555757",
          4766 => x"72812e81",
          4767 => x"e9387589",
          4768 => x"2e81f938",
          4769 => x"75892481",
          4770 => x"b9387581",
          4771 => x"2e838538",
          4772 => x"75882e82",
          4773 => x"d53884b8",
          4774 => x"803383f9",
          4775 => x"bc3383f9",
          4776 => x"bd337272",
          4777 => x"29055556",
          4778 => x"5484b888",
          4779 => x"163387a3",
          4780 => x"a0801434",
          4781 => x"84b88033",
          4782 => x"83f9bd33",
          4783 => x"83f9ba22",
          4784 => x"72712912",
          4785 => x"5a5a5653",
          4786 => x"7583f9be",
          4787 => x"183483f9",
          4788 => x"bc337371",
          4789 => x"29165854",
          4790 => x"83f9b833",
          4791 => x"87a3b080",
          4792 => x"183484b8",
          4793 => x"80337081",
          4794 => x"ff0683f9",
          4795 => x"ba2283f9",
          4796 => x"bd337272",
          4797 => x"2911575b",
          4798 => x"57555783",
          4799 => x"f9b83384",
          4800 => x"98de1434",
          4801 => x"81187081",
          4802 => x"ff065955",
          4803 => x"73782681",
          4804 => x"993884b8",
          4805 => x"81335877",
          4806 => x"81ea38ff",
          4807 => x"17537283",
          4808 => x"f9bd3484",
          4809 => x"b8833353",
          4810 => x"72802e8c",
          4811 => x"3884b884",
          4812 => x"33577680",
          4813 => x"2e80fb38",
          4814 => x"800b84ba",
          4815 => x"8c0c893d",
          4816 => x"0d04758d",
          4817 => x"2e973875",
          4818 => x"8d2480f7",
          4819 => x"38758a2e",
          4820 => x"098106fe",
          4821 => x"c1388152",
          4822 => x"8151f196",
          4823 => x"3f800b83",
          4824 => x"f9bd34ff",
          4825 => x"be3983f9",
          4826 => x"be153353",
          4827 => x"84b88813",
          4828 => x"33743475",
          4829 => x"892e0981",
          4830 => x"06fe8938",
          4831 => x"80537652",
          4832 => x"a051fdba",
          4833 => x"3f811370",
          4834 => x"81ff0654",
          4835 => x"54728326",
          4836 => x"ff913876",
          4837 => x"52a051fd",
          4838 => x"a53f8113",
          4839 => x"7081ff06",
          4840 => x"54548373",
          4841 => x"27d838fe",
          4842 => x"fa397483",
          4843 => x"f9bd34fe",
          4844 => x"f2397552",
          4845 => x"8351f9de",
          4846 => x"3f800b84",
          4847 => x"ba8c0c89",
          4848 => x"3d0d0475",
          4849 => x"80ff2e09",
          4850 => x"8106fdca",
          4851 => x"3883f9bd",
          4852 => x"337081ff",
          4853 => x"0655ff05",
          4854 => x"53738338",
          4855 => x"73537283",
          4856 => x"f9bd3476",
          4857 => x"52a051fc",
          4858 => x"d53f83f9",
          4859 => x"bd337081",
          4860 => x"ff0655ff",
          4861 => x"055373fe",
          4862 => x"a5387353",
          4863 => x"7283f9bd",
          4864 => x"34fea039",
          4865 => x"800b83f9",
          4866 => x"bd348152",
          4867 => x"8151efe2",
          4868 => x"3ffe9039",
          4869 => x"80527551",
          4870 => x"efd83ffe",
          4871 => x"8639e63d",
          4872 => x"0d0280f3",
          4873 => x"053384b9",
          4874 => x"88085759",
          4875 => x"75812e81",
          4876 => x"b8387582",
          4877 => x"2e838238",
          4878 => x"788a2e84",
          4879 => x"b538788a",
          4880 => x"2482d138",
          4881 => x"78882e84",
          4882 => x"b9387889",
          4883 => x"2e888f38",
          4884 => x"84b88033",
          4885 => x"83f9bc33",
          4886 => x"83f9bd33",
          4887 => x"72722905",
          4888 => x"585e5c84",
          4889 => x"b8881933",
          4890 => x"87a3a080",
          4891 => x"173484b8",
          4892 => x"803383f9",
          4893 => x"bd3383f9",
          4894 => x"ba227271",
          4895 => x"29125a5a",
          4896 => x"42407883",
          4897 => x"f9be1834",
          4898 => x"83f9bc33",
          4899 => x"60712962",
          4900 => x"05405a83",
          4901 => x"f9b8337f",
          4902 => x"87a3b080",
          4903 => x"053484b8",
          4904 => x"80337081",
          4905 => x"ff0683f9",
          4906 => x"ba2283f9",
          4907 => x"bd337272",
          4908 => x"29114240",
          4909 => x"5d585983",
          4910 => x"f9b83384",
          4911 => x"98de1f34",
          4912 => x"811d7081",
          4913 => x"ff064258",
          4914 => x"76612681",
          4915 => x"b83884b8",
          4916 => x"81335a79",
          4917 => x"86f138ff",
          4918 => x"19567583",
          4919 => x"f9bd3480",
          4920 => x"0b84ba8c",
          4921 => x"0c9c3d0d",
          4922 => x"0478b72e",
          4923 => x"848a38b7",
          4924 => x"792581fd",
          4925 => x"3878b82e",
          4926 => x"9bb33878",
          4927 => x"80db2e89",
          4928 => x"cc38800b",
          4929 => x"84b9880c",
          4930 => x"84b88033",
          4931 => x"83f9bc33",
          4932 => x"83f9bd33",
          4933 => x"72722905",
          4934 => x"5e404084",
          4935 => x"b8881933",
          4936 => x"87a3a080",
          4937 => x"1d3484b8",
          4938 => x"803383f9",
          4939 => x"bd3383f9",
          4940 => x"ba227271",
          4941 => x"2912415f",
          4942 => x"59567883",
          4943 => x"f9be1f34",
          4944 => x"83f9bc33",
          4945 => x"76712919",
          4946 => x"5b5783f9",
          4947 => x"b83387a3",
          4948 => x"b0801b34",
          4949 => x"84b88033",
          4950 => x"7081ff06",
          4951 => x"83f9ba22",
          4952 => x"83f9bd33",
          4953 => x"72722911",
          4954 => x"44424358",
          4955 => x"5983f9b8",
          4956 => x"33608498",
          4957 => x"de053481",
          4958 => x"1f587781",
          4959 => x"ff064160",
          4960 => x"7727feca",
          4961 => x"387783f9",
          4962 => x"bd34800b",
          4963 => x"84ba8c0c",
          4964 => x"9c3d0d04",
          4965 => x"789b2e82",
          4966 => x"b738789b",
          4967 => x"24838138",
          4968 => x"788d2e09",
          4969 => x"8106fda8",
          4970 => x"38800b83",
          4971 => x"f9bd3480",
          4972 => x"0b84ba8c",
          4973 => x"0c9c3d0d",
          4974 => x"04789b2e",
          4975 => x"82aa38d0",
          4976 => x"19567589",
          4977 => x"2684d038",
          4978 => x"84b98c33",
          4979 => x"81115957",
          4980 => x"7784b98c",
          4981 => x"347884b9",
          4982 => x"90183477",
          4983 => x"81ff0659",
          4984 => x"800b84b9",
          4985 => x"901a3480",
          4986 => x"0b84ba8c",
          4987 => x"0c9c3d0d",
          4988 => x"04789b2e",
          4989 => x"fde93880",
          4990 => x"0b84b988",
          4991 => x"0c84b880",
          4992 => x"3383f9bc",
          4993 => x"3383f9bd",
          4994 => x"33727229",
          4995 => x"055e4040",
          4996 => x"84b88819",
          4997 => x"3387a3a0",
          4998 => x"801d3484",
          4999 => x"b8803383",
          5000 => x"f9bd3383",
          5001 => x"f9ba2272",
          5002 => x"71291241",
          5003 => x"5f595678",
          5004 => x"83f9be1f",
          5005 => x"3483f9bc",
          5006 => x"33767129",
          5007 => x"195b5783",
          5008 => x"f9b83387",
          5009 => x"a3b0801b",
          5010 => x"3484b880",
          5011 => x"337081ff",
          5012 => x"0683f9ba",
          5013 => x"2283f9bd",
          5014 => x"33727229",
          5015 => x"11444243",
          5016 => x"585983f9",
          5017 => x"b8336084",
          5018 => x"98de0534",
          5019 => x"811f58fe",
          5020 => x"89398152",
          5021 => x"8151eafa",
          5022 => x"3f800b83",
          5023 => x"f9bd34fe",
          5024 => x"ae3984b8",
          5025 => x"803383f9",
          5026 => x"bd337081",
          5027 => x"ff0683f9",
          5028 => x"bc337371",
          5029 => x"291287a3",
          5030 => x"a0800583",
          5031 => x"f9ba2240",
          5032 => x"515d727e",
          5033 => x"29057083",
          5034 => x"ffff0683",
          5035 => x"f892335a",
          5036 => x"51595a5c",
          5037 => x"75812e86",
          5038 => x"a4387881",
          5039 => x"ff06ff1a",
          5040 => x"575776fc",
          5041 => x"95387656",
          5042 => x"7583f9bd",
          5043 => x"34fc9039",
          5044 => x"800b84b9",
          5045 => x"8c34800b",
          5046 => x"84b98d34",
          5047 => x"800b84b9",
          5048 => x"8e34800b",
          5049 => x"84b98f34",
          5050 => x"810b84b9",
          5051 => x"880c800b",
          5052 => x"84ba8c0c",
          5053 => x"9c3d0d04",
          5054 => x"83f9bc33",
          5055 => x"84b9f434",
          5056 => x"83f9bd33",
          5057 => x"84b9f534",
          5058 => x"83f9bb33",
          5059 => x"84b9f634",
          5060 => x"800b84b9",
          5061 => x"880c800b",
          5062 => x"84ba8c0c",
          5063 => x"9c3d0d04",
          5064 => x"7880ff2e",
          5065 => x"098106fa",
          5066 => x"a73883f9",
          5067 => x"bc3384b8",
          5068 => x"80337081",
          5069 => x"ff0683f9",
          5070 => x"bd337081",
          5071 => x"ff067275",
          5072 => x"291187a3",
          5073 => x"a0800583",
          5074 => x"f9ba225c",
          5075 => x"40727b29",
          5076 => x"057083ff",
          5077 => x"ff0683f8",
          5078 => x"9233445c",
          5079 => x"435c425b",
          5080 => x"5c7d812e",
          5081 => x"85fe3878",
          5082 => x"81ff06ff",
          5083 => x"1a585675",
          5084 => x"83387557",
          5085 => x"7683f9bd",
          5086 => x"347b81ff",
          5087 => x"067a81ff",
          5088 => x"067881ff",
          5089 => x"06727229",
          5090 => x"055f405b",
          5091 => x"84b8a833",
          5092 => x"87a3a080",
          5093 => x"1e3484b8",
          5094 => x"803383f9",
          5095 => x"bd3383f9",
          5096 => x"ba227271",
          5097 => x"29125a5e",
          5098 => x"4240a00b",
          5099 => x"83f9be18",
          5100 => x"3483f9bc",
          5101 => x"33607129",
          5102 => x"62055a56",
          5103 => x"83f9b833",
          5104 => x"87a3b080",
          5105 => x"1a3484b8",
          5106 => x"80337081",
          5107 => x"ff0683f9",
          5108 => x"ba2283f9",
          5109 => x"bd337272",
          5110 => x"2911435d",
          5111 => x"5a5e5983",
          5112 => x"f9b8337f",
          5113 => x"8498de05",
          5114 => x"34811a70",
          5115 => x"81ff065c",
          5116 => x"587c7b26",
          5117 => x"95ea3884",
          5118 => x"b881335a",
          5119 => x"7996d038",
          5120 => x"ff195877",
          5121 => x"83f9bd34",
          5122 => x"83f9bd33",
          5123 => x"7081ff06",
          5124 => x"58ff0556",
          5125 => x"fdac3978",
          5126 => x"bb2e95d8",
          5127 => x"3878bd2e",
          5128 => x"83d73878",
          5129 => x"bf2e95a8",
          5130 => x"3884b98c",
          5131 => x"335f7e83",
          5132 => x"f938ffbf",
          5133 => x"195675b4",
          5134 => x"2684c838",
          5135 => x"75101083",
          5136 => x"c6980558",
          5137 => x"77080480",
          5138 => x"0b83f9bd",
          5139 => x"34805281",
          5140 => x"51e79f3f",
          5141 => x"800b84ba",
          5142 => x"8c0c9c3d",
          5143 => x"0d0483f9",
          5144 => x"bc3384b8",
          5145 => x"80337081",
          5146 => x"ff0683f9",
          5147 => x"bd337081",
          5148 => x"ff067275",
          5149 => x"291187a3",
          5150 => x"a0800583",
          5151 => x"f9ba225c",
          5152 => x"41727b29",
          5153 => x"057083ff",
          5154 => x"ff0683f8",
          5155 => x"92334653",
          5156 => x"455c595b",
          5157 => x"5b7f812e",
          5158 => x"82ef3880",
          5159 => x"5c7a81ff",
          5160 => x"067a81ff",
          5161 => x"067a81ff",
          5162 => x"06727229",
          5163 => x"055c5840",
          5164 => x"84b8a833",
          5165 => x"87a3a080",
          5166 => x"1b3484b8",
          5167 => x"803383f9",
          5168 => x"bd3383f9",
          5169 => x"ba227271",
          5170 => x"29125e41",
          5171 => x"5e56a00b",
          5172 => x"83f9be1c",
          5173 => x"3483f9bc",
          5174 => x"33767129",
          5175 => x"1e5a5e83",
          5176 => x"f9b83387",
          5177 => x"a3b0801a",
          5178 => x"3484b880",
          5179 => x"337081ff",
          5180 => x"0683f9ba",
          5181 => x"2283f9bd",
          5182 => x"33727229",
          5183 => x"115b445a",
          5184 => x"405983f9",
          5185 => x"b8338498",
          5186 => x"de183460",
          5187 => x"81057081",
          5188 => x"ff065b58",
          5189 => x"7e7a2681",
          5190 => x"ac3884b8",
          5191 => x"81335877",
          5192 => x"92fb38ff",
          5193 => x"19567583",
          5194 => x"f9bd3481",
          5195 => x"1c7081ff",
          5196 => x"065d597b",
          5197 => x"8326f7a7",
          5198 => x"3883f9bc",
          5199 => x"3384b880",
          5200 => x"3383f9bd",
          5201 => x"337281ff",
          5202 => x"067281ff",
          5203 => x"067281ff",
          5204 => x"06727229",
          5205 => x"05545b43",
          5206 => x"5b5b5b84",
          5207 => x"b8a83387",
          5208 => x"a3a0801b",
          5209 => x"3484b880",
          5210 => x"3383f9bd",
          5211 => x"3383f9ba",
          5212 => x"22727129",
          5213 => x"125e415e",
          5214 => x"56a00b83",
          5215 => x"f9be1c34",
          5216 => x"83f9bc33",
          5217 => x"7671291e",
          5218 => x"5a5e83f9",
          5219 => x"b83387a3",
          5220 => x"b0801a34",
          5221 => x"84b88033",
          5222 => x"7081ff06",
          5223 => x"83f9ba22",
          5224 => x"83f9bd33",
          5225 => x"72722911",
          5226 => x"5b445a40",
          5227 => x"5983f9b8",
          5228 => x"338498de",
          5229 => x"18346081",
          5230 => x"057081ff",
          5231 => x"065b5879",
          5232 => x"7f27fed6",
          5233 => x"387783f9",
          5234 => x"bd34fedf",
          5235 => x"39820b84",
          5236 => x"b9880c80",
          5237 => x"0b84ba8c",
          5238 => x"0c9c3d0d",
          5239 => x"0483f9be",
          5240 => x"17335984",
          5241 => x"b8881933",
          5242 => x"7a3483f9",
          5243 => x"bd337081",
          5244 => x"ff0658ff",
          5245 => x"0556f9ca",
          5246 => x"39810b84",
          5247 => x"b98e3480",
          5248 => x"0b84ba8c",
          5249 => x"0c9c3d0d",
          5250 => x"0483f9be",
          5251 => x"17335b84",
          5252 => x"b8881b33",
          5253 => x"7c3483f9",
          5254 => x"bc3384b8",
          5255 => x"803383f9",
          5256 => x"bd335b5b",
          5257 => x"5b805cfc",
          5258 => x"f43984b9",
          5259 => x"90429c3d",
          5260 => x"dc1153d8",
          5261 => x"0551ff8a",
          5262 => x"cd3f84ba",
          5263 => x"8c08802e",
          5264 => x"fbf03884",
          5265 => x"b98d3381",
          5266 => x"11575a75",
          5267 => x"84b98d34",
          5268 => x"791083fe",
          5269 => x"06410280",
          5270 => x"ca052261",
          5271 => x"84b9e005",
          5272 => x"23fbcf39",
          5273 => x"83f9be17",
          5274 => x"335c84b8",
          5275 => x"881c337b",
          5276 => x"3483f9bc",
          5277 => x"3384b880",
          5278 => x"3383f9bd",
          5279 => x"335b5b5c",
          5280 => x"f9e53984",
          5281 => x"b8803383",
          5282 => x"f9bc3383",
          5283 => x"f9bd3372",
          5284 => x"72290541",
          5285 => x"5d5b84b8",
          5286 => x"8819337f",
          5287 => x"87a3a080",
          5288 => x"053484b8",
          5289 => x"803383f9",
          5290 => x"bd3383f9",
          5291 => x"ba227271",
          5292 => x"29125a43",
          5293 => x"5b567883",
          5294 => x"f9be1834",
          5295 => x"83f9bc33",
          5296 => x"7671291b",
          5297 => x"415e83f9",
          5298 => x"b8336087",
          5299 => x"a3b08005",
          5300 => x"3484b880",
          5301 => x"337081ff",
          5302 => x"0683f9ba",
          5303 => x"2283f9bd",
          5304 => x"33727229",
          5305 => x"11415f5a",
          5306 => x"425a83f9",
          5307 => x"b8338498",
          5308 => x"de1e3481",
          5309 => x"1c7081ff",
          5310 => x"065c5860",
          5311 => x"7b2690a2",
          5312 => x"3884b881",
          5313 => x"33587790",
          5314 => x"e238ff1a",
          5315 => x"567583f9",
          5316 => x"bd34800b",
          5317 => x"84b9880c",
          5318 => x"84b88333",
          5319 => x"407f802e",
          5320 => x"f3bd3884",
          5321 => x"b8843356",
          5322 => x"75f3b438",
          5323 => x"78528151",
          5324 => x"eae43f80",
          5325 => x"0b84ba8c",
          5326 => x"0c9c3d0d",
          5327 => x"0484b9f4",
          5328 => x"3383f9bc",
          5329 => x"3484b9f5",
          5330 => x"3383f9bd",
          5331 => x"3484b9f6",
          5332 => x"33577683",
          5333 => x"f9ba23ff",
          5334 => x"b93983f9",
          5335 => x"bc3384b9",
          5336 => x"f43483f9",
          5337 => x"bd3384b9",
          5338 => x"f53483f9",
          5339 => x"bb3384b9",
          5340 => x"f634ff9e",
          5341 => x"3984b98d",
          5342 => x"335b7a80",
          5343 => x"2eff9338",
          5344 => x"84b9e022",
          5345 => x"5d7c862e",
          5346 => x"098106ff",
          5347 => x"853883f9",
          5348 => x"bd338105",
          5349 => x"5583f9bc",
          5350 => x"33810554",
          5351 => x"9b5383e4",
          5352 => x"8c52943d",
          5353 => x"705257fe",
          5354 => x"edfe3f76",
          5355 => x"51fefef8",
          5356 => x"3f84ba8c",
          5357 => x"0881ff06",
          5358 => x"83f89033",
          5359 => x"57760541",
          5360 => x"60a024fe",
          5361 => x"cd387652",
          5362 => x"83f7f051",
          5363 => x"fefdc33f",
          5364 => x"fec03980",
          5365 => x"0b84b98d",
          5366 => x"335b5879",
          5367 => x"81ff065b",
          5368 => x"777b27fe",
          5369 => x"ad387710",
          5370 => x"84b9e005",
          5371 => x"81113357",
          5372 => x"4175b126",
          5373 => x"8aa53875",
          5374 => x"101083c7",
          5375 => x"ec055f7e",
          5376 => x"080484b9",
          5377 => x"8d335e7d",
          5378 => x"802e8fa4",
          5379 => x"3883f9bc",
          5380 => x"3384b9e1",
          5381 => x"33717131",
          5382 => x"7009709f",
          5383 => x"2c72065a",
          5384 => x"42595e5c",
          5385 => x"7583f9bc",
          5386 => x"34fde739",
          5387 => x"84b98d33",
          5388 => x"5675802e",
          5389 => x"8ee73884",
          5390 => x"b9e133ff",
          5391 => x"057081ff",
          5392 => x"0684b880",
          5393 => x"335d575f",
          5394 => x"757b27fd",
          5395 => x"c5387583",
          5396 => x"f9bd34fd",
          5397 => x"bd39800b",
          5398 => x"83f9bd34",
          5399 => x"83f9bc33",
          5400 => x"7081ff06",
          5401 => x"5d577b80",
          5402 => x"2efda738",
          5403 => x"ff175675",
          5404 => x"83f9bc34",
          5405 => x"fd9c3980",
          5406 => x"0b83f9bd",
          5407 => x"3483f9bc",
          5408 => x"3384b7ff",
          5409 => x"33ff0557",
          5410 => x"57767625",
          5411 => x"fd843881",
          5412 => x"17567583",
          5413 => x"f9bc34fc",
          5414 => x"f93984b9",
          5415 => x"8d33407f",
          5416 => x"802e8de0",
          5417 => x"3883f9bd",
          5418 => x"3384b9e1",
          5419 => x"33717131",
          5420 => x"7009709f",
          5421 => x"2c72065a",
          5422 => x"4159425a",
          5423 => x"7583f9bd",
          5424 => x"34fccf39",
          5425 => x"84b98d33",
          5426 => x"5b7a802e",
          5427 => x"fcc43884",
          5428 => x"b9e02241",
          5429 => x"60992e09",
          5430 => x"8106fcb6",
          5431 => x"3884b880",
          5432 => x"3383f9bd",
          5433 => x"3383f9bc",
          5434 => x"33727129",
          5435 => x"1287a3a0",
          5436 => x"801183f9",
          5437 => x"ba224351",
          5438 => x"5a587160",
          5439 => x"29057083",
          5440 => x"ffff0683",
          5441 => x"f8900887",
          5442 => x"fffe8006",
          5443 => x"425a5d5d",
          5444 => x"7e848280",
          5445 => x"2e92bf38",
          5446 => x"800b83f8",
          5447 => x"9134fbf2",
          5448 => x"3984b98d",
          5449 => x"335a7980",
          5450 => x"2efbe738",
          5451 => x"84b9e022",
          5452 => x"5877992e",
          5453 => x"098106fb",
          5454 => x"d938810b",
          5455 => x"83f89134",
          5456 => x"fbd03984",
          5457 => x"b98d3356",
          5458 => x"75802e90",
          5459 => x"be3884b9",
          5460 => x"e13383f9",
          5461 => x"bd335d7c",
          5462 => x"0584b880",
          5463 => x"33ff1159",
          5464 => x"5e56757d",
          5465 => x"25833875",
          5466 => x"577683f9",
          5467 => x"bd34fba2",
          5468 => x"3984b98d",
          5469 => x"33577680",
          5470 => x"2e8cc838",
          5471 => x"84b9e133",
          5472 => x"83f9bc33",
          5473 => x"42610584",
          5474 => x"b7ff33ff",
          5475 => x"11594156",
          5476 => x"75602583",
          5477 => x"38755776",
          5478 => x"83f9bc34",
          5479 => x"faf43983",
          5480 => x"e49851fe",
          5481 => x"e8e23f80",
          5482 => x"0b84b98d",
          5483 => x"33575776",
          5484 => x"76278bc7",
          5485 => x"38761084",
          5486 => x"b9e00570",
          5487 => x"22535a83",
          5488 => x"e3f851fe",
          5489 => x"e8c23f81",
          5490 => x"177081ff",
          5491 => x"0684b98d",
          5492 => x"33585858",
          5493 => x"da39820b",
          5494 => x"84b98d33",
          5495 => x"5f577d80",
          5496 => x"2e8d3884",
          5497 => x"b9e02256",
          5498 => x"75832683",
          5499 => x"38755781",
          5500 => x"527681ff",
          5501 => x"0651d5f3",
          5502 => x"3ffa9739",
          5503 => x"84b98d33",
          5504 => x"57817727",
          5505 => x"8eb73884",
          5506 => x"b9e333ff",
          5507 => x"057081ff",
          5508 => x"0684b9e1",
          5509 => x"33ff0570",
          5510 => x"81ff0684",
          5511 => x"b7ff3370",
          5512 => x"81ff06ff",
          5513 => x"11404352",
          5514 => x"5b595c5c",
          5515 => x"777e2783",
          5516 => x"38775a79",
          5517 => x"83f9ba23",
          5518 => x"7681ff06",
          5519 => x"ff18585f",
          5520 => x"777f2783",
          5521 => x"38775776",
          5522 => x"83f9bc34",
          5523 => x"84b88033",
          5524 => x"ff115740",
          5525 => x"7a6027f9",
          5526 => x"b4387a56",
          5527 => x"7583f9bd",
          5528 => x"34f9af39",
          5529 => x"84b98d33",
          5530 => x"5f7e802e",
          5531 => x"8aef3884",
          5532 => x"b9e13384",
          5533 => x"b7ff3340",
          5534 => x"5b7a7f26",
          5535 => x"f9943883",
          5536 => x"f9bc3384",
          5537 => x"b8803370",
          5538 => x"81ff0683",
          5539 => x"f9bd3371",
          5540 => x"74291187",
          5541 => x"a3a08005",
          5542 => x"83f9ba22",
          5543 => x"5f40717e",
          5544 => x"29057083",
          5545 => x"ffff0683",
          5546 => x"f8923346",
          5547 => x"5259595f",
          5548 => x"5d60812e",
          5549 => x"84f03879",
          5550 => x"83ffff06",
          5551 => x"707c315d",
          5552 => x"57807c24",
          5553 => x"8efe3884",
          5554 => x"b7ff3356",
          5555 => x"7676278e",
          5556 => x"d638ff16",
          5557 => x"567583f9",
          5558 => x"ba237c81",
          5559 => x"ff06707c",
          5560 => x"31415780",
          5561 => x"60248ee5",
          5562 => x"3884b7ff",
          5563 => x"33567676",
          5564 => x"278dee38",
          5565 => x"ff165675",
          5566 => x"83f9bc34",
          5567 => x"7e81ff06",
          5568 => x"83f9ba22",
          5569 => x"5757805a",
          5570 => x"76762690",
          5571 => x"38757731",
          5572 => x"81057e81",
          5573 => x"ff067171",
          5574 => x"295c5e5b",
          5575 => x"795887a3",
          5576 => x"a0805b87",
          5577 => x"a3b0807f",
          5578 => x"81ff067f",
          5579 => x"81ff0671",
          5580 => x"71291d42",
          5581 => x"58425c79",
          5582 => x"7f27f7d6",
          5583 => x"388498de",
          5584 => x"1a57e0e0",
          5585 => x"17335f84",
          5586 => x"b8881f33",
          5587 => x"7b708105",
          5588 => x"5d347670",
          5589 => x"81055833",
          5590 => x"7c708105",
          5591 => x"5e348118",
          5592 => x"84b88033",
          5593 => x"84b7ff33",
          5594 => x"7171291d",
          5595 => x"43405e58",
          5596 => x"776027f7",
          5597 => x"9d38e0e0",
          5598 => x"17335f84",
          5599 => x"b8881f33",
          5600 => x"7b708105",
          5601 => x"5d347670",
          5602 => x"81055833",
          5603 => x"7c708105",
          5604 => x"5e348118",
          5605 => x"84b88033",
          5606 => x"84b7ff33",
          5607 => x"7171291d",
          5608 => x"43405e58",
          5609 => x"7f7826ff",
          5610 => x"9938f6e6",
          5611 => x"3984b98d",
          5612 => x"33567580",
          5613 => x"2e87e038",
          5614 => x"805284b9",
          5615 => x"e13351d8",
          5616 => x"b13ff6ce",
          5617 => x"39800b84",
          5618 => x"b88033ff",
          5619 => x"1184b98d",
          5620 => x"335d5940",
          5621 => x"5879782e",
          5622 => x"943884b9",
          5623 => x"e0225675",
          5624 => x"782e0981",
          5625 => x"068bbe38",
          5626 => x"83f9bd33",
          5627 => x"587681ff",
          5628 => x"0683f9bc",
          5629 => x"3379435c",
          5630 => x"5c76ff2e",
          5631 => x"81ed3884",
          5632 => x"b7ff3340",
          5633 => x"7a6026f6",
          5634 => x"89387e81",
          5635 => x"ff065660",
          5636 => x"7626f5fe",
          5637 => x"387b7626",
          5638 => x"617d2707",
          5639 => x"5776f5f2",
          5640 => x"387a1010",
          5641 => x"1b709029",
          5642 => x"620587a3",
          5643 => x"a0801170",
          5644 => x"1f5d5a87",
          5645 => x"a3b08005",
          5646 => x"79830658",
          5647 => x"515d758b",
          5648 => x"ac387983",
          5649 => x"0657768b",
          5650 => x"a43883f9",
          5651 => x"b8337098",
          5652 => x"2b71902b",
          5653 => x"0771882b",
          5654 => x"07710779",
          5655 => x"7f59525f",
          5656 => x"57777a27",
          5657 => x"9e388077",
          5658 => x"70840559",
          5659 => x"0c7d7670",
          5660 => x"8405580c",
          5661 => x"797726ee",
          5662 => x"3884b880",
          5663 => x"3384b7ff",
          5664 => x"33415f7e",
          5665 => x"81ff0660",
          5666 => x"81ff0683",
          5667 => x"f9ba227d",
          5668 => x"73296405",
          5669 => x"5959595a",
          5670 => x"7777268c",
          5671 => x"38767831",
          5672 => x"1b707b29",
          5673 => x"62055740",
          5674 => x"75761d57",
          5675 => x"57767626",
          5676 => x"f4e03883",
          5677 => x"f9b83384",
          5678 => x"98de1859",
          5679 => x"5aa00be0",
          5680 => x"e0193479",
          5681 => x"78708105",
          5682 => x"5a348117",
          5683 => x"57767626",
          5684 => x"f4c038a0",
          5685 => x"0be0e019",
          5686 => x"34797870",
          5687 => x"81055a34",
          5688 => x"81175775",
          5689 => x"7727d638",
          5690 => x"f4a839ff",
          5691 => x"1f7081ff",
          5692 => x"065d58fe",
          5693 => x"8a3983f9",
          5694 => x"b8337080",
          5695 => x"f0067184",
          5696 => x"2b80f006",
          5697 => x"71842a07",
          5698 => x"585d577b",
          5699 => x"80f02e09",
          5700 => x"8106be38",
          5701 => x"80f20b83",
          5702 => x"f9b83481",
          5703 => x"187081ff",
          5704 => x"065956f5",
          5705 => x"b63983f9",
          5706 => x"be17335e",
          5707 => x"84b8881e",
          5708 => x"337c3483",
          5709 => x"f9bc3384",
          5710 => x"b8803383",
          5711 => x"f9ba2284",
          5712 => x"b7ff3342",
          5713 => x"5c5f5dfa",
          5714 => x"ee3983f9",
          5715 => x"b8338707",
          5716 => x"567583f9",
          5717 => x"b8348118",
          5718 => x"7081ff06",
          5719 => x"5956f4fb",
          5720 => x"3983f9b8",
          5721 => x"3381fd06",
          5722 => x"85075675",
          5723 => x"83f9b834",
          5724 => x"e53983f9",
          5725 => x"b83381fb",
          5726 => x"06830756",
          5727 => x"7583f9b8",
          5728 => x"34d43983",
          5729 => x"f9b83381",
          5730 => x"f9068107",
          5731 => x"567583f9",
          5732 => x"b834c339",
          5733 => x"83f9b833",
          5734 => x"819f0690",
          5735 => x"07567583",
          5736 => x"f9b834ff",
          5737 => x"b13980f1",
          5738 => x"0b83f9b8",
          5739 => x"34811870",
          5740 => x"81ff0659",
          5741 => x"56f4a439",
          5742 => x"83f9b833",
          5743 => x"818f0656",
          5744 => x"7583f9b8",
          5745 => x"34ff8f39",
          5746 => x"83f9b833",
          5747 => x"819f0690",
          5748 => x"07567583",
          5749 => x"f9b834fe",
          5750 => x"fd3983f9",
          5751 => x"b83381ef",
          5752 => x"0680e007",
          5753 => x"567583f9",
          5754 => x"b834feea",
          5755 => x"3983f9b8",
          5756 => x"3381cf06",
          5757 => x"80c00756",
          5758 => x"7583f9b8",
          5759 => x"34fed739",
          5760 => x"83f9b833",
          5761 => x"81af06a0",
          5762 => x"07567583",
          5763 => x"f9b834fe",
          5764 => x"c53983f9",
          5765 => x"b83381fe",
          5766 => x"06860756",
          5767 => x"7583f9b8",
          5768 => x"34feb339",
          5769 => x"83f9b833",
          5770 => x"81fc0684",
          5771 => x"07567583",
          5772 => x"f9b834fe",
          5773 => x"a13983f9",
          5774 => x"b83381fa",
          5775 => x"06820756",
          5776 => x"7583f9b8",
          5777 => x"34fe8f39",
          5778 => x"83f9b833",
          5779 => x"81f80656",
          5780 => x"7583f9b8",
          5781 => x"34fdff39",
          5782 => x"83f9b833",
          5783 => x"80f00756",
          5784 => x"7583f9b8",
          5785 => x"34fdef39",
          5786 => x"83f9b833",
          5787 => x"80f00756",
          5788 => x"7583f9b8",
          5789 => x"34fddf39",
          5790 => x"83f9b833",
          5791 => x"81df0680",
          5792 => x"d0075675",
          5793 => x"83f9b834",
          5794 => x"fdcc3983",
          5795 => x"f9b83381",
          5796 => x"bf06b007",
          5797 => x"567583f9",
          5798 => x"b834fdba",
          5799 => x"39800b83",
          5800 => x"f9bd3480",
          5801 => x"528151d2",
          5802 => x"c93fecff",
          5803 => x"3984b9f4",
          5804 => x"3383f9bc",
          5805 => x"3484b9f5",
          5806 => x"3383f9bd",
          5807 => x"3484b9f6",
          5808 => x"33597883",
          5809 => x"f9ba2380",
          5810 => x"0b84b988",
          5811 => x"0ce8c739",
          5812 => x"810b84b9",
          5813 => x"8f34800b",
          5814 => x"84ba8c0c",
          5815 => x"9c3d0d04",
          5816 => x"7783f9bd",
          5817 => x"3483f9bd",
          5818 => x"337081ff",
          5819 => x"0658ff05",
          5820 => x"56e7cf39",
          5821 => x"84b99042",
          5822 => x"9c3ddc11",
          5823 => x"53d80551",
          5824 => x"fef9833f",
          5825 => x"84ba8c08",
          5826 => x"a13884ba",
          5827 => x"8c0884b9",
          5828 => x"880c800b",
          5829 => x"84b98c34",
          5830 => x"800b84ba",
          5831 => x"8c0c9c3d",
          5832 => x"0d047783",
          5833 => x"f9bd34ef",
          5834 => x"e93984b9",
          5835 => x"8d338111",
          5836 => x"5c5c7a84",
          5837 => x"b98d347b",
          5838 => x"1083fe06",
          5839 => x"5d0280ca",
          5840 => x"052284b9",
          5841 => x"e01e2380",
          5842 => x"0b84b98c",
          5843 => x"34ca3980",
          5844 => x"0b83f9bd",
          5845 => x"34805281",
          5846 => x"51d1973f",
          5847 => x"83f9bd33",
          5848 => x"7081ff06",
          5849 => x"58ff0556",
          5850 => x"e6d83980",
          5851 => x"0b83f9bd",
          5852 => x"34805281",
          5853 => x"51d0fb3f",
          5854 => x"ef98398a",
          5855 => x"51feebde",
          5856 => x"3fef8f39",
          5857 => x"83f9bd33",
          5858 => x"ff057009",
          5859 => x"709f2c72",
          5860 => x"06585f57",
          5861 => x"f2a63975",
          5862 => x"528151d9",
          5863 => x"3984b880",
          5864 => x"33407560",
          5865 => x"27eeeb38",
          5866 => x"7583f9bd",
          5867 => x"34eee339",
          5868 => x"83f9bc33",
          5869 => x"ff057009",
          5870 => x"709f2c72",
          5871 => x"06584057",
          5872 => x"f0e23983",
          5873 => x"f9bc3381",
          5874 => x"0584b7ff",
          5875 => x"33ff1159",
          5876 => x"59567578",
          5877 => x"25f3c038",
          5878 => x"7557f3bb",
          5879 => x"3984b7ff",
          5880 => x"337081ff",
          5881 => x"06585c81",
          5882 => x"7726eea6",
          5883 => x"3883f9bc",
          5884 => x"3384b880",
          5885 => x"337081ff",
          5886 => x"0683f9bd",
          5887 => x"33717429",
          5888 => x"1187a3a0",
          5889 => x"800583f9",
          5890 => x"ba225f5f",
          5891 => x"717e2905",
          5892 => x"7083ffff",
          5893 => x"0683f892",
          5894 => x"335d5b44",
          5895 => x"425f5d77",
          5896 => x"812e81f5",
          5897 => x"387983ff",
          5898 => x"ff06ff11",
          5899 => x"5c57807b",
          5900 => x"24848938",
          5901 => x"84b7ff33",
          5902 => x"56767627",
          5903 => x"839838ff",
          5904 => x"16567583",
          5905 => x"f9ba237c",
          5906 => x"81ff06ff",
          5907 => x"11575780",
          5908 => x"762483df",
          5909 => x"3884b7ff",
          5910 => x"33567676",
          5911 => x"2782ec38",
          5912 => x"ff165675",
          5913 => x"83f9bc34",
          5914 => x"7b81ff06",
          5915 => x"83f9ba22",
          5916 => x"5757805a",
          5917 => x"76762690",
          5918 => x"38757731",
          5919 => x"81057e81",
          5920 => x"ff067171",
          5921 => x"295c5e5f",
          5922 => x"795887a3",
          5923 => x"a0805b87",
          5924 => x"a3b0807c",
          5925 => x"81ff067f",
          5926 => x"81ff0671",
          5927 => x"71291d41",
          5928 => x"42425d79",
          5929 => x"7e27ecea",
          5930 => x"388498de",
          5931 => x"1a57e0e0",
          5932 => x"17335e84",
          5933 => x"b8881e33",
          5934 => x"7b708105",
          5935 => x"5d347670",
          5936 => x"81055833",
          5937 => x"7d708105",
          5938 => x"5f348118",
          5939 => x"84b88033",
          5940 => x"84b7ff33",
          5941 => x"7171291d",
          5942 => x"59415d58",
          5943 => x"777627ec",
          5944 => x"b138e0e0",
          5945 => x"17335e84",
          5946 => x"b8881e33",
          5947 => x"7b708105",
          5948 => x"5d347670",
          5949 => x"81055833",
          5950 => x"7d708105",
          5951 => x"5f348118",
          5952 => x"84b88033",
          5953 => x"84b7ff33",
          5954 => x"7171291d",
          5955 => x"59415d58",
          5956 => x"757826ff",
          5957 => x"9938ebfa",
          5958 => x"3983f9be",
          5959 => x"17335c84",
          5960 => x"b8881c33",
          5961 => x"7b3483f9",
          5962 => x"bc3384b8",
          5963 => x"803383f9",
          5964 => x"ba2284b7",
          5965 => x"ff335f5c",
          5966 => x"5f5dfde9",
          5967 => x"3976ebd2",
          5968 => x"3884b7ff",
          5969 => x"337081ff",
          5970 => x"06ff115c",
          5971 => x"42587661",
          5972 => x"27833876",
          5973 => x"5a7983f9",
          5974 => x"ba237781",
          5975 => x"ff06ff19",
          5976 => x"585a807a",
          5977 => x"27833880",
          5978 => x"577683f9",
          5979 => x"bc3484b8",
          5980 => x"80337081",
          5981 => x"ff06ff12",
          5982 => x"52595680",
          5983 => x"7827eb8d",
          5984 => x"38805675",
          5985 => x"83f9bd34",
          5986 => x"eb883983",
          5987 => x"f9bd3381",
          5988 => x"0584b880",
          5989 => x"33ff1159",
          5990 => x"4056757f",
          5991 => x"25efca38",
          5992 => x"7557efc5",
          5993 => x"3975812e",
          5994 => x"098106f4",
          5995 => x"c03883f9",
          5996 => x"bd337081",
          5997 => x"ff0683f9",
          5998 => x"bc337a44",
          5999 => x"5d5d5776",
          6000 => x"ff2e0981",
          6001 => x"06f4b838",
          6002 => x"f6a139ff",
          6003 => x"1d567583",
          6004 => x"f9bc34fd",
          6005 => x"9339ff1a",
          6006 => x"567583f9",
          6007 => x"ba23fce7",
          6008 => x"397c7b31",
          6009 => x"567583f9",
          6010 => x"bc34f290",
          6011 => x"39777d58",
          6012 => x"56777a26",
          6013 => x"f58d3880",
          6014 => x"76708105",
          6015 => x"583483f9",
          6016 => x"b8337770",
          6017 => x"81055934",
          6018 => x"757a26f4",
          6019 => x"ec388076",
          6020 => x"70810558",
          6021 => x"3483f9b8",
          6022 => x"33777081",
          6023 => x"05593479",
          6024 => x"7627d438",
          6025 => x"f4d33979",
          6026 => x"7b315675",
          6027 => x"83f9ba23",
          6028 => x"f1a83980",
          6029 => x"0b83f9bc",
          6030 => x"34fcad39",
          6031 => x"7e83f9ba",
          6032 => x"23fc8439",
          6033 => x"800b83f9",
          6034 => x"ba23f18e",
          6035 => x"39800b83",
          6036 => x"f9bc34f1",
          6037 => x"a73983f9",
          6038 => x"be18335a",
          6039 => x"84b8881a",
          6040 => x"33773480",
          6041 => x"0b83f891",
          6042 => x"34e9a739",
          6043 => x"fd3d0d02",
          6044 => x"97053384",
          6045 => x"b8823354",
          6046 => x"5472802e",
          6047 => x"90387351",
          6048 => x"db9c3f80",
          6049 => x"0b84ba8c",
          6050 => x"0c853d0d",
          6051 => x"04765273",
          6052 => x"51d7ab3f",
          6053 => x"800b84ba",
          6054 => x"8c0c853d",
          6055 => x"0d04f33d",
          6056 => x"0d02bf05",
          6057 => x"335cff0b",
          6058 => x"83f89033",
          6059 => x"7081ff06",
          6060 => x"83f7f011",
          6061 => x"33585555",
          6062 => x"5974802e",
          6063 => x"80d63881",
          6064 => x"14567583",
          6065 => x"f8903474",
          6066 => x"597884ba",
          6067 => x"8c0c8f3d",
          6068 => x"0d0483f7",
          6069 => x"ec085482",
          6070 => x"5373802e",
          6071 => x"91387373",
          6072 => x"32703071",
          6073 => x"07700970",
          6074 => x"9f2a565d",
          6075 => x"5e587283",
          6076 => x"f7ec0cff",
          6077 => x"5980547b",
          6078 => x"812e0981",
          6079 => x"0683387b",
          6080 => x"547b8332",
          6081 => x"70307080",
          6082 => x"2576075c",
          6083 => x"5c5d7980",
          6084 => x"2e85c438",
          6085 => x"84b88033",
          6086 => x"83f9bd33",
          6087 => x"83f9bc33",
          6088 => x"72712912",
          6089 => x"87a3a080",
          6090 => x"0583f9ba",
          6091 => x"225b595d",
          6092 => x"71792905",
          6093 => x"7083ffff",
          6094 => x"0683f891",
          6095 => x"33585955",
          6096 => x"5874812e",
          6097 => x"838c3881",
          6098 => x"f0547386",
          6099 => x"ee808034",
          6100 => x"800b87c0",
          6101 => x"98880c87",
          6102 => x"c0988808",
          6103 => x"5675802e",
          6104 => x"f63886ee",
          6105 => x"80840857",
          6106 => x"7683f5bc",
          6107 => x"15348114",
          6108 => x"7081ff06",
          6109 => x"555581f9",
          6110 => x"7427cf38",
          6111 => x"805483f7",
          6112 => x"ac143370",
          6113 => x"81ff0683",
          6114 => x"f7b61633",
          6115 => x"58545572",
          6116 => x"762e85c1",
          6117 => x"387281ff",
          6118 => x"2e86b438",
          6119 => x"7483f7c0",
          6120 => x"15347581",
          6121 => x"ff065a79",
          6122 => x"81ff2e85",
          6123 => x"cd387583",
          6124 => x"f7ca1534",
          6125 => x"83f7ac14",
          6126 => x"3383f7b6",
          6127 => x"15348114",
          6128 => x"7081ff06",
          6129 => x"555e8974",
          6130 => x"27ffb338",
          6131 => x"83f7b433",
          6132 => x"70982b70",
          6133 => x"80255856",
          6134 => x"547583f7",
          6135 => x"e4347381",
          6136 => x"ff067086",
          6137 => x"2a813270",
          6138 => x"81065154",
          6139 => x"5872802e",
          6140 => x"85e73881",
          6141 => x"0b83f7e5",
          6142 => x"34730981",
          6143 => x"06537280",
          6144 => x"2e85e438",
          6145 => x"810b83f7",
          6146 => x"e634800b",
          6147 => x"83f7e533",
          6148 => x"83f7ec08",
          6149 => x"83f7e633",
          6150 => x"7083f7e8",
          6151 => x"3383f7e7",
          6152 => x"335d5d42",
          6153 => x"5e5c5e56",
          6154 => x"83f7c016",
          6155 => x"33557481",
          6156 => x"ff2e8d38",
          6157 => x"83f7d416",
          6158 => x"33547380",
          6159 => x"2e828238",
          6160 => x"83f7ca16",
          6161 => x"33537281",
          6162 => x"ff2e8b38",
          6163 => x"83f7d416",
          6164 => x"33547381",
          6165 => x"ec387481",
          6166 => x"ff065473",
          6167 => x"81ff2e8d",
          6168 => x"3883f7d4",
          6169 => x"16335372",
          6170 => x"812e81da",
          6171 => x"387481ff",
          6172 => x"06537281",
          6173 => x"ff2e848c",
          6174 => x"3883f7d4",
          6175 => x"16335481",
          6176 => x"74278480",
          6177 => x"3883f7e0",
          6178 => x"0887e805",
          6179 => x"87c0989c",
          6180 => x"08545473",
          6181 => x"732783ec",
          6182 => x"38810b87",
          6183 => x"c0989c08",
          6184 => x"83f7e00c",
          6185 => x"58811670",
          6186 => x"81ff0657",
          6187 => x"54897627",
          6188 => x"fef63876",
          6189 => x"83f7e734",
          6190 => x"7783f7e8",
          6191 => x"34fe9e19",
          6192 => x"53729c26",
          6193 => x"828b3872",
          6194 => x"101083c9",
          6195 => x"b4055a79",
          6196 => x"080483f8",
          6197 => x"94085473",
          6198 => x"802e9138",
          6199 => x"83f41487",
          6200 => x"c0989c08",
          6201 => x"5e5e7d7d",
          6202 => x"27fcdc38",
          6203 => x"800b83f8",
          6204 => x"92335454",
          6205 => x"72812e83",
          6206 => x"38745473",
          6207 => x"83f89234",
          6208 => x"87c0989c",
          6209 => x"0883f894",
          6210 => x"0c7381ff",
          6211 => x"06587781",
          6212 => x"2e943883",
          6213 => x"f9be1733",
          6214 => x"5484b888",
          6215 => x"14337634",
          6216 => x"81f054fc",
          6217 => x"a53983f7",
          6218 => x"ec085372",
          6219 => x"802e829c",
          6220 => x"3872812e",
          6221 => x"83f43880",
          6222 => x"c3763481",
          6223 => x"f054fc8a",
          6224 => x"398058fe",
          6225 => x"e0398074",
          6226 => x"56578359",
          6227 => x"7c812e9b",
          6228 => x"3879772e",
          6229 => x"09810683",
          6230 => x"b4387d81",
          6231 => x"2e80ed38",
          6232 => x"79812e80",
          6233 => x"d7387981",
          6234 => x"ff065987",
          6235 => x"77277598",
          6236 => x"2b545472",
          6237 => x"8025a138",
          6238 => x"73802e9c",
          6239 => x"38811770",
          6240 => x"81ff0676",
          6241 => x"1081fe06",
          6242 => x"87722771",
          6243 => x"982b5753",
          6244 => x"57585480",
          6245 => x"7324e138",
          6246 => x"78101010",
          6247 => x"79100576",
          6248 => x"11832b78",
          6249 => x"0583f49c",
          6250 => x"0570335b",
          6251 => x"56547887",
          6252 => x"c0989c08",
          6253 => x"83f7e00c",
          6254 => x"57fdea39",
          6255 => x"80597d81",
          6256 => x"2effa838",
          6257 => x"7981ff06",
          6258 => x"59ffa039",
          6259 => x"8259ff9b",
          6260 => x"3978ff2e",
          6261 => x"fa9f3880",
          6262 => x"0b84b882",
          6263 => x"33545472",
          6264 => x"812e83e8",
          6265 => x"387b8232",
          6266 => x"70307080",
          6267 => x"25760740",
          6268 => x"59567d8a",
          6269 => x"387b832e",
          6270 => x"098106f9",
          6271 => x"cc3878ff",
          6272 => x"2ef9c638",
          6273 => x"80537210",
          6274 => x"101083f8",
          6275 => x"98057033",
          6276 => x"5d54787c",
          6277 => x"2e83ba38",
          6278 => x"81137081",
          6279 => x"ff065457",
          6280 => x"937327e2",
          6281 => x"3884b883",
          6282 => x"33537280",
          6283 => x"2ef99a38",
          6284 => x"84b88433",
          6285 => x"5574f991",
          6286 => x"387881ff",
          6287 => x"06528251",
          6288 => x"ccd43f78",
          6289 => x"84ba8c0c",
          6290 => x"8f3d0d04",
          6291 => x"be763481",
          6292 => x"f054f9f6",
          6293 => x"397281ff",
          6294 => x"2e923883",
          6295 => x"f7d41433",
          6296 => x"81055b7a",
          6297 => x"83f7d415",
          6298 => x"34fac939",
          6299 => x"800b83f7",
          6300 => x"d41534ff",
          6301 => x"0b83f7c0",
          6302 => x"1534ff0b",
          6303 => x"83f7ca15",
          6304 => x"34fab139",
          6305 => x"7481ff06",
          6306 => x"537281ff",
          6307 => x"2efc9638",
          6308 => x"83f7d416",
          6309 => x"33558175",
          6310 => x"27fc8a38",
          6311 => x"7781ff06",
          6312 => x"5473812e",
          6313 => x"098106fb",
          6314 => x"fc3883f7",
          6315 => x"e00881fa",
          6316 => x"0587c098",
          6317 => x"9c085455",
          6318 => x"747327fb",
          6319 => x"e83887c0",
          6320 => x"989c0883",
          6321 => x"f7e00c76",
          6322 => x"81ff0659",
          6323 => x"fbd739ff",
          6324 => x"0b83f7c0",
          6325 => x"1534f9ca",
          6326 => x"397283f7",
          6327 => x"e5347309",
          6328 => x"81065372",
          6329 => x"fa9e3872",
          6330 => x"83f7e634",
          6331 => x"800b83f7",
          6332 => x"e53383f7",
          6333 => x"ec0883f7",
          6334 => x"e6337083",
          6335 => x"f7e83383",
          6336 => x"f7e7335d",
          6337 => x"5d425e5c",
          6338 => x"5e56fa9c",
          6339 => x"3979822e",
          6340 => x"098106fc",
          6341 => x"cb387a59",
          6342 => x"7a812efc",
          6343 => x"ce387981",
          6344 => x"2e098106",
          6345 => x"fcc038fd",
          6346 => x"9339ef76",
          6347 => x"3481f054",
          6348 => x"f8983980",
          6349 => x"0b84b883",
          6350 => x"33575475",
          6351 => x"83388154",
          6352 => x"7384b883",
          6353 => x"34ff59f7",
          6354 => x"ac39800b",
          6355 => x"84b88233",
          6356 => x"58547683",
          6357 => x"38815473",
          6358 => x"84b88234",
          6359 => x"ff59f795",
          6360 => x"39815383",
          6361 => x"f7ec0884",
          6362 => x"2ef78338",
          6363 => x"840b83f7",
          6364 => x"ec0cf6ff",
          6365 => x"3984b7ff",
          6366 => x"337081ff",
          6367 => x"06ff1157",
          6368 => x"5a548079",
          6369 => x"27833880",
          6370 => x"557483f9",
          6371 => x"ba237381",
          6372 => x"ff06ff15",
          6373 => x"55538073",
          6374 => x"27833880",
          6375 => x"547383f9",
          6376 => x"bc3484b8",
          6377 => x"80337081",
          6378 => x"ff0656ff",
          6379 => x"05538075",
          6380 => x"27833880",
          6381 => x"537283f9",
          6382 => x"bd34ff59",
          6383 => x"f6b73981",
          6384 => x"528351ff",
          6385 => x"baa53fff",
          6386 => x"59f6aa39",
          6387 => x"7254fc95",
          6388 => x"39841408",
          6389 => x"5283f7f0",
          6390 => x"51fedeeb",
          6391 => x"3f810b83",
          6392 => x"f8903483",
          6393 => x"f7f03359",
          6394 => x"fcbb3980",
          6395 => x"3d0d8151",
          6396 => x"f5ac3f82",
          6397 => x"3d0d04f9",
          6398 => x"3d0d800b",
          6399 => x"83f49808",
          6400 => x"545802a7",
          6401 => x"05338214",
          6402 => x"3483f498",
          6403 => x"085280e0",
          6404 => x"7234850b",
          6405 => x"83f49808",
          6406 => x"5657fe0b",
          6407 => x"81163480",
          6408 => x"0b86f080",
          6409 => x"e83487c0",
          6410 => x"989c0883",
          6411 => x"f4980856",
          6412 => x"80ce9005",
          6413 => x"5487c098",
          6414 => x"9c085387",
          6415 => x"c0989c08",
          6416 => x"5271732e",
          6417 => x"f6388115",
          6418 => x"3387c098",
          6419 => x"9c085753",
          6420 => x"75742787",
          6421 => x"387281fe",
          6422 => x"2edb3887",
          6423 => x"c098a408",
          6424 => x"52ff5671",
          6425 => x"742780cd",
          6426 => x"38725672",
          6427 => x"ff2e80c5",
          6428 => x"3887c098",
          6429 => x"9c0880ce",
          6430 => x"90055487",
          6431 => x"c0989c08",
          6432 => x"5387c098",
          6433 => x"9c085675",
          6434 => x"732ef638",
          6435 => x"81153387",
          6436 => x"c0989c08",
          6437 => x"53537174",
          6438 => x"27873872",
          6439 => x"81ff2edb",
          6440 => x"3887c098",
          6441 => x"a40852ff",
          6442 => x"56717427",
          6443 => x"a4387256",
          6444 => x"72ff2e9d",
          6445 => x"3876802e",
          6446 => x"a3387581",
          6447 => x"ff065372",
          6448 => x"fed83875",
          6449 => x"ff2e9538",
          6450 => x"7784ba8c",
          6451 => x"0c893d0d",
          6452 => x"04ff1770",
          6453 => x"81ff0658",
          6454 => x"5476df38",
          6455 => x"810b83e4",
          6456 => x"d45258fe",
          6457 => x"d78d3f77",
          6458 => x"84ba8c0c",
          6459 => x"893d0d04",
          6460 => x"f93d0d7a",
          6461 => x"028405a7",
          6462 => x"05335753",
          6463 => x"800b83f4",
          6464 => x"98087488",
          6465 => x"2b87fc80",
          6466 => x"80067076",
          6467 => x"982a0751",
          6468 => x"56565872",
          6469 => x"83163473",
          6470 => x"902a5271",
          6471 => x"84163472",
          6472 => x"902a5776",
          6473 => x"85163473",
          6474 => x"86163483",
          6475 => x"f4980853",
          6476 => x"75821434",
          6477 => x"83f49808",
          6478 => x"5280e172",
          6479 => x"34850b83",
          6480 => x"f4980856",
          6481 => x"57fe0b81",
          6482 => x"1634800b",
          6483 => x"86f080e8",
          6484 => x"3487c098",
          6485 => x"9c0883f4",
          6486 => x"98085680",
          6487 => x"ce900554",
          6488 => x"87c0989c",
          6489 => x"085387c0",
          6490 => x"989c0852",
          6491 => x"71732ef6",
          6492 => x"38811533",
          6493 => x"87c0989c",
          6494 => x"08575375",
          6495 => x"74278738",
          6496 => x"7281fe2e",
          6497 => x"db3887c0",
          6498 => x"98a40852",
          6499 => x"ff567174",
          6500 => x"2780cf38",
          6501 => x"725672ff",
          6502 => x"2e80c738",
          6503 => x"87c0989c",
          6504 => x"0880ce90",
          6505 => x"055487c0",
          6506 => x"989c0853",
          6507 => x"87c0989c",
          6508 => x"08567573",
          6509 => x"2ef63881",
          6510 => x"153387c0",
          6511 => x"989c0853",
          6512 => x"53717427",
          6513 => x"87387281",
          6514 => x"ff2edb38",
          6515 => x"87c098a4",
          6516 => x"0852ff56",
          6517 => x"71742780",
          6518 => x"df387256",
          6519 => x"72ff2e80",
          6520 => x"d7387680",
          6521 => x"2e80dd38",
          6522 => x"7581ff06",
          6523 => x"5372fed5",
          6524 => x"38755271",
          6525 => x"81ff0657",
          6526 => x"76aa3880",
          6527 => x"c6157c84",
          6528 => x"80115653",
          6529 => x"53717427",
          6530 => x"92387270",
          6531 => x"81055433",
          6532 => x"72708105",
          6533 => x"54347372",
          6534 => x"26f03877",
          6535 => x"84ba8c0c",
          6536 => x"893d0d04",
          6537 => x"810b83e4",
          6538 => x"e85258fe",
          6539 => x"d4c53f77",
          6540 => x"84ba8c0c",
          6541 => x"893d0d04",
          6542 => x"ff177081",
          6543 => x"ff065854",
          6544 => x"76ffa538",
          6545 => x"ff52ffab",
          6546 => x"39f93d0d",
          6547 => x"7a028405",
          6548 => x"a7053357",
          6549 => x"57800b83",
          6550 => x"f4980878",
          6551 => x"882b87fc",
          6552 => x"80800670",
          6553 => x"7a982a07",
          6554 => x"51565658",
          6555 => x"76831634",
          6556 => x"73902a52",
          6557 => x"71841634",
          6558 => x"76902a53",
          6559 => x"72851634",
          6560 => x"73861634",
          6561 => x"7b83f498",
          6562 => x"0880c611",
          6563 => x"84801357",
          6564 => x"55565271",
          6565 => x"74279738",
          6566 => x"71708105",
          6567 => x"53337370",
          6568 => x"81055534",
          6569 => x"737226f0",
          6570 => x"3883f498",
          6571 => x"08557582",
          6572 => x"163483f4",
          6573 => x"98085680",
          6574 => x"e2763485",
          6575 => x"0b83f498",
          6576 => x"085657fe",
          6577 => x"0b811634",
          6578 => x"800b86f0",
          6579 => x"80e83487",
          6580 => x"c0989c08",
          6581 => x"83f49808",
          6582 => x"5680ce90",
          6583 => x"055487c0",
          6584 => x"989c0853",
          6585 => x"87c0989c",
          6586 => x"08527173",
          6587 => x"2ef63881",
          6588 => x"153387c0",
          6589 => x"989c0857",
          6590 => x"53757427",
          6591 => x"87387281",
          6592 => x"fe2edb38",
          6593 => x"87c098a4",
          6594 => x"0852ff56",
          6595 => x"71742780",
          6596 => x"cd387256",
          6597 => x"72ff2e80",
          6598 => x"c53887c0",
          6599 => x"989c0880",
          6600 => x"ce900554",
          6601 => x"87c0989c",
          6602 => x"085387c0",
          6603 => x"989c0856",
          6604 => x"75732ef6",
          6605 => x"38811533",
          6606 => x"87c0989c",
          6607 => x"08535371",
          6608 => x"74278738",
          6609 => x"7281ff2e",
          6610 => x"db3887c0",
          6611 => x"98a40852",
          6612 => x"ff567174",
          6613 => x"27a93872",
          6614 => x"5672ff2e",
          6615 => x"a2387680",
          6616 => x"2ea83875",
          6617 => x"81ff0653",
          6618 => x"72fed838",
          6619 => x"757081ff",
          6620 => x"06565274",
          6621 => x"a1387784",
          6622 => x"ba8c0c89",
          6623 => x"3d0d04ff",
          6624 => x"177081ff",
          6625 => x"06585476",
          6626 => x"da38ff70",
          6627 => x"81ff0656",
          6628 => x"5274802e",
          6629 => x"e138810b",
          6630 => x"83e4fc52",
          6631 => x"58fed1d3",
          6632 => x"3f7784ba",
          6633 => x"8c0c893d",
          6634 => x"0d04fb3d",
          6635 => x"0d83f498",
          6636 => x"085180d0",
          6637 => x"7134850b",
          6638 => x"83f49808",
          6639 => x"5656fe0b",
          6640 => x"81163480",
          6641 => x"0b86f080",
          6642 => x"e83487c0",
          6643 => x"989c0883",
          6644 => x"f4980856",
          6645 => x"80ce9005",
          6646 => x"5487c098",
          6647 => x"9c085287",
          6648 => x"c0989c08",
          6649 => x"5372722e",
          6650 => x"f6388115",
          6651 => x"3387c098",
          6652 => x"9c085252",
          6653 => x"70742787",
          6654 => x"387181fe",
          6655 => x"2edb3887",
          6656 => x"c098a408",
          6657 => x"51ff5370",
          6658 => x"742780cd",
          6659 => x"38715371",
          6660 => x"ff2e80c5",
          6661 => x"3887c098",
          6662 => x"9c0880ce",
          6663 => x"90055487",
          6664 => x"c0989c08",
          6665 => x"5287c098",
          6666 => x"9c085372",
          6667 => x"722ef638",
          6668 => x"81153387",
          6669 => x"c0989c08",
          6670 => x"52527074",
          6671 => x"27873871",
          6672 => x"81ff2edb",
          6673 => x"3887c098",
          6674 => x"a40851ff",
          6675 => x"53707427",
          6676 => x"98387153",
          6677 => x"71ff2e91",
          6678 => x"3875802e",
          6679 => x"8a387281",
          6680 => x"ff065271",
          6681 => x"fed838ff",
          6682 => x"39ff1670",
          6683 => x"81ff0657",
          6684 => x"54e73980",
          6685 => x"3d0d83e5",
          6686 => x"9051fecf",
          6687 => x"f63f823d",
          6688 => x"0d04f93d",
          6689 => x"0d84b9fc",
          6690 => x"087a7131",
          6691 => x"832a7083",
          6692 => x"ffff0670",
          6693 => x"832b7311",
          6694 => x"70338112",
          6695 => x"33718b2b",
          6696 => x"71832b07",
          6697 => x"77117033",
          6698 => x"81123371",
          6699 => x"982b7190",
          6700 => x"2b075c54",
          6701 => x"4153535d",
          6702 => x"57595256",
          6703 => x"57538071",
          6704 => x"2481af38",
          6705 => x"72168211",
          6706 => x"33831233",
          6707 => x"718b2b71",
          6708 => x"832b0776",
          6709 => x"05703381",
          6710 => x"12337198",
          6711 => x"2b71902b",
          6712 => x"0757535c",
          6713 => x"52595652",
          6714 => x"80712483",
          6715 => x"9e388413",
          6716 => x"33851433",
          6717 => x"718b2b71",
          6718 => x"832b0775",
          6719 => x"0576882a",
          6720 => x"52545657",
          6721 => x"74861334",
          6722 => x"7381ff06",
          6723 => x"54738713",
          6724 => x"3484b9fc",
          6725 => x"08701784",
          6726 => x"12338513",
          6727 => x"3371882b",
          6728 => x"0770882a",
          6729 => x"5c555954",
          6730 => x"51778414",
          6731 => x"34718514",
          6732 => x"3484b9fc",
          6733 => x"08165280",
          6734 => x"0b861334",
          6735 => x"800b8713",
          6736 => x"3484b9fc",
          6737 => x"08537484",
          6738 => x"14347385",
          6739 => x"143484b9",
          6740 => x"fc081670",
          6741 => x"33811233",
          6742 => x"71882b07",
          6743 => x"82808007",
          6744 => x"70882a58",
          6745 => x"58525274",
          6746 => x"72347581",
          6747 => x"1334893d",
          6748 => x"0d048612",
          6749 => x"33871333",
          6750 => x"718b2b71",
          6751 => x"832b0775",
          6752 => x"11841633",
          6753 => x"85173371",
          6754 => x"882b0770",
          6755 => x"882a5858",
          6756 => x"54515358",
          6757 => x"58718412",
          6758 => x"34728512",
          6759 => x"3484b9fc",
          6760 => x"08701684",
          6761 => x"11338512",
          6762 => x"33718b2b",
          6763 => x"71832b07",
          6764 => x"565a5a52",
          6765 => x"72058612",
          6766 => x"33871333",
          6767 => x"71882b07",
          6768 => x"70882a52",
          6769 => x"55595277",
          6770 => x"86133472",
          6771 => x"87133484",
          6772 => x"b9fc0815",
          6773 => x"70338112",
          6774 => x"3371882b",
          6775 => x"0781ffff",
          6776 => x"0670882a",
          6777 => x"5a5a5452",
          6778 => x"76723477",
          6779 => x"81133484",
          6780 => x"b9fc0870",
          6781 => x"17703381",
          6782 => x"1233718b",
          6783 => x"2b71832b",
          6784 => x"07740570",
          6785 => x"33811233",
          6786 => x"71882b07",
          6787 => x"70832b8f",
          6788 => x"fff80677",
          6789 => x"057b882a",
          6790 => x"54525354",
          6791 => x"5c5a5754",
          6792 => x"52778214",
          6793 => x"34738314",
          6794 => x"3484b9fc",
          6795 => x"08701770",
          6796 => x"33811233",
          6797 => x"718b2b71",
          6798 => x"832b0774",
          6799 => x"05703381",
          6800 => x"12337188",
          6801 => x"2b0781ff",
          6802 => x"ff067088",
          6803 => x"2a5f5253",
          6804 => x"555a5754",
          6805 => x"52777334",
          6806 => x"70811434",
          6807 => x"84b9fc08",
          6808 => x"70178211",
          6809 => x"33831233",
          6810 => x"718b2b71",
          6811 => x"832b0774",
          6812 => x"05703381",
          6813 => x"12337198",
          6814 => x"2b71902b",
          6815 => x"0758535d",
          6816 => x"525a5753",
          6817 => x"53708025",
          6818 => x"fce43871",
          6819 => x"33811333",
          6820 => x"71882b07",
          6821 => x"82808007",
          6822 => x"70882a59",
          6823 => x"59547675",
          6824 => x"34778116",
          6825 => x"3484b9fc",
          6826 => x"08701770",
          6827 => x"33811233",
          6828 => x"718b2b71",
          6829 => x"832b0774",
          6830 => x"05821433",
          6831 => x"83153371",
          6832 => x"882b0770",
          6833 => x"882a575c",
          6834 => x"5c525856",
          6835 => x"52537282",
          6836 => x"15347583",
          6837 => x"1534893d",
          6838 => x"0d04f93d",
          6839 => x"0d7984b9",
          6840 => x"fc085858",
          6841 => x"76802e8f",
          6842 => x"3877802e",
          6843 => x"86387751",
          6844 => x"fb903f89",
          6845 => x"3d0d0484",
          6846 => x"fff40b84",
          6847 => x"b9fc0ca0",
          6848 => x"800b84b9",
          6849 => x"f8238280",
          6850 => x"80537652",
          6851 => x"84fff451",
          6852 => x"fed2ec3f",
          6853 => x"84b9fc08",
          6854 => x"55767534",
          6855 => x"810b8116",
          6856 => x"3484b9fc",
          6857 => x"08547684",
          6858 => x"1534810b",
          6859 => x"85153484",
          6860 => x"b9fc0856",
          6861 => x"76861734",
          6862 => x"810b8717",
          6863 => x"3484b9fc",
          6864 => x"0884b9f8",
          6865 => x"22ff05fe",
          6866 => x"80800770",
          6867 => x"83ffff06",
          6868 => x"70882a58",
          6869 => x"51555674",
          6870 => x"88173473",
          6871 => x"89173484",
          6872 => x"b9f82270",
          6873 => x"10101084",
          6874 => x"b9fc0805",
          6875 => x"f8055555",
          6876 => x"76821534",
          6877 => x"810b8315",
          6878 => x"34feee39",
          6879 => x"f73d0d7b",
          6880 => x"52805381",
          6881 => x"51847227",
          6882 => x"8e38fb12",
          6883 => x"832a8205",
          6884 => x"7083ffff",
          6885 => x"06515170",
          6886 => x"83ffff06",
          6887 => x"84b9fc08",
          6888 => x"84113385",
          6889 => x"12337188",
          6890 => x"2b077052",
          6891 => x"595a5855",
          6892 => x"81ffff54",
          6893 => x"75802e80",
          6894 => x"cc387510",
          6895 => x"10101770",
          6896 => x"33811233",
          6897 => x"71882b07",
          6898 => x"7081ffff",
          6899 => x"06793170",
          6900 => x"83ffff06",
          6901 => x"707a2756",
          6902 => x"535c5c54",
          6903 => x"52727427",
          6904 => x"8a387080",
          6905 => x"2e853875",
          6906 => x"73555884",
          6907 => x"12338513",
          6908 => x"3371882b",
          6909 => x"07575a75",
          6910 => x"c1387381",
          6911 => x"ffff2e85",
          6912 => x"38777454",
          6913 => x"56807683",
          6914 => x"2b781170",
          6915 => x"33811233",
          6916 => x"71882b07",
          6917 => x"7081ffff",
          6918 => x"0656565d",
          6919 => x"56595970",
          6920 => x"792e8338",
          6921 => x"81598051",
          6922 => x"74732682",
          6923 => x"8d387851",
          6924 => x"78802e82",
          6925 => x"85387275",
          6926 => x"2e828838",
          6927 => x"74167083",
          6928 => x"2b781174",
          6929 => x"82808007",
          6930 => x"70882a5b",
          6931 => x"5c56565a",
          6932 => x"76743478",
          6933 => x"81153484",
          6934 => x"b9fc0815",
          6935 => x"76882a53",
          6936 => x"53718214",
          6937 => x"34758314",
          6938 => x"3484b9fc",
          6939 => x"08701970",
          6940 => x"33811233",
          6941 => x"71882b07",
          6942 => x"70832b8f",
          6943 => x"fff80674",
          6944 => x"057e83ff",
          6945 => x"ff067088",
          6946 => x"2a5c5853",
          6947 => x"57595252",
          6948 => x"75821234",
          6949 => x"7281ff06",
          6950 => x"53728312",
          6951 => x"3484b9fc",
          6952 => x"08185475",
          6953 => x"74347281",
          6954 => x"153484b9",
          6955 => x"fc087019",
          6956 => x"86113387",
          6957 => x"1233718b",
          6958 => x"2b71832b",
          6959 => x"07740558",
          6960 => x"5c5c5357",
          6961 => x"75841534",
          6962 => x"72851534",
          6963 => x"84b9fc08",
          6964 => x"70165578",
          6965 => x"05861133",
          6966 => x"87123371",
          6967 => x"882b0770",
          6968 => x"882a5454",
          6969 => x"58597086",
          6970 => x"15347187",
          6971 => x"153484b9",
          6972 => x"fc087019",
          6973 => x"84113385",
          6974 => x"1233718b",
          6975 => x"2b71832b",
          6976 => x"07740558",
          6977 => x"5a5c5a52",
          6978 => x"75861534",
          6979 => x"72871534",
          6980 => x"84b9fc08",
          6981 => x"70165578",
          6982 => x"05841133",
          6983 => x"85123371",
          6984 => x"882b0770",
          6985 => x"882a545c",
          6986 => x"57597084",
          6987 => x"15347985",
          6988 => x"153484b9",
          6989 => x"fc081884",
          6990 => x"05517084",
          6991 => x"ba8c0c8b",
          6992 => x"3d0d0486",
          6993 => x"14338715",
          6994 => x"33718b2b",
          6995 => x"71832b07",
          6996 => x"79058417",
          6997 => x"33851833",
          6998 => x"71882b07",
          6999 => x"70882a5a",
          7000 => x"5b595354",
          7001 => x"52748412",
          7002 => x"34768512",
          7003 => x"3484b9fc",
          7004 => x"08701984",
          7005 => x"11338512",
          7006 => x"33718b2b",
          7007 => x"71832b07",
          7008 => x"74058614",
          7009 => x"33871533",
          7010 => x"71882b07",
          7011 => x"70882a58",
          7012 => x"5d5f5256",
          7013 => x"5b575270",
          7014 => x"861a3476",
          7015 => x"871a3484",
          7016 => x"b9fc0818",
          7017 => x"70338112",
          7018 => x"3371882b",
          7019 => x"0781ffff",
          7020 => x"0670882a",
          7021 => x"59575457",
          7022 => x"75773474",
          7023 => x"81183484",
          7024 => x"b9fc0818",
          7025 => x"840551fe",
          7026 => x"f139f93d",
          7027 => x"0d7984b9",
          7028 => x"fc085858",
          7029 => x"76802ea0",
          7030 => x"38775477",
          7031 => x"8a387384",
          7032 => x"ba8c0c89",
          7033 => x"3d0d0477",
          7034 => x"51fb913f",
          7035 => x"84ba8c08",
          7036 => x"84ba8c0c",
          7037 => x"893d0d04",
          7038 => x"84fff40b",
          7039 => x"84b9fc0c",
          7040 => x"a0800b84",
          7041 => x"b9f82382",
          7042 => x"80805376",
          7043 => x"5284fff4",
          7044 => x"51fecceb",
          7045 => x"3f84b9fc",
          7046 => x"08557675",
          7047 => x"34810b81",
          7048 => x"163484b9",
          7049 => x"fc085476",
          7050 => x"84153481",
          7051 => x"0b851534",
          7052 => x"84b9fc08",
          7053 => x"56768617",
          7054 => x"34810b87",
          7055 => x"173484b9",
          7056 => x"fc0884b9",
          7057 => x"f822ff05",
          7058 => x"fe808007",
          7059 => x"7083ffff",
          7060 => x"0670882a",
          7061 => x"58515556",
          7062 => x"74881734",
          7063 => x"73891734",
          7064 => x"84b9f822",
          7065 => x"70101010",
          7066 => x"84b9fc08",
          7067 => x"05f80555",
          7068 => x"55768215",
          7069 => x"34810b83",
          7070 => x"15347754",
          7071 => x"77802efe",
          7072 => x"dd38fee3",
          7073 => x"39ed3d0d",
          7074 => x"6567415f",
          7075 => x"807084b9",
          7076 => x"fc085945",
          7077 => x"4176612e",
          7078 => x"84aa387e",
          7079 => x"802e85af",
          7080 => x"387f802e",
          7081 => x"88d73881",
          7082 => x"54846027",
          7083 => x"8f387ffb",
          7084 => x"05832a82",
          7085 => x"057083ff",
          7086 => x"ff065558",
          7087 => x"7383ffff",
          7088 => x"067f7831",
          7089 => x"832a7083",
          7090 => x"ffff0670",
          7091 => x"832b7a11",
          7092 => x"70338112",
          7093 => x"3371882b",
          7094 => x"07707531",
          7095 => x"7083ffff",
          7096 => x"06701010",
          7097 => x"10fc0573",
          7098 => x"832b6111",
          7099 => x"70338112",
          7100 => x"3371882b",
          7101 => x"0770902b",
          7102 => x"70902c53",
          7103 => x"42454644",
          7104 => x"53544344",
          7105 => x"5c485952",
          7106 => x"5e5f4280",
          7107 => x"7a2485fd",
          7108 => x"38821533",
          7109 => x"83163371",
          7110 => x"882b0770",
          7111 => x"10101019",
          7112 => x"70338112",
          7113 => x"3371982b",
          7114 => x"71902b07",
          7115 => x"535c5356",
          7116 => x"56568074",
          7117 => x"2485c938",
          7118 => x"7a622782",
          7119 => x"f638631b",
          7120 => x"5877622e",
          7121 => x"87a23860",
          7122 => x"802e85f9",
          7123 => x"38601b58",
          7124 => x"77622587",
          7125 => x"be386318",
          7126 => x"59617924",
          7127 => x"92f73876",
          7128 => x"1e703381",
          7129 => x"1233718b",
          7130 => x"2b71832b",
          7131 => x"077a1170",
          7132 => x"33811233",
          7133 => x"71982b71",
          7134 => x"902b0747",
          7135 => x"43595253",
          7136 => x"575b5880",
          7137 => x"60248cba",
          7138 => x"38761e82",
          7139 => x"11338312",
          7140 => x"33718b2b",
          7141 => x"71832b07",
          7142 => x"7a118611",
          7143 => x"33871233",
          7144 => x"718b2b71",
          7145 => x"832b077e",
          7146 => x"05841433",
          7147 => x"85153371",
          7148 => x"882b0770",
          7149 => x"882a5957",
          7150 => x"48525b41",
          7151 => x"58535c59",
          7152 => x"5677841d",
          7153 => x"3479851d",
          7154 => x"3484b9fc",
          7155 => x"08701784",
          7156 => x"11338512",
          7157 => x"33718b2b",
          7158 => x"71832b07",
          7159 => x"74058614",
          7160 => x"33871533",
          7161 => x"71882b07",
          7162 => x"70882a5f",
          7163 => x"425e5240",
          7164 => x"57415777",
          7165 => x"8616347b",
          7166 => x"87163484",
          7167 => x"b9fc0816",
          7168 => x"70338112",
          7169 => x"3371882b",
          7170 => x"0781ffff",
          7171 => x"0670882a",
          7172 => x"5a5c5e59",
          7173 => x"76793479",
          7174 => x"811a3484",
          7175 => x"b9fc0870",
          7176 => x"1f821133",
          7177 => x"83123371",
          7178 => x"8b2b7183",
          7179 => x"2b077405",
          7180 => x"73338115",
          7181 => x"3371882b",
          7182 => x"0770882a",
          7183 => x"415c455d",
          7184 => x"5f5a5555",
          7185 => x"79793475",
          7186 => x"811a3484",
          7187 => x"b9fc0870",
          7188 => x"1f703381",
          7189 => x"1233718b",
          7190 => x"2b71832b",
          7191 => x"07740582",
          7192 => x"14338315",
          7193 => x"3371882b",
          7194 => x"0770882a",
          7195 => x"415c455d",
          7196 => x"5f5a5555",
          7197 => x"79821a34",
          7198 => x"75831a34",
          7199 => x"84b9fc08",
          7200 => x"701f8211",
          7201 => x"33831233",
          7202 => x"71882b07",
          7203 => x"66576256",
          7204 => x"70832b42",
          7205 => x"525a5d7e",
          7206 => x"05840551",
          7207 => x"fec4a33f",
          7208 => x"84b9fc08",
          7209 => x"1e840561",
          7210 => x"65051c70",
          7211 => x"83ffff06",
          7212 => x"5d445f7a",
          7213 => x"622681b6",
          7214 => x"387e5473",
          7215 => x"84ba8c0c",
          7216 => x"953d0d04",
          7217 => x"84fff40b",
          7218 => x"84b9fc0c",
          7219 => x"a0800b84",
          7220 => x"b9f82382",
          7221 => x"80805360",
          7222 => x"5284fff4",
          7223 => x"51fec79f",
          7224 => x"3f84b9fc",
          7225 => x"085e607e",
          7226 => x"34810b81",
          7227 => x"1f3484b9",
          7228 => x"fc085d60",
          7229 => x"841e3481",
          7230 => x"0b851e34",
          7231 => x"84b9fc08",
          7232 => x"5c60861d",
          7233 => x"34810b87",
          7234 => x"1d3484b9",
          7235 => x"fc0884b9",
          7236 => x"f822ff05",
          7237 => x"fe808007",
          7238 => x"7083ffff",
          7239 => x"0670882a",
          7240 => x"5c5a5b57",
          7241 => x"78881834",
          7242 => x"77891834",
          7243 => x"84b9f822",
          7244 => x"70101010",
          7245 => x"84b9fc08",
          7246 => x"05f80555",
          7247 => x"56608215",
          7248 => x"34810b83",
          7249 => x"153484b9",
          7250 => x"fc08577e",
          7251 => x"fad33876",
          7252 => x"802e828c",
          7253 => x"387e547f",
          7254 => x"802efedf",
          7255 => x"387f51f4",
          7256 => x"9b3f84ba",
          7257 => x"8c0884ba",
          7258 => x"8c0c953d",
          7259 => x"0d04611c",
          7260 => x"84b9fc08",
          7261 => x"71832b71",
          7262 => x"115e447f",
          7263 => x"05703381",
          7264 => x"12337188",
          7265 => x"2b0781ff",
          7266 => x"ff067088",
          7267 => x"2a48445b",
          7268 => x"5e40637b",
          7269 => x"3460811c",
          7270 => x"346184b9",
          7271 => x"fc08057c",
          7272 => x"882a5758",
          7273 => x"75821934",
          7274 => x"7b831934",
          7275 => x"84b9fc08",
          7276 => x"701f7033",
          7277 => x"81123371",
          7278 => x"882b0770",
          7279 => x"832b8fff",
          7280 => x"f8067405",
          7281 => x"6483ffff",
          7282 => x"0670882a",
          7283 => x"4a5c4757",
          7284 => x"5e5b5d63",
          7285 => x"63820534",
          7286 => x"7681ff06",
          7287 => x"41606383",
          7288 => x"053484b9",
          7289 => x"fc081e5b",
          7290 => x"637b3460",
          7291 => x"811c3461",
          7292 => x"84b9fc08",
          7293 => x"05840551",
          7294 => x"ed883f7e",
          7295 => x"54fdbc39",
          7296 => x"7b753170",
          7297 => x"83ffff06",
          7298 => x"4254faac",
          7299 => x"397781ff",
          7300 => x"ff067631",
          7301 => x"7083ffff",
          7302 => x"06821733",
          7303 => x"83183371",
          7304 => x"882b0770",
          7305 => x"1010101b",
          7306 => x"70338112",
          7307 => x"3371982b",
          7308 => x"71902b07",
          7309 => x"535e5354",
          7310 => x"58584554",
          7311 => x"738025f9",
          7312 => x"f738ffbc",
          7313 => x"39617824",
          7314 => x"fa833880",
          7315 => x"7a248b8f",
          7316 => x"387783ff",
          7317 => x"ff065b61",
          7318 => x"7b27fcdd",
          7319 => x"38fe8f39",
          7320 => x"84fff40b",
          7321 => x"84b9fc0c",
          7322 => x"a0800b84",
          7323 => x"b9f82382",
          7324 => x"8080537e",
          7325 => x"5284fff4",
          7326 => x"51fec483",
          7327 => x"3f84b9fc",
          7328 => x"085a7e7a",
          7329 => x"34810b81",
          7330 => x"1b3484b9",
          7331 => x"fc08597e",
          7332 => x"841a3481",
          7333 => x"0b851a34",
          7334 => x"84b9fc08",
          7335 => x"587e8619",
          7336 => x"34810b87",
          7337 => x"193484b9",
          7338 => x"fc0884b9",
          7339 => x"f822ff05",
          7340 => x"fe808007",
          7341 => x"7083ffff",
          7342 => x"0670882a",
          7343 => x"58565744",
          7344 => x"74648805",
          7345 => x"34736489",
          7346 => x"053484b9",
          7347 => x"f8227010",
          7348 => x"101084b9",
          7349 => x"fc0805f8",
          7350 => x"0542437e",
          7351 => x"61820534",
          7352 => x"81618305",
          7353 => x"34fcee39",
          7354 => x"807a2483",
          7355 => x"de386183",
          7356 => x"ffff065b",
          7357 => x"617b27fb",
          7358 => x"c038fcf2",
          7359 => x"3976802e",
          7360 => x"82bd387e",
          7361 => x"51eafb3f",
          7362 => x"7f547384",
          7363 => x"ba8c0c95",
          7364 => x"3d0d0476",
          7365 => x"1e821133",
          7366 => x"83123371",
          7367 => x"8b2b7183",
          7368 => x"2b077a11",
          7369 => x"86113387",
          7370 => x"1233718b",
          7371 => x"2b71832b",
          7372 => x"077e0584",
          7373 => x"14338515",
          7374 => x"3371882b",
          7375 => x"0770882a",
          7376 => x"43444556",
          7377 => x"5b465853",
          7378 => x"5c455678",
          7379 => x"64840534",
          7380 => x"7a648505",
          7381 => x"3484b9fc",
          7382 => x"08701784",
          7383 => x"11338512",
          7384 => x"33718b2b",
          7385 => x"71832b07",
          7386 => x"74058614",
          7387 => x"33871533",
          7388 => x"71882b07",
          7389 => x"70882a5b",
          7390 => x"4142485d",
          7391 => x"595d4173",
          7392 => x"64860534",
          7393 => x"7a648705",
          7394 => x"3484b9fc",
          7395 => x"08167033",
          7396 => x"81123371",
          7397 => x"882b0781",
          7398 => x"ffff0670",
          7399 => x"882a5f5c",
          7400 => x"5a5d7b7d",
          7401 => x"3479811e",
          7402 => x"3484b9fc",
          7403 => x"08701f82",
          7404 => x"11338312",
          7405 => x"33718b2b",
          7406 => x"71832b07",
          7407 => x"74057333",
          7408 => x"81153371",
          7409 => x"882b0770",
          7410 => x"882a5e5c",
          7411 => x"5e404357",
          7412 => x"4554767c",
          7413 => x"3475811d",
          7414 => x"3484b9fc",
          7415 => x"08701f70",
          7416 => x"33811233",
          7417 => x"718b2b71",
          7418 => x"832b0774",
          7419 => x"05821433",
          7420 => x"83153371",
          7421 => x"882b0770",
          7422 => x"882a4047",
          7423 => x"405b405c",
          7424 => x"55557882",
          7425 => x"18346083",
          7426 => x"183484b9",
          7427 => x"fc08701f",
          7428 => x"82113383",
          7429 => x"12337188",
          7430 => x"2b076657",
          7431 => x"62567083",
          7432 => x"2b425258",
          7433 => x"5d7e0584",
          7434 => x"0551febd",
          7435 => x"953f84b9",
          7436 => x"fc081e84",
          7437 => x"057883ff",
          7438 => x"ff065c5f",
          7439 => x"fc993984",
          7440 => x"fff40b84",
          7441 => x"b9fc0ca0",
          7442 => x"800b84b9",
          7443 => x"f8238280",
          7444 => x"80537f52",
          7445 => x"84fff451",
          7446 => x"fec0a43f",
          7447 => x"84b9fc08",
          7448 => x"567f7634",
          7449 => x"810b8117",
          7450 => x"3484b9fc",
          7451 => x"08557f84",
          7452 => x"1634810b",
          7453 => x"85163484",
          7454 => x"b9fc0854",
          7455 => x"7f861534",
          7456 => x"810b8715",
          7457 => x"3484b9fc",
          7458 => x"0884b9f8",
          7459 => x"22ff05fe",
          7460 => x"80800770",
          7461 => x"83ffff06",
          7462 => x"70882a45",
          7463 => x"43445e61",
          7464 => x"881f3460",
          7465 => x"891f3484",
          7466 => x"b9f82270",
          7467 => x"10101084",
          7468 => x"b9fc0805",
          7469 => x"f8055c5d",
          7470 => x"7f821c34",
          7471 => x"810b831c",
          7472 => x"347e51e7",
          7473 => x"bd3f7f54",
          7474 => x"fcc03986",
          7475 => x"1933871a",
          7476 => x"33718b2b",
          7477 => x"71832b07",
          7478 => x"7905841c",
          7479 => x"33851d33",
          7480 => x"71882b07",
          7481 => x"70882a5c",
          7482 => x"485e4359",
          7483 => x"55766184",
          7484 => x"05346361",
          7485 => x"85053484",
          7486 => x"b9fc0870",
          7487 => x"1e841133",
          7488 => x"85123371",
          7489 => x"8b2b7183",
          7490 => x"2b077405",
          7491 => x"86143387",
          7492 => x"15337188",
          7493 => x"2b077088",
          7494 => x"2a415f48",
          7495 => x"48595659",
          7496 => x"40796486",
          7497 => x"05347864",
          7498 => x"87053484",
          7499 => x"b9fc081d",
          7500 => x"70338112",
          7501 => x"3371882b",
          7502 => x"0781ffff",
          7503 => x"0670882a",
          7504 => x"59425858",
          7505 => x"7578347f",
          7506 => x"81193484",
          7507 => x"b9fc0870",
          7508 => x"1f703381",
          7509 => x"1233718b",
          7510 => x"2b71832b",
          7511 => x"07740570",
          7512 => x"33811233",
          7513 => x"71882b07",
          7514 => x"70832b8f",
          7515 => x"fff80677",
          7516 => x"0563882a",
          7517 => x"485d5d5a",
          7518 => x"5d405d44",
          7519 => x"417f8217",
          7520 => x"347b8317",
          7521 => x"3484b9fc",
          7522 => x"08701f70",
          7523 => x"33811233",
          7524 => x"718b2b71",
          7525 => x"832b0774",
          7526 => x"05703381",
          7527 => x"12337188",
          7528 => x"2b0781ff",
          7529 => x"ff067088",
          7530 => x"2a485d5e",
          7531 => x"5e465a41",
          7532 => x"5b606034",
          7533 => x"76608105",
          7534 => x"346183ff",
          7535 => x"ff065bfa",
          7536 => x"b3398615",
          7537 => x"33871633",
          7538 => x"718b2b71",
          7539 => x"832b0779",
          7540 => x"05841833",
          7541 => x"85193371",
          7542 => x"882b0770",
          7543 => x"882a5e5e",
          7544 => x"5a52415d",
          7545 => x"78841e34",
          7546 => x"79851e34",
          7547 => x"84b9fc08",
          7548 => x"70198411",
          7549 => x"33851233",
          7550 => x"718b2b71",
          7551 => x"832b0774",
          7552 => x"05861433",
          7553 => x"87153371",
          7554 => x"882b0770",
          7555 => x"882a4456",
          7556 => x"5e525a42",
          7557 => x"55567c60",
          7558 => x"86053475",
          7559 => x"60870534",
          7560 => x"84b9fc08",
          7561 => x"18703381",
          7562 => x"12337188",
          7563 => x"2b0781ff",
          7564 => x"ff067088",
          7565 => x"2a5b5b58",
          7566 => x"55777534",
          7567 => x"78811634",
          7568 => x"84b9fc08",
          7569 => x"701f7033",
          7570 => x"81123371",
          7571 => x"8b2b7183",
          7572 => x"2b077405",
          7573 => x"70338112",
          7574 => x"3371882b",
          7575 => x"0770832b",
          7576 => x"8ffff806",
          7577 => x"77056388",
          7578 => x"2a56545f",
          7579 => x"5f585942",
          7580 => x"5e557f82",
          7581 => x"17347b83",
          7582 => x"173484b9",
          7583 => x"fc08701f",
          7584 => x"70338112",
          7585 => x"33718b2b",
          7586 => x"71832b07",
          7587 => x"74057033",
          7588 => x"81123371",
          7589 => x"882b0781",
          7590 => x"ffff0670",
          7591 => x"882a5d54",
          7592 => x"5e585b59",
          7593 => x"5d55757c",
          7594 => x"3476811d",
          7595 => x"3484b9fc",
          7596 => x"08701f82",
          7597 => x"11338312",
          7598 => x"33718b2b",
          7599 => x"71832b07",
          7600 => x"74118611",
          7601 => x"33871233",
          7602 => x"718b2b71",
          7603 => x"832b0778",
          7604 => x"05841433",
          7605 => x"85153371",
          7606 => x"882b0770",
          7607 => x"882a5957",
          7608 => x"49525c42",
          7609 => x"59535d5a",
          7610 => x"57577784",
          7611 => x"1d347985",
          7612 => x"1d3484b9",
          7613 => x"fc087017",
          7614 => x"84113385",
          7615 => x"1233718b",
          7616 => x"2b71832b",
          7617 => x"07740586",
          7618 => x"14338715",
          7619 => x"3371882b",
          7620 => x"0770882a",
          7621 => x"5f425e52",
          7622 => x"40574157",
          7623 => x"77861634",
          7624 => x"7b871634",
          7625 => x"84b9fc08",
          7626 => x"16703381",
          7627 => x"12337188",
          7628 => x"2b0781ff",
          7629 => x"ff067088",
          7630 => x"2a5a5c5e",
          7631 => x"59767934",
          7632 => x"79811a34",
          7633 => x"84b9fc08",
          7634 => x"701f8211",
          7635 => x"33831233",
          7636 => x"718b2b71",
          7637 => x"832b0774",
          7638 => x"05733381",
          7639 => x"15337188",
          7640 => x"2b077088",
          7641 => x"2a415c45",
          7642 => x"5d5f5a55",
          7643 => x"55797934",
          7644 => x"75811a34",
          7645 => x"84b9fc08",
          7646 => x"701f7033",
          7647 => x"81123371",
          7648 => x"8b2b7183",
          7649 => x"2b077405",
          7650 => x"82143383",
          7651 => x"15337188",
          7652 => x"2b077088",
          7653 => x"2a415c45",
          7654 => x"5d5f5a55",
          7655 => x"5579821a",
          7656 => x"3475831a",
          7657 => x"3484b9fc",
          7658 => x"08701f82",
          7659 => x"11338312",
          7660 => x"3371882b",
          7661 => x"07665762",
          7662 => x"5670832b",
          7663 => x"42525a5d",
          7664 => x"7e058405",
          7665 => x"51feb5fa",
          7666 => x"3f84b9fc",
          7667 => x"081e8405",
          7668 => x"6165051c",
          7669 => x"7083ffff",
          7670 => x"065d445f",
          7671 => x"f1d53986",
          7672 => x"1933871a",
          7673 => x"33718b2b",
          7674 => x"71832b07",
          7675 => x"7905841c",
          7676 => x"33851d33",
          7677 => x"71882b07",
          7678 => x"70882a40",
          7679 => x"485d4341",
          7680 => x"557a6184",
          7681 => x"05346361",
          7682 => x"85053484",
          7683 => x"b9fc0870",
          7684 => x"1e841133",
          7685 => x"85123371",
          7686 => x"8b2b7183",
          7687 => x"2b077405",
          7688 => x"86143387",
          7689 => x"15337188",
          7690 => x"2b077088",
          7691 => x"2a5b415f",
          7692 => x"485c5941",
          7693 => x"56736486",
          7694 => x"05347a64",
          7695 => x"87053484",
          7696 => x"b9fc081d",
          7697 => x"70338112",
          7698 => x"3371882b",
          7699 => x"0781ffff",
          7700 => x"0670882a",
          7701 => x"5c5f4255",
          7702 => x"7875347c",
          7703 => x"81163484",
          7704 => x"b9fc0870",
          7705 => x"1f703381",
          7706 => x"1233718b",
          7707 => x"2b71832b",
          7708 => x"07740570",
          7709 => x"33811233",
          7710 => x"71882b07",
          7711 => x"70832b8f",
          7712 => x"fff80677",
          7713 => x"0563882a",
          7714 => x"5d445c49",
          7715 => x"585e4558",
          7716 => x"4074821e",
          7717 => x"347b831e",
          7718 => x"3484b9fc",
          7719 => x"08701f70",
          7720 => x"33811233",
          7721 => x"718b2b71",
          7722 => x"832b0774",
          7723 => x"05703381",
          7724 => x"12337188",
          7725 => x"2b0781ff",
          7726 => x"ff067088",
          7727 => x"2a475f49",
          7728 => x"5846595e",
          7729 => x"5b7f7d34",
          7730 => x"78811e34",
          7731 => x"7783ffff",
          7732 => x"065bf383",
          7733 => x"397e6052",
          7734 => x"54e5a13f",
          7735 => x"84ba8c08",
          7736 => x"5f84ba8c",
          7737 => x"08802e93",
          7738 => x"38625373",
          7739 => x"5284ba8c",
          7740 => x"0851feb4",
          7741 => x"f53f7351",
          7742 => x"df883f61",
          7743 => x"5b617b27",
          7744 => x"efb738f0",
          7745 => x"e939f93d",
          7746 => x"0d7a7a29",
          7747 => x"84b9fc08",
          7748 => x"58587680",
          7749 => x"2eb73877",
          7750 => x"54778a38",
          7751 => x"7384ba8c",
          7752 => x"0c893d0d",
          7753 => x"047751e4",
          7754 => x"d33f84ba",
          7755 => x"8c085484",
          7756 => x"ba8c0880",
          7757 => x"2ee63877",
          7758 => x"53805284",
          7759 => x"ba8c0851",
          7760 => x"feb6bc3f",
          7761 => x"7384ba8c",
          7762 => x"0c893d0d",
          7763 => x"0484fff4",
          7764 => x"0b84b9fc",
          7765 => x"0ca0800b",
          7766 => x"84b9f823",
          7767 => x"82808053",
          7768 => x"765284ff",
          7769 => x"f451feb6",
          7770 => x"963f84b9",
          7771 => x"fc085576",
          7772 => x"7534810b",
          7773 => x"81163484",
          7774 => x"b9fc0854",
          7775 => x"76841534",
          7776 => x"810b8515",
          7777 => x"3484b9fc",
          7778 => x"08567686",
          7779 => x"1734810b",
          7780 => x"87173484",
          7781 => x"b9fc0884",
          7782 => x"b9f822ff",
          7783 => x"05fe8080",
          7784 => x"077083ff",
          7785 => x"ff067088",
          7786 => x"2a585155",
          7787 => x"56748817",
          7788 => x"34738917",
          7789 => x"3484b9f8",
          7790 => x"22701010",
          7791 => x"1084b9fc",
          7792 => x"0805f805",
          7793 => x"55557682",
          7794 => x"1534810b",
          7795 => x"83153477",
          7796 => x"5477802e",
          7797 => x"fec638fe",
          7798 => x"cc39ff3d",
          7799 => x"0d028f05",
          7800 => x"33518152",
          7801 => x"70722687",
          7802 => x"3884ba88",
          7803 => x"11335271",
          7804 => x"84ba8c0c",
          7805 => x"833d0d04",
          7806 => x"fe3d0d02",
          7807 => x"93053352",
          7808 => x"83537181",
          7809 => x"269d3871",
          7810 => x"51d3ec3f",
          7811 => x"84ba8c08",
          7812 => x"81ff0653",
          7813 => x"72873872",
          7814 => x"84ba8813",
          7815 => x"3484ba88",
          7816 => x"12335372",
          7817 => x"84ba8c0c",
          7818 => x"843d0d04",
          7819 => x"f73d0d7c",
          7820 => x"7e60028c",
          7821 => x"05af0533",
          7822 => x"5a5c5759",
          7823 => x"81547674",
          7824 => x"26873884",
          7825 => x"ba881733",
          7826 => x"54738106",
          7827 => x"54835573",
          7828 => x"bd387358",
          7829 => x"850b87c0",
          7830 => x"988c0c78",
          7831 => x"53755276",
          7832 => x"51d58d3f",
          7833 => x"84ba8c08",
          7834 => x"81ff0655",
          7835 => x"74802ea7",
          7836 => x"3887c098",
          7837 => x"8c085473",
          7838 => x"e2387978",
          7839 => x"26d63874",
          7840 => x"fc808006",
          7841 => x"5473802e",
          7842 => x"83388154",
          7843 => x"73557484",
          7844 => x"ba8c0c8b",
          7845 => x"3d0d0484",
          7846 => x"80168119",
          7847 => x"7081ff06",
          7848 => x"5a555679",
          7849 => x"7826ffac",
          7850 => x"38d539f7",
          7851 => x"3d0d7c7e",
          7852 => x"60028c05",
          7853 => x"af05335a",
          7854 => x"5c575981",
          7855 => x"54767426",
          7856 => x"873884ba",
          7857 => x"88173354",
          7858 => x"73810654",
          7859 => x"835573bd",
          7860 => x"38735885",
          7861 => x"0b87c098",
          7862 => x"8c0c7853",
          7863 => x"75527651",
          7864 => x"d6e73f84",
          7865 => x"ba8c0881",
          7866 => x"ff065574",
          7867 => x"802ea738",
          7868 => x"87c0988c",
          7869 => x"085473e2",
          7870 => x"38797826",
          7871 => x"d63874fc",
          7872 => x"80800654",
          7873 => x"73802e83",
          7874 => x"38815473",
          7875 => x"557484ba",
          7876 => x"8c0c8b3d",
          7877 => x"0d048480",
          7878 => x"16811970",
          7879 => x"81ff065a",
          7880 => x"55567978",
          7881 => x"26ffac38",
          7882 => x"d539fc3d",
          7883 => x"0d780284",
          7884 => x"059b0533",
          7885 => x"0288059f",
          7886 => x"05335353",
          7887 => x"55815371",
          7888 => x"73268738",
          7889 => x"84ba8812",
          7890 => x"33537281",
          7891 => x"06548353",
          7892 => x"739b3885",
          7893 => x"0b87c098",
          7894 => x"8c0c8153",
          7895 => x"70732e96",
          7896 => x"38727125",
          7897 => x"ad387083",
          7898 => x"2e9a3884",
          7899 => x"537284ba",
          7900 => x"8c0c863d",
          7901 => x"0d048880",
          7902 => x"0a750c73",
          7903 => x"84ba8c0c",
          7904 => x"863d0d04",
          7905 => x"8180750c",
          7906 => x"800b84ba",
          7907 => x"8c0c863d",
          7908 => x"0d047184",
          7909 => x"2b87c092",
          7910 => x"8c115354",
          7911 => x"70cd3871",
          7912 => x"0870812a",
          7913 => x"81065151",
          7914 => x"70802e8a",
          7915 => x"3887c098",
          7916 => x"8c085574",
          7917 => x"ea3887c0",
          7918 => x"988c0851",
          7919 => x"70ca3881",
          7920 => x"720c87c0",
          7921 => x"928c1452",
          7922 => x"71088206",
          7923 => x"5473802e",
          7924 => x"ff9b3871",
          7925 => x"08820654",
          7926 => x"73ee38ff",
          7927 => x"9039f63d",
          7928 => x"0d7c5880",
          7929 => x"0b831933",
          7930 => x"715b5657",
          7931 => x"74772e09",
          7932 => x"8106a838",
          7933 => x"77335675",
          7934 => x"832e8187",
          7935 => x"38805380",
          7936 => x"52811833",
          7937 => x"51fea33f",
          7938 => x"84ba8c08",
          7939 => x"802e8338",
          7940 => x"81597884",
          7941 => x"ba8c0c8c",
          7942 => x"3d0d0481",
          7943 => x"54b41808",
          7944 => x"53b81870",
          7945 => x"53811933",
          7946 => x"525afcff",
          7947 => x"3f815984",
          7948 => x"ba8c0877",
          7949 => x"2e098106",
          7950 => x"d93884ba",
          7951 => x"8c088319",
          7952 => x"34b41808",
          7953 => x"70a81a08",
          7954 => x"31a01a08",
          7955 => x"84ba8c08",
          7956 => x"5c58565b",
          7957 => x"747627ff",
          7958 => x"9b388218",
          7959 => x"33557482",
          7960 => x"2e098106",
          7961 => x"ff8e3881",
          7962 => x"54751b53",
          7963 => x"79528118",
          7964 => x"3351fcb7",
          7965 => x"3f767833",
          7966 => x"57597583",
          7967 => x"2e098106",
          7968 => x"fefb3884",
          7969 => x"18335776",
          7970 => x"812e0981",
          7971 => x"06feee38",
          7972 => x"b8185a84",
          7973 => x"807a5657",
          7974 => x"80757081",
          7975 => x"055734ff",
          7976 => x"175776f4",
          7977 => x"3880d50b",
          7978 => x"84b61934",
          7979 => x"ffaa0b84",
          7980 => x"b7193480",
          7981 => x"d27a3480",
          7982 => x"d20bb919",
          7983 => x"3480e10b",
          7984 => x"ba193480",
          7985 => x"c10bbb19",
          7986 => x"3480f20b",
          7987 => x"849c1934",
          7988 => x"80f20b84",
          7989 => x"9d193480",
          7990 => x"c10b849e",
          7991 => x"193480e1",
          7992 => x"0b849f19",
          7993 => x"34941808",
          7994 => x"557484a0",
          7995 => x"19347488",
          7996 => x"2a5b7a84",
          7997 => x"a1193474",
          7998 => x"902a5675",
          7999 => x"84a21934",
          8000 => x"74982a5b",
          8001 => x"7a84a319",
          8002 => x"34901808",
          8003 => x"5b7a84a4",
          8004 => x"19347a88",
          8005 => x"2a557484",
          8006 => x"a519347a",
          8007 => x"902a5675",
          8008 => x"84a61934",
          8009 => x"7a982a55",
          8010 => x"7484a719",
          8011 => x"34a41808",
          8012 => x"810570b4",
          8013 => x"1a0c5b81",
          8014 => x"547a5379",
          8015 => x"52811833",
          8016 => x"51fae83f",
          8017 => x"76841934",
          8018 => x"80538052",
          8019 => x"81183351",
          8020 => x"fbd83f84",
          8021 => x"ba8c0880",
          8022 => x"2efdb738",
          8023 => x"fdb239f3",
          8024 => x"3d0d6060",
          8025 => x"70085956",
          8026 => x"56817627",
          8027 => x"88389c17",
          8028 => x"0876268c",
          8029 => x"38815877",
          8030 => x"84ba8c0c",
          8031 => x"8f3d0d04",
          8032 => x"ff773356",
          8033 => x"5874822e",
          8034 => x"81cc3874",
          8035 => x"822482a5",
          8036 => x"3874812e",
          8037 => x"098106dd",
          8038 => x"3875812a",
          8039 => x"1670892a",
          8040 => x"a8190805",
          8041 => x"5a5a805b",
          8042 => x"b4170879",
          8043 => x"2eb03883",
          8044 => x"17335c7b",
          8045 => x"7b2e0981",
          8046 => x"0683de38",
          8047 => x"81547853",
          8048 => x"b8175281",
          8049 => x"173351f8",
          8050 => x"e33f84ba",
          8051 => x"8c08802e",
          8052 => x"8538ff59",
          8053 => x"815b78b4",
          8054 => x"180c7aff",
          8055 => x"9a387983",
          8056 => x"ff0617b8",
          8057 => x"1133811c",
          8058 => x"70892aa8",
          8059 => x"1b080553",
          8060 => x"5d5d59b4",
          8061 => x"1708792e",
          8062 => x"b538800b",
          8063 => x"83183371",
          8064 => x"5c565d74",
          8065 => x"7d2e0981",
          8066 => x"0684b538",
          8067 => x"81547853",
          8068 => x"b8175281",
          8069 => x"173351f8",
          8070 => x"933f84ba",
          8071 => x"8c08802e",
          8072 => x"8538ff59",
          8073 => x"815a78b4",
          8074 => x"180c79fe",
          8075 => x"ca387a83",
          8076 => x"ff0617b8",
          8077 => x"11337088",
          8078 => x"2b7e0778",
          8079 => x"81067184",
          8080 => x"2a535d59",
          8081 => x"595d79fe",
          8082 => x"ae38769f",
          8083 => x"ff0684ba",
          8084 => x"8c0c8f3d",
          8085 => x"0d047588",
          8086 => x"2aa81808",
          8087 => x"0559b417",
          8088 => x"08792eb5",
          8089 => x"38800b83",
          8090 => x"1833715c",
          8091 => x"5d5b7b7b",
          8092 => x"2e098106",
          8093 => x"81c23881",
          8094 => x"547853b8",
          8095 => x"17528117",
          8096 => x"3351f7a8",
          8097 => x"3f84ba8c",
          8098 => x"08802e85",
          8099 => x"38ff5981",
          8100 => x"5a78b418",
          8101 => x"0c79fddf",
          8102 => x"38751083",
          8103 => x"fe067705",
          8104 => x"b8058111",
          8105 => x"33713371",
          8106 => x"882b0784",
          8107 => x"ba8c0c57",
          8108 => x"5b8f3d0d",
          8109 => x"0474832e",
          8110 => x"098106fd",
          8111 => x"b8387587",
          8112 => x"2aa81808",
          8113 => x"0559b417",
          8114 => x"08792eb5",
          8115 => x"38800b83",
          8116 => x"1833715c",
          8117 => x"5e5b7c7b",
          8118 => x"2e098106",
          8119 => x"82813881",
          8120 => x"547853b8",
          8121 => x"17528117",
          8122 => x"3351f6c0",
          8123 => x"3f84ba8c",
          8124 => x"08802e85",
          8125 => x"38ff5981",
          8126 => x"5a78b418",
          8127 => x"0c79fcf7",
          8128 => x"3875822b",
          8129 => x"83fc0677",
          8130 => x"05b80583",
          8131 => x"11338212",
          8132 => x"3371902b",
          8133 => x"71882b07",
          8134 => x"81143370",
          8135 => x"7207882b",
          8136 => x"75337180",
          8137 => x"fffffe80",
          8138 => x"060784ba",
          8139 => x"8c0c415c",
          8140 => x"5e595a56",
          8141 => x"8f3d0d04",
          8142 => x"8154b417",
          8143 => x"0853b817",
          8144 => x"70538118",
          8145 => x"33525cf6",
          8146 => x"e23f815a",
          8147 => x"84ba8c08",
          8148 => x"7b2e0981",
          8149 => x"06febe38",
          8150 => x"84ba8c08",
          8151 => x"831834b4",
          8152 => x"1708a818",
          8153 => x"083184ba",
          8154 => x"8c085b5e",
          8155 => x"7da01808",
          8156 => x"27fe8438",
          8157 => x"82173355",
          8158 => x"74822e09",
          8159 => x"8106fdf7",
          8160 => x"388154b4",
          8161 => x"1708a018",
          8162 => x"0805537b",
          8163 => x"52811733",
          8164 => x"51f6983f",
          8165 => x"7a5afddf",
          8166 => x"398154b4",
          8167 => x"170853b8",
          8168 => x"17705381",
          8169 => x"1833525c",
          8170 => x"f6813f84",
          8171 => x"ba8c087b",
          8172 => x"2e098106",
          8173 => x"82813884",
          8174 => x"ba8c0883",
          8175 => x"1834b417",
          8176 => x"08a81808",
          8177 => x"315d7ca0",
          8178 => x"1808278b",
          8179 => x"38821733",
          8180 => x"5e7d822e",
          8181 => x"81cb3884",
          8182 => x"ba8c085b",
          8183 => x"fbde3981",
          8184 => x"54b41708",
          8185 => x"53b81770",
          8186 => x"53811833",
          8187 => x"525cf5bb",
          8188 => x"3f815a84",
          8189 => x"ba8c087b",
          8190 => x"2e098106",
          8191 => x"fdff3884",
          8192 => x"ba8c0883",
          8193 => x"1834b417",
          8194 => x"08a81808",
          8195 => x"3184ba8c",
          8196 => x"085b5e7d",
          8197 => x"a0180827",
          8198 => x"fdc53882",
          8199 => x"17335574",
          8200 => x"822e0981",
          8201 => x"06fdb838",
          8202 => x"8154b417",
          8203 => x"08a01808",
          8204 => x"05537b52",
          8205 => x"81173351",
          8206 => x"f4f13f7a",
          8207 => x"5afda039",
          8208 => x"8154b417",
          8209 => x"0853b817",
          8210 => x"70538118",
          8211 => x"33525ef4",
          8212 => x"da3f815a",
          8213 => x"84ba8c08",
          8214 => x"7d2e0981",
          8215 => x"06fbcb38",
          8216 => x"84ba8c08",
          8217 => x"831834b4",
          8218 => x"1708a818",
          8219 => x"083184ba",
          8220 => x"8c085b55",
          8221 => x"74a01808",
          8222 => x"27fb9138",
          8223 => x"82173355",
          8224 => x"74822e09",
          8225 => x"8106fb84",
          8226 => x"388154b4",
          8227 => x"1708a018",
          8228 => x"0805537d",
          8229 => x"52811733",
          8230 => x"51f4903f",
          8231 => x"7c5afaec",
          8232 => x"398154b4",
          8233 => x"1708a018",
          8234 => x"0805537b",
          8235 => x"52811733",
          8236 => x"51f3f83f",
          8237 => x"fa863981",
          8238 => x"5b7af9bb",
          8239 => x"38fa9f39",
          8240 => x"f23d0d60",
          8241 => x"62645d57",
          8242 => x"59825881",
          8243 => x"76279c38",
          8244 => x"759c1a08",
          8245 => x"27953878",
          8246 => x"33557478",
          8247 => x"2e963874",
          8248 => x"78248180",
          8249 => x"3874812e",
          8250 => x"828a3877",
          8251 => x"84ba8c0c",
          8252 => x"903d0d04",
          8253 => x"75882aa8",
          8254 => x"1a080558",
          8255 => x"800bb41a",
          8256 => x"08585c76",
          8257 => x"782e86b6",
          8258 => x"38831933",
          8259 => x"7c5b5d7c",
          8260 => x"7c2e0981",
          8261 => x"0683fa38",
          8262 => x"81547753",
          8263 => x"b8195281",
          8264 => x"193351f2",
          8265 => x"873f84ba",
          8266 => x"8c08802e",
          8267 => x"8538ff58",
          8268 => x"815a77b4",
          8269 => x"1a0c7958",
          8270 => x"79ffb038",
          8271 => x"751083fe",
          8272 => x"0679057b",
          8273 => x"83ffff06",
          8274 => x"585e76b8",
          8275 => x"1f347688",
          8276 => x"2a5a79b9",
          8277 => x"1f34810b",
          8278 => x"831a3477",
          8279 => x"84ba8c0c",
          8280 => x"903d0d04",
          8281 => x"74832e09",
          8282 => x"8106feff",
          8283 => x"3875872a",
          8284 => x"a81a0805",
          8285 => x"58800bb4",
          8286 => x"1a08585c",
          8287 => x"76782e85",
          8288 => x"e1388319",
          8289 => x"337c5b5d",
          8290 => x"7c7c2e09",
          8291 => x"810684bd",
          8292 => x"38815477",
          8293 => x"53b81952",
          8294 => x"81193351",
          8295 => x"f18e3f84",
          8296 => x"ba8c0880",
          8297 => x"2e8538ff",
          8298 => x"58815a77",
          8299 => x"b41a0c79",
          8300 => x"5879feb7",
          8301 => x"3875822b",
          8302 => x"83fc0679",
          8303 => x"05b81183",
          8304 => x"11337098",
          8305 => x"2b8f0a06",
          8306 => x"7ef00a06",
          8307 => x"0741575e",
          8308 => x"5c7d7d34",
          8309 => x"7d882a56",
          8310 => x"75b91d34",
          8311 => x"7d902a5a",
          8312 => x"79ba1d34",
          8313 => x"7d982a5b",
          8314 => x"7abb1d34",
          8315 => x"810b831a",
          8316 => x"34fee839",
          8317 => x"75812a16",
          8318 => x"70892aa8",
          8319 => x"1b0805b4",
          8320 => x"1b085959",
          8321 => x"5a76782e",
          8322 => x"b738800b",
          8323 => x"831a3371",
          8324 => x"5e565d74",
          8325 => x"7d2e0981",
          8326 => x"0682d438",
          8327 => x"81547753",
          8328 => x"b8195281",
          8329 => x"193351f0",
          8330 => x"833f84ba",
          8331 => x"8c08802e",
          8332 => x"8538ff58",
          8333 => x"815c77b4",
          8334 => x"1a0c7b58",
          8335 => x"7bfdac38",
          8336 => x"7983ff06",
          8337 => x"19b80581",
          8338 => x"1b778106",
          8339 => x"5f5f577a",
          8340 => x"557c802e",
          8341 => x"8f387a84",
          8342 => x"2b9ff006",
          8343 => x"77338f06",
          8344 => x"7107565a",
          8345 => x"74773481",
          8346 => x"0b831a34",
          8347 => x"7d892aa8",
          8348 => x"1a080556",
          8349 => x"800bb41a",
          8350 => x"08565f74",
          8351 => x"762e83dd",
          8352 => x"38815474",
          8353 => x"53b81970",
          8354 => x"53811a33",
          8355 => x"5257f09b",
          8356 => x"3f815884",
          8357 => x"ba8c087f",
          8358 => x"2e098106",
          8359 => x"80c73884",
          8360 => x"ba8c0883",
          8361 => x"1a34b419",
          8362 => x"0870a81b",
          8363 => x"0831a01b",
          8364 => x"0884ba8c",
          8365 => x"085b5c56",
          8366 => x"5c747a27",
          8367 => x"8b388219",
          8368 => x"33557482",
          8369 => x"2e82e438",
          8370 => x"81547553",
          8371 => x"76528119",
          8372 => x"3351eed8",
          8373 => x"3f84ba8c",
          8374 => x"08802e85",
          8375 => x"38ff5681",
          8376 => x"5875b41a",
          8377 => x"0c77fc83",
          8378 => x"387d83ff",
          8379 => x"0619b805",
          8380 => x"7b842a56",
          8381 => x"567c8f38",
          8382 => x"7a882a76",
          8383 => x"3381f006",
          8384 => x"718f0607",
          8385 => x"565c7476",
          8386 => x"34810b83",
          8387 => x"1a34fccb",
          8388 => x"39815476",
          8389 => x"53b81970",
          8390 => x"53811a33",
          8391 => x"525def8b",
          8392 => x"3f815a84",
          8393 => x"ba8c087c",
          8394 => x"2e098106",
          8395 => x"fc883884",
          8396 => x"ba8c0883",
          8397 => x"1a34b419",
          8398 => x"0870a81b",
          8399 => x"0831a01b",
          8400 => x"0884ba8c",
          8401 => x"085d5940",
          8402 => x"5e7e7727",
          8403 => x"fbca3882",
          8404 => x"19335574",
          8405 => x"822e0981",
          8406 => x"06fbbd38",
          8407 => x"8154761e",
          8408 => x"537c5281",
          8409 => x"193351ee",
          8410 => x"c23f7b5a",
          8411 => x"fbaa3981",
          8412 => x"547653b8",
          8413 => x"19705381",
          8414 => x"1a335257",
          8415 => x"eead3f81",
          8416 => x"5c84ba8c",
          8417 => x"087d2e09",
          8418 => x"8106fdae",
          8419 => x"3884ba8c",
          8420 => x"08831a34",
          8421 => x"b4190870",
          8422 => x"a81b0831",
          8423 => x"a01b0884",
          8424 => x"ba8c085f",
          8425 => x"40565f74",
          8426 => x"7e27fcf0",
          8427 => x"38821933",
          8428 => x"5574822e",
          8429 => x"098106fc",
          8430 => x"e3388154",
          8431 => x"7d1f5376",
          8432 => x"52811933",
          8433 => x"51ede43f",
          8434 => x"7c5cfcd0",
          8435 => x"39815476",
          8436 => x"53b81970",
          8437 => x"53811a33",
          8438 => x"5257edcf",
          8439 => x"3f815a84",
          8440 => x"ba8c087c",
          8441 => x"2e098106",
          8442 => x"fbc53884",
          8443 => x"ba8c0883",
          8444 => x"1a34b419",
          8445 => x"0870a81b",
          8446 => x"0831a01b",
          8447 => x"0884ba8c",
          8448 => x"085d5f40",
          8449 => x"5e7e7d27",
          8450 => x"fb873882",
          8451 => x"19335574",
          8452 => x"822e0981",
          8453 => x"06fafa38",
          8454 => x"81547c1e",
          8455 => x"53765281",
          8456 => x"193351ed",
          8457 => x"863f7b5a",
          8458 => x"fae73981",
          8459 => x"54791c53",
          8460 => x"76528119",
          8461 => x"3351ecf3",
          8462 => x"3f7e58fd",
          8463 => x"8b397b76",
          8464 => x"1083fe06",
          8465 => x"7a057c83",
          8466 => x"ffff0659",
          8467 => x"5f5876b8",
          8468 => x"1f347688",
          8469 => x"2a5a79b9",
          8470 => x"1f34f9fa",
          8471 => x"397e58fd",
          8472 => x"88397b76",
          8473 => x"822b83fc",
          8474 => x"067a05b8",
          8475 => x"11831133",
          8476 => x"70982b8f",
          8477 => x"0a067ff0",
          8478 => x"0a060742",
          8479 => x"585f5d58",
          8480 => x"7d7d347d",
          8481 => x"882a5675",
          8482 => x"b91d347d",
          8483 => x"902a5a79",
          8484 => x"ba1d347d",
          8485 => x"982a5b7a",
          8486 => x"bb1d34fa",
          8487 => x"cf39f63d",
          8488 => x"0d7c7e71",
          8489 => x"085b5c5a",
          8490 => x"7a818a38",
          8491 => x"90190857",
          8492 => x"76802e80",
          8493 => x"f438769c",
          8494 => x"1a082780",
          8495 => x"ec389419",
          8496 => x"08705654",
          8497 => x"73802e80",
          8498 => x"d738767b",
          8499 => x"2e819338",
          8500 => x"76568116",
          8501 => x"569c1908",
          8502 => x"76268938",
          8503 => x"82567577",
          8504 => x"2682b238",
          8505 => x"75527951",
          8506 => x"f0f53f84",
          8507 => x"ba8c0880",
          8508 => x"2e81d038",
          8509 => x"805884ba",
          8510 => x"8c08812e",
          8511 => x"b13884ba",
          8512 => x"8c080970",
          8513 => x"30707207",
          8514 => x"8025707b",
          8515 => x"07515155",
          8516 => x"557382aa",
          8517 => x"3875772e",
          8518 => x"098106ff",
          8519 => x"b5387355",
          8520 => x"7484ba8c",
          8521 => x"0c8c3d0d",
          8522 => x"048157ff",
          8523 => x"913984ba",
          8524 => x"8c0858ca",
          8525 => x"397a5279",
          8526 => x"51f0a43f",
          8527 => x"81557484",
          8528 => x"ba8c0827",
          8529 => x"db3884ba",
          8530 => x"8c085584",
          8531 => x"ba8c08ff",
          8532 => x"2ece389c",
          8533 => x"190884ba",
          8534 => x"8c0826c4",
          8535 => x"387a57fe",
          8536 => x"dd39811b",
          8537 => x"569c1908",
          8538 => x"76268338",
          8539 => x"82567552",
          8540 => x"7951efeb",
          8541 => x"3f805884",
          8542 => x"ba8c0881",
          8543 => x"2e81a038",
          8544 => x"84ba8c08",
          8545 => x"09703070",
          8546 => x"72078025",
          8547 => x"707b0784",
          8548 => x"ba8c0854",
          8549 => x"51515555",
          8550 => x"73ff8538",
          8551 => x"84ba8c08",
          8552 => x"802e9a38",
          8553 => x"90190854",
          8554 => x"817427fe",
          8555 => x"a338739c",
          8556 => x"1a0827fe",
          8557 => x"9b387370",
          8558 => x"5757fe96",
          8559 => x"3975802e",
          8560 => x"fe8e38ff",
          8561 => x"53755278",
          8562 => x"51f5f53f",
          8563 => x"84ba8c08",
          8564 => x"84ba8c08",
          8565 => x"307084ba",
          8566 => x"8c080780",
          8567 => x"25565855",
          8568 => x"7a80c438",
          8569 => x"7480e338",
          8570 => x"75901a0c",
          8571 => x"9c1908fe",
          8572 => x"05941a08",
          8573 => x"56587478",
          8574 => x"268638ff",
          8575 => x"15941a0c",
          8576 => x"84193381",
          8577 => x"075a7984",
          8578 => x"1a347555",
          8579 => x"7484ba8c",
          8580 => x"0c8c3d0d",
          8581 => x"04800b84",
          8582 => x"ba8c0c8c",
          8583 => x"3d0d0484",
          8584 => x"ba8c0858",
          8585 => x"feda3973",
          8586 => x"802effb8",
          8587 => x"3875537a",
          8588 => x"527851f5",
          8589 => x"8b3f84ba",
          8590 => x"8c0855ff",
          8591 => x"a73984ba",
          8592 => x"8c0884ba",
          8593 => x"8c0c8c3d",
          8594 => x"0d04ff56",
          8595 => x"74812eff",
          8596 => x"b9388155",
          8597 => x"ffb639f8",
          8598 => x"3d0d7a7c",
          8599 => x"71085955",
          8600 => x"5873f080",
          8601 => x"0a2680df",
          8602 => x"38739f06",
          8603 => x"537280d7",
          8604 => x"38739019",
          8605 => x"0c881808",
          8606 => x"557480df",
          8607 => x"38763356",
          8608 => x"75822680",
          8609 => x"cc387385",
          8610 => x"2a53820b",
          8611 => x"8818225a",
          8612 => x"56727927",
          8613 => x"a938ac17",
          8614 => x"0898190c",
          8615 => x"7494190c",
          8616 => x"98180853",
          8617 => x"82567280",
          8618 => x"2e943873",
          8619 => x"892a1398",
          8620 => x"190c7383",
          8621 => x"ff0617b8",
          8622 => x"059c190c",
          8623 => x"80567584",
          8624 => x"ba8c0c8a",
          8625 => x"3d0d0482",
          8626 => x"0b84ba8c",
          8627 => x"0c8a3d0d",
          8628 => x"04ac1708",
          8629 => x"5574802e",
          8630 => x"ffac388a",
          8631 => x"17227089",
          8632 => x"2b575973",
          8633 => x"7627a538",
          8634 => x"9c170853",
          8635 => x"fe15fe14",
          8636 => x"54568059",
          8637 => x"7573278d",
          8638 => x"388a1722",
          8639 => x"767129b0",
          8640 => x"1908055a",
          8641 => x"53789819",
          8642 => x"0cff9139",
          8643 => x"74527751",
          8644 => x"eccd3f84",
          8645 => x"ba8c0855",
          8646 => x"84ba8c08",
          8647 => x"ff2ea438",
          8648 => x"810b84ba",
          8649 => x"8c0827ff",
          8650 => x"9e389c17",
          8651 => x"085384ba",
          8652 => x"8c087327",
          8653 => x"ff913873",
          8654 => x"76315473",
          8655 => x"7627cd38",
          8656 => x"ffaa3981",
          8657 => x"0b84ba8c",
          8658 => x"0c8a3d0d",
          8659 => x"04f33d0d",
          8660 => x"7f700890",
          8661 => x"1208a005",
          8662 => x"5c5a57f0",
          8663 => x"800a7a27",
          8664 => x"8638800b",
          8665 => x"98180c98",
          8666 => x"17085584",
          8667 => x"5674802e",
          8668 => x"b2387983",
          8669 => x"ff065b7a",
          8670 => x"9d388115",
          8671 => x"94180857",
          8672 => x"5875a938",
          8673 => x"79852a88",
          8674 => x"1a225755",
          8675 => x"74762781",
          8676 => x"f5387798",
          8677 => x"180c7990",
          8678 => x"180c781b",
          8679 => x"b8059c18",
          8680 => x"0c805675",
          8681 => x"84ba8c0c",
          8682 => x"8f3d0d04",
          8683 => x"7798180c",
          8684 => x"8a1922ff",
          8685 => x"057a892a",
          8686 => x"065c7bda",
          8687 => x"38755276",
          8688 => x"51eb9c3f",
          8689 => x"84ba8c08",
          8690 => x"5d825681",
          8691 => x"0b84ba8c",
          8692 => x"0827d038",
          8693 => x"815684ba",
          8694 => x"8c08ff2e",
          8695 => x"c6389c19",
          8696 => x"0884ba8c",
          8697 => x"08268291",
          8698 => x"3860802e",
          8699 => x"81983894",
          8700 => x"17085276",
          8701 => x"51f9a73f",
          8702 => x"84ba8c08",
          8703 => x"5d875684",
          8704 => x"ba8c0880",
          8705 => x"2eff9c38",
          8706 => x"825684ba",
          8707 => x"8c08812e",
          8708 => x"ff913881",
          8709 => x"5684ba8c",
          8710 => x"08ff2eff",
          8711 => x"863884ba",
          8712 => x"8c08831a",
          8713 => x"335f587d",
          8714 => x"80ea38fe",
          8715 => x"189c1a08",
          8716 => x"fe055956",
          8717 => x"805c7578",
          8718 => x"278d388a",
          8719 => x"19227671",
          8720 => x"29b01b08",
          8721 => x"055d5e7b",
          8722 => x"b41a0cb8",
          8723 => x"19588480",
          8724 => x"78575580",
          8725 => x"76708105",
          8726 => x"5834ff15",
          8727 => x"5574f438",
          8728 => x"74568a19",
          8729 => x"22557575",
          8730 => x"27818038",
          8731 => x"8154751c",
          8732 => x"53775281",
          8733 => x"193351e4",
          8734 => x"b23f84ba",
          8735 => x"8c0880e7",
          8736 => x"38811656",
          8737 => x"dd397a98",
          8738 => x"180c840b",
          8739 => x"84ba8c0c",
          8740 => x"8f3d0d04",
          8741 => x"7554b419",
          8742 => x"0853b819",
          8743 => x"7053811a",
          8744 => x"335256e4",
          8745 => x"863f84ba",
          8746 => x"8c0880f3",
          8747 => x"3884ba8c",
          8748 => x"08831a34",
          8749 => x"b41908a8",
          8750 => x"1a083155",
          8751 => x"74a01a08",
          8752 => x"27fee838",
          8753 => x"8219335c",
          8754 => x"7b822e09",
          8755 => x"8106fedb",
          8756 => x"388154b4",
          8757 => x"1908a01a",
          8758 => x"08055375",
          8759 => x"52811933",
          8760 => x"51e3c83f",
          8761 => x"fec5398a",
          8762 => x"19225574",
          8763 => x"83ffff06",
          8764 => x"5574762e",
          8765 => x"098106a7",
          8766 => x"387c9418",
          8767 => x"0cfe1d9c",
          8768 => x"1a08fe05",
          8769 => x"5e568058",
          8770 => x"757d27fd",
          8771 => x"85388a19",
          8772 => x"22767129",
          8773 => x"b01b0805",
          8774 => x"98190c5c",
          8775 => x"fcf83981",
          8776 => x"0b84ba8c",
          8777 => x"0c8f3d0d",
          8778 => x"04ee3d0d",
          8779 => x"6466415c",
          8780 => x"847c085a",
          8781 => x"5b81ff70",
          8782 => x"981e0858",
          8783 => x"5e5e7580",
          8784 => x"2e82d238",
          8785 => x"b8195f75",
          8786 => x"5a8058b4",
          8787 => x"1908762e",
          8788 => x"82d13883",
          8789 => x"19337858",
          8790 => x"5574782e",
          8791 => x"09810681",
          8792 => x"94388154",
          8793 => x"7553b819",
          8794 => x"52811933",
          8795 => x"51e1bd3f",
          8796 => x"84ba8c08",
          8797 => x"802e8538",
          8798 => x"ff5a8157",
          8799 => x"79b41a0c",
          8800 => x"765b7682",
          8801 => x"90389c1c",
          8802 => x"08703358",
          8803 => x"5876802e",
          8804 => x"8281388b",
          8805 => x"1833bf06",
          8806 => x"7081ff06",
          8807 => x"5b416086",
          8808 => x"1d347681",
          8809 => x"e5327030",
          8810 => x"78ae3270",
          8811 => x"30728025",
          8812 => x"71802507",
          8813 => x"54454557",
          8814 => x"55749338",
          8815 => x"747adf06",
          8816 => x"43566188",
          8817 => x"2e81bf38",
          8818 => x"75602e81",
          8819 => x"863881ff",
          8820 => x"5d80527b",
          8821 => x"51faf63f",
          8822 => x"84ba8c08",
          8823 => x"5b84ba8c",
          8824 => x"0881b238",
          8825 => x"981c0856",
          8826 => x"75fedc38",
          8827 => x"7a84ba8c",
          8828 => x"0c943d0d",
          8829 => x"048154b4",
          8830 => x"1908537e",
          8831 => x"52811933",
          8832 => x"51e1a83f",
          8833 => x"815784ba",
          8834 => x"8c08782e",
          8835 => x"098106fe",
          8836 => x"ef3884ba",
          8837 => x"8c08831a",
          8838 => x"34b41908",
          8839 => x"a81a0831",
          8840 => x"84ba8c08",
          8841 => x"585b7aa0",
          8842 => x"1a0827fe",
          8843 => x"b5388219",
          8844 => x"33416082",
          8845 => x"2e098106",
          8846 => x"fea83881",
          8847 => x"54b41908",
          8848 => x"a01a0805",
          8849 => x"537e5281",
          8850 => x"193351e0",
          8851 => x"de3f7757",
          8852 => x"fe903979",
          8853 => x"8f2e0981",
          8854 => x"0681e738",
          8855 => x"76862a81",
          8856 => x"065b7a80",
          8857 => x"2e93388d",
          8858 => x"18337781",
          8859 => x"bf067090",
          8860 => x"1f087fac",
          8861 => x"050c595e",
          8862 => x"5e767d2e",
          8863 => x"ab3881ff",
          8864 => x"55745dfe",
          8865 => x"cc398156",
          8866 => x"75602e09",
          8867 => x"8106febe",
          8868 => x"38c13984",
          8869 => x"5b800b98",
          8870 => x"1d0c7a84",
          8871 => x"ba8c0c94",
          8872 => x"3d0d0477",
          8873 => x"5bfddf39",
          8874 => x"8d183357",
          8875 => x"7d772e09",
          8876 => x"8106cb38",
          8877 => x"8c19089b",
          8878 => x"19339a1a",
          8879 => x"3371882b",
          8880 => x"07585641",
          8881 => x"75ffb738",
          8882 => x"77337081",
          8883 => x"bf068d29",
          8884 => x"f305515a",
          8885 => x"8176585b",
          8886 => x"83e68c17",
          8887 => x"33780581",
          8888 => x"11337133",
          8889 => x"71882b07",
          8890 => x"5244567a",
          8891 => x"802e80c5",
          8892 => x"387981fe",
          8893 => x"26ff8738",
          8894 => x"79106105",
          8895 => x"765c4275",
          8896 => x"6223811a",
          8897 => x"5a811757",
          8898 => x"8c7727cc",
          8899 => x"38773370",
          8900 => x"862a8106",
          8901 => x"59577780",
          8902 => x"2e903879",
          8903 => x"81fe26fe",
          8904 => x"dd387910",
          8905 => x"61054380",
          8906 => x"6323ff1d",
          8907 => x"7081ff06",
          8908 => x"5e41fd9d",
          8909 => x"397583ff",
          8910 => x"ff2eca38",
          8911 => x"81ff55fe",
          8912 => x"c0397ca8",
          8913 => x"387c558b",
          8914 => x"5774812a",
          8915 => x"75818029",
          8916 => x"05787081",
          8917 => x"055a3340",
          8918 => x"7f057081",
          8919 => x"ff06ff19",
          8920 => x"59565976",
          8921 => x"e438747e",
          8922 => x"2efd8138",
          8923 => x"ff0bac1d",
          8924 => x"0c7a84ba",
          8925 => x"8c0c943d",
          8926 => x"0d04ef3d",
          8927 => x"0d637008",
          8928 => x"5c5c8052",
          8929 => x"7b51f5cf",
          8930 => x"3f84ba8c",
          8931 => x"085a84ba",
          8932 => x"8c088280",
          8933 => x"3881ff70",
          8934 => x"405dff0b",
          8935 => x"ac1d0cb8",
          8936 => x"1b5e981c",
          8937 => x"08568058",
          8938 => x"b41b0876",
          8939 => x"2e82cc38",
          8940 => x"831b3378",
          8941 => x"58557478",
          8942 => x"2e098106",
          8943 => x"81df3881",
          8944 => x"547553b8",
          8945 => x"1b52811b",
          8946 => x"3351dce0",
          8947 => x"3f84ba8c",
          8948 => x"08802e85",
          8949 => x"38ff5681",
          8950 => x"5775b41c",
          8951 => x"0c765a76",
          8952 => x"81b2389c",
          8953 => x"1c087033",
          8954 => x"58597680",
          8955 => x"2e849938",
          8956 => x"8b1933bf",
          8957 => x"067081ff",
          8958 => x"06575877",
          8959 => x"861d3476",
          8960 => x"81e52e80",
          8961 => x"f2387583",
          8962 => x"2a810655",
          8963 => x"758f2e81",
          8964 => x"ef387480",
          8965 => x"e238758f",
          8966 => x"2e81e538",
          8967 => x"7caa3878",
          8968 => x"7d56588b",
          8969 => x"5774812a",
          8970 => x"75818029",
          8971 => x"05787081",
          8972 => x"055a3357",
          8973 => x"76057081",
          8974 => x"ff06ff19",
          8975 => x"59565d76",
          8976 => x"e438747f",
          8977 => x"2e80cd38",
          8978 => x"ab1c3381",
          8979 => x"065776a7",
          8980 => x"388b0ba0",
          8981 => x"1d595778",
          8982 => x"7081055a",
          8983 => x"33787081",
          8984 => x"055a3371",
          8985 => x"7131ff1a",
          8986 => x"5a584240",
          8987 => x"76802e81",
          8988 => x"dc387580",
          8989 => x"2ee13881",
          8990 => x"ff5dff0b",
          8991 => x"ac1d0c80",
          8992 => x"527b51f5",
          8993 => x"c83f84ba",
          8994 => x"8c085a84",
          8995 => x"ba8c0880",
          8996 => x"2efe8f38",
          8997 => x"7984ba8c",
          8998 => x"0c933d0d",
          8999 => x"048154b4",
          9000 => x"1b08537d",
          9001 => x"52811b33",
          9002 => x"51dc803f",
          9003 => x"815784ba",
          9004 => x"8c08782e",
          9005 => x"098106fe",
          9006 => x"a43884ba",
          9007 => x"8c08831c",
          9008 => x"34b41b08",
          9009 => x"a81c0831",
          9010 => x"84ba8c08",
          9011 => x"585978a0",
          9012 => x"1c0827fd",
          9013 => x"ea38821b",
          9014 => x"335a7982",
          9015 => x"2e098106",
          9016 => x"fddd3881",
          9017 => x"54b41b08",
          9018 => x"a01c0805",
          9019 => x"537d5281",
          9020 => x"1b3351db",
          9021 => x"b63f7757",
          9022 => x"fdc53977",
          9023 => x"5afde439",
          9024 => x"ab1c3370",
          9025 => x"862a8106",
          9026 => x"425560fe",
          9027 => x"f2387686",
          9028 => x"2a81065a",
          9029 => x"79802e93",
          9030 => x"388d1933",
          9031 => x"7781bf06",
          9032 => x"70901f08",
          9033 => x"7fac050c",
          9034 => x"595e5f76",
          9035 => x"7d2eaf38",
          9036 => x"81ff5574",
          9037 => x"5d80527b",
          9038 => x"51f4923f",
          9039 => x"84ba8c08",
          9040 => x"5a84ba8c",
          9041 => x"08802efc",
          9042 => x"d938fec8",
          9043 => x"3975802e",
          9044 => x"fec23881",
          9045 => x"ff5dff0b",
          9046 => x"ac1d0cfe",
          9047 => x"a2398d19",
          9048 => x"33577e77",
          9049 => x"2e098106",
          9050 => x"c7388c1b",
          9051 => x"089b1a33",
          9052 => x"9a1b3371",
          9053 => x"882b0759",
          9054 => x"424076ff",
          9055 => x"b3387833",
          9056 => x"70bf068d",
          9057 => x"29f3055b",
          9058 => x"55817759",
          9059 => x"5683e68c",
          9060 => x"18337905",
          9061 => x"81113371",
          9062 => x"3371882b",
          9063 => x"07524257",
          9064 => x"75802e80",
          9065 => x"ed387981",
          9066 => x"fe26ff84",
          9067 => x"38765181",
          9068 => x"a18a3f84",
          9069 => x"ba8c087a",
          9070 => x"10610570",
          9071 => x"22534381",
          9072 => x"1b5b5681",
          9073 => x"a0f63f75",
          9074 => x"84ba8c08",
          9075 => x"2e098106",
          9076 => x"fede3876",
          9077 => x"56811858",
          9078 => x"8c7827ff",
          9079 => x"b0387833",
          9080 => x"70862a81",
          9081 => x"06565975",
          9082 => x"802e9238",
          9083 => x"74802e8d",
          9084 => x"38791060",
          9085 => x"05702241",
          9086 => x"417ffeb4",
          9087 => x"38ff1d70",
          9088 => x"81ff065e",
          9089 => x"5afeae39",
          9090 => x"840b84ba",
          9091 => x"8c0c933d",
          9092 => x"0d047683",
          9093 => x"ffff2eff",
          9094 => x"bc3881ff",
          9095 => x"55fe9439",
          9096 => x"ea3d0d68",
          9097 => x"700870ab",
          9098 => x"133381a0",
          9099 => x"06585a5d",
          9100 => x"5e865674",
          9101 => x"85b53874",
          9102 => x"8c1d0870",
          9103 => x"2257575d",
          9104 => x"74802e8e",
          9105 => x"38811d70",
          9106 => x"10177022",
          9107 => x"51565d74",
          9108 => x"f438953d",
          9109 => x"a01f5b40",
          9110 => x"8c607b58",
          9111 => x"58557570",
          9112 => x"81055733",
          9113 => x"77708105",
          9114 => x"5934ff15",
          9115 => x"5574ef38",
          9116 => x"0280db05",
          9117 => x"33708106",
          9118 => x"58567680",
          9119 => x"2e82aa38",
          9120 => x"80c00bab",
          9121 => x"1f34810b",
          9122 => x"943d405b",
          9123 => x"8c1c087b",
          9124 => x"58598b7a",
          9125 => x"615a5755",
          9126 => x"77708105",
          9127 => x"59337670",
          9128 => x"81055834",
          9129 => x"ff155574",
          9130 => x"ef38857b",
          9131 => x"2780c238",
          9132 => x"7a792256",
          9133 => x"5774802e",
          9134 => x"b8387482",
          9135 => x"1a5a568f",
          9136 => x"58758106",
          9137 => x"77100776",
          9138 => x"812a7083",
          9139 => x"ffff0672",
          9140 => x"902a8106",
          9141 => x"44585657",
          9142 => x"60802e87",
          9143 => x"387684a0",
          9144 => x"a13257ff",
          9145 => x"18587780",
          9146 => x"25d73878",
          9147 => x"225574ca",
          9148 => x"38870284",
          9149 => x"0580cf05",
          9150 => x"575876b0",
          9151 => x"07bf0655",
          9152 => x"b9752784",
          9153 => x"38871555",
          9154 => x"747634ff",
          9155 => x"16ff1978",
          9156 => x"842a5959",
          9157 => x"5676e338",
          9158 => x"771f5980",
          9159 => x"fe793476",
          9160 => x"7a585680",
          9161 => x"7827a038",
          9162 => x"79335574",
          9163 => x"a02e9838",
          9164 => x"81165675",
          9165 => x"782788a2",
          9166 => x"38751a70",
          9167 => x"33565774",
          9168 => x"a02e0981",
          9169 => x"06ea3881",
          9170 => x"1656a055",
          9171 => x"7787268e",
          9172 => x"38983d78",
          9173 => x"05ec0581",
          9174 => x"19713357",
          9175 => x"59417477",
          9176 => x"34877627",
          9177 => x"87f4387d",
          9178 => x"51f88f3f",
          9179 => x"84ba8c08",
          9180 => x"8b38811b",
          9181 => x"5b80e37b",
          9182 => x"27fe9138",
          9183 => x"87567a80",
          9184 => x"e42e82e7",
          9185 => x"3884ba8c",
          9186 => x"085684ba",
          9187 => x"8c08842e",
          9188 => x"09810682",
          9189 => x"d6380280",
          9190 => x"db0533ab",
          9191 => x"1f347d08",
          9192 => x"02840580",
          9193 => x"db053357",
          9194 => x"5875812a",
          9195 => x"81065f81",
          9196 => x"5b7e802e",
          9197 => x"90388d52",
          9198 => x"8c1d51fe",
          9199 => x"89e73f84",
          9200 => x"ba8c081b",
          9201 => x"5b80527d",
          9202 => x"51ed8c3f",
          9203 => x"84ba8c08",
          9204 => x"5684ba8c",
          9205 => x"08818238",
          9206 => x"84ba8c08",
          9207 => x"b8195e59",
          9208 => x"981e0856",
          9209 => x"8057b418",
          9210 => x"08762e85",
          9211 => x"f3388318",
          9212 => x"33407f77",
          9213 => x"2e098106",
          9214 => x"82a33881",
          9215 => x"547553b8",
          9216 => x"18528118",
          9217 => x"3351d4a4",
          9218 => x"3f84ba8c",
          9219 => x"08802e85",
          9220 => x"38ff5681",
          9221 => x"5775b419",
          9222 => x"0c765676",
          9223 => x"bc389c1e",
          9224 => x"08703356",
          9225 => x"427481e5",
          9226 => x"2e81c938",
          9227 => x"74307080",
          9228 => x"25780756",
          9229 => x"5f74802e",
          9230 => x"81c93881",
          9231 => x"1959787b",
          9232 => x"2e868938",
          9233 => x"81527d51",
          9234 => x"ee833f84",
          9235 => x"ba8c0856",
          9236 => x"84ba8c08",
          9237 => x"802eff88",
          9238 => x"38875875",
          9239 => x"842e8189",
          9240 => x"38755875",
          9241 => x"818338ff",
          9242 => x"1b407f81",
          9243 => x"f338981e",
          9244 => x"0857b41c",
          9245 => x"08772eaf",
          9246 => x"38831c33",
          9247 => x"7857407f",
          9248 => x"84823881",
          9249 => x"547653b8",
          9250 => x"1c52811c",
          9251 => x"3351d39c",
          9252 => x"3f84ba8c",
          9253 => x"08802e85",
          9254 => x"38ff5781",
          9255 => x"5676b41d",
          9256 => x"0c755875",
          9257 => x"80c338a0",
          9258 => x"0b9c1f08",
          9259 => x"57558076",
          9260 => x"70810558",
          9261 => x"34ff1555",
          9262 => x"74f4388b",
          9263 => x"0b9c1f08",
          9264 => x"7b585855",
          9265 => x"75708105",
          9266 => x"57337770",
          9267 => x"81055934",
          9268 => x"ff155574",
          9269 => x"ef389c1e",
          9270 => x"08ab1f33",
          9271 => x"98065e5a",
          9272 => x"7c8c1b34",
          9273 => x"810b831d",
          9274 => x"34775675",
          9275 => x"84ba8c0c",
          9276 => x"983d0d04",
          9277 => x"81753070",
          9278 => x"80257207",
          9279 => x"57405774",
          9280 => x"feb93874",
          9281 => x"5981527d",
          9282 => x"51ecc23f",
          9283 => x"84ba8c08",
          9284 => x"5684ba8c",
          9285 => x"08802efd",
          9286 => x"c738febd",
          9287 => x"398154b4",
          9288 => x"1808537c",
          9289 => x"52811833",
          9290 => x"51d3803f",
          9291 => x"84ba8c08",
          9292 => x"772e0981",
          9293 => x"0683bf38",
          9294 => x"84ba8c08",
          9295 => x"831934b4",
          9296 => x"1808a819",
          9297 => x"08315574",
          9298 => x"a0190827",
          9299 => x"8b388218",
          9300 => x"33416082",
          9301 => x"2e84ac38",
          9302 => x"84ba8c08",
          9303 => x"57fd9c39",
          9304 => x"7f852b90",
          9305 => x"1f087131",
          9306 => x"53587d51",
          9307 => x"e9e93f84",
          9308 => x"ba8c0858",
          9309 => x"84ba8c08",
          9310 => x"feef3879",
          9311 => x"84ba8c08",
          9312 => x"56588b57",
          9313 => x"74812a75",
          9314 => x"81802905",
          9315 => x"78708105",
          9316 => x"5a335776",
          9317 => x"057081ff",
          9318 => x"06ff1959",
          9319 => x"565d76e4",
          9320 => x"387481ff",
          9321 => x"06b81d43",
          9322 => x"41981e08",
          9323 => x"578056b4",
          9324 => x"1c08772e",
          9325 => x"b238831c",
          9326 => x"335b7a76",
          9327 => x"2e098106",
          9328 => x"82c93881",
          9329 => x"547653b8",
          9330 => x"1c52811c",
          9331 => x"3351d0dc",
          9332 => x"3f84ba8c",
          9333 => x"08802e85",
          9334 => x"38ff5781",
          9335 => x"5676b41d",
          9336 => x"0c755875",
          9337 => x"fe83388c",
          9338 => x"1c089c1f",
          9339 => x"086181ff",
          9340 => x"065f5c5f",
          9341 => x"608d1c34",
          9342 => x"8f0b8b1c",
          9343 => x"34758c1c",
          9344 => x"34759a1c",
          9345 => x"34759b1c",
          9346 => x"347c8d29",
          9347 => x"f3057677",
          9348 => x"5a585976",
          9349 => x"83ffff2e",
          9350 => x"8b387810",
          9351 => x"1f702281",
          9352 => x"1b5b5856",
          9353 => x"83e68c18",
          9354 => x"337b0555",
          9355 => x"76757081",
          9356 => x"05573476",
          9357 => x"882a5675",
          9358 => x"75347685",
          9359 => x"3883ffff",
          9360 => x"57811858",
          9361 => x"8c7827cb",
          9362 => x"387683ff",
          9363 => x"ff2e81b3",
          9364 => x"3878101f",
          9365 => x"70225858",
          9366 => x"76802e81",
          9367 => x"a6387c7b",
          9368 => x"34810b83",
          9369 => x"1d348052",
          9370 => x"7d51e9e1",
          9371 => x"3f84ba8c",
          9372 => x"085884ba",
          9373 => x"8c08fcf1",
          9374 => x"387fff05",
          9375 => x"407ffea9",
          9376 => x"38fbeb39",
          9377 => x"8154b41c",
          9378 => x"0853b81c",
          9379 => x"7053811d",
          9380 => x"335259d0",
          9381 => x"963f8156",
          9382 => x"84ba8c08",
          9383 => x"fc833884",
          9384 => x"ba8c0883",
          9385 => x"1d34b41c",
          9386 => x"08a81d08",
          9387 => x"3184ba8c",
          9388 => x"08574160",
          9389 => x"a01d0827",
          9390 => x"fbc93882",
          9391 => x"1c334261",
          9392 => x"822e0981",
          9393 => x"06fbbc38",
          9394 => x"8154b41c",
          9395 => x"08a01d08",
          9396 => x"05537852",
          9397 => x"811c3351",
          9398 => x"cfd13f77",
          9399 => x"56fba439",
          9400 => x"769c1f08",
          9401 => x"70335743",
          9402 => x"567481e5",
          9403 => x"2e098106",
          9404 => x"faba38fb",
          9405 => x"ff398170",
          9406 => x"57577680",
          9407 => x"2efa9f38",
          9408 => x"fad7397c",
          9409 => x"80c0075d",
          9410 => x"fed43981",
          9411 => x"54b41c08",
          9412 => x"53615281",
          9413 => x"1c3351cf",
          9414 => x"923f84ba",
          9415 => x"8c08762e",
          9416 => x"098106bc",
          9417 => x"3884ba8c",
          9418 => x"08831d34",
          9419 => x"b41c08a8",
          9420 => x"1d083155",
          9421 => x"74a01d08",
          9422 => x"278a3882",
          9423 => x"1c335f7e",
          9424 => x"822eaa38",
          9425 => x"84ba8c08",
          9426 => x"56fcf839",
          9427 => x"75ff1c41",
          9428 => x"587f802e",
          9429 => x"fa9838fc",
          9430 => x"8739751a",
          9431 => x"57f7e839",
          9432 => x"81705956",
          9433 => x"75802efc",
          9434 => x"fe38fafd",
          9435 => x"398154b4",
          9436 => x"1c08a01d",
          9437 => x"08055361",
          9438 => x"52811c33",
          9439 => x"51ceac3f",
          9440 => x"fcc13981",
          9441 => x"54b41808",
          9442 => x"a0190805",
          9443 => x"537c5281",
          9444 => x"183351ce",
          9445 => x"963ff8e3",
          9446 => x"39f33d0d",
          9447 => x"7f617108",
          9448 => x"405e5c80",
          9449 => x"0b961e34",
          9450 => x"981c0880",
          9451 => x"2e82b538",
          9452 => x"ac1c08ff",
          9453 => x"2e80d938",
          9454 => x"80707160",
          9455 => x"8c050870",
          9456 => x"2257585b",
          9457 => x"5c587278",
          9458 => x"2ebc3877",
          9459 => x"54741470",
          9460 => x"22811b5b",
          9461 => x"55567a82",
          9462 => x"953880d0",
          9463 => x"80147083",
          9464 => x"ffff0658",
          9465 => x"5a768fff",
          9466 => x"26828338",
          9467 => x"73791a76",
          9468 => x"1170225d",
          9469 => x"58555b79",
          9470 => x"d4387a30",
          9471 => x"70802570",
          9472 => x"307a065a",
          9473 => x"5c5e7c18",
          9474 => x"94055780",
          9475 => x"0b821834",
          9476 => x"8070891f",
          9477 => x"5957589c",
          9478 => x"1c081670",
          9479 => x"33811858",
          9480 => x"565374a0",
          9481 => x"2eb23874",
          9482 => x"852e81bc",
          9483 => x"38758932",
          9484 => x"70307072",
          9485 => x"07802555",
          9486 => x"5b54778b",
          9487 => x"26903872",
          9488 => x"802e8b38",
          9489 => x"ae777081",
          9490 => x"05593481",
          9491 => x"18587477",
          9492 => x"70810559",
          9493 => x"34811858",
          9494 => x"8a7627ff",
          9495 => x"ba387c18",
          9496 => x"88055580",
          9497 => x"0b811634",
          9498 => x"961d3353",
          9499 => x"72a53877",
          9500 => x"81f338bf",
          9501 => x"0b961e34",
          9502 => x"81577c17",
          9503 => x"94055680",
          9504 => x"0b821734",
          9505 => x"9c1c088c",
          9506 => x"11335553",
          9507 => x"73893873",
          9508 => x"891e349c",
          9509 => x"1c08538b",
          9510 => x"1333881e",
          9511 => x"349c1c08",
          9512 => x"9c118311",
          9513 => x"33821233",
          9514 => x"71902b71",
          9515 => x"882b0781",
          9516 => x"14337072",
          9517 => x"07882b75",
          9518 => x"33710764",
          9519 => x"0c599716",
          9520 => x"33961733",
          9521 => x"71882b07",
          9522 => x"5f415b40",
          9523 => x"5a565b55",
          9524 => x"77861e23",
          9525 => x"99153398",
          9526 => x"16337188",
          9527 => x"2b075d54",
          9528 => x"7b841e23",
          9529 => x"8f3d0d04",
          9530 => x"81e555fe",
          9531 => x"c039771d",
          9532 => x"961181ff",
          9533 => x"7a31585b",
          9534 => x"5783b552",
          9535 => x"7a902b74",
          9536 => x"07518191",
          9537 => x"893f84ba",
          9538 => x"8c0883ff",
          9539 => x"ff065581",
          9540 => x"ff7527ad",
          9541 => x"38817627",
          9542 => x"81b33874",
          9543 => x"882a5473",
          9544 => x"7a347497",
          9545 => x"18348278",
          9546 => x"0558800b",
          9547 => x"8c1f0856",
          9548 => x"5b781975",
          9549 => x"1170225c",
          9550 => x"575479fd",
          9551 => x"9038fdba",
          9552 => x"39743076",
          9553 => x"30707807",
          9554 => x"80257280",
          9555 => x"25075855",
          9556 => x"577580f9",
          9557 => x"38747a34",
          9558 => x"81780558",
          9559 => x"800b8c1f",
          9560 => x"08565bcd",
          9561 => x"39727389",
          9562 => x"1f335a57",
          9563 => x"5777802e",
          9564 => x"fe88387c",
          9565 => x"961e7e57",
          9566 => x"59548914",
          9567 => x"33ffbf11",
          9568 => x"5a547899",
          9569 => x"26a4389c",
          9570 => x"1c088c11",
          9571 => x"33545b88",
          9572 => x"7627b438",
          9573 => x"72842a53",
          9574 => x"7281065e",
          9575 => x"7d802e8a",
          9576 => x"38a01470",
          9577 => x"83ffff06",
          9578 => x"55537378",
          9579 => x"7081055a",
          9580 => x"34811681",
          9581 => x"16811971",
          9582 => x"8913335e",
          9583 => x"57595656",
          9584 => x"79ffb738",
          9585 => x"fdb43972",
          9586 => x"832a53cc",
          9587 => x"39807b30",
          9588 => x"70802570",
          9589 => x"30730653",
          9590 => x"5d5f58fc",
          9591 => x"a939ef3d",
          9592 => x"0d637008",
          9593 => x"7042575c",
          9594 => x"80657033",
          9595 => x"57555374",
          9596 => x"af2e8338",
          9597 => x"81537480",
          9598 => x"dc2e81df",
          9599 => x"3872802e",
          9600 => x"81d93898",
          9601 => x"1608881d",
          9602 => x"0c733396",
          9603 => x"3d943d41",
          9604 => x"42559f75",
          9605 => x"2782a738",
          9606 => x"73428c16",
          9607 => x"08588057",
          9608 => x"61707081",
          9609 => x"05523355",
          9610 => x"537381df",
          9611 => x"38727f0c",
          9612 => x"73ff2e81",
          9613 => x"ec3883ff",
          9614 => x"ff74278b",
          9615 => x"38761018",
          9616 => x"56807623",
          9617 => x"81175773",
          9618 => x"83ffff06",
          9619 => x"70af3270",
          9620 => x"309f7327",
          9621 => x"71802507",
          9622 => x"575b5b55",
          9623 => x"73829038",
          9624 => x"7480dc2e",
          9625 => x"82893874",
          9626 => x"80ff26b2",
          9627 => x"3883e5a8",
          9628 => x"0b83e5a8",
          9629 => x"337081ff",
          9630 => x"06565456",
          9631 => x"73802e81",
          9632 => x"ab387375",
          9633 => x"2e8f3881",
          9634 => x"16703370",
          9635 => x"81ff0656",
          9636 => x"545673ee",
          9637 => x"387281ff",
          9638 => x"065b7a81",
          9639 => x"84387681",
          9640 => x"fe2680fd",
          9641 => x"38761018",
          9642 => x"5d747d23",
          9643 => x"81176270",
          9644 => x"70810552",
          9645 => x"33565457",
          9646 => x"73802efe",
          9647 => x"f03880cb",
          9648 => x"39817380",
          9649 => x"dc327030",
          9650 => x"70802573",
          9651 => x"07515558",
          9652 => x"5572802e",
          9653 => x"a1388114",
          9654 => x"70465480",
          9655 => x"74335455",
          9656 => x"72af2edd",
          9657 => x"387280dc",
          9658 => x"32703070",
          9659 => x"80257707",
          9660 => x"51545772",
          9661 => x"e1387288",
          9662 => x"1d0c7333",
          9663 => x"963d943d",
          9664 => x"41425574",
          9665 => x"9f26fe90",
          9666 => x"38b43983",
          9667 => x"b5527351",
          9668 => x"818de73f",
          9669 => x"84ba8c08",
          9670 => x"83ffff06",
          9671 => x"5473fe8d",
          9672 => x"38865473",
          9673 => x"84ba8c0c",
          9674 => x"933d0d04",
          9675 => x"83e5a833",
          9676 => x"7081ff06",
          9677 => x"5c537a80",
          9678 => x"2efee338",
          9679 => x"e439ff80",
          9680 => x"0bab1d34",
          9681 => x"80527b51",
          9682 => x"de8d3f84",
          9683 => x"ba8c0884",
          9684 => x"ba8c0c93",
          9685 => x"3d0d0481",
          9686 => x"7380dc32",
          9687 => x"70307080",
          9688 => x"25730741",
          9689 => x"555a567d",
          9690 => x"802ea138",
          9691 => x"81144280",
          9692 => x"62703355",
          9693 => x"555672af",
          9694 => x"2edd3872",
          9695 => x"80dc3270",
          9696 => x"30708025",
          9697 => x"78074054",
          9698 => x"597de138",
          9699 => x"73610c9f",
          9700 => x"7527822b",
          9701 => x"5a76812e",
          9702 => x"84f83876",
          9703 => x"822e83d1",
          9704 => x"38761759",
          9705 => x"76802ea7",
          9706 => x"38761778",
          9707 => x"11fe0570",
          9708 => x"2270a032",
          9709 => x"7030709f",
          9710 => x"2a524256",
          9711 => x"5f56597c",
          9712 => x"ae2e8438",
          9713 => x"728938ff",
          9714 => x"175776dd",
          9715 => x"38765977",
          9716 => x"19568076",
          9717 => x"2376802e",
          9718 => x"fec73880",
          9719 => x"78227083",
          9720 => x"ffff0672",
          9721 => x"585d5556",
          9722 => x"7aa02e82",
          9723 => x"e6387383",
          9724 => x"ffff0653",
          9725 => x"72ae2e82",
          9726 => x"f1387680",
          9727 => x"2eaa3877",
          9728 => x"19fe0570",
          9729 => x"225a5478",
          9730 => x"ae2e9d38",
          9731 => x"761018fe",
          9732 => x"0554ff17",
          9733 => x"5776802e",
          9734 => x"8f38fe14",
          9735 => x"70225e54",
          9736 => x"7cae2e09",
          9737 => x"8106eb38",
          9738 => x"8b0ba01d",
          9739 => x"5553a074",
          9740 => x"70810556",
          9741 => x"34ff1353",
          9742 => x"72f43872",
          9743 => x"735c5e88",
          9744 => x"78167022",
          9745 => x"81195957",
          9746 => x"545d7480",
          9747 => x"2e80ed38",
          9748 => x"74a02e83",
          9749 => x"d03874ae",
          9750 => x"32703070",
          9751 => x"8025555a",
          9752 => x"5475772e",
          9753 => x"85ce3872",
          9754 => x"83bb3872",
          9755 => x"597c7b26",
          9756 => x"83388159",
          9757 => x"75773270",
          9758 => x"30707207",
          9759 => x"8025707c",
          9760 => x"07515154",
          9761 => x"5472802e",
          9762 => x"83e0387c",
          9763 => x"8b2e8683",
          9764 => x"3875772e",
          9765 => x"8a387983",
          9766 => x"075a7577",
          9767 => x"269e3876",
          9768 => x"56885b8b",
          9769 => x"7e822b81",
          9770 => x"fc067718",
          9771 => x"575f5d77",
          9772 => x"15702281",
          9773 => x"18585653",
          9774 => x"74ff9538",
          9775 => x"a01c3357",
          9776 => x"7681e52e",
          9777 => x"8384387c",
          9778 => x"882e82e3",
          9779 => x"387d8c06",
          9780 => x"58778c2e",
          9781 => x"82ed387d",
          9782 => x"83065574",
          9783 => x"832e82e3",
          9784 => x"3879812a",
          9785 => x"81065675",
          9786 => x"9d387d81",
          9787 => x"065d7c80",
          9788 => x"2e853879",
          9789 => x"90075a7d",
          9790 => x"822a8106",
          9791 => x"5e7d802e",
          9792 => x"85387988",
          9793 => x"075a79ab",
          9794 => x"1d347b51",
          9795 => x"e4ec3f84",
          9796 => x"ba8c08ab",
          9797 => x"1d335654",
          9798 => x"84ba8c08",
          9799 => x"802e81ac",
          9800 => x"3884ba8c",
          9801 => x"08842e09",
          9802 => x"8106fbf7",
          9803 => x"3874852a",
          9804 => x"81065a79",
          9805 => x"802e84f0",
          9806 => x"3874822a",
          9807 => x"81065978",
          9808 => x"8298387b",
          9809 => x"08655556",
          9810 => x"73428c16",
          9811 => x"08588057",
          9812 => x"f9ce3981",
          9813 => x"16701179",
          9814 => x"11702240",
          9815 => x"4056567c",
          9816 => x"a02ef038",
          9817 => x"75802efd",
          9818 => x"85387983",
          9819 => x"075afd8a",
          9820 => x"39821822",
          9821 => x"5675ae2e",
          9822 => x"098106fc",
          9823 => x"ac387722",
          9824 => x"5473ae2e",
          9825 => x"098106fc",
          9826 => x"a0387610",
          9827 => x"185b807b",
          9828 => x"23800ba0",
          9829 => x"1d5653ae",
          9830 => x"54767326",
          9831 => x"8338a054",
          9832 => x"73757081",
          9833 => x"05573481",
          9834 => x"13538a73",
          9835 => x"27e93879",
          9836 => x"a0075877",
          9837 => x"ab1d347b",
          9838 => x"51e3bf3f",
          9839 => x"84ba8c08",
          9840 => x"ab1d3356",
          9841 => x"5484ba8c",
          9842 => x"08fed638",
          9843 => x"74822a81",
          9844 => x"065877fa",
          9845 => x"ce38861c",
          9846 => x"3370842a",
          9847 => x"8106565d",
          9848 => x"74802e83",
          9849 => x"cd38901c",
          9850 => x"0883ff06",
          9851 => x"600580d3",
          9852 => x"113380d2",
          9853 => x"12337188",
          9854 => x"2b076233",
          9855 => x"41575454",
          9856 => x"7d832e82",
          9857 => x"d8387488",
          9858 => x"1d0c7b08",
          9859 => x"655556fe",
          9860 => x"b7397722",
          9861 => x"5574ae2e",
          9862 => x"fef03876",
          9863 => x"175976fb",
          9864 => x"8838fbab",
          9865 => x"39798307",
          9866 => x"7617565a",
          9867 => x"fd81397d",
          9868 => x"822b81fc",
          9869 => x"06708c06",
          9870 => x"595e778c",
          9871 => x"2e098106",
          9872 => x"fd953879",
          9873 => x"82075afd",
          9874 => x"9839850b",
          9875 => x"a01d347c",
          9876 => x"882e0981",
          9877 => x"06fcf638",
          9878 => x"d639ff80",
          9879 => x"0bab1d34",
          9880 => x"800b84ba",
          9881 => x"8c0c933d",
          9882 => x"0d047480",
          9883 => x"ff269d38",
          9884 => x"81ff7527",
          9885 => x"80c938ff",
          9886 => x"1d59787b",
          9887 => x"2681f738",
          9888 => x"7983077d",
          9889 => x"7718575c",
          9890 => x"5afca439",
          9891 => x"7982075a",
          9892 => x"83b55274",
          9893 => x"518185f6",
          9894 => x"3f84ba8c",
          9895 => x"0883ffff",
          9896 => x"0670872a",
          9897 => x"81065a55",
          9898 => x"78802ec4",
          9899 => x"387480ff",
          9900 => x"0683e69c",
          9901 => x"11335654",
          9902 => x"7481ff26",
          9903 => x"ffb93874",
          9904 => x"802e8185",
          9905 => x"3883e5b4",
          9906 => x"0b83e5b4",
          9907 => x"337081ff",
          9908 => x"06565459",
          9909 => x"73802e80",
          9910 => x"e0387375",
          9911 => x"2e8f3881",
          9912 => x"19703370",
          9913 => x"81ff0656",
          9914 => x"545973ee",
          9915 => x"387281ff",
          9916 => x"06597880",
          9917 => x"d438ffbf",
          9918 => x"15547399",
          9919 => x"268a387d",
          9920 => x"82077081",
          9921 => x"ff065f53",
          9922 => x"ff9f1559",
          9923 => x"78992693",
          9924 => x"387d8107",
          9925 => x"7081ff06",
          9926 => x"e0177083",
          9927 => x"ffff0658",
          9928 => x"565f537b",
          9929 => x"1ba00559",
          9930 => x"74793481",
          9931 => x"1b5b7516",
          9932 => x"55fafc39",
          9933 => x"8053fab3",
          9934 => x"3983e5b4",
          9935 => x"337081ff",
          9936 => x"065a5378",
          9937 => x"802effae",
          9938 => x"3880df7a",
          9939 => x"83077d1d",
          9940 => x"a0055b5b",
          9941 => x"55747934",
          9942 => x"811b5bd2",
          9943 => x"3980cd14",
          9944 => x"3380cc15",
          9945 => x"3371982b",
          9946 => x"71902b07",
          9947 => x"7707881f",
          9948 => x"0c5a57fd",
          9949 => x"95397b1b",
          9950 => x"a0057588",
          9951 => x"2a545472",
          9952 => x"7434811b",
          9953 => x"7c11a005",
          9954 => x"5a5b7479",
          9955 => x"34811b5b",
          9956 => x"ff9c3979",
          9957 => x"8307a01d",
          9958 => x"33585a76",
          9959 => x"81e52e09",
          9960 => x"8106faa3",
          9961 => x"38fda339",
          9962 => x"74822a81",
          9963 => x"065c7bf6",
          9964 => x"f238850b",
          9965 => x"84ba8c0c",
          9966 => x"933d0d04",
          9967 => x"eb3d0d67",
          9968 => x"69028805",
          9969 => x"80e70533",
          9970 => x"42425e80",
          9971 => x"610cff7e",
          9972 => x"0870595b",
          9973 => x"4279802e",
          9974 => x"85d73879",
          9975 => x"7081055b",
          9976 => x"33709f26",
          9977 => x"565675ba",
          9978 => x"2e85d038",
          9979 => x"74ed3875",
          9980 => x"ba2e85c7",
          9981 => x"3884d1e8",
          9982 => x"33568076",
          9983 => x"2485b238",
          9984 => x"75101084",
          9985 => x"d1d40570",
          9986 => x"08585a8c",
          9987 => x"5876802e",
          9988 => x"85963876",
          9989 => x"610c7f81",
          9990 => x"fe067733",
          9991 => x"5d597b80",
          9992 => x"2e9b3881",
          9993 => x"173351ff",
          9994 => x"bbb03f84",
          9995 => x"ba8c0881",
          9996 => x"ff067081",
          9997 => x"065e587c",
          9998 => x"802e8696",
          9999 => x"38807734",
         10000 => x"75165d84",
         10001 => x"ba801d33",
         10002 => x"81183481",
         10003 => x"52811733",
         10004 => x"51ffbba4",
         10005 => x"3f84ba8c",
         10006 => x"0881ff06",
         10007 => x"70810641",
         10008 => x"5683587f",
         10009 => x"84c23878",
         10010 => x"802e8d38",
         10011 => x"75822a81",
         10012 => x"06418a58",
         10013 => x"6084b138",
         10014 => x"805b7a83",
         10015 => x"1834ff0b",
         10016 => x"b4180c7a",
         10017 => x"7b5a5581",
         10018 => x"547a53b8",
         10019 => x"17705381",
         10020 => x"18335258",
         10021 => x"ffbb953f",
         10022 => x"84ba8c08",
         10023 => x"7b2e8538",
         10024 => x"ff558159",
         10025 => x"74b4180c",
         10026 => x"84567899",
         10027 => x"3884b717",
         10028 => x"3384b618",
         10029 => x"3371882b",
         10030 => x"07565683",
         10031 => x"567482d4",
         10032 => x"d52e85a5",
         10033 => x"38758126",
         10034 => x"8b3884ba",
         10035 => x"811d3342",
         10036 => x"6185bf38",
         10037 => x"81587584",
         10038 => x"2e83cd38",
         10039 => x"8d587581",
         10040 => x"2683c538",
         10041 => x"80c41733",
         10042 => x"80c31833",
         10043 => x"71882b07",
         10044 => x"5e597c84",
         10045 => x"802e0981",
         10046 => x"0683ad38",
         10047 => x"80cf1733",
         10048 => x"80ce1833",
         10049 => x"71882b07",
         10050 => x"575a75a4",
         10051 => x"3880dc17",
         10052 => x"83113382",
         10053 => x"12337190",
         10054 => x"2b71882b",
         10055 => x"07811433",
         10056 => x"70720788",
         10057 => x"2b753371",
         10058 => x"07565a45",
         10059 => x"435e5f56",
         10060 => x"75a0180c",
         10061 => x"80c81733",
         10062 => x"82183480",
         10063 => x"c81733ff",
         10064 => x"117081ff",
         10065 => x"065f4059",
         10066 => x"8d587c81",
         10067 => x"2682d938",
         10068 => x"7881ff06",
         10069 => x"76712980",
         10070 => x"c519335a",
         10071 => x"5f5a778a",
         10072 => x"18237759",
         10073 => x"77802e87",
         10074 => x"c438ff18",
         10075 => x"78064261",
         10076 => x"87bb3880",
         10077 => x"ca173380",
         10078 => x"c9183371",
         10079 => x"882b0756",
         10080 => x"40748818",
         10081 => x"2374758f",
         10082 => x"065e5a8d",
         10083 => x"587c8298",
         10084 => x"3880cc17",
         10085 => x"3380cb18",
         10086 => x"3371882b",
         10087 => x"07565c74",
         10088 => x"a43880d8",
         10089 => x"17831133",
         10090 => x"82123371",
         10091 => x"902b7188",
         10092 => x"2b078114",
         10093 => x"33707207",
         10094 => x"882b7533",
         10095 => x"71075344",
         10096 => x"5a584242",
         10097 => x"4280c717",
         10098 => x"3380c618",
         10099 => x"3371882b",
         10100 => x"075d588d",
         10101 => x"587b802e",
         10102 => x"81ce387d",
         10103 => x"1c7a842a",
         10104 => x"055a7975",
         10105 => x"2681c138",
         10106 => x"7852747a",
         10107 => x"3151fded",
         10108 => x"b43f84ba",
         10109 => x"8c085684",
         10110 => x"ba8c0880",
         10111 => x"2e81a938",
         10112 => x"84ba8c08",
         10113 => x"80ffffff",
         10114 => x"f5268338",
         10115 => x"835d7583",
         10116 => x"fff52683",
         10117 => x"38825d75",
         10118 => x"9ff52685",
         10119 => x"eb38815d",
         10120 => x"8216709c",
         10121 => x"190c7ba4",
         10122 => x"190c7b1d",
         10123 => x"70a81a0c",
         10124 => x"7b1db01a",
         10125 => x"0c57597c",
         10126 => x"832e8a87",
         10127 => x"38881722",
         10128 => x"5c8d587b",
         10129 => x"802e80e0",
         10130 => x"387d16ac",
         10131 => x"180c7819",
         10132 => x"557c822e",
         10133 => x"8d387810",
         10134 => x"1970812a",
         10135 => x"7a810605",
         10136 => x"565a83ff",
         10137 => x"15892a59",
         10138 => x"8d5878a0",
         10139 => x"180826b8",
         10140 => x"38ff0b94",
         10141 => x"180cff0b",
         10142 => x"90180cff",
         10143 => x"800b8418",
         10144 => x"347c832e",
         10145 => x"8696387c",
         10146 => x"773484d1",
         10147 => x"e4228105",
         10148 => x"5d7c84d1",
         10149 => x"e4237c86",
         10150 => x"182384d1",
         10151 => x"ec0b8c18",
         10152 => x"0c800b98",
         10153 => x"180c8058",
         10154 => x"7784ba8c",
         10155 => x"0c973d0d",
         10156 => x"048b0b84",
         10157 => x"ba8c0c97",
         10158 => x"3d0d0476",
         10159 => x"33d01170",
         10160 => x"81ff0657",
         10161 => x"57587489",
         10162 => x"26913882",
         10163 => x"177881ff",
         10164 => x"06d0055d",
         10165 => x"59787a2e",
         10166 => x"87fe3880",
         10167 => x"7e0883e5",
         10168 => x"fc5f405c",
         10169 => x"7c087f5a",
         10170 => x"5b7a7081",
         10171 => x"055c3379",
         10172 => x"7081055b",
         10173 => x"33ff9f12",
         10174 => x"5a585677",
         10175 => x"99268938",
         10176 => x"e0167081",
         10177 => x"ff065755",
         10178 => x"ff9f1758",
         10179 => x"77992689",
         10180 => x"38e01770",
         10181 => x"81ff0658",
         10182 => x"55753070",
         10183 => x"9f2a5955",
         10184 => x"75772e09",
         10185 => x"81068538",
         10186 => x"77ffbe38",
         10187 => x"787a3270",
         10188 => x"30707207",
         10189 => x"9f2a7a07",
         10190 => x"5d58557a",
         10191 => x"802e8798",
         10192 => x"38811c84",
         10193 => x"1e5e5c83",
         10194 => x"7c25ff98",
         10195 => x"386156f9",
         10196 => x"a9397880",
         10197 => x"2efecf38",
         10198 => x"77822a81",
         10199 => x"065e8a58",
         10200 => x"7dfec538",
         10201 => x"8058fec0",
         10202 => x"397a7833",
         10203 => x"57597581",
         10204 => x"e92e0981",
         10205 => x"06833881",
         10206 => x"597581eb",
         10207 => x"32703070",
         10208 => x"80257b07",
         10209 => x"5a5b5c77",
         10210 => x"83ad3875",
         10211 => x"81e82e83",
         10212 => x"a638933d",
         10213 => x"77575a83",
         10214 => x"5983fa16",
         10215 => x"3370595b",
         10216 => x"7a802ea5",
         10217 => x"38848116",
         10218 => x"33848017",
         10219 => x"3371902b",
         10220 => x"71882b07",
         10221 => x"83ff1933",
         10222 => x"70720788",
         10223 => x"2b83fe1b",
         10224 => x"33710752",
         10225 => x"595b4040",
         10226 => x"40777a70",
         10227 => x"84055c0c",
         10228 => x"ff199017",
         10229 => x"57597880",
         10230 => x"25ffbe38",
         10231 => x"84ba811d",
         10232 => x"33703070",
         10233 => x"9f2a7271",
         10234 => x"319b3d71",
         10235 => x"101005f0",
         10236 => x"0584b61c",
         10237 => x"445d5243",
         10238 => x"5b427808",
         10239 => x"5b83567a",
         10240 => x"802e80fb",
         10241 => x"38800b83",
         10242 => x"1834ff0b",
         10243 => x"b4180c7a",
         10244 => x"5580567a",
         10245 => x"ff2ea538",
         10246 => x"81547a53",
         10247 => x"b8175281",
         10248 => x"173351ff",
         10249 => x"b4863f84",
         10250 => x"ba8c0876",
         10251 => x"2e8538ff",
         10252 => x"55815674",
         10253 => x"b4180c84",
         10254 => x"5875bf38",
         10255 => x"811f337f",
         10256 => x"3371882b",
         10257 => x"075d5e83",
         10258 => x"587b82d4",
         10259 => x"d52e0981",
         10260 => x"06a83880",
         10261 => x"0bb81833",
         10262 => x"57587581",
         10263 => x"e92e82b7",
         10264 => x"387581eb",
         10265 => x"32703070",
         10266 => x"80257a07",
         10267 => x"4242427f",
         10268 => x"bc387581",
         10269 => x"e82eb638",
         10270 => x"82587781",
         10271 => x"ff065680",
         10272 => x"0b84ba81",
         10273 => x"1e335d58",
         10274 => x"7b782e09",
         10275 => x"81068338",
         10276 => x"81588176",
         10277 => x"27f8bd38",
         10278 => x"77802ef8",
         10279 => x"b738811a",
         10280 => x"841a5a5a",
         10281 => x"837a27fe",
         10282 => x"d138f8a8",
         10283 => x"39830b80",
         10284 => x"ee1883e5",
         10285 => x"bc405d58",
         10286 => x"7b708105",
         10287 => x"5d337e70",
         10288 => x"81054033",
         10289 => x"717131ff",
         10290 => x"1b5b5256",
         10291 => x"5677802e",
         10292 => x"80c53875",
         10293 => x"802ee138",
         10294 => x"850b818a",
         10295 => x"1883e5c0",
         10296 => x"405d587b",
         10297 => x"7081055d",
         10298 => x"337e7081",
         10299 => x"05403371",
         10300 => x"7131ff1b",
         10301 => x"5b584240",
         10302 => x"77802e85",
         10303 => x"8e387580",
         10304 => x"2ee13882",
         10305 => x"58fef339",
         10306 => x"8d587cfa",
         10307 => x"93387784",
         10308 => x"ba8c0c97",
         10309 => x"3d0d0475",
         10310 => x"5875802e",
         10311 => x"fedc3885",
         10312 => x"0b818a18",
         10313 => x"83e5c040",
         10314 => x"5d58ffb7",
         10315 => x"398d0b84",
         10316 => x"ba8c0c97",
         10317 => x"3d0d0483",
         10318 => x"0b80ee18",
         10319 => x"83e5bc5c",
         10320 => x"5a587870",
         10321 => x"81055a33",
         10322 => x"7a708105",
         10323 => x"5c337171",
         10324 => x"31ff1b5b",
         10325 => x"575f5f77",
         10326 => x"802e83d1",
         10327 => x"3874802e",
         10328 => x"e138850b",
         10329 => x"818a1883",
         10330 => x"e5c05c5a",
         10331 => x"58787081",
         10332 => x"055a337a",
         10333 => x"7081055c",
         10334 => x"33717131",
         10335 => x"ff1b5b58",
         10336 => x"42407780",
         10337 => x"2e849138",
         10338 => x"75802ee1",
         10339 => x"38933d77",
         10340 => x"575a8359",
         10341 => x"fc833981",
         10342 => x"58fdc639",
         10343 => x"80e91733",
         10344 => x"80e81833",
         10345 => x"71882b07",
         10346 => x"57557581",
         10347 => x"2e098106",
         10348 => x"f9d53881",
         10349 => x"1b58805a",
         10350 => x"b4170878",
         10351 => x"2eb13883",
         10352 => x"17335b7a",
         10353 => x"7a2e0981",
         10354 => x"06829b38",
         10355 => x"81547753",
         10356 => x"b8175281",
         10357 => x"173351ff",
         10358 => x"b0d23f84",
         10359 => x"ba8c0880",
         10360 => x"2e8538ff",
         10361 => x"58815a77",
         10362 => x"b4180c79",
         10363 => x"f9993879",
         10364 => x"84183484",
         10365 => x"b7173384",
         10366 => x"b6183371",
         10367 => x"882b0757",
         10368 => x"5e7582d4",
         10369 => x"d52e0981",
         10370 => x"06f8fc38",
         10371 => x"b8178311",
         10372 => x"33821233",
         10373 => x"71902b71",
         10374 => x"882b0781",
         10375 => x"14337072",
         10376 => x"07882b75",
         10377 => x"3371075e",
         10378 => x"41594542",
         10379 => x"5c597784",
         10380 => x"8b85a4d2",
         10381 => x"2e098106",
         10382 => x"f8cd3884",
         10383 => x"9c178311",
         10384 => x"33821233",
         10385 => x"71902b71",
         10386 => x"882b0781",
         10387 => x"14337072",
         10388 => x"07882b75",
         10389 => x"33710747",
         10390 => x"44405b5c",
         10391 => x"5a5e6086",
         10392 => x"8a85e4f2",
         10393 => x"2e098106",
         10394 => x"f89d3884",
         10395 => x"a0178311",
         10396 => x"33821233",
         10397 => x"71902b71",
         10398 => x"882b0781",
         10399 => x"14337072",
         10400 => x"07882b75",
         10401 => x"33710794",
         10402 => x"1e0c5d84",
         10403 => x"a41c8311",
         10404 => x"33821233",
         10405 => x"71902b71",
         10406 => x"882b0781",
         10407 => x"14337072",
         10408 => x"07882b75",
         10409 => x"33710762",
         10410 => x"90050c59",
         10411 => x"4449465c",
         10412 => x"4540455b",
         10413 => x"565a7c77",
         10414 => x"3484d1e4",
         10415 => x"2281055d",
         10416 => x"7c84d1e4",
         10417 => x"237c8618",
         10418 => x"2384d1ec",
         10419 => x"0b8c180c",
         10420 => x"800b9818",
         10421 => x"0cf7cf39",
         10422 => x"7b8324f8",
         10423 => x"f0387b7a",
         10424 => x"7f0c56f2",
         10425 => x"95397554",
         10426 => x"b4170853",
         10427 => x"b8177053",
         10428 => x"81183352",
         10429 => x"59ffafb3",
         10430 => x"3f84ba8c",
         10431 => x"087a2e09",
         10432 => x"810681a4",
         10433 => x"3884ba8c",
         10434 => x"08831834",
         10435 => x"b41708a8",
         10436 => x"18083140",
         10437 => x"7fa01808",
         10438 => x"278b3882",
         10439 => x"17334160",
         10440 => x"822e818d",
         10441 => x"3884ba8c",
         10442 => x"085afda0",
         10443 => x"39745674",
         10444 => x"802ef391",
         10445 => x"38850b81",
         10446 => x"8a1883e5",
         10447 => x"c05c5a58",
         10448 => x"fcab3980",
         10449 => x"e3173380",
         10450 => x"e2183371",
         10451 => x"882b075f",
         10452 => x"5a8d587d",
         10453 => x"f6d23888",
         10454 => x"17224261",
         10455 => x"f6ca3880",
         10456 => x"e4178311",
         10457 => x"33821233",
         10458 => x"71902b71",
         10459 => x"882b0781",
         10460 => x"14337072",
         10461 => x"07882b75",
         10462 => x"337107ac",
         10463 => x"1e0c5a7d",
         10464 => x"822b5a43",
         10465 => x"44405940",
         10466 => x"f5d83975",
         10467 => x"5875802e",
         10468 => x"f9e83882",
         10469 => x"58f9e339",
         10470 => x"75802ef2",
         10471 => x"a838933d",
         10472 => x"77575a83",
         10473 => x"59f7f239",
         10474 => x"755a79f5",
         10475 => x"da38fcbf",
         10476 => x"397554b4",
         10477 => x"1708a018",
         10478 => x"08055378",
         10479 => x"52811733",
         10480 => x"51ffade7",
         10481 => x"3ffc8539",
         10482 => x"f03d0d02",
         10483 => x"80d30533",
         10484 => x"64704393",
         10485 => x"3d41575d",
         10486 => x"ff765a40",
         10487 => x"75802e80",
         10488 => x"e9387870",
         10489 => x"81055a33",
         10490 => x"709f2655",
         10491 => x"5574ba2e",
         10492 => x"80e23873",
         10493 => x"ed3874ba",
         10494 => x"2e80d938",
         10495 => x"84d1e833",
         10496 => x"54807424",
         10497 => x"80c43873",
         10498 => x"101084d1",
         10499 => x"d4057008",
         10500 => x"55557380",
         10501 => x"2e843880",
         10502 => x"74346254",
         10503 => x"73802e86",
         10504 => x"38807434",
         10505 => x"62547375",
         10506 => x"0c7c547c",
         10507 => x"802e9238",
         10508 => x"8053933d",
         10509 => x"70538405",
         10510 => x"51ef813f",
         10511 => x"84ba8c08",
         10512 => x"547384ba",
         10513 => x"8c0c923d",
         10514 => x"0d048b0b",
         10515 => x"84ba8c0c",
         10516 => x"923d0d04",
         10517 => x"7533d011",
         10518 => x"7081ff06",
         10519 => x"56565773",
         10520 => x"89269138",
         10521 => x"82167781",
         10522 => x"ff06d005",
         10523 => x"5c587779",
         10524 => x"2e80f738",
         10525 => x"807f0883",
         10526 => x"e5fc5e5f",
         10527 => x"5b7b087e",
         10528 => x"595a7970",
         10529 => x"81055b33",
         10530 => x"78708105",
         10531 => x"5a33ff9f",
         10532 => x"12595755",
         10533 => x"76992689",
         10534 => x"38e01570",
         10535 => x"81ff0656",
         10536 => x"54ff9f16",
         10537 => x"57769926",
         10538 => x"8938e016",
         10539 => x"7081ff06",
         10540 => x"57547430",
         10541 => x"709f2a58",
         10542 => x"5474762e",
         10543 => x"09810685",
         10544 => x"3876ffbe",
         10545 => x"38777932",
         10546 => x"70307072",
         10547 => x"079f2a79",
         10548 => x"075c5754",
         10549 => x"79802e92",
         10550 => x"38811b84",
         10551 => x"1d5d5b83",
         10552 => x"7b25ff99",
         10553 => x"387f54fe",
         10554 => x"98397a83",
         10555 => x"24f7387a",
         10556 => x"79600c54",
         10557 => x"fe8b39e6",
         10558 => x"3d0d6c02",
         10559 => x"840580fb",
         10560 => x"05335659",
         10561 => x"89567880",
         10562 => x"2ea63874",
         10563 => x"bf067054",
         10564 => x"9d3dcc05",
         10565 => x"539e3d84",
         10566 => x"055258ed",
         10567 => x"9f3f84ba",
         10568 => x"8c085784",
         10569 => x"ba8c0880",
         10570 => x"2e8f3880",
         10571 => x"790c7656",
         10572 => x"7584ba8c",
         10573 => x"0c9c3d0d",
         10574 => x"047e406d",
         10575 => x"52903d70",
         10576 => x"525ae19a",
         10577 => x"3f84ba8c",
         10578 => x"085784ba",
         10579 => x"8c08802e",
         10580 => x"81ba3877",
         10581 => x"9c065d7c",
         10582 => x"802e81ca",
         10583 => x"3876802e",
         10584 => x"83c13876",
         10585 => x"842e83ea",
         10586 => x"38778807",
         10587 => x"5876ffbb",
         10588 => x"3877832a",
         10589 => x"81065b7a",
         10590 => x"802e81d1",
         10591 => x"38669b11",
         10592 => x"339a1233",
         10593 => x"71882b07",
         10594 => x"61703342",
         10595 => x"585e5e56",
         10596 => x"7d832e84",
         10597 => x"e938800b",
         10598 => x"8e173480",
         10599 => x"0b8f1734",
         10600 => x"a10b9017",
         10601 => x"3480cc0b",
         10602 => x"91173466",
         10603 => x"56a00b8b",
         10604 => x"17347e67",
         10605 => x"575e800b",
         10606 => x"9a173480",
         10607 => x"0b9b1734",
         10608 => x"7d335d7c",
         10609 => x"832e84a9",
         10610 => x"38665b80",
         10611 => x"0b9c1c34",
         10612 => x"800b9d1c",
         10613 => x"34800b9e",
         10614 => x"1c34800b",
         10615 => x"9f1c347e",
         10616 => x"55810b83",
         10617 => x"16347b80",
         10618 => x"2e80e238",
         10619 => x"7eb41108",
         10620 => x"7d7c0853",
         10621 => x"575f5781",
         10622 => x"7c278938",
         10623 => x"9c17087c",
         10624 => x"26838a38",
         10625 => x"82578079",
         10626 => x"0cfea339",
         10627 => x"0280e705",
         10628 => x"3370982b",
         10629 => x"5d5b7b80",
         10630 => x"25feb838",
         10631 => x"86789c06",
         10632 => x"5e577cfe",
         10633 => x"b83876fe",
         10634 => x"82380280",
         10635 => x"c2053370",
         10636 => x"842a8106",
         10637 => x"5d567b82",
         10638 => x"91387781",
         10639 => x"2a81065e",
         10640 => x"7d802e89",
         10641 => x"38758106",
         10642 => x"5a7981f6",
         10643 => x"3877832a",
         10644 => x"81065675",
         10645 => x"802e8638",
         10646 => x"7780c007",
         10647 => x"587eb411",
         10648 => x"08a01b0c",
         10649 => x"67a41b0c",
         10650 => x"679b1133",
         10651 => x"9a123371",
         10652 => x"882b0773",
         10653 => x"33405e40",
         10654 => x"575a7b83",
         10655 => x"2e81f138",
         10656 => x"7a881a0c",
         10657 => x"9c168311",
         10658 => x"33821233",
         10659 => x"71902b71",
         10660 => x"882b0781",
         10661 => x"14337072",
         10662 => x"07882b75",
         10663 => x"33710770",
         10664 => x"608c050c",
         10665 => x"60600c51",
         10666 => x"52415957",
         10667 => x"5d5e861a",
         10668 => x"22841a23",
         10669 => x"77901a34",
         10670 => x"800b911a",
         10671 => x"34800b9c",
         10672 => x"1a0c7785",
         10673 => x"2a810655",
         10674 => x"74802e84",
         10675 => x"ac387580",
         10676 => x"2e84f138",
         10677 => x"75941a0c",
         10678 => x"8a1a2270",
         10679 => x"892b7c52",
         10680 => x"5b587630",
         10681 => x"70780780",
         10682 => x"25565b79",
         10683 => x"76278492",
         10684 => x"38817076",
         10685 => x"065f5b7d",
         10686 => x"802e8486",
         10687 => x"38775278",
         10688 => x"51ffacdb",
         10689 => x"3f84ba8c",
         10690 => x"085884ba",
         10691 => x"8c088126",
         10692 => x"83388257",
         10693 => x"84ba8c08",
         10694 => x"ff2e80cb",
         10695 => x"38757a31",
         10696 => x"56c03902",
         10697 => x"80c20533",
         10698 => x"91065e7d",
         10699 => x"95387782",
         10700 => x"2a810655",
         10701 => x"74802efc",
         10702 => x"b8388857",
         10703 => x"80790cfb",
         10704 => x"ed398757",
         10705 => x"80790cfb",
         10706 => x"e5398457",
         10707 => x"80790cfb",
         10708 => x"dd397951",
         10709 => x"cdca3f84",
         10710 => x"ba8c0878",
         10711 => x"88075957",
         10712 => x"76fbc838",
         10713 => x"fc8b397a",
         10714 => x"767b3157",
         10715 => x"57fef339",
         10716 => x"95163394",
         10717 => x"17337198",
         10718 => x"2b71902b",
         10719 => x"077d075d",
         10720 => x"5e5cfdfc",
         10721 => x"397c557c",
         10722 => x"7b2781bd",
         10723 => x"38745279",
         10724 => x"51ffabcb",
         10725 => x"3f84ba8c",
         10726 => x"085d84ba",
         10727 => x"8c08802e",
         10728 => x"81a73884",
         10729 => x"ba8c0881",
         10730 => x"2efcd938",
         10731 => x"84ba8c08",
         10732 => x"ff2e8399",
         10733 => x"38805374",
         10734 => x"527651ff",
         10735 => x"b2823f84",
         10736 => x"ba8c0883",
         10737 => x"90389c17",
         10738 => x"08fe1194",
         10739 => x"19085856",
         10740 => x"5b757527",
         10741 => x"ffaf3881",
         10742 => x"1694180c",
         10743 => x"84173381",
         10744 => x"07557484",
         10745 => x"18347c55",
         10746 => x"7a7d26ff",
         10747 => x"a03880d9",
         10748 => x"39800b94",
         10749 => x"1734800b",
         10750 => x"951734fb",
         10751 => x"cc399516",
         10752 => x"33941733",
         10753 => x"71982b71",
         10754 => x"902b077e",
         10755 => x"075e565b",
         10756 => x"800b8e17",
         10757 => x"34800b8f",
         10758 => x"1734a10b",
         10759 => x"90173480",
         10760 => x"cc0b9117",
         10761 => x"346656a0",
         10762 => x"0b8b1734",
         10763 => x"7e67575e",
         10764 => x"800b9a17",
         10765 => x"34800b9b",
         10766 => x"17347d33",
         10767 => x"5d7c832e",
         10768 => x"098106fb",
         10769 => x"8438ffa9",
         10770 => x"39807f7f",
         10771 => x"725e5957",
         10772 => x"5db41608",
         10773 => x"7e2eae38",
         10774 => x"8316335a",
         10775 => x"797d2e09",
         10776 => x"8106b538",
         10777 => x"81547d53",
         10778 => x"b8165281",
         10779 => x"163351ff",
         10780 => x"a3ba3f84",
         10781 => x"ba8c0880",
         10782 => x"2e8538ff",
         10783 => x"57815b76",
         10784 => x"b4170c7e",
         10785 => x"567aff1d",
         10786 => x"90180c57",
         10787 => x"7a802efb",
         10788 => x"bc388079",
         10789 => x"0cf99739",
         10790 => x"8154b416",
         10791 => x"0853b816",
         10792 => x"70538117",
         10793 => x"33525aff",
         10794 => x"a4813f84",
         10795 => x"ba8c087d",
         10796 => x"2e098106",
         10797 => x"81aa3884",
         10798 => x"ba8c0883",
         10799 => x"1734b416",
         10800 => x"08a81708",
         10801 => x"3184ba8c",
         10802 => x"085c5574",
         10803 => x"a0170827",
         10804 => x"ff923882",
         10805 => x"16335574",
         10806 => x"822e0981",
         10807 => x"06ff8538",
         10808 => x"8154b416",
         10809 => x"08a01708",
         10810 => x"05537952",
         10811 => x"81163351",
         10812 => x"ffa3b83f",
         10813 => x"7c5bfeec",
         10814 => x"3974941a",
         10815 => x"0c7656f8",
         10816 => x"af397798",
         10817 => x"1a0c76f8",
         10818 => x"a2387583",
         10819 => x"ff065a79",
         10820 => x"802ef89a",
         10821 => x"387efe19",
         10822 => x"9c1208fe",
         10823 => x"055f595a",
         10824 => x"777d27f9",
         10825 => x"df388a1a",
         10826 => x"22787129",
         10827 => x"b01c0805",
         10828 => x"565c7480",
         10829 => x"2ef9cd38",
         10830 => x"75892a15",
         10831 => x"9c1a0c76",
         10832 => x"56f7ed39",
         10833 => x"75941a0c",
         10834 => x"7656f7e4",
         10835 => x"39815780",
         10836 => x"790cf7da",
         10837 => x"3984ba8c",
         10838 => x"08578079",
         10839 => x"0cf7cf39",
         10840 => x"817f575b",
         10841 => x"fe9f39f0",
         10842 => x"3d0d6265",
         10843 => x"67664040",
         10844 => x"5d5a807e",
         10845 => x"0c895779",
         10846 => x"802e9f38",
         10847 => x"79085675",
         10848 => x"802e9738",
         10849 => x"75335574",
         10850 => x"802e8f38",
         10851 => x"86162284",
         10852 => x"1b225959",
         10853 => x"78782e84",
         10854 => x"b7388055",
         10855 => x"74417655",
         10856 => x"76828c38",
         10857 => x"911a3355",
         10858 => x"74828438",
         10859 => x"901a3381",
         10860 => x"06578756",
         10861 => x"76802e81",
         10862 => x"ed38941a",
         10863 => x"088c1b08",
         10864 => x"71315656",
         10865 => x"7b752681",
         10866 => x"ef387b80",
         10867 => x"2e81d538",
         10868 => x"60597583",
         10869 => x"ff065b7a",
         10870 => x"81e3388a",
         10871 => x"1922ff05",
         10872 => x"76892a06",
         10873 => x"5b7a9b38",
         10874 => x"7583d338",
         10875 => x"881a0855",
         10876 => x"81752784",
         10877 => x"853874ff",
         10878 => x"2e83f038",
         10879 => x"74981b0c",
         10880 => x"6059981a",
         10881 => x"08fe059c",
         10882 => x"1a08fe05",
         10883 => x"41577660",
         10884 => x"2783e738",
         10885 => x"8a192270",
         10886 => x"7829b01b",
         10887 => x"08055656",
         10888 => x"74802e83",
         10889 => x"d5387a15",
         10890 => x"7c892a59",
         10891 => x"5777802e",
         10892 => x"83813877",
         10893 => x"1b557575",
         10894 => x"27853875",
         10895 => x"7b315877",
         10896 => x"5476537c",
         10897 => x"52811933",
         10898 => x"51ff9fe0",
         10899 => x"3f84ba8c",
         10900 => x"08839838",
         10901 => x"60831133",
         10902 => x"57597580",
         10903 => x"2ea938b4",
         10904 => x"19087731",
         10905 => x"56757827",
         10906 => x"9e388480",
         10907 => x"7671291e",
         10908 => x"b81b5858",
         10909 => x"55757081",
         10910 => x"05573377",
         10911 => x"70810559",
         10912 => x"34ff1555",
         10913 => x"74ef3877",
         10914 => x"892b587b",
         10915 => x"78317e08",
         10916 => x"197f0c78",
         10917 => x"1e941c08",
         10918 => x"1a705994",
         10919 => x"1d0c5e5c",
         10920 => x"7bfeaf38",
         10921 => x"80567584",
         10922 => x"ba8c0c92",
         10923 => x"3d0d0474",
         10924 => x"84ba8c0c",
         10925 => x"923d0d04",
         10926 => x"745cfe8e",
         10927 => x"399c1a08",
         10928 => x"577583ff",
         10929 => x"06848071",
         10930 => x"31595b7b",
         10931 => x"78278338",
         10932 => x"7b587656",
         10933 => x"b4190877",
         10934 => x"2eb63880",
         10935 => x"0b831a33",
         10936 => x"715d415f",
         10937 => x"7f7f2e09",
         10938 => x"810680e4",
         10939 => x"38815476",
         10940 => x"53b81952",
         10941 => x"81193351",
         10942 => x"ff9eb13f",
         10943 => x"84ba8c08",
         10944 => x"802e8538",
         10945 => x"ff56815b",
         10946 => x"75b41a0c",
         10947 => x"7a81dc38",
         10948 => x"60941b08",
         10949 => x"83ff0611",
         10950 => x"797f5a58",
         10951 => x"b8055659",
         10952 => x"77802efe",
         10953 => x"e6387470",
         10954 => x"81055633",
         10955 => x"77708105",
         10956 => x"5934ff16",
         10957 => x"5675802e",
         10958 => x"fed13874",
         10959 => x"70810556",
         10960 => x"33777081",
         10961 => x"055934ff",
         10962 => x"165675da",
         10963 => x"38febc39",
         10964 => x"8154b419",
         10965 => x"0853b819",
         10966 => x"7053811a",
         10967 => x"335240ff",
         10968 => x"9ec93f81",
         10969 => x"5b84ba8c",
         10970 => x"087f2e09",
         10971 => x"8106ff9c",
         10972 => x"3884ba8c",
         10973 => x"08831a34",
         10974 => x"b41908a8",
         10975 => x"1a083184",
         10976 => x"ba8c085c",
         10977 => x"5574a01a",
         10978 => x"0827fee1",
         10979 => x"38821933",
         10980 => x"5574822e",
         10981 => x"098106fe",
         10982 => x"d4388154",
         10983 => x"b41908a0",
         10984 => x"1a080553",
         10985 => x"7f528119",
         10986 => x"3351ff9d",
         10987 => x"fe3f7e5b",
         10988 => x"febb3976",
         10989 => x"9c1b0c94",
         10990 => x"1a0856fe",
         10991 => x"8439981a",
         10992 => x"08527951",
         10993 => x"ffa3983f",
         10994 => x"84ba8c08",
         10995 => x"55fca139",
         10996 => x"81163351",
         10997 => x"ff9c833f",
         10998 => x"84ba8c08",
         10999 => x"81065574",
         11000 => x"fbb83874",
         11001 => x"7a085657",
         11002 => x"fbb23981",
         11003 => x"0b911b34",
         11004 => x"810b84ba",
         11005 => x"8c0c923d",
         11006 => x"0d04820b",
         11007 => x"911b3482",
         11008 => x"0b84ba8c",
         11009 => x"0c923d0d",
         11010 => x"04f03d0d",
         11011 => x"62656766",
         11012 => x"40405c5a",
         11013 => x"807e0c89",
         11014 => x"5779802e",
         11015 => x"9f387908",
         11016 => x"5675802e",
         11017 => x"97387533",
         11018 => x"5574802e",
         11019 => x"8f388616",
         11020 => x"22841b22",
         11021 => x"59597878",
         11022 => x"2e85fd38",
         11023 => x"80557441",
         11024 => x"76557682",
         11025 => x"c438911a",
         11026 => x"33557482",
         11027 => x"bc38901a",
         11028 => x"3370812a",
         11029 => x"81065858",
         11030 => x"87567680",
         11031 => x"2e82a138",
         11032 => x"941a087b",
         11033 => x"115d577b",
         11034 => x"77278438",
         11035 => x"76095b7a",
         11036 => x"802e8281",
         11037 => x"387683ff",
         11038 => x"065f7e82",
         11039 => x"a238608a",
         11040 => x"1122ff05",
         11041 => x"78892a06",
         11042 => x"5a5678aa",
         11043 => x"3876849e",
         11044 => x"38881a08",
         11045 => x"5574802e",
         11046 => x"84b13874",
         11047 => x"812e86a1",
         11048 => x"3874ff2e",
         11049 => x"868c3874",
         11050 => x"981b0c88",
         11051 => x"1a088538",
         11052 => x"74881b0c",
         11053 => x"6056b416",
         11054 => x"089c1b08",
         11055 => x"2e81d338",
         11056 => x"981a08fe",
         11057 => x"059c1708",
         11058 => x"fe055858",
         11059 => x"77772785",
         11060 => x"f0388a16",
         11061 => x"22707929",
         11062 => x"b0180805",
         11063 => x"56577480",
         11064 => x"2e85de38",
         11065 => x"78157b89",
         11066 => x"2a595c77",
         11067 => x"802e8398",
         11068 => x"3877195f",
         11069 => x"767f2785",
         11070 => x"38767931",
         11071 => x"5877547b",
         11072 => x"537c5281",
         11073 => x"163351ff",
         11074 => x"9ba13f84",
         11075 => x"ba8c0885",
         11076 => x"a13860b4",
         11077 => x"11087d31",
         11078 => x"56577478",
         11079 => x"27a53884",
         11080 => x"800bb818",
         11081 => x"7672291f",
         11082 => x"57585674",
         11083 => x"70810556",
         11084 => x"33777081",
         11085 => x"055934ff",
         11086 => x"165675ef",
         11087 => x"38605975",
         11088 => x"831a3477",
         11089 => x"892b597a",
         11090 => x"79317e08",
         11091 => x"1a7f0c79",
         11092 => x"1e941c08",
         11093 => x"1b707194",
         11094 => x"1f0c8c1e",
         11095 => x"085a5a57",
         11096 => x"5e5b7575",
         11097 => x"27833874",
         11098 => x"56758c1b",
         11099 => x"0c7afe85",
         11100 => x"38901a33",
         11101 => x"587780c0",
         11102 => x"075b7a90",
         11103 => x"1b348056",
         11104 => x"7584ba8c",
         11105 => x"0c923d0d",
         11106 => x"047484ba",
         11107 => x"8c0c923d",
         11108 => x"0d048316",
         11109 => x"33557482",
         11110 => x"c8386056",
         11111 => x"fea23960",
         11112 => x"9c1b0859",
         11113 => x"567683ff",
         11114 => x"06848071",
         11115 => x"315a5c7a",
         11116 => x"79278338",
         11117 => x"7a597757",
         11118 => x"b4160878",
         11119 => x"2eb63880",
         11120 => x"0b831733",
         11121 => x"715e415f",
         11122 => x"7f7f2e09",
         11123 => x"810680d5",
         11124 => x"38815477",
         11125 => x"53b81652",
         11126 => x"81163351",
         11127 => x"ff98cd3f",
         11128 => x"84ba8c08",
         11129 => x"802e8538",
         11130 => x"ff57815c",
         11131 => x"76b4170c",
         11132 => x"7b83bf38",
         11133 => x"60941b08",
         11134 => x"83ff0611",
         11135 => x"7a58b805",
         11136 => x"7e595658",
         11137 => x"78802e95",
         11138 => x"38767081",
         11139 => x"05583375",
         11140 => x"70810557",
         11141 => x"34ff1656",
         11142 => x"75ef3860",
         11143 => x"58810b83",
         11144 => x"1934fea3",
         11145 => x"398154b4",
         11146 => x"160853b8",
         11147 => x"16705381",
         11148 => x"17335240",
         11149 => x"ff98f43f",
         11150 => x"815c84ba",
         11151 => x"8c087f2e",
         11152 => x"098106ff",
         11153 => x"ab3884ba",
         11154 => x"8c088317",
         11155 => x"34b41608",
         11156 => x"a8170831",
         11157 => x"84ba8c08",
         11158 => x"5d5574a0",
         11159 => x"170827fe",
         11160 => x"f0388216",
         11161 => x"33557482",
         11162 => x"2e098106",
         11163 => x"fee33881",
         11164 => x"54b41608",
         11165 => x"a0170805",
         11166 => x"537f5281",
         11167 => x"163351ff",
         11168 => x"98a93f7e",
         11169 => x"5cfeca39",
         11170 => x"941a0857",
         11171 => x"8c1a0877",
         11172 => x"26933883",
         11173 => x"1633407f",
         11174 => x"81b93860",
         11175 => x"7cb4120c",
         11176 => x"941b0858",
         11177 => x"567b7c9c",
         11178 => x"1c0c58fd",
         11179 => x"f839981a",
         11180 => x"08527951",
         11181 => x"ffabe73f",
         11182 => x"84ba8c08",
         11183 => x"5584ba8c",
         11184 => x"08fbd838",
         11185 => x"901a3358",
         11186 => x"fdab3976",
         11187 => x"527951ff",
         11188 => x"abcc3f84",
         11189 => x"ba8c0855",
         11190 => x"84ba8c08",
         11191 => x"fbbd38e4",
         11192 => x"398154b4",
         11193 => x"160853b8",
         11194 => x"16705381",
         11195 => x"17335257",
         11196 => x"ff97b83f",
         11197 => x"84ba8c08",
         11198 => x"81b83884",
         11199 => x"ba8c0883",
         11200 => x"1734b416",
         11201 => x"08a81708",
         11202 => x"315877a0",
         11203 => x"170827fd",
         11204 => x"89388216",
         11205 => x"335c7b82",
         11206 => x"2e098106",
         11207 => x"fcfc3881",
         11208 => x"54b41608",
         11209 => x"a0170805",
         11210 => x"53765281",
         11211 => x"163351ff",
         11212 => x"96f93f60",
         11213 => x"56fb8939",
         11214 => x"81163351",
         11215 => x"ff959b3f",
         11216 => x"84ba8c08",
         11217 => x"81065574",
         11218 => x"f9f23874",
         11219 => x"7a085657",
         11220 => x"f9ec3981",
         11221 => x"54b41608",
         11222 => x"53b81670",
         11223 => x"53811733",
         11224 => x"5257ff96",
         11225 => x"c63f84ba",
         11226 => x"8c0880c6",
         11227 => x"3884ba8c",
         11228 => x"08831734",
         11229 => x"b41608a8",
         11230 => x"17083155",
         11231 => x"74a01708",
         11232 => x"27fe9838",
         11233 => x"82163358",
         11234 => x"77822e09",
         11235 => x"8106fe8b",
         11236 => x"388154b4",
         11237 => x"1608a017",
         11238 => x"08055376",
         11239 => x"52811633",
         11240 => x"51ff9687",
         11241 => x"3f607cb4",
         11242 => x"120c941b",
         11243 => x"085856fd",
         11244 => x"f439810b",
         11245 => x"911b3481",
         11246 => x"0b84ba8c",
         11247 => x"0c923d0d",
         11248 => x"04820b91",
         11249 => x"1b34820b",
         11250 => x"84ba8c0c",
         11251 => x"923d0d04",
         11252 => x"f53d0d7d",
         11253 => x"58895a77",
         11254 => x"802e9f38",
         11255 => x"77085675",
         11256 => x"802e9738",
         11257 => x"75335574",
         11258 => x"802e8f38",
         11259 => x"86162284",
         11260 => x"19225859",
         11261 => x"78772e83",
         11262 => x"b5388055",
         11263 => x"745c7956",
         11264 => x"7981d838",
         11265 => x"90183370",
         11266 => x"862a8106",
         11267 => x"5c577a80",
         11268 => x"2e81c838",
         11269 => x"7ba01908",
         11270 => x"5a57b417",
         11271 => x"08792eac",
         11272 => x"38831733",
         11273 => x"5b7a81bc",
         11274 => x"38815478",
         11275 => x"53b81752",
         11276 => x"81173351",
         11277 => x"ff93f53f",
         11278 => x"84ba8c08",
         11279 => x"802e8538",
         11280 => x"ff598156",
         11281 => x"78b4180c",
         11282 => x"75819038",
         11283 => x"a418088b",
         11284 => x"1133a007",
         11285 => x"5a57788b",
         11286 => x"18347708",
         11287 => x"88190870",
         11288 => x"83ffff06",
         11289 => x"5d5a567a",
         11290 => x"9a18347a",
         11291 => x"882a5a79",
         11292 => x"9b18349c",
         11293 => x"17763396",
         11294 => x"195c565b",
         11295 => x"74832e81",
         11296 => x"c1388c18",
         11297 => x"0855747b",
         11298 => x"3474882a",
         11299 => x"5b7a9d18",
         11300 => x"3474902a",
         11301 => x"56759e18",
         11302 => x"3474982a",
         11303 => x"59789f18",
         11304 => x"34807a34",
         11305 => x"800b9718",
         11306 => x"34a10b98",
         11307 => x"183480cc",
         11308 => x"0b991834",
         11309 => x"800b9218",
         11310 => x"34800b93",
         11311 => x"18347b5b",
         11312 => x"810b831c",
         11313 => x"347b51ff",
         11314 => x"96943f84",
         11315 => x"ba8c0890",
         11316 => x"193381bf",
         11317 => x"065b5679",
         11318 => x"90193475",
         11319 => x"84ba8c0c",
         11320 => x"8d3d0d04",
         11321 => x"8154b417",
         11322 => x"0853b817",
         11323 => x"70538118",
         11324 => x"33525bff",
         11325 => x"93b53f81",
         11326 => x"5684ba8c",
         11327 => x"08fec938",
         11328 => x"84ba8c08",
         11329 => x"831834b4",
         11330 => x"1708a818",
         11331 => x"083184ba",
         11332 => x"8c085755",
         11333 => x"74a01808",
         11334 => x"27fe8e38",
         11335 => x"82173355",
         11336 => x"74822e09",
         11337 => x"8106fe81",
         11338 => x"388154b4",
         11339 => x"1708a018",
         11340 => x"0805537a",
         11341 => x"52811733",
         11342 => x"51ff92ef",
         11343 => x"3f7956fd",
         11344 => x"e8397890",
         11345 => x"2a557494",
         11346 => x"18347488",
         11347 => x"2a567595",
         11348 => x"18348c18",
         11349 => x"0855747b",
         11350 => x"3474882a",
         11351 => x"5b7a9d18",
         11352 => x"3474902a",
         11353 => x"56759e18",
         11354 => x"3474982a",
         11355 => x"59789f18",
         11356 => x"34807a34",
         11357 => x"800b9718",
         11358 => x"34a10b98",
         11359 => x"183480cc",
         11360 => x"0b991834",
         11361 => x"800b9218",
         11362 => x"34800b93",
         11363 => x"18347b5b",
         11364 => x"810b831c",
         11365 => x"347b51ff",
         11366 => x"94c43f84",
         11367 => x"ba8c0890",
         11368 => x"193381bf",
         11369 => x"065b5679",
         11370 => x"901934fe",
         11371 => x"ae398116",
         11372 => x"3351ff90",
         11373 => x"a53f84ba",
         11374 => x"8c088106",
         11375 => x"5574fcba",
         11376 => x"38747808",
         11377 => x"565afcb4",
         11378 => x"39f93d0d",
         11379 => x"79705255",
         11380 => x"fbfe3f84",
         11381 => x"ba8c0854",
         11382 => x"84ba8c08",
         11383 => x"b1388956",
         11384 => x"74802e9e",
         11385 => x"38740853",
         11386 => x"72802e96",
         11387 => x"38723352",
         11388 => x"71802e8e",
         11389 => x"38861322",
         11390 => x"84162258",
         11391 => x"5271772e",
         11392 => x"96388052",
         11393 => x"71587554",
         11394 => x"75843875",
         11395 => x"750c7384",
         11396 => x"ba8c0c89",
         11397 => x"3d0d0481",
         11398 => x"133351ff",
         11399 => x"8fbc3f84",
         11400 => x"ba8c0881",
         11401 => x"065372da",
         11402 => x"38737508",
         11403 => x"5356d539",
         11404 => x"f63d0dff",
         11405 => x"7d705b57",
         11406 => x"5b75802e",
         11407 => x"b2387570",
         11408 => x"81055733",
         11409 => x"709f2652",
         11410 => x"5271ba2e",
         11411 => x"ac3870ee",
         11412 => x"3871ba2e",
         11413 => x"a43884d1",
         11414 => x"e8335180",
         11415 => x"71249038",
         11416 => x"7084d1e8",
         11417 => x"34800b84",
         11418 => x"ba8c0c8c",
         11419 => x"3d0d048b",
         11420 => x"0b84ba8c",
         11421 => x"0c8c3d0d",
         11422 => x"047833d0",
         11423 => x"117081ff",
         11424 => x"06535353",
         11425 => x"70892691",
         11426 => x"38821973",
         11427 => x"81ff06d0",
         11428 => x"05595473",
         11429 => x"762e80f5",
         11430 => x"38800b83",
         11431 => x"e5fc5b58",
         11432 => x"79087956",
         11433 => x"57767081",
         11434 => x"05583375",
         11435 => x"70810557",
         11436 => x"33ff9f12",
         11437 => x"53545270",
         11438 => x"99268938",
         11439 => x"e0127081",
         11440 => x"ff065354",
         11441 => x"ff9f1351",
         11442 => x"70992689",
         11443 => x"38e01370",
         11444 => x"81ff0654",
         11445 => x"54713070",
         11446 => x"9f2a5551",
         11447 => x"71732e09",
         11448 => x"81068538",
         11449 => x"73ffbe38",
         11450 => x"74763270",
         11451 => x"30707207",
         11452 => x"9f2a7607",
         11453 => x"59525276",
         11454 => x"802e9238",
         11455 => x"8118841b",
         11456 => x"5b588378",
         11457 => x"25ff9938",
         11458 => x"7a51fecf",
         11459 => x"39778324",
         11460 => x"f7387776",
         11461 => x"5e51fec3",
         11462 => x"39ea3d0d",
         11463 => x"8053983d",
         11464 => x"cc055299",
         11465 => x"3d51d194",
         11466 => x"3f84ba8c",
         11467 => x"085584ba",
         11468 => x"8c08802e",
         11469 => x"8a387484",
         11470 => x"ba8c0c98",
         11471 => x"3d0d047a",
         11472 => x"5c685298",
         11473 => x"3dd00551",
         11474 => x"c5943f84",
         11475 => x"ba8c0855",
         11476 => x"84ba8c08",
         11477 => x"80c63802",
         11478 => x"80d70533",
         11479 => x"70982b58",
         11480 => x"5a807724",
         11481 => x"80e23802",
         11482 => x"b2053370",
         11483 => x"842a8106",
         11484 => x"57597580",
         11485 => x"2eb2387a",
         11486 => x"639b1133",
         11487 => x"9a123371",
         11488 => x"882b0773",
         11489 => x"335e5a5b",
         11490 => x"57587983",
         11491 => x"2ea43876",
         11492 => x"98190c74",
         11493 => x"84ba8c0c",
         11494 => x"983d0d04",
         11495 => x"84ba8c08",
         11496 => x"842e0981",
         11497 => x"06ff8f38",
         11498 => x"850b84ba",
         11499 => x"8c0c983d",
         11500 => x"0d049516",
         11501 => x"33941733",
         11502 => x"71982b71",
         11503 => x"902b0779",
         11504 => x"07981b0c",
         11505 => x"5b54cc39",
         11506 => x"7a7e9812",
         11507 => x"0c587484",
         11508 => x"ba8c0c98",
         11509 => x"3d0d04ff",
         11510 => x"9e3d0d80",
         11511 => x"e63d0880",
         11512 => x"e63d085d",
         11513 => x"40807c34",
         11514 => x"805380e4",
         11515 => x"3dfdb405",
         11516 => x"5280e53d",
         11517 => x"51cfc53f",
         11518 => x"84ba8c08",
         11519 => x"5984ba8c",
         11520 => x"0883c838",
         11521 => x"6080d93d",
         11522 => x"0c7f6198",
         11523 => x"110880dd",
         11524 => x"3d0c5880",
         11525 => x"db3d085b",
         11526 => x"5879802e",
         11527 => x"82cc3880",
         11528 => x"d83d983d",
         11529 => x"405ba052",
         11530 => x"7a51ffa4",
         11531 => x"aa3f84ba",
         11532 => x"8c085984",
         11533 => x"ba8c0883",
         11534 => x"92386080",
         11535 => x"df3d0858",
         11536 => x"56b41608",
         11537 => x"772eb138",
         11538 => x"84ba8c08",
         11539 => x"8317335f",
         11540 => x"5d7d83c7",
         11541 => x"38815476",
         11542 => x"53b81652",
         11543 => x"81163351",
         11544 => x"ff8bc93f",
         11545 => x"84ba8c08",
         11546 => x"802e8538",
         11547 => x"ff578159",
         11548 => x"76b4170c",
         11549 => x"7882d438",
         11550 => x"80df3d08",
         11551 => x"9b11339a",
         11552 => x"12337188",
         11553 => x"2b076370",
         11554 => x"335d4059",
         11555 => x"56567883",
         11556 => x"2e82da38",
         11557 => x"7680db3d",
         11558 => x"0c80527a",
         11559 => x"51ffa3b7",
         11560 => x"3f84ba8c",
         11561 => x"085984ba",
         11562 => x"8c08829f",
         11563 => x"3880527a",
         11564 => x"51ffa8f5",
         11565 => x"3f84ba8c",
         11566 => x"085984ba",
         11567 => x"8c08bb38",
         11568 => x"80df3d08",
         11569 => x"9b11339a",
         11570 => x"12337188",
         11571 => x"2b076370",
         11572 => x"33425859",
         11573 => x"5e567d83",
         11574 => x"2e81fd38",
         11575 => x"767a2ea4",
         11576 => x"3884ba8c",
         11577 => x"08527a51",
         11578 => x"ffa4e23f",
         11579 => x"84ba8c08",
         11580 => x"5984ba8c",
         11581 => x"08802eff",
         11582 => x"b4387884",
         11583 => x"2e83d838",
         11584 => x"7881c838",
         11585 => x"80e43dfd",
         11586 => x"b805527a",
         11587 => x"51ffbd89",
         11588 => x"3f787f82",
         11589 => x"05335b57",
         11590 => x"79802e90",
         11591 => x"38821f56",
         11592 => x"81178117",
         11593 => x"70335f57",
         11594 => x"577cf538",
         11595 => x"81175675",
         11596 => x"78268195",
         11597 => x"3876802e",
         11598 => x"9c387e17",
         11599 => x"820556ff",
         11600 => x"1880e63d",
         11601 => x"0811ff19",
         11602 => x"ff195959",
         11603 => x"56587533",
         11604 => x"753476eb",
         11605 => x"38ff1880",
         11606 => x"e63d0811",
         11607 => x"5f58af7e",
         11608 => x"3480da3d",
         11609 => x"085a79fd",
         11610 => x"bd387760",
         11611 => x"2e828a38",
         11612 => x"800b84d1",
         11613 => x"e8337010",
         11614 => x"1083e5fc",
         11615 => x"05700870",
         11616 => x"33435959",
         11617 => x"5e5a7e7a",
         11618 => x"2e8d3881",
         11619 => x"1a701770",
         11620 => x"33575f5a",
         11621 => x"74f53882",
         11622 => x"1a5b7a78",
         11623 => x"26ab3880",
         11624 => x"57767a27",
         11625 => x"94387616",
         11626 => x"5f7e337c",
         11627 => x"7081055e",
         11628 => x"34811757",
         11629 => x"797726ee",
         11630 => x"38ba7c70",
         11631 => x"81055e34",
         11632 => x"76ff2e09",
         11633 => x"810681df",
         11634 => x"38915980",
         11635 => x"7c347884",
         11636 => x"ba8c0c80",
         11637 => x"e43d0d04",
         11638 => x"95163394",
         11639 => x"17337198",
         11640 => x"2b71902b",
         11641 => x"07790759",
         11642 => x"565efdf0",
         11643 => x"39951633",
         11644 => x"94173371",
         11645 => x"982b7190",
         11646 => x"2b077907",
         11647 => x"80dd3d0c",
         11648 => x"5a5d8052",
         11649 => x"7a51ffa0",
         11650 => x"ce3f84ba",
         11651 => x"8c085984",
         11652 => x"ba8c0880",
         11653 => x"2efd9638",
         11654 => x"ffb13981",
         11655 => x"54b41608",
         11656 => x"53b81670",
         11657 => x"53811733",
         11658 => x"525eff88",
         11659 => x"fe3f8159",
         11660 => x"84ba8c08",
         11661 => x"fcbe3884",
         11662 => x"ba8c0883",
         11663 => x"1734b416",
         11664 => x"08a81708",
         11665 => x"3184ba8c",
         11666 => x"085a5574",
         11667 => x"a0170827",
         11668 => x"fc833882",
         11669 => x"16335574",
         11670 => x"822e0981",
         11671 => x"06fbf638",
         11672 => x"8154b416",
         11673 => x"08a01708",
         11674 => x"05537d52",
         11675 => x"81163351",
         11676 => x"ff88b83f",
         11677 => x"7c59fbdd",
         11678 => x"39ff1880",
         11679 => x"e63d0811",
         11680 => x"5c58af7b",
         11681 => x"34800b84",
         11682 => x"d1e83370",
         11683 => x"101083e5",
         11684 => x"fc057008",
         11685 => x"70334359",
         11686 => x"595e5a7e",
         11687 => x"7a2e0981",
         11688 => x"06fde838",
         11689 => x"fdf13980",
         11690 => x"e53d0818",
         11691 => x"8119595a",
         11692 => x"79337c70",
         11693 => x"81055e34",
         11694 => x"776027fe",
         11695 => x"8e3880e5",
         11696 => x"3d081881",
         11697 => x"19595a79",
         11698 => x"337c7081",
         11699 => x"055e347f",
         11700 => x"7826d438",
         11701 => x"fdf53982",
         11702 => x"59807c34",
         11703 => x"7884ba8c",
         11704 => x"0c80e43d",
         11705 => x"0d04f73d",
         11706 => x"0d7b7d58",
         11707 => x"55895674",
         11708 => x"802e9f38",
         11709 => x"74085473",
         11710 => x"802e9738",
         11711 => x"73335372",
         11712 => x"802e8f38",
         11713 => x"86142284",
         11714 => x"16225959",
         11715 => x"78782e83",
         11716 => x"a0388053",
         11717 => x"725a7553",
         11718 => x"7581c238",
         11719 => x"91153353",
         11720 => x"7281ba38",
         11721 => x"8c150856",
         11722 => x"76762681",
         11723 => x"b9389415",
         11724 => x"08548058",
         11725 => x"76782e81",
         11726 => x"cc38798a",
         11727 => x"11227089",
         11728 => x"2b525a56",
         11729 => x"73782e81",
         11730 => x"f7387552",
         11731 => x"ff1751fd",
         11732 => x"bad33f84",
         11733 => x"ba8c08ff",
         11734 => x"15775470",
         11735 => x"535553fd",
         11736 => x"bac33f84",
         11737 => x"ba8c0873",
         11738 => x"2681d538",
         11739 => x"75307406",
         11740 => x"7094170c",
         11741 => x"77713198",
         11742 => x"17085658",
         11743 => x"5973802e",
         11744 => x"82983875",
         11745 => x"772781d9",
         11746 => x"38767631",
         11747 => x"94160817",
         11748 => x"94170c90",
         11749 => x"16337081",
         11750 => x"2a810651",
         11751 => x"5a577880",
         11752 => x"2e81fe38",
         11753 => x"73527451",
         11754 => x"ff99f33f",
         11755 => x"84ba8c08",
         11756 => x"5484ba8c",
         11757 => x"08802e81",
         11758 => x"a33873ff",
         11759 => x"2e983881",
         11760 => x"742782b4",
         11761 => x"38795373",
         11762 => x"9c140827",
         11763 => x"82aa3873",
         11764 => x"98160cff",
         11765 => x"ae39810b",
         11766 => x"91163481",
         11767 => x"537284ba",
         11768 => x"8c0c8b3d",
         11769 => x"0d049015",
         11770 => x"3370812a",
         11771 => x"81065558",
         11772 => x"73febb38",
         11773 => x"75941608",
         11774 => x"55578058",
         11775 => x"76782e09",
         11776 => x"8106feb6",
         11777 => x"38779416",
         11778 => x"0c941508",
         11779 => x"54757427",
         11780 => x"9038738c",
         11781 => x"160c9015",
         11782 => x"3380c007",
         11783 => x"57769016",
         11784 => x"347383ff",
         11785 => x"06597880",
         11786 => x"2e8c389c",
         11787 => x"1508782e",
         11788 => x"8538779c",
         11789 => x"160c800b",
         11790 => x"84ba8c0c",
         11791 => x"8b3d0d04",
         11792 => x"800b9416",
         11793 => x"0c881508",
         11794 => x"5473802e",
         11795 => x"80fe3873",
         11796 => x"98160c73",
         11797 => x"802e80c2",
         11798 => x"38fea839",
         11799 => x"84ba8c08",
         11800 => x"57941508",
         11801 => x"1794160c",
         11802 => x"7683ff06",
         11803 => x"5675802e",
         11804 => x"a93879fe",
         11805 => x"159c1208",
         11806 => x"fe055a55",
         11807 => x"56737827",
         11808 => x"80f6388a",
         11809 => x"16227471",
         11810 => x"29b01808",
         11811 => x"0578892a",
         11812 => x"115a5a53",
         11813 => x"78802e80",
         11814 => x"df388c15",
         11815 => x"0856fee9",
         11816 => x"39735274",
         11817 => x"51ff89b7",
         11818 => x"3f84ba8c",
         11819 => x"0854fe8a",
         11820 => x"39811433",
         11821 => x"51ff82a2",
         11822 => x"3f84ba8c",
         11823 => x"08810653",
         11824 => x"72fccf38",
         11825 => x"72750854",
         11826 => x"56fcc939",
         11827 => x"73527451",
         11828 => x"ff97cb3f",
         11829 => x"84ba8c08",
         11830 => x"5484ba8c",
         11831 => x"08812e98",
         11832 => x"3884ba8c",
         11833 => x"08ff2efd",
         11834 => x"ed3884ba",
         11835 => x"8c088816",
         11836 => x"0c739816",
         11837 => x"0cfedc39",
         11838 => x"820b9116",
         11839 => x"34820b84",
         11840 => x"ba8c0c8b",
         11841 => x"3d0d04f6",
         11842 => x"3d0d7c56",
         11843 => x"89547580",
         11844 => x"2ea23880",
         11845 => x"538c3dfc",
         11846 => x"05528d3d",
         11847 => x"840551c5",
         11848 => x"9b3f84ba",
         11849 => x"8c085584",
         11850 => x"ba8c0880",
         11851 => x"2e8f3880",
         11852 => x"760c7454",
         11853 => x"7384ba8c",
         11854 => x"0c8c3d0d",
         11855 => x"047a760c",
         11856 => x"7d527551",
         11857 => x"ffb9973f",
         11858 => x"84ba8c08",
         11859 => x"5584ba8c",
         11860 => x"0880d138",
         11861 => x"ab163370",
         11862 => x"982b5959",
         11863 => x"807824af",
         11864 => x"38861633",
         11865 => x"70842a81",
         11866 => x"065b5479",
         11867 => x"802e80c5",
         11868 => x"389c1608",
         11869 => x"9b11339a",
         11870 => x"12337188",
         11871 => x"2b077d70",
         11872 => x"335d5d5a",
         11873 => x"55577883",
         11874 => x"2eb33877",
         11875 => x"88170c7a",
         11876 => x"58861822",
         11877 => x"84172374",
         11878 => x"527551ff",
         11879 => x"99b93f84",
         11880 => x"ba8c0855",
         11881 => x"74842e8d",
         11882 => x"3874802e",
         11883 => x"ff843880",
         11884 => x"760cfefe",
         11885 => x"39855580",
         11886 => x"760cfef6",
         11887 => x"39951733",
         11888 => x"94183371",
         11889 => x"982b7190",
         11890 => x"2b077a07",
         11891 => x"88190c5a",
         11892 => x"5affbc39",
         11893 => x"fa3d0d78",
         11894 => x"55895474",
         11895 => x"802e9e38",
         11896 => x"74085372",
         11897 => x"802e9638",
         11898 => x"72335271",
         11899 => x"802e8e38",
         11900 => x"86132284",
         11901 => x"16225752",
         11902 => x"71762e94",
         11903 => x"38805271",
         11904 => x"57738438",
         11905 => x"73750c73",
         11906 => x"84ba8c0c",
         11907 => x"883d0d04",
         11908 => x"81133351",
         11909 => x"feffc33f",
         11910 => x"84ba8c08",
         11911 => x"81065271",
         11912 => x"dc387175",
         11913 => x"085354d7",
         11914 => x"39f83d0d",
         11915 => x"7a7c5855",
         11916 => x"89567480",
         11917 => x"2e9f3874",
         11918 => x"08547380",
         11919 => x"2e973873",
         11920 => x"33537280",
         11921 => x"2e8f3886",
         11922 => x"14228416",
         11923 => x"22595372",
         11924 => x"782e8197",
         11925 => x"38805372",
         11926 => x"59755375",
         11927 => x"80c73876",
         11928 => x"802e80f3",
         11929 => x"38755274",
         11930 => x"51ff9dbd",
         11931 => x"3f84ba8c",
         11932 => x"085384ba",
         11933 => x"8c08842e",
         11934 => x"b53884ba",
         11935 => x"8c08a638",
         11936 => x"76527451",
         11937 => x"ffb2923f",
         11938 => x"72527451",
         11939 => x"ff99be3f",
         11940 => x"84ba8c08",
         11941 => x"84327030",
         11942 => x"7072079f",
         11943 => x"2c84ba8c",
         11944 => x"08065557",
         11945 => x"547284ba",
         11946 => x"8c0c8a3d",
         11947 => x"0d047577",
         11948 => x"53755253",
         11949 => x"ffb1e23f",
         11950 => x"72527451",
         11951 => x"ff998e3f",
         11952 => x"84ba8c08",
         11953 => x"84327030",
         11954 => x"7072079f",
         11955 => x"2c84ba8c",
         11956 => x"08065557",
         11957 => x"54cf3975",
         11958 => x"527451ff",
         11959 => x"96f93f84",
         11960 => x"ba8c0884",
         11961 => x"ba8c0c8a",
         11962 => x"3d0d0481",
         11963 => x"143351fe",
         11964 => x"fde83f84",
         11965 => x"ba8c0881",
         11966 => x"065372fe",
         11967 => x"d8387275",
         11968 => x"085456fe",
         11969 => x"d239ed3d",
         11970 => x"0d665780",
         11971 => x"53893d70",
         11972 => x"53973d52",
         11973 => x"56c1a53f",
         11974 => x"84ba8c08",
         11975 => x"5584ba8c",
         11976 => x"08802e8a",
         11977 => x"387484ba",
         11978 => x"8c0c953d",
         11979 => x"0d046552",
         11980 => x"7551ffb5",
         11981 => x"a93f84ba",
         11982 => x"8c085584",
         11983 => x"ba8c08e5",
         11984 => x"380280cb",
         11985 => x"05337098",
         11986 => x"2b555880",
         11987 => x"74249738",
         11988 => x"76802ed1",
         11989 => x"38765275",
         11990 => x"51ffb0bd",
         11991 => x"3f7484ba",
         11992 => x"8c0c953d",
         11993 => x"0d04860b",
         11994 => x"84ba8c0c",
         11995 => x"953d0d04",
         11996 => x"ed3d0d66",
         11997 => x"68565f80",
         11998 => x"53953dec",
         11999 => x"0552963d",
         12000 => x"51c0b93f",
         12001 => x"84ba8c08",
         12002 => x"5a84ba8c",
         12003 => x"089a387f",
         12004 => x"750c7408",
         12005 => x"9c1108fe",
         12006 => x"11941308",
         12007 => x"59575957",
         12008 => x"7575268d",
         12009 => x"38757f0c",
         12010 => x"7984ba8c",
         12011 => x"0c953d0d",
         12012 => x"0484ba8c",
         12013 => x"0877335a",
         12014 => x"5b78812e",
         12015 => x"82933877",
         12016 => x"a8180884",
         12017 => x"ba8c085a",
         12018 => x"5d597780",
         12019 => x"c1387b81",
         12020 => x"1d715c5d",
         12021 => x"56b41708",
         12022 => x"762e82ef",
         12023 => x"38831733",
         12024 => x"785f5d7c",
         12025 => x"818d3881",
         12026 => x"547553b8",
         12027 => x"17528117",
         12028 => x"3351fefc",
         12029 => x"b73f84ba",
         12030 => x"8c08802e",
         12031 => x"8538ff5a",
         12032 => x"815e79b4",
         12033 => x"180c7f7e",
         12034 => x"5b577d80",
         12035 => x"cc387633",
         12036 => x"5e7d822e",
         12037 => x"828d3877",
         12038 => x"17b80583",
         12039 => x"11338212",
         12040 => x"3371902b",
         12041 => x"71882b07",
         12042 => x"81143370",
         12043 => x"7207882b",
         12044 => x"75337180",
         12045 => x"fffffe80",
         12046 => x"06077030",
         12047 => x"70802563",
         12048 => x"05608405",
         12049 => x"83ff0662",
         12050 => x"ff054341",
         12051 => x"43535452",
         12052 => x"5358405e",
         12053 => x"5678fef2",
         12054 => x"387a7f0c",
         12055 => x"7a94180c",
         12056 => x"84173381",
         12057 => x"07587784",
         12058 => x"18347984",
         12059 => x"ba8c0c95",
         12060 => x"3d0d0481",
         12061 => x"54b41708",
         12062 => x"53b81770",
         12063 => x"53811833",
         12064 => x"525dfefc",
         12065 => x"a63f815e",
         12066 => x"84ba8c08",
         12067 => x"fef83884",
         12068 => x"ba8c0883",
         12069 => x"1834b417",
         12070 => x"08a81808",
         12071 => x"3184ba8c",
         12072 => x"085f5574",
         12073 => x"a0180827",
         12074 => x"febd3882",
         12075 => x"17335574",
         12076 => x"822e0981",
         12077 => x"06feb038",
         12078 => x"8154b417",
         12079 => x"08a01808",
         12080 => x"05537c52",
         12081 => x"81173351",
         12082 => x"fefbe03f",
         12083 => x"775efe97",
         12084 => x"39827742",
         12085 => x"923d5956",
         12086 => x"75527751",
         12087 => x"ff81803f",
         12088 => x"84ba8c08",
         12089 => x"ff2e80e8",
         12090 => x"3884ba8c",
         12091 => x"08812e80",
         12092 => x"f73884ba",
         12093 => x"8c083070",
         12094 => x"84ba8c08",
         12095 => x"0780257c",
         12096 => x"05811862",
         12097 => x"5a585c5c",
         12098 => x"9c170876",
         12099 => x"26ca387a",
         12100 => x"7f0c7a94",
         12101 => x"180c8417",
         12102 => x"33810758",
         12103 => x"77841834",
         12104 => x"fec83977",
         12105 => x"17b80581",
         12106 => x"11337133",
         12107 => x"71882b07",
         12108 => x"70307080",
         12109 => x"251f821d",
         12110 => x"83ff06ff",
         12111 => x"1f5f5d5f",
         12112 => x"595f5f55",
         12113 => x"78fd8338",
         12114 => x"fe8f3977",
         12115 => x"5afdbf39",
         12116 => x"8160585a",
         12117 => x"7a7f0c7a",
         12118 => x"94180c84",
         12119 => x"17338107",
         12120 => x"58778418",
         12121 => x"34fe8339",
         12122 => x"8260585a",
         12123 => x"e739f73d",
         12124 => x"0d7b5789",
         12125 => x"5676802e",
         12126 => x"9f387608",
         12127 => x"5574802e",
         12128 => x"97387433",
         12129 => x"5473802e",
         12130 => x"8f388615",
         12131 => x"22841822",
         12132 => x"59597878",
         12133 => x"2e81da38",
         12134 => x"8054735a",
         12135 => x"7580dc38",
         12136 => x"91173356",
         12137 => x"7580d438",
         12138 => x"90173370",
         12139 => x"812a8106",
         12140 => x"55588755",
         12141 => x"73802e80",
         12142 => x"c4389417",
         12143 => x"0854738c",
         12144 => x"180827b7",
         12145 => x"387381d5",
         12146 => x"38881708",
         12147 => x"77085754",
         12148 => x"81742788",
         12149 => x"389c1608",
         12150 => x"7426b338",
         12151 => x"8256800b",
         12152 => x"88180c94",
         12153 => x"17088c18",
         12154 => x"0c7780c0",
         12155 => x"07597890",
         12156 => x"18347580",
         12157 => x"2e853875",
         12158 => x"91183475",
         12159 => x"557484ba",
         12160 => x"8c0c8b3d",
         12161 => x"0d047854",
         12162 => x"78782780",
         12163 => x"ff387352",
         12164 => x"7651fefe",
         12165 => x"ca3f84ba",
         12166 => x"8c085984",
         12167 => x"ba8c0880",
         12168 => x"2e80e938",
         12169 => x"84ba8c08",
         12170 => x"812e82d8",
         12171 => x"3884ba8c",
         12172 => x"08ff2e82",
         12173 => x"e5388053",
         12174 => x"73527551",
         12175 => x"ff85813f",
         12176 => x"84ba8c08",
         12177 => x"82c8389c",
         12178 => x"1608fe11",
         12179 => x"94180857",
         12180 => x"55587474",
         12181 => x"27ffaf38",
         12182 => x"81159417",
         12183 => x"0c841633",
         12184 => x"81075473",
         12185 => x"84173478",
         12186 => x"54777926",
         12187 => x"ffa0389c",
         12188 => x"39811533",
         12189 => x"51fef6e2",
         12190 => x"3f84ba8c",
         12191 => x"08810654",
         12192 => x"73fe9538",
         12193 => x"73770855",
         12194 => x"56fe8f39",
         12195 => x"800b9018",
         12196 => x"33595473",
         12197 => x"56800b88",
         12198 => x"180cfec7",
         12199 => x"39981708",
         12200 => x"527651fe",
         12201 => x"fdb93f84",
         12202 => x"ba8c08ff",
         12203 => x"2e81c238",
         12204 => x"84ba8c08",
         12205 => x"812e81be",
         12206 => x"387581ae",
         12207 => x"38795884",
         12208 => x"ba8c089c",
         12209 => x"19082781",
         12210 => x"a13884ba",
         12211 => x"8c089818",
         12212 => x"08780858",
         12213 => x"5654810b",
         12214 => x"84ba8c08",
         12215 => x"2781a138",
         12216 => x"84ba8c08",
         12217 => x"9c170827",
         12218 => x"81963874",
         12219 => x"802e9738",
         12220 => x"ff537452",
         12221 => x"7551ff83",
         12222 => x"c73f84ba",
         12223 => x"8c085584",
         12224 => x"ba8c0880",
         12225 => x"e3387352",
         12226 => x"7651fefc",
         12227 => x"d23f84ba",
         12228 => x"8c085984",
         12229 => x"ba8c0880",
         12230 => x"2e80cb38",
         12231 => x"84ba8c08",
         12232 => x"812e80dc",
         12233 => x"3884ba8c",
         12234 => x"08ff2e80",
         12235 => x"fe388053",
         12236 => x"73527551",
         12237 => x"ff83893f",
         12238 => x"84ba8c08",
         12239 => x"80e6389c",
         12240 => x"1608fe11",
         12241 => x"94180857",
         12242 => x"55587474",
         12243 => x"27903881",
         12244 => x"1594170c",
         12245 => x"84163381",
         12246 => x"07547384",
         12247 => x"17347854",
         12248 => x"777926ff",
         12249 => x"a1388055",
         12250 => x"74569017",
         12251 => x"3358fcf3",
         12252 => x"398156fe",
         12253 => x"bb39820b",
         12254 => x"90183359",
         12255 => x"56fce439",
         12256 => x"8256e739",
         12257 => x"820b9018",
         12258 => x"335954fe",
         12259 => x"863984ba",
         12260 => x"8c089018",
         12261 => x"335954fd",
         12262 => x"fa39810b",
         12263 => x"90183359",
         12264 => x"54fdf039",
         12265 => x"84ba8c08",
         12266 => x"56c03981",
         12267 => x"56ffbb39",
         12268 => x"db3d0d82",
         12269 => x"53a73dff",
         12270 => x"9c0552a8",
         12271 => x"3d51ffb7",
         12272 => x"fb3f84ba",
         12273 => x"8c085684",
         12274 => x"ba8c0880",
         12275 => x"2e8a3875",
         12276 => x"84ba8c0c",
         12277 => x"a73d0d04",
         12278 => x"7d4ba83d",
         12279 => x"08529b3d",
         12280 => x"705259ff",
         12281 => x"abf83f84",
         12282 => x"ba8c0856",
         12283 => x"84ba8c08",
         12284 => x"de380281",
         12285 => x"93053370",
         12286 => x"852a8106",
         12287 => x"59578656",
         12288 => x"77cd3876",
         12289 => x"982b5b80",
         12290 => x"7b24c438",
         12291 => x"0280ee05",
         12292 => x"33708106",
         12293 => x"5d578756",
         12294 => x"7bffb438",
         12295 => x"7da33d08",
         12296 => x"9b11339a",
         12297 => x"12337188",
         12298 => x"2b077333",
         12299 => x"415e5c57",
         12300 => x"587c832e",
         12301 => x"80d53876",
         12302 => x"842a8106",
         12303 => x"5776802e",
         12304 => x"80ed3887",
         12305 => x"56981808",
         12306 => x"7b2eff83",
         12307 => x"38775f7a",
         12308 => x"4184ba8c",
         12309 => x"08528f3d",
         12310 => x"705255ff",
         12311 => x"8bf93f84",
         12312 => x"ba8c0856",
         12313 => x"84ba8c08",
         12314 => x"fee53884",
         12315 => x"ba8c0852",
         12316 => x"7451ff91",
         12317 => x"b43f84ba",
         12318 => x"8c085684",
         12319 => x"ba8c08a0",
         12320 => x"38870b84",
         12321 => x"ba8c0ca7",
         12322 => x"3d0d0495",
         12323 => x"16339417",
         12324 => x"3371982b",
         12325 => x"71902b07",
         12326 => x"7d075d5d",
         12327 => x"5dff9839",
         12328 => x"84ba8c08",
         12329 => x"842e8838",
         12330 => x"84ba8c08",
         12331 => x"fea13878",
         12332 => x"086fa83d",
         12333 => x"08575d57",
         12334 => x"74ff2e80",
         12335 => x"d3387452",
         12336 => x"7851ff8b",
         12337 => x"923f84ba",
         12338 => x"8c085684",
         12339 => x"ba8c0880",
         12340 => x"2ebe3875",
         12341 => x"30707707",
         12342 => x"8025565a",
         12343 => x"7a802e9a",
         12344 => x"3874802e",
         12345 => x"95387a79",
         12346 => x"08585581",
         12347 => x"7b278938",
         12348 => x"9c17087b",
         12349 => x"2681fd38",
         12350 => x"825675fd",
         12351 => x"d2387d51",
         12352 => x"fef5db3f",
         12353 => x"84ba8c08",
         12354 => x"84ba8c0c",
         12355 => x"a73d0d04",
         12356 => x"b8175d98",
         12357 => x"19085680",
         12358 => x"5ab41708",
         12359 => x"762e82b9",
         12360 => x"38831733",
         12361 => x"7a595574",
         12362 => x"7a2e0981",
         12363 => x"0680dd38",
         12364 => x"81547553",
         12365 => x"b8175281",
         12366 => x"173351fe",
         12367 => x"f1ee3f84",
         12368 => x"ba8c0880",
         12369 => x"2e8538ff",
         12370 => x"56815875",
         12371 => x"b4180c77",
         12372 => x"5677ab38",
         12373 => x"9c190858",
         12374 => x"e5783481",
         12375 => x"0b831834",
         12376 => x"9019087c",
         12377 => x"27feec38",
         12378 => x"80527851",
         12379 => x"ff8bde3f",
         12380 => x"84ba8c08",
         12381 => x"5684ba8c",
         12382 => x"08802eff",
         12383 => x"96387584",
         12384 => x"2e098106",
         12385 => x"fecd3882",
         12386 => x"56fec839",
         12387 => x"8154b417",
         12388 => x"08537c52",
         12389 => x"81173351",
         12390 => x"fef2903f",
         12391 => x"815884ba",
         12392 => x"8c087a2e",
         12393 => x"098106ff",
         12394 => x"a63884ba",
         12395 => x"8c088318",
         12396 => x"34b41708",
         12397 => x"a8180831",
         12398 => x"84ba8c08",
         12399 => x"595574a0",
         12400 => x"180827fe",
         12401 => x"eb388217",
         12402 => x"33557482",
         12403 => x"2e098106",
         12404 => x"fede3881",
         12405 => x"54b41708",
         12406 => x"a0180805",
         12407 => x"537c5281",
         12408 => x"173351fe",
         12409 => x"f1c53f79",
         12410 => x"58fec539",
         12411 => x"79557978",
         12412 => x"2780e138",
         12413 => x"74527851",
         12414 => x"fef6e43f",
         12415 => x"84ba8c08",
         12416 => x"5a84ba8c",
         12417 => x"08802e80",
         12418 => x"cb3884ba",
         12419 => x"8c08812e",
         12420 => x"fde63884",
         12421 => x"ba8c08ff",
         12422 => x"2e80cb38",
         12423 => x"80537452",
         12424 => x"7651fefd",
         12425 => x"9b3f84ba",
         12426 => x"8c08b338",
         12427 => x"9c1708fe",
         12428 => x"11941908",
         12429 => x"585c5875",
         12430 => x"7b27ffb0",
         12431 => x"38811694",
         12432 => x"180c8417",
         12433 => x"3381075c",
         12434 => x"7b841834",
         12435 => x"7955777a",
         12436 => x"26ffa138",
         12437 => x"8056fda2",
         12438 => x"397956fd",
         12439 => x"f73984ba",
         12440 => x"8c0856fd",
         12441 => x"95398156",
         12442 => x"fd9039e3",
         12443 => x"3d0d8253",
         12444 => x"9f3dffbc",
         12445 => x"0552a03d",
         12446 => x"51ffb2c0",
         12447 => x"3f84ba8c",
         12448 => x"085684ba",
         12449 => x"8c08802e",
         12450 => x"8a387584",
         12451 => x"ba8c0c9f",
         12452 => x"3d0d047d",
         12453 => x"436f5293",
         12454 => x"3d70525a",
         12455 => x"ffa6bf3f",
         12456 => x"84ba8c08",
         12457 => x"5684ba8c",
         12458 => x"088b3888",
         12459 => x"0b84ba8c",
         12460 => x"0c9f3d0d",
         12461 => x"0484ba8c",
         12462 => x"08842e09",
         12463 => x"8106cb38",
         12464 => x"0280f305",
         12465 => x"3370852a",
         12466 => x"81065658",
         12467 => x"865674ff",
         12468 => x"b9387d5f",
         12469 => x"74528f3d",
         12470 => x"70525dff",
         12471 => x"83c03f84",
         12472 => x"ba8c0875",
         12473 => x"575c84ba",
         12474 => x"8c088338",
         12475 => x"875684ba",
         12476 => x"8c08812e",
         12477 => x"80f93884",
         12478 => x"ba8c08ff",
         12479 => x"2e81cb38",
         12480 => x"7581c938",
         12481 => x"7d84ba8c",
         12482 => x"08831233",
         12483 => x"5d5a577a",
         12484 => x"80e238fe",
         12485 => x"199c1808",
         12486 => x"fe055a56",
         12487 => x"805b7579",
         12488 => x"278d388a",
         12489 => x"17227671",
         12490 => x"29b01908",
         12491 => x"055c587a",
         12492 => x"b4180cb8",
         12493 => x"17598480",
         12494 => x"79575580",
         12495 => x"76708105",
         12496 => x"5834ff15",
         12497 => x"5574f438",
         12498 => x"74588a17",
         12499 => x"22557775",
         12500 => x"2781f938",
         12501 => x"8154771b",
         12502 => x"53785281",
         12503 => x"173351fe",
         12504 => x"eec93f84",
         12505 => x"ba8c0881",
         12506 => x"df388118",
         12507 => x"58dc3982",
         12508 => x"56ff8439",
         12509 => x"8154b417",
         12510 => x"0853b817",
         12511 => x"70538118",
         12512 => x"335258fe",
         12513 => x"eea53f81",
         12514 => x"5684ba8c",
         12515 => x"08be3884",
         12516 => x"ba8c0883",
         12517 => x"1834b417",
         12518 => x"08a81808",
         12519 => x"315574a0",
         12520 => x"180827fe",
         12521 => x"ee388217",
         12522 => x"335b7a82",
         12523 => x"2e098106",
         12524 => x"fee13875",
         12525 => x"54b41708",
         12526 => x"a0180805",
         12527 => x"53775281",
         12528 => x"173351fe",
         12529 => x"ede53ffe",
         12530 => x"ca398156",
         12531 => x"7b7d0858",
         12532 => x"55817c27",
         12533 => x"fdb4387b",
         12534 => x"9c180827",
         12535 => x"fdac3874",
         12536 => x"527c51fe",
         12537 => x"f2f93f84",
         12538 => x"ba8c085a",
         12539 => x"84ba8c08",
         12540 => x"802efd96",
         12541 => x"3884ba8c",
         12542 => x"08812efd",
         12543 => x"8d3884ba",
         12544 => x"8c08ff2e",
         12545 => x"fd843880",
         12546 => x"53745276",
         12547 => x"51fef9b0",
         12548 => x"3f84ba8c",
         12549 => x"08fcf338",
         12550 => x"9c1708fe",
         12551 => x"11941908",
         12552 => x"5a5c5977",
         12553 => x"7b279038",
         12554 => x"81189418",
         12555 => x"0c841733",
         12556 => x"81075c7b",
         12557 => x"84183479",
         12558 => x"55787a26",
         12559 => x"ffa13875",
         12560 => x"84ba8c0c",
         12561 => x"9f3d0d04",
         12562 => x"8a172255",
         12563 => x"7483ffff",
         12564 => x"06578156",
         12565 => x"76782e09",
         12566 => x"8106fef0",
         12567 => x"388b0bb8",
         12568 => x"1f5656a0",
         12569 => x"75708105",
         12570 => x"5734ff16",
         12571 => x"5675f438",
         12572 => x"7d57ae0b",
         12573 => x"b818347d",
         12574 => x"58900b80",
         12575 => x"c319347d",
         12576 => x"597580ce",
         12577 => x"1a347580",
         12578 => x"cf1a34a1",
         12579 => x"0b80d01a",
         12580 => x"3480cc0b",
         12581 => x"80d11a34",
         12582 => x"7d7c83ff",
         12583 => x"ff065956",
         12584 => x"7780d217",
         12585 => x"3477882a",
         12586 => x"5b7a80d3",
         12587 => x"17347533",
         12588 => x"5574832e",
         12589 => x"81cc387d",
         12590 => x"59a00b80",
         12591 => x"d81ab81b",
         12592 => x"57585674",
         12593 => x"70810556",
         12594 => x"33777081",
         12595 => x"055934ff",
         12596 => x"165675ef",
         12597 => x"387d56ae",
         12598 => x"0b80d917",
         12599 => x"34647e71",
         12600 => x"83ffff06",
         12601 => x"5b575778",
         12602 => x"80f21734",
         12603 => x"78882a5b",
         12604 => x"7a80f317",
         12605 => x"34753355",
         12606 => x"74832e80",
         12607 => x"f0387d5b",
         12608 => x"810b831c",
         12609 => x"347951ff",
         12610 => x"92963f84",
         12611 => x"ba8c0856",
         12612 => x"84ba8c08",
         12613 => x"fdb63869",
         12614 => x"5684ba8c",
         12615 => x"08961734",
         12616 => x"84ba8c08",
         12617 => x"971734a1",
         12618 => x"0b981734",
         12619 => x"80cc0b99",
         12620 => x"17347d6a",
         12621 => x"585d779a",
         12622 => x"18347788",
         12623 => x"2a59789b",
         12624 => x"18347c33",
         12625 => x"5a79832e",
         12626 => x"80d93869",
         12627 => x"55900b8b",
         12628 => x"16347d57",
         12629 => x"810b8318",
         12630 => x"347d51fe",
         12631 => x"ed803f84",
         12632 => x"ba8c0856",
         12633 => x"7584ba8c",
         12634 => x"0c9f3d0d",
         12635 => x"0476902a",
         12636 => x"557480ec",
         12637 => x"17347488",
         12638 => x"2a577680",
         12639 => x"ed1734fe",
         12640 => x"fd397b90",
         12641 => x"2a5b7a80",
         12642 => x"cc17347a",
         12643 => x"882a5574",
         12644 => x"80cd1734",
         12645 => x"7d59a00b",
         12646 => x"80d81ab8",
         12647 => x"1b575856",
         12648 => x"fea1397b",
         12649 => x"902a5877",
         12650 => x"94183477",
         12651 => x"882a5c7b",
         12652 => x"95183469",
         12653 => x"55900b8b",
         12654 => x"16347d57",
         12655 => x"810b8318",
         12656 => x"347d51fe",
         12657 => x"ec983f84",
         12658 => x"ba8c0856",
         12659 => x"ff9639d1",
         12660 => x"3d0db33d",
         12661 => x"b43d0870",
         12662 => x"595b5f79",
         12663 => x"802e9b38",
         12664 => x"79708105",
         12665 => x"5b33709f",
         12666 => x"26565675",
         12667 => x"ba2e81b8",
         12668 => x"3874ed38",
         12669 => x"75ba2e81",
         12670 => x"af388253",
         12671 => x"b13dfefc",
         12672 => x"0552b23d",
         12673 => x"51ffabb4",
         12674 => x"3f84ba8c",
         12675 => x"085684ba",
         12676 => x"8c08802e",
         12677 => x"8a387584",
         12678 => x"ba8c0cb1",
         12679 => x"3d0d047f",
         12680 => x"a63d0cb2",
         12681 => x"3d0852a5",
         12682 => x"3d705259",
         12683 => x"ff9faf3f",
         12684 => x"84ba8c08",
         12685 => x"5684ba8c",
         12686 => x"08dc3802",
         12687 => x"81bb0533",
         12688 => x"81a0065d",
         12689 => x"86567cce",
         12690 => x"38a00b92",
         12691 => x"3dae3d08",
         12692 => x"58585575",
         12693 => x"70810557",
         12694 => x"33777081",
         12695 => x"055934ff",
         12696 => x"155574ef",
         12697 => x"38993d58",
         12698 => x"b0787a58",
         12699 => x"58557570",
         12700 => x"81055733",
         12701 => x"77708105",
         12702 => x"5934ff15",
         12703 => x"5574ef38",
         12704 => x"b33d0852",
         12705 => x"7751ff9e",
         12706 => x"d53f84ba",
         12707 => x"8c085684",
         12708 => x"ba8c0885",
         12709 => x"d8386aa8",
         12710 => x"3d082e81",
         12711 => x"cb38880b",
         12712 => x"84ba8c0c",
         12713 => x"b13d0d04",
         12714 => x"7633d011",
         12715 => x"7081ff06",
         12716 => x"57575874",
         12717 => x"89269138",
         12718 => x"82177881",
         12719 => x"ff06d005",
         12720 => x"5d59787a",
         12721 => x"2e80fa38",
         12722 => x"807f0883",
         12723 => x"e5fc7008",
         12724 => x"725d5e5f",
         12725 => x"5f5c7a70",
         12726 => x"81055c33",
         12727 => x"79708105",
         12728 => x"5b33ff9f",
         12729 => x"125a5856",
         12730 => x"77992689",
         12731 => x"38e01670",
         12732 => x"81ff0657",
         12733 => x"55ff9f17",
         12734 => x"58779926",
         12735 => x"8938e017",
         12736 => x"7081ff06",
         12737 => x"58557530",
         12738 => x"709f2a59",
         12739 => x"5575772e",
         12740 => x"09810685",
         12741 => x"3877ffbe",
         12742 => x"38787a32",
         12743 => x"70307072",
         12744 => x"079f2a7a",
         12745 => x"075d5855",
         12746 => x"7a802e95",
         12747 => x"38811c84",
         12748 => x"1e5e5c7b",
         12749 => x"8324fdc2",
         12750 => x"387c087e",
         12751 => x"5a5bff96",
         12752 => x"397b8324",
         12753 => x"fdb43879",
         12754 => x"7f0c8253",
         12755 => x"b13dfefc",
         12756 => x"0552b23d",
         12757 => x"51ffa8e4",
         12758 => x"3f84ba8c",
         12759 => x"085684ba",
         12760 => x"8c08fdb2",
         12761 => x"38fdb839",
         12762 => x"6caa3d08",
         12763 => x"2e098106",
         12764 => x"feac3877",
         12765 => x"51ff8da8",
         12766 => x"3f84ba8c",
         12767 => x"085684ba",
         12768 => x"8c08fd92",
         12769 => x"386f5893",
         12770 => x"0b8d1902",
         12771 => x"880580cd",
         12772 => x"0558565a",
         12773 => x"75708105",
         12774 => x"57337570",
         12775 => x"81055734",
         12776 => x"ff1a5a79",
         12777 => x"ef380280",
         12778 => x"cb05338b",
         12779 => x"19348b18",
         12780 => x"3370842a",
         12781 => x"81064056",
         12782 => x"7e893875",
         12783 => x"a0075776",
         12784 => x"8b19347f",
         12785 => x"5d810b83",
         12786 => x"1e348b18",
         12787 => x"3370842a",
         12788 => x"8106575c",
         12789 => x"75802e81",
         12790 => x"c538a73d",
         12791 => x"086b2e81",
         12792 => x"bd387f9b",
         12793 => x"19339a1a",
         12794 => x"3371882b",
         12795 => x"07723341",
         12796 => x"585c577d",
         12797 => x"832e82e0",
         12798 => x"38fe169c",
         12799 => x"1808fe05",
         12800 => x"5e56757d",
         12801 => x"2782c738",
         12802 => x"8a172276",
         12803 => x"7129b019",
         12804 => x"0805575e",
         12805 => x"75802e82",
         12806 => x"b538757a",
         12807 => x"5d58b417",
         12808 => x"08762eaa",
         12809 => x"38831733",
         12810 => x"5f7e83bc",
         12811 => x"38815475",
         12812 => x"53b81752",
         12813 => x"81173351",
         12814 => x"fee3f13f",
         12815 => x"84ba8c08",
         12816 => x"802e8538",
         12817 => x"ff58815c",
         12818 => x"77b4180c",
         12819 => x"7f577b80",
         12820 => x"d8185656",
         12821 => x"7bfbbf38",
         12822 => x"8115335a",
         12823 => x"79ae2e09",
         12824 => x"8106bb38",
         12825 => x"6a7083ff",
         12826 => x"ff065d56",
         12827 => x"7b80f218",
         12828 => x"347b882a",
         12829 => x"587780f3",
         12830 => x"18347633",
         12831 => x"5b7a832e",
         12832 => x"09810693",
         12833 => x"3875902a",
         12834 => x"5e7d80ec",
         12835 => x"18347d88",
         12836 => x"2a567580",
         12837 => x"ed18347f",
         12838 => x"57810b83",
         12839 => x"18347808",
         12840 => x"aa3d08b2",
         12841 => x"3d08575c",
         12842 => x"5674ff2e",
         12843 => x"95387452",
         12844 => x"7851fefb",
         12845 => x"a23f84ba",
         12846 => x"8c085584",
         12847 => x"ba8c0880",
         12848 => x"f538b816",
         12849 => x"5c981908",
         12850 => x"57805ab4",
         12851 => x"1608772e",
         12852 => x"b4388316",
         12853 => x"337a595f",
         12854 => x"7e7a2e09",
         12855 => x"810681a8",
         12856 => x"38815476",
         12857 => x"53b81652",
         12858 => x"81163351",
         12859 => x"fee2bd3f",
         12860 => x"84ba8c08",
         12861 => x"802e8538",
         12862 => x"ff578158",
         12863 => x"76b4170c",
         12864 => x"775577aa",
         12865 => x"389c1908",
         12866 => x"5ae57a34",
         12867 => x"810b8317",
         12868 => x"34901908",
         12869 => x"7b27a538",
         12870 => x"80527851",
         12871 => x"fefcae3f",
         12872 => x"84ba8c08",
         12873 => x"5584ba8c",
         12874 => x"08802eff",
         12875 => x"98388256",
         12876 => x"74842ef9",
         12877 => x"e1387456",
         12878 => x"74f9db38",
         12879 => x"7f51fee5",
         12880 => x"9d3f84ba",
         12881 => x"8c0884ba",
         12882 => x"8c0cb13d",
         12883 => x"0d04820b",
         12884 => x"84ba8c0c",
         12885 => x"b13d0d04",
         12886 => x"95183394",
         12887 => x"19337198",
         12888 => x"2b71902b",
         12889 => x"07780758",
         12890 => x"565cfd8d",
         12891 => x"3984ba8c",
         12892 => x"08842efb",
         12893 => x"fe3884ba",
         12894 => x"8c08802e",
         12895 => x"fea03875",
         12896 => x"84ba8c0c",
         12897 => x"b13d0d04",
         12898 => x"8154b416",
         12899 => x"08537b52",
         12900 => x"81163351",
         12901 => x"fee2943f",
         12902 => x"815884ba",
         12903 => x"8c087a2e",
         12904 => x"098106fe",
         12905 => x"db3884ba",
         12906 => x"8c088317",
         12907 => x"34b41608",
         12908 => x"a8170831",
         12909 => x"84ba8c08",
         12910 => x"595574a0",
         12911 => x"170827fe",
         12912 => x"a0388216",
         12913 => x"335d7c82",
         12914 => x"2e098106",
         12915 => x"fe933881",
         12916 => x"54b41608",
         12917 => x"a0170805",
         12918 => x"537b5281",
         12919 => x"163351fe",
         12920 => x"e1c93f79",
         12921 => x"58fdfa39",
         12922 => x"8154b417",
         12923 => x"0853b817",
         12924 => x"70538118",
         12925 => x"33525bfe",
         12926 => x"e1b13f81",
         12927 => x"5c84ba8c",
         12928 => x"08fcc938",
         12929 => x"84ba8c08",
         12930 => x"831834b4",
         12931 => x"1708a818",
         12932 => x"083184ba",
         12933 => x"8c085d55",
         12934 => x"74a01808",
         12935 => x"27fc8e38",
         12936 => x"8217335d",
         12937 => x"7c822e09",
         12938 => x"8106fc81",
         12939 => x"388154b4",
         12940 => x"1708a018",
         12941 => x"0805537a",
         12942 => x"52811733",
         12943 => x"51fee0eb",
         12944 => x"3f795cfb",
         12945 => x"e839ec3d",
         12946 => x"0d0280df",
         12947 => x"05330284",
         12948 => x"0580e305",
         12949 => x"33565782",
         12950 => x"53963dcc",
         12951 => x"0552973d",
         12952 => x"51ffa2d8",
         12953 => x"3f84ba8c",
         12954 => x"085684ba",
         12955 => x"8c08802e",
         12956 => x"8a387584",
         12957 => x"ba8c0c96",
         12958 => x"3d0d0478",
         12959 => x"5a665296",
         12960 => x"3dd00551",
         12961 => x"ff96d73f",
         12962 => x"84ba8c08",
         12963 => x"5684ba8c",
         12964 => x"08e03802",
         12965 => x"80cf0533",
         12966 => x"81a00654",
         12967 => x"865673d2",
         12968 => x"3874a706",
         12969 => x"6171098b",
         12970 => x"12337106",
         12971 => x"7a740607",
         12972 => x"51565755",
         12973 => x"738b1734",
         12974 => x"7855810b",
         12975 => x"83163478",
         12976 => x"51fee29a",
         12977 => x"3f84ba8c",
         12978 => x"0884ba8c",
         12979 => x"0c963d0d",
         12980 => x"04ec3d0d",
         12981 => x"67578253",
         12982 => x"963dcc05",
         12983 => x"52973d51",
         12984 => x"ffa1d93f",
         12985 => x"84ba8c08",
         12986 => x"5584ba8c",
         12987 => x"08802e8a",
         12988 => x"387484ba",
         12989 => x"8c0c963d",
         12990 => x"0d04785a",
         12991 => x"6652963d",
         12992 => x"d00551ff",
         12993 => x"95d83f84",
         12994 => x"ba8c0855",
         12995 => x"84ba8c08",
         12996 => x"e0380280",
         12997 => x"cf053381",
         12998 => x"a0065686",
         12999 => x"5575d238",
         13000 => x"60841822",
         13001 => x"86192271",
         13002 => x"902b0759",
         13003 => x"59567696",
         13004 => x"17347688",
         13005 => x"2a557497",
         13006 => x"17347690",
         13007 => x"2a587798",
         13008 => x"17347698",
         13009 => x"2a547399",
         13010 => x"17347857",
         13011 => x"810b8318",
         13012 => x"347851fe",
         13013 => x"e1883f84",
         13014 => x"ba8c0884",
         13015 => x"ba8c0c96",
         13016 => x"3d0d04e8",
         13017 => x"3d0d6b6d",
         13018 => x"5d5b8053",
         13019 => x"9a3dcc05",
         13020 => x"529b3d51",
         13021 => x"ffa0c53f",
         13022 => x"84ba8c08",
         13023 => x"84ba8c08",
         13024 => x"307084ba",
         13025 => x"8c080780",
         13026 => x"25515657",
         13027 => x"7a802e8b",
         13028 => x"38817076",
         13029 => x"065a5678",
         13030 => x"81a43876",
         13031 => x"30707807",
         13032 => x"8025565b",
         13033 => x"7b802e81",
         13034 => x"8c388170",
         13035 => x"76065a58",
         13036 => x"78802e81",
         13037 => x"80387ca4",
         13038 => x"11085856",
         13039 => x"805ab416",
         13040 => x"08772e82",
         13041 => x"f6388316",
         13042 => x"337a5a55",
         13043 => x"747a2e09",
         13044 => x"81068198",
         13045 => x"38815476",
         13046 => x"53b81652",
         13047 => x"81163351",
         13048 => x"fedcc93f",
         13049 => x"84ba8c08",
         13050 => x"802e8538",
         13051 => x"ff578159",
         13052 => x"76b4170c",
         13053 => x"785778bd",
         13054 => x"387c7033",
         13055 => x"565880c3",
         13056 => x"5674832e",
         13057 => x"8b3880e4",
         13058 => x"5674842e",
         13059 => x"8338a756",
         13060 => x"7518b805",
         13061 => x"83113382",
         13062 => x"12337190",
         13063 => x"2b71882b",
         13064 => x"07811433",
         13065 => x"70720788",
         13066 => x"2b753371",
         13067 => x"07620c5f",
         13068 => x"5d5e5759",
         13069 => x"567684ba",
         13070 => x"8c0c9a3d",
         13071 => x"0d047c5e",
         13072 => x"80408052",
         13073 => x"8e3d7052",
         13074 => x"55fef48b",
         13075 => x"3f84ba8c",
         13076 => x"085784ba",
         13077 => x"8c08802e",
         13078 => x"818d3876",
         13079 => x"842e0981",
         13080 => x"06feb838",
         13081 => x"807b3480",
         13082 => x"57feb039",
         13083 => x"7754b416",
         13084 => x"0853b816",
         13085 => x"70538117",
         13086 => x"33525bfe",
         13087 => x"dcad3f77",
         13088 => x"5984ba8c",
         13089 => x"087a2e09",
         13090 => x"8106fee8",
         13091 => x"3884ba8c",
         13092 => x"08831734",
         13093 => x"b41608a8",
         13094 => x"17083184",
         13095 => x"ba8c085a",
         13096 => x"5574a017",
         13097 => x"0827fead",
         13098 => x"38821633",
         13099 => x"5574822e",
         13100 => x"098106fe",
         13101 => x"a0387754",
         13102 => x"b41608a0",
         13103 => x"17080553",
         13104 => x"7a528116",
         13105 => x"3351fedb",
         13106 => x"e23f7959",
         13107 => x"81547653",
         13108 => x"b8165281",
         13109 => x"163351fe",
         13110 => x"dad23f84",
         13111 => x"ba8c0880",
         13112 => x"2efe8d38",
         13113 => x"fe863975",
         13114 => x"527451fe",
         13115 => x"f8bb3f84",
         13116 => x"ba8c0857",
         13117 => x"84ba8c08",
         13118 => x"fee13884",
         13119 => x"ba8c0884",
         13120 => x"ba8c0866",
         13121 => x"5c595979",
         13122 => x"1881197c",
         13123 => x"1b575956",
         13124 => x"75337534",
         13125 => x"8119598a",
         13126 => x"7827ec38",
         13127 => x"8b701c57",
         13128 => x"58807634",
         13129 => x"77802efc",
         13130 => x"f238ff18",
         13131 => x"7b117033",
         13132 => x"5c575879",
         13133 => x"a02eea38",
         13134 => x"fce13979",
         13135 => x"57fdba39",
         13136 => x"e13d0d82",
         13137 => x"53a13dff",
         13138 => x"b40552a2",
         13139 => x"3d51ff9c",
         13140 => x"eb3f84ba",
         13141 => x"8c085684",
         13142 => x"ba8c0882",
         13143 => x"a6388f3d",
         13144 => x"5d8b7d57",
         13145 => x"55a07670",
         13146 => x"81055834",
         13147 => x"ff155574",
         13148 => x"f43874a3",
         13149 => x"3d087033",
         13150 => x"7081ff06",
         13151 => x"5b58585a",
         13152 => x"9f782781",
         13153 => x"b738a23d",
         13154 => x"903d5c5c",
         13155 => x"7581ff06",
         13156 => x"81185755",
         13157 => x"7481f538",
         13158 => x"757c0c74",
         13159 => x"83ffff26",
         13160 => x"81ff3874",
         13161 => x"51a1953f",
         13162 => x"83b55284",
         13163 => x"ba8c0851",
         13164 => x"9fdc3f84",
         13165 => x"ba8c0883",
         13166 => x"ffff0657",
         13167 => x"76802e81",
         13168 => x"e03883e7",
         13169 => x"9c0b83e7",
         13170 => x"9c337081",
         13171 => x"ff065b56",
         13172 => x"5878802e",
         13173 => x"81d63874",
         13174 => x"5678772e",
         13175 => x"99388118",
         13176 => x"70337081",
         13177 => x"ff065757",
         13178 => x"5874802e",
         13179 => x"89387477",
         13180 => x"2e098106",
         13181 => x"e9387581",
         13182 => x"ff065978",
         13183 => x"81a33881",
         13184 => x"ff772781",
         13185 => x"f8387989",
         13186 => x"26819638",
         13187 => x"81ff7727",
         13188 => x"8f387688",
         13189 => x"2a55747b",
         13190 => x"7081055d",
         13191 => x"34811a5a",
         13192 => x"767b7081",
         13193 => x"055d3481",
         13194 => x"1aa33d08",
         13195 => x"70337081",
         13196 => x"ff065b58",
         13197 => x"585a779f",
         13198 => x"26fed138",
         13199 => x"8f3d3357",
         13200 => x"86567681",
         13201 => x"e52ebc38",
         13202 => x"79802e99",
         13203 => x"3802b705",
         13204 => x"56791670",
         13205 => x"335c5c7a",
         13206 => x"a02e0981",
         13207 => x"068738ff",
         13208 => x"1a5a79ed",
         13209 => x"387d4580",
         13210 => x"47805295",
         13211 => x"3d705256",
         13212 => x"feefe43f",
         13213 => x"84ba8c08",
         13214 => x"5584ba8c",
         13215 => x"08802eb4",
         13216 => x"38745675",
         13217 => x"84ba8c0c",
         13218 => x"a13d0d04",
         13219 => x"83b55274",
         13220 => x"519ee73f",
         13221 => x"84ba8c08",
         13222 => x"83ffff06",
         13223 => x"5574fdf8",
         13224 => x"38865675",
         13225 => x"84ba8c0c",
         13226 => x"a13d0d04",
         13227 => x"83e79c33",
         13228 => x"56fec339",
         13229 => x"81527551",
         13230 => x"fef4ee3f",
         13231 => x"84ba8c08",
         13232 => x"5584ba8c",
         13233 => x"0880c138",
         13234 => x"79802e82",
         13235 => x"c4388b6c",
         13236 => x"7e595755",
         13237 => x"76708105",
         13238 => x"58337670",
         13239 => x"81055834",
         13240 => x"ff155574",
         13241 => x"ef387d5d",
         13242 => x"810b831e",
         13243 => x"347d51fe",
         13244 => x"d9ec3f84",
         13245 => x"ba8c0855",
         13246 => x"7456ff87",
         13247 => x"398a7a27",
         13248 => x"fe8a3886",
         13249 => x"56ff9c39",
         13250 => x"84ba8c08",
         13251 => x"842e0981",
         13252 => x"06feee38",
         13253 => x"80557975",
         13254 => x"2efee638",
         13255 => x"75087553",
         13256 => x"765258fe",
         13257 => x"eeb13f84",
         13258 => x"ba8c0857",
         13259 => x"84ba8c08",
         13260 => x"752e0981",
         13261 => x"06818438",
         13262 => x"84ba8c08",
         13263 => x"b8195c5a",
         13264 => x"98160857",
         13265 => x"8059b418",
         13266 => x"08772eb2",
         13267 => x"38831833",
         13268 => x"5574792e",
         13269 => x"09810681",
         13270 => x"d7388154",
         13271 => x"7653b818",
         13272 => x"52811833",
         13273 => x"51fed5c4",
         13274 => x"3f84ba8c",
         13275 => x"08802e85",
         13276 => x"38ff5781",
         13277 => x"5976b419",
         13278 => x"0c785778",
         13279 => x"be38789c",
         13280 => x"17087033",
         13281 => x"575a5774",
         13282 => x"81e52e81",
         13283 => x"9e387430",
         13284 => x"70802578",
         13285 => x"07565c74",
         13286 => x"802e81d7",
         13287 => x"38811a5a",
         13288 => x"79812ea5",
         13289 => x"38815275",
         13290 => x"51feefa1",
         13291 => x"3f84ba8c",
         13292 => x"085784ba",
         13293 => x"8c08802e",
         13294 => x"ff863887",
         13295 => x"5576842e",
         13296 => x"fdbf3876",
         13297 => x"5576fdb9",
         13298 => x"38a06c57",
         13299 => x"55807670",
         13300 => x"81055834",
         13301 => x"ff155574",
         13302 => x"f4386b56",
         13303 => x"880b8b17",
         13304 => x"348b6c7e",
         13305 => x"59575576",
         13306 => x"70810558",
         13307 => x"33767081",
         13308 => x"055834ff",
         13309 => x"15557480",
         13310 => x"2efdeb38",
         13311 => x"76708105",
         13312 => x"58337670",
         13313 => x"81055834",
         13314 => x"ff155574",
         13315 => x"da38fdd6",
         13316 => x"396b5ae5",
         13317 => x"7a347d5d",
         13318 => x"810b831e",
         13319 => x"347d51fe",
         13320 => x"d7bc3f84",
         13321 => x"ba8c0855",
         13322 => x"fdce3981",
         13323 => x"57fedf39",
         13324 => x"8154b418",
         13325 => x"08537a52",
         13326 => x"81183351",
         13327 => x"fed4ec3f",
         13328 => x"84ba8c08",
         13329 => x"792e0981",
         13330 => x"0680c338",
         13331 => x"84ba8c08",
         13332 => x"831934b4",
         13333 => x"1808a819",
         13334 => x"08315c7b",
         13335 => x"a0190827",
         13336 => x"8a388218",
         13337 => x"33557482",
         13338 => x"2eb13884",
         13339 => x"ba8c0859",
         13340 => x"fde83974",
         13341 => x"5a815275",
         13342 => x"51feedd1",
         13343 => x"3f84ba8c",
         13344 => x"085784ba",
         13345 => x"8c08802e",
         13346 => x"fdb638fe",
         13347 => x"ae398170",
         13348 => x"58597880",
         13349 => x"2efde738",
         13350 => x"fea13981",
         13351 => x"54b41808",
         13352 => x"a0190805",
         13353 => x"537a5281",
         13354 => x"183351fe",
         13355 => x"d3fd3ffd",
         13356 => x"a939f23d",
         13357 => x"0d606202",
         13358 => x"880580cb",
         13359 => x"05335e5b",
         13360 => x"57895676",
         13361 => x"802e9f38",
         13362 => x"76085574",
         13363 => x"802e9738",
         13364 => x"74335473",
         13365 => x"802e8f38",
         13366 => x"86152284",
         13367 => x"18225959",
         13368 => x"78782e81",
         13369 => x"c2388054",
         13370 => x"735f7581",
         13371 => x"a5389117",
         13372 => x"33567581",
         13373 => x"9d387980",
         13374 => x"2e81a238",
         13375 => x"8c170881",
         13376 => x"9c389017",
         13377 => x"3370812a",
         13378 => x"8106565d",
         13379 => x"74802e81",
         13380 => x"8c387e8a",
         13381 => x"11227089",
         13382 => x"2b70557c",
         13383 => x"54575c59",
         13384 => x"fd87823f",
         13385 => x"ff157a06",
         13386 => x"70307072",
         13387 => x"079f2a84",
         13388 => x"ba8c0805",
         13389 => x"901c0879",
         13390 => x"42535f55",
         13391 => x"58817827",
         13392 => x"88389c19",
         13393 => x"08782683",
         13394 => x"38825877",
         13395 => x"78565b80",
         13396 => x"59745276",
         13397 => x"51fed887",
         13398 => x"3f81157f",
         13399 => x"55559c14",
         13400 => x"08752683",
         13401 => x"38825584",
         13402 => x"ba8c0881",
         13403 => x"2e81dc38",
         13404 => x"84ba8c08",
         13405 => x"ff2e81d8",
         13406 => x"3884ba8c",
         13407 => x"0881c538",
         13408 => x"81195978",
         13409 => x"7d2ebb38",
         13410 => x"74782e09",
         13411 => x"8106c238",
         13412 => x"87567554",
         13413 => x"7384ba8c",
         13414 => x"0c903d0d",
         13415 => x"04870b84",
         13416 => x"ba8c0c90",
         13417 => x"3d0d0481",
         13418 => x"153351fe",
         13419 => x"d0ac3f84",
         13420 => x"ba8c0881",
         13421 => x"065473fe",
         13422 => x"ad387377",
         13423 => x"085556fe",
         13424 => x"a7397b80",
         13425 => x"2e818e38",
         13426 => x"7a7d5658",
         13427 => x"7c802eab",
         13428 => x"38811854",
         13429 => x"74812e80",
         13430 => x"e6387353",
         13431 => x"77527e51",
         13432 => x"fedddd3f",
         13433 => x"84ba8c08",
         13434 => x"5684ba8c",
         13435 => x"08ffa338",
         13436 => x"778119ff",
         13437 => x"1757595e",
         13438 => x"74d7387e",
         13439 => x"7e90120c",
         13440 => x"557b802e",
         13441 => x"ff8c387a",
         13442 => x"88180c79",
         13443 => x"8c180c90",
         13444 => x"173380c0",
         13445 => x"075c7b90",
         13446 => x"18349c15",
         13447 => x"08fe0594",
         13448 => x"1608585a",
         13449 => x"767a26fe",
         13450 => x"e938767d",
         13451 => x"3194160c",
         13452 => x"84153381",
         13453 => x"075d7c84",
         13454 => x"16347554",
         13455 => x"fed639ff",
         13456 => x"54ff9739",
         13457 => x"745b8059",
         13458 => x"febe3982",
         13459 => x"54fec539",
         13460 => x"8154fec0",
         13461 => x"39ff1b5e",
         13462 => x"ffa13984",
         13463 => x"ba9808e3",
         13464 => x"3d0da33d",
         13465 => x"08a53d08",
         13466 => x"02880581",
         13467 => x"87053344",
         13468 => x"425fff0b",
         13469 => x"a23d0870",
         13470 => x"5f5b4079",
         13471 => x"802e858a",
         13472 => x"38797081",
         13473 => x"055b3370",
         13474 => x"9f265656",
         13475 => x"75ba2e85",
         13476 => x"9b3874ed",
         13477 => x"3875ba2e",
         13478 => x"85923884",
         13479 => x"d1e83356",
         13480 => x"80762484",
         13481 => x"e5387510",
         13482 => x"1084d1d4",
         13483 => x"05700856",
         13484 => x"5a74802e",
         13485 => x"84388075",
         13486 => x"34751684",
         13487 => x"ba801133",
         13488 => x"84ba8112",
         13489 => x"33405b5d",
         13490 => x"81527951",
         13491 => x"fecea93f",
         13492 => x"84ba8c08",
         13493 => x"81ff0670",
         13494 => x"81065d56",
         13495 => x"83577b84",
         13496 => x"ab387582",
         13497 => x"2a810640",
         13498 => x"8a577f84",
         13499 => x"9f389f3d",
         13500 => x"fc055383",
         13501 => x"527951fe",
         13502 => x"d0b03f84",
         13503 => x"ba8c0884",
         13504 => x"98386d55",
         13505 => x"74802e84",
         13506 => x"90387482",
         13507 => x"80802684",
         13508 => x"8838ff15",
         13509 => x"75065574",
         13510 => x"83ff387e",
         13511 => x"802e8838",
         13512 => x"84807f26",
         13513 => x"83f8387e",
         13514 => x"81800a26",
         13515 => x"83f038ff",
         13516 => x"1f7f0655",
         13517 => x"7483e738",
         13518 => x"7e892aa6",
         13519 => x"3d08892a",
         13520 => x"70892b77",
         13521 => x"594c475b",
         13522 => x"60802e85",
         13523 => x"ab386530",
         13524 => x"70802577",
         13525 => x"07565f91",
         13526 => x"577483b0",
         13527 => x"387d802e",
         13528 => x"84df3881",
         13529 => x"54745360",
         13530 => x"527951fe",
         13531 => x"cdbe3f81",
         13532 => x"5784ba8c",
         13533 => x"08839538",
         13534 => x"6083ff05",
         13535 => x"336183fe",
         13536 => x"05337188",
         13537 => x"2b075956",
         13538 => x"8e577782",
         13539 => x"d4d52e09",
         13540 => x"810682f8",
         13541 => x"387d9029",
         13542 => x"610583b2",
         13543 => x"11334458",
         13544 => x"62802e82",
         13545 => x"e73883b6",
         13546 => x"18831133",
         13547 => x"82123371",
         13548 => x"902b7188",
         13549 => x"2b078114",
         13550 => x"33707207",
         13551 => x"882b7533",
         13552 => x"710783ba",
         13553 => x"1f831133",
         13554 => x"82123371",
         13555 => x"902b7188",
         13556 => x"2b078114",
         13557 => x"33707207",
         13558 => x"882b7533",
         13559 => x"71075ca2",
         13560 => x"3d0c42a3",
         13561 => x"3d0ca33d",
         13562 => x"0c444e54",
         13563 => x"45594f41",
         13564 => x"5a4b784d",
         13565 => x"8e5780ff",
         13566 => x"79278290",
         13567 => x"3893577a",
         13568 => x"81802682",
         13569 => x"87386181",
         13570 => x"2a708106",
         13571 => x"45496380",
         13572 => x"2e83f938",
         13573 => x"61870645",
         13574 => x"64822e89",
         13575 => x"38618106",
         13576 => x"476683f4",
         13577 => x"38836e70",
         13578 => x"304a4643",
         13579 => x"7a586283",
         13580 => x"2e8ac238",
         13581 => x"7aae3878",
         13582 => x"8c2a5781",
         13583 => x"0b83e7b0",
         13584 => x"22565874",
         13585 => x"802e9d38",
         13586 => x"74772698",
         13587 => x"3883e7b0",
         13588 => x"56771082",
         13589 => x"17702257",
         13590 => x"57587480",
         13591 => x"2e863876",
         13592 => x"7527ee38",
         13593 => x"77527851",
         13594 => x"fd80ba3f",
         13595 => x"84ba8c08",
         13596 => x"10840555",
         13597 => x"84ba8c08",
         13598 => x"9ff52696",
         13599 => x"38810b84",
         13600 => x"ba8c0810",
         13601 => x"84ba8c08",
         13602 => x"05711172",
         13603 => x"2a830557",
         13604 => x"4c4383ff",
         13605 => x"15892a5d",
         13606 => x"815ca047",
         13607 => x"7b1f7d11",
         13608 => x"68056611",
         13609 => x"ff05706b",
         13610 => x"06723158",
         13611 => x"4e574462",
         13612 => x"832e89b8",
         13613 => x"38741d5d",
         13614 => x"77902916",
         13615 => x"70603156",
         13616 => x"57747926",
         13617 => x"82f23878",
         13618 => x"7c317d31",
         13619 => x"78537068",
         13620 => x"315256fc",
         13621 => x"ffcf3f84",
         13622 => x"ba8c0840",
         13623 => x"62832e89",
         13624 => x"f6386282",
         13625 => x"2e098106",
         13626 => x"82dd3883",
         13627 => x"fff50b84",
         13628 => x"ba8c0827",
         13629 => x"82ac387a",
         13630 => x"89f93877",
         13631 => x"18557480",
         13632 => x"c02689ef",
         13633 => x"38745bfe",
         13634 => x"a3398b57",
         13635 => x"7684ba8c",
         13636 => x"0c9f3d0d",
         13637 => x"84ba980c",
         13638 => x"04814efb",
         13639 => x"fe39930b",
         13640 => x"84ba8c0c",
         13641 => x"9f3d0d84",
         13642 => x"ba980c04",
         13643 => x"7c33d011",
         13644 => x"7081ff06",
         13645 => x"57575774",
         13646 => x"89269138",
         13647 => x"821d7781",
         13648 => x"ff06d005",
         13649 => x"5d58777a",
         13650 => x"2e81b238",
         13651 => x"800b83e5",
         13652 => x"fc5f5c7d",
         13653 => x"087d575b",
         13654 => x"7a708105",
         13655 => x"5c337670",
         13656 => x"81055833",
         13657 => x"ff9f1245",
         13658 => x"59576299",
         13659 => x"268938e0",
         13660 => x"177081ff",
         13661 => x"065844ff",
         13662 => x"9f184564",
         13663 => x"99268938",
         13664 => x"e0187081",
         13665 => x"ff065946",
         13666 => x"7630709f",
         13667 => x"2a5a4776",
         13668 => x"782e0981",
         13669 => x"06853878",
         13670 => x"ffbe3875",
         13671 => x"7a327030",
         13672 => x"7072079f",
         13673 => x"2a7b075d",
         13674 => x"4a4a7a80",
         13675 => x"2e80ce38",
         13676 => x"811c841f",
         13677 => x"5f5c837c",
         13678 => x"25ff9838",
         13679 => x"7f56f9e0",
         13680 => x"399f3df8",
         13681 => x"05538152",
         13682 => x"7951feca",
         13683 => x"dd3f8157",
         13684 => x"84ba8c08",
         13685 => x"feb63861",
         13686 => x"832a7706",
         13687 => x"84ba8c08",
         13688 => x"40567583",
         13689 => x"38bf5f6c",
         13690 => x"558e577e",
         13691 => x"7526fe9c",
         13692 => x"38747f31",
         13693 => x"59fbfb39",
         13694 => x"8156fad2",
         13695 => x"397b8324",
         13696 => x"ffba387b",
         13697 => x"7aa33d0c",
         13698 => x"56f99539",
         13699 => x"61810648",
         13700 => x"93576780",
         13701 => x"2efdf538",
         13702 => x"826e7030",
         13703 => x"4a4643fc",
         13704 => x"8b3984ba",
         13705 => x"8c089ff5",
         13706 => x"269d387a",
         13707 => x"8b387718",
         13708 => x"5b81807b",
         13709 => x"27fbf538",
         13710 => x"8e577684",
         13711 => x"ba8c0c9f",
         13712 => x"3d0d84ba",
         13713 => x"980c0480",
         13714 => x"5562812e",
         13715 => x"8699389f",
         13716 => x"f560278b",
         13717 => x"38748106",
         13718 => x"5b8e577a",
         13719 => x"fdae3884",
         13720 => x"80615755",
         13721 => x"80767081",
         13722 => x"055834ff",
         13723 => x"155574f4",
         13724 => x"388b6183",
         13725 => x"e5c85957",
         13726 => x"55767081",
         13727 => x"05583376",
         13728 => x"70810558",
         13729 => x"34ff1555",
         13730 => x"74ef3860",
         13731 => x"8b054574",
         13732 => x"65348261",
         13733 => x"8c053477",
         13734 => x"618d0534",
         13735 => x"7b83ffff",
         13736 => x"064b6a61",
         13737 => x"8e05346a",
         13738 => x"882a5c7b",
         13739 => x"618f0534",
         13740 => x"81619005",
         13741 => x"34628332",
         13742 => x"70305a48",
         13743 => x"80619105",
         13744 => x"34789e2a",
         13745 => x"82064968",
         13746 => x"61920534",
         13747 => x"6c567583",
         13748 => x"ffff2686",
         13749 => x"ad387583",
         13750 => x"ffff0655",
         13751 => x"74619305",
         13752 => x"3474882a",
         13753 => x"4c6b6194",
         13754 => x"0534f861",
         13755 => x"950534bf",
         13756 => x"61980534",
         13757 => x"80619905",
         13758 => x"34ff619a",
         13759 => x"05348061",
         13760 => x"9b05347e",
         13761 => x"619c0534",
         13762 => x"7e882a48",
         13763 => x"67619d05",
         13764 => x"347e902a",
         13765 => x"4c6b619e",
         13766 => x"05347e98",
         13767 => x"2a84ba98",
         13768 => x"0c84ba98",
         13769 => x"08619f05",
         13770 => x"3462832e",
         13771 => x"85f73880",
         13772 => x"61a70534",
         13773 => x"8061a805",
         13774 => x"34a161a9",
         13775 => x"053480cc",
         13776 => x"61aa0534",
         13777 => x"7c83ffff",
         13778 => x"06557461",
         13779 => x"96053474",
         13780 => x"882a4b6a",
         13781 => x"61970534",
         13782 => x"ff8061a4",
         13783 => x"0534a961",
         13784 => x"a6053493",
         13785 => x"61ab0583",
         13786 => x"e5d45957",
         13787 => x"55767081",
         13788 => x"05583376",
         13789 => x"70810558",
         13790 => x"34ff1555",
         13791 => x"74ef3860",
         13792 => x"83fe0549",
         13793 => x"80d56934",
         13794 => x"6083ff05",
         13795 => x"4bffaa6b",
         13796 => x"3481547e",
         13797 => x"53605279",
         13798 => x"51fec68f",
         13799 => x"3f815784",
         13800 => x"ba8c08fa",
         13801 => x"e7386017",
         13802 => x"5c62832e",
         13803 => x"879c3869",
         13804 => x"61575580",
         13805 => x"76708105",
         13806 => x"5834ff15",
         13807 => x"5574f438",
         13808 => x"6375415b",
         13809 => x"62832e86",
         13810 => x"c03887ff",
         13811 => x"fff85762",
         13812 => x"812e8338",
         13813 => x"f8577661",
         13814 => x"3476882a",
         13815 => x"7c455574",
         13816 => x"64708105",
         13817 => x"46347690",
         13818 => x"2a597864",
         13819 => x"70810546",
         13820 => x"3476982a",
         13821 => x"56756434",
         13822 => x"7c576559",
         13823 => x"76662683",
         13824 => x"38765978",
         13825 => x"547a5360",
         13826 => x"527951fe",
         13827 => x"c59d3f84",
         13828 => x"ba8c0885",
         13829 => x"e6388480",
         13830 => x"61575580",
         13831 => x"76708105",
         13832 => x"5834ff15",
         13833 => x"5574f438",
         13834 => x"781b777a",
         13835 => x"31585b76",
         13836 => x"c9387f81",
         13837 => x"05407f80",
         13838 => x"2eff8938",
         13839 => x"77566283",
         13840 => x"2e833866",
         13841 => x"56655575",
         13842 => x"66268338",
         13843 => x"75557454",
         13844 => x"7a536052",
         13845 => x"7951fec4",
         13846 => x"d23f84ba",
         13847 => x"8c08859b",
         13848 => x"38741b76",
         13849 => x"7631575b",
         13850 => x"75db388c",
         13851 => x"5862832e",
         13852 => x"93388658",
         13853 => x"6c83ffff",
         13854 => x"268a3884",
         13855 => x"5862822e",
         13856 => x"83388158",
         13857 => x"7d84c138",
         13858 => x"61832a81",
         13859 => x"065e7d81",
         13860 => x"b3388480",
         13861 => x"61565980",
         13862 => x"75708105",
         13863 => x"5734ff19",
         13864 => x"5978f438",
         13865 => x"80d56934",
         13866 => x"ffaa6b34",
         13867 => x"6083be05",
         13868 => x"47786734",
         13869 => x"81678105",
         13870 => x"34816782",
         13871 => x"05347867",
         13872 => x"83053477",
         13873 => x"67840534",
         13874 => x"6c4380fd",
         13875 => x"c152621f",
         13876 => x"51fcf7d1",
         13877 => x"3ffe6785",
         13878 => x"053484ba",
         13879 => x"8c08822a",
         13880 => x"bf075776",
         13881 => x"67860534",
         13882 => x"84ba8c08",
         13883 => x"67870534",
         13884 => x"7e6183c6",
         13885 => x"05346761",
         13886 => x"83c70534",
         13887 => x"6b6183c8",
         13888 => x"053484ba",
         13889 => x"98086183",
         13890 => x"c9053462",
         13891 => x"6183ca05",
         13892 => x"3462882a",
         13893 => x"45646183",
         13894 => x"cb053462",
         13895 => x"902a5877",
         13896 => x"6183cc05",
         13897 => x"3462982a",
         13898 => x"5f7e6183",
         13899 => x"cd053481",
         13900 => x"54785360",
         13901 => x"527951fe",
         13902 => x"c2f13f81",
         13903 => x"5784ba8c",
         13904 => x"08f7c938",
         13905 => x"80538052",
         13906 => x"7951fec3",
         13907 => x"dd3f8157",
         13908 => x"84ba8c08",
         13909 => x"f7b63884",
         13910 => x"ba8c0884",
         13911 => x"ba8c0c9f",
         13912 => x"3d0d84ba",
         13913 => x"980c0462",
         13914 => x"55f9e439",
         13915 => x"741c6416",
         13916 => x"455cf6c4",
         13917 => x"397aae38",
         13918 => x"78912a57",
         13919 => x"810b83e7",
         13920 => x"c0225658",
         13921 => x"74802e9d",
         13922 => x"38747726",
         13923 => x"983883e7",
         13924 => x"c0567710",
         13925 => x"82177022",
         13926 => x"57575874",
         13927 => x"802e8638",
         13928 => x"767527ee",
         13929 => x"38775278",
         13930 => x"51fcf5f9",
         13931 => x"3f84ba8c",
         13932 => x"08101084",
         13933 => x"87057089",
         13934 => x"2a5e5ca0",
         13935 => x"5c800b84",
         13936 => x"ba8c08fc",
         13937 => x"808a0558",
         13938 => x"47fdfff0",
         13939 => x"0a7727f5",
         13940 => x"cb388e57",
         13941 => x"f8e43984",
         13942 => x"ba8c0883",
         13943 => x"fff526f8",
         13944 => x"e6387af8",
         13945 => x"d3387781",
         13946 => x"2a5b7af4",
         13947 => x"bf388e57",
         13948 => x"f8c83968",
         13949 => x"81064463",
         13950 => x"802ef8af",
         13951 => x"388343f4",
         13952 => x"ab397561",
         13953 => x"a0053475",
         13954 => x"882a4968",
         13955 => x"61a10534",
         13956 => x"75902a5b",
         13957 => x"7a61a205",
         13958 => x"3475982a",
         13959 => x"577661a3",
         13960 => x"0534f9c6",
         13961 => x"39806180",
         13962 => x"c3053480",
         13963 => x"6180c405",
         13964 => x"34a16180",
         13965 => x"c5053480",
         13966 => x"cc6180c6",
         13967 => x"05347c61",
         13968 => x"a405347c",
         13969 => x"882a5c7b",
         13970 => x"61a50534",
         13971 => x"7c902a59",
         13972 => x"7861a605",
         13973 => x"347c982a",
         13974 => x"567561a7",
         13975 => x"05348261",
         13976 => x"ac053480",
         13977 => x"61ad0534",
         13978 => x"8061ae05",
         13979 => x"348061af",
         13980 => x"05348161",
         13981 => x"b0053480",
         13982 => x"61b10534",
         13983 => x"8661b205",
         13984 => x"348061b3",
         13985 => x"0534ff80",
         13986 => x"6180c005",
         13987 => x"34a96180",
         13988 => x"c2053493",
         13989 => x"6180c705",
         13990 => x"83e5e859",
         13991 => x"57557670",
         13992 => x"81055833",
         13993 => x"76708105",
         13994 => x"5834ff15",
         13995 => x"5574802e",
         13996 => x"f9cd3876",
         13997 => x"70810558",
         13998 => x"33767081",
         13999 => x"055834ff",
         14000 => x"155574da",
         14001 => x"38f9b839",
         14002 => x"81548053",
         14003 => x"60527951",
         14004 => x"febed93f",
         14005 => x"815784ba",
         14006 => x"8c08f4b0",
         14007 => x"387d9029",
         14008 => x"61054277",
         14009 => x"6283b205",
         14010 => x"34765484",
         14011 => x"ba8c0853",
         14012 => x"60527951",
         14013 => x"febfb43f",
         14014 => x"fcc33981",
         14015 => x"0b84ba8c",
         14016 => x"0c9f3d0d",
         14017 => x"84ba980c",
         14018 => x"04f86134",
         14019 => x"7b4aff6a",
         14020 => x"7081054c",
         14021 => x"34ff6a70",
         14022 => x"81054c34",
         14023 => x"ff6a34ff",
         14024 => x"61840534",
         14025 => x"ff618505",
         14026 => x"34ff6186",
         14027 => x"0534ff61",
         14028 => x"870534ff",
         14029 => x"61880534",
         14030 => x"ff618905",
         14031 => x"34ff618a",
         14032 => x"05348f65",
         14033 => x"347c57f9",
         14034 => x"b1397654",
         14035 => x"861f5360",
         14036 => x"527951fe",
         14037 => x"bed53f84",
         14038 => x"80615657",
         14039 => x"80757081",
         14040 => x"055734ff",
         14041 => x"175776f4",
         14042 => x"38605c80",
         14043 => x"d27c7081",
         14044 => x"055e347b",
         14045 => x"5580d275",
         14046 => x"70810557",
         14047 => x"3480e175",
         14048 => x"70810557",
         14049 => x"3480c175",
         14050 => x"3480f261",
         14051 => x"83e40534",
         14052 => x"80f26183",
         14053 => x"e5053480",
         14054 => x"c16183e6",
         14055 => x"053480e1",
         14056 => x"6183e705",
         14057 => x"347fff05",
         14058 => x"5b7a6183",
         14059 => x"e805347a",
         14060 => x"882a5978",
         14061 => x"6183e905",
         14062 => x"347a902a",
         14063 => x"56756183",
         14064 => x"ea05347a",
         14065 => x"982a407f",
         14066 => x"6183eb05",
         14067 => x"34826183",
         14068 => x"ec053476",
         14069 => x"6183ed05",
         14070 => x"34766183",
         14071 => x"ee053476",
         14072 => x"6183ef05",
         14073 => x"3480d569",
         14074 => x"34ffaa6b",
         14075 => x"34815487",
         14076 => x"1f536052",
         14077 => x"7951febd",
         14078 => x"b23f8154",
         14079 => x"811f5360",
         14080 => x"527951fe",
         14081 => x"bda53f69",
         14082 => x"615755f7",
         14083 => x"a639f43d",
         14084 => x"0d7e615b",
         14085 => x"5b807b61",
         14086 => x"ff055a57",
         14087 => x"57767825",
         14088 => x"b8388d3d",
         14089 => x"598e3df8",
         14090 => x"05548153",
         14091 => x"78527951",
         14092 => x"ff9ab43f",
         14093 => x"7b812e09",
         14094 => x"81069e38",
         14095 => x"8d3d3355",
         14096 => x"748d2e90",
         14097 => x"38747670",
         14098 => x"81055834",
         14099 => x"81175774",
         14100 => x"8a2e8638",
         14101 => x"777724cd",
         14102 => x"38807634",
         14103 => x"7a557683",
         14104 => x"38765574",
         14105 => x"84ba8c0c",
         14106 => x"8e3d0d04",
         14107 => x"f73d0d7b",
         14108 => x"028405b3",
         14109 => x"05335957",
         14110 => x"778a2e80",
         14111 => x"d5388417",
         14112 => x"08568076",
         14113 => x"249e3888",
         14114 => x"17087717",
         14115 => x"8c055659",
         14116 => x"77753481",
         14117 => x"165574bb",
         14118 => x"248e3874",
         14119 => x"84180c81",
         14120 => x"1988180c",
         14121 => x"8b3d0d04",
         14122 => x"8b3dfc05",
         14123 => x"5474538c",
         14124 => x"17527608",
         14125 => x"51ff9ed1",
         14126 => x"3f747a32",
         14127 => x"70307072",
         14128 => x"079f2a70",
         14129 => x"30841b0c",
         14130 => x"811c881b",
         14131 => x"0c5a5656",
         14132 => x"d3398d52",
         14133 => x"7651ff94",
         14134 => x"3fffa339",
         14135 => x"e33d0d02",
         14136 => x"80ff0533",
         14137 => x"8d3d5858",
         14138 => x"80cc7757",
         14139 => x"55807670",
         14140 => x"81055834",
         14141 => x"ff155574",
         14142 => x"f438a13d",
         14143 => x"08770c77",
         14144 => x"8a2e80f7",
         14145 => x"387c5680",
         14146 => x"762480c0",
         14147 => x"387d7717",
         14148 => x"8c055659",
         14149 => x"77753481",
         14150 => x"165574bb",
         14151 => x"24b83874",
         14152 => x"84180c81",
         14153 => x"1988180c",
         14154 => x"7c558075",
         14155 => x"249e389f",
         14156 => x"3dffac11",
         14157 => x"557554c0",
         14158 => x"05527608",
         14159 => x"51ff9dc9",
         14160 => x"3f84ba8c",
         14161 => x"0886387c",
         14162 => x"7a2eba38",
         14163 => x"ff0b84ba",
         14164 => x"8c0c9f3d",
         14165 => x"0d049f3d",
         14166 => x"ffb01155",
         14167 => x"7554c005",
         14168 => x"52760851",
         14169 => x"ff9da23f",
         14170 => x"747b3270",
         14171 => x"30707207",
         14172 => x"9f2a7030",
         14173 => x"525a5656",
         14174 => x"ffa5398d",
         14175 => x"527651fd",
         14176 => x"eb3fff81",
         14177 => x"397d84ba",
         14178 => x"8c0c9f3d",
         14179 => x"0d04fd3d",
         14180 => x"0d750284",
         14181 => x"059a0522",
         14182 => x"52538052",
         14183 => x"7280ff26",
         14184 => x"90387283",
         14185 => x"ffff0652",
         14186 => x"7184ba8c",
         14187 => x"0c853d0d",
         14188 => x"0483ffff",
         14189 => x"73275470",
         14190 => x"83b52e09",
         14191 => x"8106e938",
         14192 => x"73802ee4",
         14193 => x"3883e7d0",
         14194 => x"22517271",
         14195 => x"2e9c3881",
         14196 => x"127083ff",
         14197 => x"ff065354",
         14198 => x"7180ff26",
         14199 => x"8d387110",
         14200 => x"83e7d005",
         14201 => x"70225151",
         14202 => x"e1398180",
         14203 => x"127081ff",
         14204 => x"0684ba8c",
         14205 => x"0c53853d",
         14206 => x"0d04fe3d",
         14207 => x"0d029205",
         14208 => x"22028405",
         14209 => x"96052253",
         14210 => x"51805370",
         14211 => x"80ff268c",
         14212 => x"38705372",
         14213 => x"84ba8c0c",
         14214 => x"843d0d04",
         14215 => x"7183b52e",
         14216 => x"098106ef",
         14217 => x"387081ff",
         14218 => x"26e93870",
         14219 => x"1083e5d0",
         14220 => x"05702284",
         14221 => x"ba8c0c51",
         14222 => x"843d0d04",
         14223 => x"fb3d0d77",
         14224 => x"517083ff",
         14225 => x"ff2680e1",
         14226 => x"387083ff",
         14227 => x"ff0683e9",
         14228 => x"d0565675",
         14229 => x"9fff2680",
         14230 => x"d9387470",
         14231 => x"82055622",
         14232 => x"75713070",
         14233 => x"8025737a",
         14234 => x"26075456",
         14235 => x"535370b7",
         14236 => x"38717082",
         14237 => x"05532272",
         14238 => x"71882a54",
         14239 => x"5681ff06",
         14240 => x"70145254",
         14241 => x"707624b1",
         14242 => x"3871cf38",
         14243 => x"73101570",
         14244 => x"70820552",
         14245 => x"22547330",
         14246 => x"70802575",
         14247 => x"79260753",
         14248 => x"55527080",
         14249 => x"2ecb3875",
         14250 => x"517084ba",
         14251 => x"8c0c873d",
         14252 => x"0d0483ed",
         14253 => x"c455ffa2",
         14254 => x"39718826",
         14255 => x"ea387110",
         14256 => x"1083caa8",
         14257 => x"05547308",
         14258 => x"04c7a016",
         14259 => x"7083ffff",
         14260 => x"06575175",
         14261 => x"51d339ff",
         14262 => x"b0167083",
         14263 => x"ffff0657",
         14264 => x"51f13988",
         14265 => x"167083ff",
         14266 => x"ff065751",
         14267 => x"e639e616",
         14268 => x"7083ffff",
         14269 => x"065751db",
         14270 => x"39d01670",
         14271 => x"83ffff06",
         14272 => x"5751d039",
         14273 => x"e0167083",
         14274 => x"ffff0657",
         14275 => x"51c539f0",
         14276 => x"167083ff",
         14277 => x"ff065751",
         14278 => x"ffb93975",
         14279 => x"73318106",
         14280 => x"76713170",
         14281 => x"83ffff06",
         14282 => x"585255ff",
         14283 => x"a6397573",
         14284 => x"31107505",
         14285 => x"70225252",
         14286 => x"feef3900",
         14287 => x"00ffffff",
         14288 => x"ff00ffff",
         14289 => x"ffff00ff",
         14290 => x"ffffff00",
         14291 => x"0000198b",
         14292 => x"00001980",
         14293 => x"00001975",
         14294 => x"0000196a",
         14295 => x"0000195f",
         14296 => x"00001954",
         14297 => x"00001949",
         14298 => x"0000193e",
         14299 => x"00001933",
         14300 => x"00001928",
         14301 => x"0000191d",
         14302 => x"00001912",
         14303 => x"00001907",
         14304 => x"000018fc",
         14305 => x"000018f1",
         14306 => x"000018e6",
         14307 => x"000018db",
         14308 => x"000018d0",
         14309 => x"000018c5",
         14310 => x"000018ba",
         14311 => x"00001ebf",
         14312 => x"00001f59",
         14313 => x"00001f59",
         14314 => x"00001f59",
         14315 => x"00001f59",
         14316 => x"00001f59",
         14317 => x"00001f59",
         14318 => x"00001f59",
         14319 => x"00001f59",
         14320 => x"00001f59",
         14321 => x"00001f59",
         14322 => x"00001f59",
         14323 => x"00001f59",
         14324 => x"00001f59",
         14325 => x"00001f59",
         14326 => x"00001f59",
         14327 => x"00001f59",
         14328 => x"00001f59",
         14329 => x"00001f59",
         14330 => x"00001f59",
         14331 => x"00001f59",
         14332 => x"00001f59",
         14333 => x"00001f59",
         14334 => x"00001f59",
         14335 => x"00001f59",
         14336 => x"00001f59",
         14337 => x"00001f59",
         14338 => x"00001f59",
         14339 => x"00001f59",
         14340 => x"00001f59",
         14341 => x"00001f59",
         14342 => x"00001f59",
         14343 => x"00001f59",
         14344 => x"00001f59",
         14345 => x"00001f59",
         14346 => x"00001f59",
         14347 => x"00001f59",
         14348 => x"00001f59",
         14349 => x"00001f59",
         14350 => x"00001f59",
         14351 => x"00001f59",
         14352 => x"00001f59",
         14353 => x"00001f59",
         14354 => x"0000247b",
         14355 => x"00001f59",
         14356 => x"00001f59",
         14357 => x"00001f59",
         14358 => x"00001f59",
         14359 => x"00001f59",
         14360 => x"00001f59",
         14361 => x"00001f59",
         14362 => x"00001f59",
         14363 => x"00001f59",
         14364 => x"00001f59",
         14365 => x"00001f59",
         14366 => x"00001f59",
         14367 => x"00001f59",
         14368 => x"00001f59",
         14369 => x"00001f59",
         14370 => x"00001f59",
         14371 => x"00002411",
         14372 => x"00002310",
         14373 => x"00001f59",
         14374 => x"00002294",
         14375 => x"000024b2",
         14376 => x"00002371",
         14377 => x"00002236",
         14378 => x"000021d8",
         14379 => x"00001f59",
         14380 => x"00001f59",
         14381 => x"00001f59",
         14382 => x"00001f59",
         14383 => x"00001f59",
         14384 => x"00001f59",
         14385 => x"00001f59",
         14386 => x"00001f59",
         14387 => x"00001f59",
         14388 => x"00001f59",
         14389 => x"00001f59",
         14390 => x"00001f59",
         14391 => x"00001f59",
         14392 => x"00001f59",
         14393 => x"00001f59",
         14394 => x"00001f59",
         14395 => x"00001f59",
         14396 => x"00001f59",
         14397 => x"00001f59",
         14398 => x"00001f59",
         14399 => x"00001f59",
         14400 => x"00001f59",
         14401 => x"00001f59",
         14402 => x"00001f59",
         14403 => x"00001f59",
         14404 => x"00001f59",
         14405 => x"00001f59",
         14406 => x"00001f59",
         14407 => x"00001f59",
         14408 => x"00001f59",
         14409 => x"00001f59",
         14410 => x"00001f59",
         14411 => x"00001f59",
         14412 => x"00001f59",
         14413 => x"00001f59",
         14414 => x"00001f59",
         14415 => x"00001f59",
         14416 => x"00001f59",
         14417 => x"00001f59",
         14418 => x"00001f59",
         14419 => x"00001f59",
         14420 => x"00001f59",
         14421 => x"00001f59",
         14422 => x"00001f59",
         14423 => x"00001f59",
         14424 => x"00001f59",
         14425 => x"00001f59",
         14426 => x"00001f59",
         14427 => x"00001f59",
         14428 => x"00001f59",
         14429 => x"00001f59",
         14430 => x"00001f59",
         14431 => x"000021b5",
         14432 => x"0000217a",
         14433 => x"00001f59",
         14434 => x"00001f59",
         14435 => x"00001f59",
         14436 => x"00001f59",
         14437 => x"00001f59",
         14438 => x"00001f59",
         14439 => x"00001f59",
         14440 => x"00001f59",
         14441 => x"0000216d",
         14442 => x"00002162",
         14443 => x"00001f59",
         14444 => x"0000214b",
         14445 => x"00001f59",
         14446 => x"0000215b",
         14447 => x"00002151",
         14448 => x"00002144",
         14449 => x"0000321c",
         14450 => x"00003234",
         14451 => x"00003240",
         14452 => x"0000324c",
         14453 => x"00003258",
         14454 => x"00003228",
         14455 => x"00003b91",
         14456 => x"00003a7f",
         14457 => x"000038fb",
         14458 => x"00003649",
         14459 => x"00003a1b",
         14460 => x"000034d8",
         14461 => x"00003795",
         14462 => x"0000366e",
         14463 => x"000039c5",
         14464 => x"0000369d",
         14465 => x"0000370c",
         14466 => x"00003924",
         14467 => x"000034d8",
         14468 => x"000038fb",
         14469 => x"00003805",
         14470 => x"00003795",
         14471 => x"000034d8",
         14472 => x"000034d8",
         14473 => x"0000370c",
         14474 => x"0000369d",
         14475 => x"0000366e",
         14476 => x"00003649",
         14477 => x"00004676",
         14478 => x"0000468f",
         14479 => x"000046b4",
         14480 => x"000046d5",
         14481 => x"00004636",
         14482 => x"000046fa",
         14483 => x"0000464f",
         14484 => x"0000479f",
         14485 => x"0000475c",
         14486 => x"0000475c",
         14487 => x"0000475c",
         14488 => x"0000475c",
         14489 => x"0000475c",
         14490 => x"0000475c",
         14491 => x"00004735",
         14492 => x"0000475c",
         14493 => x"0000475c",
         14494 => x"0000475c",
         14495 => x"0000475c",
         14496 => x"0000475c",
         14497 => x"0000475c",
         14498 => x"0000475c",
         14499 => x"0000475c",
         14500 => x"0000475c",
         14501 => x"0000475c",
         14502 => x"0000475c",
         14503 => x"0000475c",
         14504 => x"0000475c",
         14505 => x"0000475c",
         14506 => x"0000475c",
         14507 => x"0000475c",
         14508 => x"0000475c",
         14509 => x"0000475c",
         14510 => x"0000475c",
         14511 => x"0000475c",
         14512 => x"0000475c",
         14513 => x"0000475c",
         14514 => x"00004874",
         14515 => x"00004862",
         14516 => x"0000484f",
         14517 => x"0000483c",
         14518 => x"00004766",
         14519 => x"0000482a",
         14520 => x"00004817",
         14521 => x"0000477f",
         14522 => x"0000475c",
         14523 => x"0000477f",
         14524 => x"00004807",
         14525 => x"00004884",
         14526 => x"000047b0",
         14527 => x"0000478e",
         14528 => x"000047f5",
         14529 => x"000047e3",
         14530 => x"000047d1",
         14531 => x"000047c2",
         14532 => x"0000475c",
         14533 => x"00004766",
         14534 => x"00005402",
         14535 => x"00005571",
         14536 => x"00005543",
         14537 => x"0000549a",
         14538 => x"00005477",
         14539 => x"00005456",
         14540 => x"0000542c",
         14541 => x"000055fc",
         14542 => x"00005283",
         14543 => x"000055d6",
         14544 => x"000057c5",
         14545 => x"00005283",
         14546 => x"00005283",
         14547 => x"00005283",
         14548 => x"00005283",
         14549 => x"00005283",
         14550 => x"00005283",
         14551 => x"0000559f",
         14552 => x"000057ad",
         14553 => x"00005664",
         14554 => x"00005283",
         14555 => x"00005283",
         14556 => x"00005283",
         14557 => x"00005283",
         14558 => x"00005283",
         14559 => x"00005283",
         14560 => x"00005283",
         14561 => x"00005283",
         14562 => x"00005283",
         14563 => x"00005283",
         14564 => x"00005283",
         14565 => x"00005283",
         14566 => x"00005283",
         14567 => x"00005283",
         14568 => x"00005283",
         14569 => x"00005283",
         14570 => x"00005283",
         14571 => x"00005283",
         14572 => x"00005283",
         14573 => x"00005521",
         14574 => x"00005283",
         14575 => x"00005283",
         14576 => x"00005283",
         14577 => x"000054c4",
         14578 => x"000053d3",
         14579 => x"00005375",
         14580 => x"00005283",
         14581 => x"00005283",
         14582 => x"00005283",
         14583 => x"00005283",
         14584 => x"0000535a",
         14585 => x"00005283",
         14586 => x"0000533d",
         14587 => x"000059a6",
         14588 => x"0000591b",
         14589 => x"0000591b",
         14590 => x"0000591b",
         14591 => x"0000591b",
         14592 => x"0000591b",
         14593 => x"0000591b",
         14594 => x"000058f6",
         14595 => x"0000591b",
         14596 => x"0000591b",
         14597 => x"0000591b",
         14598 => x"0000591b",
         14599 => x"0000591b",
         14600 => x"0000591b",
         14601 => x"0000591b",
         14602 => x"0000591b",
         14603 => x"0000591b",
         14604 => x"0000591b",
         14605 => x"0000591b",
         14606 => x"0000591b",
         14607 => x"0000591b",
         14608 => x"0000591b",
         14609 => x"0000591b",
         14610 => x"0000591b",
         14611 => x"0000591b",
         14612 => x"0000591b",
         14613 => x"0000591b",
         14614 => x"0000591b",
         14615 => x"0000591b",
         14616 => x"0000591b",
         14617 => x"000059b8",
         14618 => x"00005a00",
         14619 => x"000059ed",
         14620 => x"000059da",
         14621 => x"000059c8",
         14622 => x"00005a8b",
         14623 => x"00005a78",
         14624 => x"00005a68",
         14625 => x"0000591b",
         14626 => x"00005a58",
         14627 => x"00005a48",
         14628 => x"00005a36",
         14629 => x"00005a24",
         14630 => x"00005a12",
         14631 => x"00005983",
         14632 => x"00005972",
         14633 => x"00005961",
         14634 => x"0000594a",
         14635 => x"0000591b",
         14636 => x"00005994",
         14637 => x"00006375",
         14638 => x"000061d1",
         14639 => x"000061d1",
         14640 => x"000061d1",
         14641 => x"000061d1",
         14642 => x"000061d1",
         14643 => x"000061d1",
         14644 => x"000061d1",
         14645 => x"000061d1",
         14646 => x"000061d1",
         14647 => x"000061d1",
         14648 => x"000061d1",
         14649 => x"000061d1",
         14650 => x"000061d1",
         14651 => x"00005ef3",
         14652 => x"000061d1",
         14653 => x"000061d1",
         14654 => x"000061d1",
         14655 => x"000061d1",
         14656 => x"000061d1",
         14657 => x"000061d1",
         14658 => x"000063bf",
         14659 => x"000061d1",
         14660 => x"000061d1",
         14661 => x"0000634a",
         14662 => x"000061d1",
         14663 => x"00006361",
         14664 => x"00005ed2",
         14665 => x"00006333",
         14666 => x"0000df2e",
         14667 => x"0000df1b",
         14668 => x"0000df0f",
         14669 => x"0000df04",
         14670 => x"0000def9",
         14671 => x"0000deee",
         14672 => x"0000dee3",
         14673 => x"0000ded7",
         14674 => x"0000dec9",
         14675 => x"00000e01",
         14676 => x"00000bfd",
         14677 => x"00000bfd",
         14678 => x"00000f49",
         14679 => x"00000bfd",
         14680 => x"00000bfd",
         14681 => x"00000bfd",
         14682 => x"00000bfd",
         14683 => x"00000bfd",
         14684 => x"00000bfd",
         14685 => x"00000bfd",
         14686 => x"00000dfd",
         14687 => x"00000bfd",
         14688 => x"00000f7f",
         14689 => x"00000f0d",
         14690 => x"00000bfd",
         14691 => x"00000bfd",
         14692 => x"00000bfd",
         14693 => x"00000bfd",
         14694 => x"00000bfd",
         14695 => x"00000bfd",
         14696 => x"00000bfd",
         14697 => x"00000bfd",
         14698 => x"00000bfd",
         14699 => x"00000bfd",
         14700 => x"00000bfd",
         14701 => x"00000bfd",
         14702 => x"00000bfd",
         14703 => x"00000bfd",
         14704 => x"00000bfd",
         14705 => x"00000bfd",
         14706 => x"00000bfd",
         14707 => x"00000bfd",
         14708 => x"00000bfd",
         14709 => x"00000bfd",
         14710 => x"00000bfd",
         14711 => x"00000bfd",
         14712 => x"00000bfd",
         14713 => x"00000bfd",
         14714 => x"00000bfd",
         14715 => x"00000bfd",
         14716 => x"00000bfd",
         14717 => x"00000bfd",
         14718 => x"00000bfd",
         14719 => x"00000bfd",
         14720 => x"00000bfd",
         14721 => x"00000bfd",
         14722 => x"00000bfd",
         14723 => x"00000bfd",
         14724 => x"00000bfd",
         14725 => x"00000bfd",
         14726 => x"00000f1d",
         14727 => x"00000bfd",
         14728 => x"00000bfd",
         14729 => x"00000bfd",
         14730 => x"00000bfd",
         14731 => x"00000e17",
         14732 => x"00000bfd",
         14733 => x"00000bfd",
         14734 => x"00000bfd",
         14735 => x"00000bfd",
         14736 => x"00000bfd",
         14737 => x"00000bfd",
         14738 => x"00000bfd",
         14739 => x"00000bfd",
         14740 => x"00000bfd",
         14741 => x"00000bfd",
         14742 => x"00000e2b",
         14743 => x"00000ee1",
         14744 => x"00000eb8",
         14745 => x"00000eb8",
         14746 => x"00000eb8",
         14747 => x"00000bfd",
         14748 => x"00000ee1",
         14749 => x"00000bfd",
         14750 => x"00000bfd",
         14751 => x"00000eff",
         14752 => x"00000bfd",
         14753 => x"00000bfd",
         14754 => x"00000c16",
         14755 => x"00000e0f",
         14756 => x"00000bfd",
         14757 => x"00000bfd",
         14758 => x"00000f58",
         14759 => x"00000bfd",
         14760 => x"00000c18",
         14761 => x"00000bfd",
         14762 => x"00000bfd",
         14763 => x"00000e17",
         14764 => x"64696e69",
         14765 => x"74000000",
         14766 => x"64696f63",
         14767 => x"746c0000",
         14768 => x"66696e69",
         14769 => x"74000000",
         14770 => x"666c6f61",
         14771 => x"64000000",
         14772 => x"66657865",
         14773 => x"63000000",
         14774 => x"6d636c65",
         14775 => x"61720000",
         14776 => x"6d636f70",
         14777 => x"79000000",
         14778 => x"6d646966",
         14779 => x"66000000",
         14780 => x"6d64756d",
         14781 => x"70000000",
         14782 => x"6d656200",
         14783 => x"6d656800",
         14784 => x"6d657700",
         14785 => x"68696400",
         14786 => x"68696500",
         14787 => x"68666400",
         14788 => x"68666500",
         14789 => x"63616c6c",
         14790 => x"00000000",
         14791 => x"6a6d7000",
         14792 => x"72657374",
         14793 => x"61727400",
         14794 => x"72657365",
         14795 => x"74000000",
         14796 => x"696e666f",
         14797 => x"00000000",
         14798 => x"74657374",
         14799 => x"00000000",
         14800 => x"636c7300",
         14801 => x"7a383000",
         14802 => x"74626173",
         14803 => x"69630000",
         14804 => x"6d626173",
         14805 => x"69630000",
         14806 => x"6b696c6f",
         14807 => x"00000000",
         14808 => x"65640000",
         14809 => x"556e6b6e",
         14810 => x"6f776e20",
         14811 => x"6572726f",
         14812 => x"722e0000",
         14813 => x"50617261",
         14814 => x"6d657465",
         14815 => x"72732069",
         14816 => x"6e636f72",
         14817 => x"72656374",
         14818 => x"2e000000",
         14819 => x"546f6f20",
         14820 => x"6d616e79",
         14821 => x"206f7065",
         14822 => x"6e206669",
         14823 => x"6c65732e",
         14824 => x"00000000",
         14825 => x"496e7375",
         14826 => x"66666963",
         14827 => x"69656e74",
         14828 => x"206d656d",
         14829 => x"6f72792e",
         14830 => x"00000000",
         14831 => x"46696c65",
         14832 => x"20697320",
         14833 => x"6c6f636b",
         14834 => x"65642e00",
         14835 => x"54696d65",
         14836 => x"6f75742c",
         14837 => x"206f7065",
         14838 => x"72617469",
         14839 => x"6f6e2063",
         14840 => x"616e6365",
         14841 => x"6c6c6564",
         14842 => x"2e000000",
         14843 => x"466f726d",
         14844 => x"61742061",
         14845 => x"626f7274",
         14846 => x"65642e00",
         14847 => x"4e6f2063",
         14848 => x"6f6d7061",
         14849 => x"7469626c",
         14850 => x"65206669",
         14851 => x"6c657379",
         14852 => x"7374656d",
         14853 => x"20666f75",
         14854 => x"6e64206f",
         14855 => x"6e206469",
         14856 => x"736b2e00",
         14857 => x"4469736b",
         14858 => x"206e6f74",
         14859 => x"20656e61",
         14860 => x"626c6564",
         14861 => x"2e000000",
         14862 => x"44726976",
         14863 => x"65206e75",
         14864 => x"6d626572",
         14865 => x"20697320",
         14866 => x"696e7661",
         14867 => x"6c69642e",
         14868 => x"00000000",
         14869 => x"53442069",
         14870 => x"73207772",
         14871 => x"69746520",
         14872 => x"70726f74",
         14873 => x"65637465",
         14874 => x"642e0000",
         14875 => x"46696c65",
         14876 => x"2068616e",
         14877 => x"646c6520",
         14878 => x"696e7661",
         14879 => x"6c69642e",
         14880 => x"00000000",
         14881 => x"46696c65",
         14882 => x"20616c72",
         14883 => x"65616479",
         14884 => x"20657869",
         14885 => x"7374732e",
         14886 => x"00000000",
         14887 => x"41636365",
         14888 => x"73732064",
         14889 => x"656e6965",
         14890 => x"642e0000",
         14891 => x"496e7661",
         14892 => x"6c696420",
         14893 => x"66696c65",
         14894 => x"6e616d65",
         14895 => x"2e000000",
         14896 => x"4e6f2070",
         14897 => x"61746820",
         14898 => x"666f756e",
         14899 => x"642e0000",
         14900 => x"4e6f2066",
         14901 => x"696c6520",
         14902 => x"666f756e",
         14903 => x"642e0000",
         14904 => x"4469736b",
         14905 => x"206e6f74",
         14906 => x"20726561",
         14907 => x"64792e00",
         14908 => x"496e7465",
         14909 => x"726e616c",
         14910 => x"20657272",
         14911 => x"6f722e00",
         14912 => x"4469736b",
         14913 => x"20457272",
         14914 => x"6f720000",
         14915 => x"53756363",
         14916 => x"6573732e",
         14917 => x"00000000",
         14918 => x"0a256c75",
         14919 => x"20627974",
         14920 => x"65732025",
         14921 => x"73206174",
         14922 => x"20256c75",
         14923 => x"20627974",
         14924 => x"65732f73",
         14925 => x"65632e0a",
         14926 => x"00000000",
         14927 => x"72656164",
         14928 => x"00000000",
         14929 => x"2530386c",
         14930 => x"58000000",
         14931 => x"3a202000",
         14932 => x"25303258",
         14933 => x"00000000",
         14934 => x"207c0000",
         14935 => x"7c000000",
         14936 => x"20200000",
         14937 => x"25303458",
         14938 => x"00000000",
         14939 => x"20202020",
         14940 => x"20202020",
         14941 => x"00000000",
         14942 => x"7a4f5300",
         14943 => x"2a2a2025",
         14944 => x"73202800",
         14945 => x"31312f31",
         14946 => x"322f3230",
         14947 => x"32300000",
         14948 => x"76312e31",
         14949 => x"64000000",
         14950 => x"205a5055",
         14951 => x"2c207265",
         14952 => x"76202530",
         14953 => x"32782920",
         14954 => x"25732025",
         14955 => x"73202a2a",
         14956 => x"0a0a0000",
         14957 => x"5a505520",
         14958 => x"496e7465",
         14959 => x"72727570",
         14960 => x"74204861",
         14961 => x"6e646c65",
         14962 => x"72000000",
         14963 => x"55415254",
         14964 => x"31205458",
         14965 => x"20696e74",
         14966 => x"65727275",
         14967 => x"70740000",
         14968 => x"55415254",
         14969 => x"31205258",
         14970 => x"20696e74",
         14971 => x"65727275",
         14972 => x"70740000",
         14973 => x"55415254",
         14974 => x"30205458",
         14975 => x"20696e74",
         14976 => x"65727275",
         14977 => x"70740000",
         14978 => x"55415254",
         14979 => x"30205258",
         14980 => x"20696e74",
         14981 => x"65727275",
         14982 => x"70740000",
         14983 => x"494f4354",
         14984 => x"4c205752",
         14985 => x"20696e74",
         14986 => x"65727275",
         14987 => x"70740000",
         14988 => x"494f4354",
         14989 => x"4c205244",
         14990 => x"20696e74",
         14991 => x"65727275",
         14992 => x"70740000",
         14993 => x"50533220",
         14994 => x"696e7465",
         14995 => x"72727570",
         14996 => x"74000000",
         14997 => x"54696d65",
         14998 => x"7220696e",
         14999 => x"74657272",
         15000 => x"75707400",
         15001 => x"53657474",
         15002 => x"696e6720",
         15003 => x"75702074",
         15004 => x"696d6572",
         15005 => x"2e2e2e00",
         15006 => x"456e6162",
         15007 => x"6c696e67",
         15008 => x"2074696d",
         15009 => x"65722e2e",
         15010 => x"2e000000",
         15011 => x"6175746f",
         15012 => x"65786563",
         15013 => x"2e626174",
         15014 => x"00000000",
         15015 => x"7a4f535f",
         15016 => x"7a70752e",
         15017 => x"68737400",
         15018 => x"4661696c",
         15019 => x"65642074",
         15020 => x"6f20696e",
         15021 => x"69746961",
         15022 => x"6c697365",
         15023 => x"20736420",
         15024 => x"63617264",
         15025 => x"20302c20",
         15026 => x"706c6561",
         15027 => x"73652069",
         15028 => x"6e697420",
         15029 => x"6d616e75",
         15030 => x"616c6c79",
         15031 => x"2e000000",
         15032 => x"2a200000",
         15033 => x"25643a5c",
         15034 => x"25730000",
         15035 => x"4469736b",
         15036 => x"20696e69",
         15037 => x"7469616c",
         15038 => x"69736564",
         15039 => x"00000000",
         15040 => x"303a0000",
         15041 => x"42616420",
         15042 => x"636f6d6d",
         15043 => x"616e642e",
         15044 => x"00000000",
         15045 => x"5a505500",
         15046 => x"62696e00",
         15047 => x"25643a5c",
         15048 => x"25735c25",
         15049 => x"732e2573",
         15050 => x"00000000",
         15051 => x"436f6c64",
         15052 => x"20726562",
         15053 => x"6f6f7469",
         15054 => x"6e672e2e",
         15055 => x"2e000000",
         15056 => x"52657374",
         15057 => x"61727469",
         15058 => x"6e672061",
         15059 => x"70706c69",
         15060 => x"63617469",
         15061 => x"6f6e2e2e",
         15062 => x"2e000000",
         15063 => x"43616c6c",
         15064 => x"696e6720",
         15065 => x"636f6465",
         15066 => x"20402025",
         15067 => x"30386c78",
         15068 => x"202e2e2e",
         15069 => x"0a000000",
         15070 => x"43616c6c",
         15071 => x"20726574",
         15072 => x"75726e65",
         15073 => x"6420636f",
         15074 => x"64652028",
         15075 => x"2564292e",
         15076 => x"0a000000",
         15077 => x"45786563",
         15078 => x"7574696e",
         15079 => x"6720636f",
         15080 => x"64652040",
         15081 => x"20253038",
         15082 => x"6c78202e",
         15083 => x"2e2e0a00",
         15084 => x"2530386c",
         15085 => x"58202530",
         15086 => x"386c582d",
         15087 => x"00000000",
         15088 => x"2530386c",
         15089 => x"58202530",
         15090 => x"34582d00",
         15091 => x"436f6d70",
         15092 => x"6172696e",
         15093 => x"672e2e2e",
         15094 => x"00000000",
         15095 => x"2530386c",
         15096 => x"78282530",
         15097 => x"3878292d",
         15098 => x"3e253038",
         15099 => x"6c782825",
         15100 => x"30387829",
         15101 => x"0a000000",
         15102 => x"436f7079",
         15103 => x"696e672e",
         15104 => x"2e2e0000",
         15105 => x"2530386c",
         15106 => x"58202530",
         15107 => x"32582d00",
         15108 => x"436c6561",
         15109 => x"72696e67",
         15110 => x"2e2e2e2e",
         15111 => x"00000000",
         15112 => x"44756d70",
         15113 => x"204d656d",
         15114 => x"6f727900",
         15115 => x"0a436f6d",
         15116 => x"706c6574",
         15117 => x"652e0000",
         15118 => x"25643a5c",
         15119 => x"25735c25",
         15120 => x"73000000",
         15121 => x"4d656d6f",
         15122 => x"72792065",
         15123 => x"78686175",
         15124 => x"73746564",
         15125 => x"2c206361",
         15126 => x"6e6e6f74",
         15127 => x"2070726f",
         15128 => x"63657373",
         15129 => x"20636f6d",
         15130 => x"6d616e64",
         15131 => x"2e000000",
         15132 => x"3f3f3f00",
         15133 => x"25642f25",
         15134 => x"642f2564",
         15135 => x"2025643a",
         15136 => x"25643a25",
         15137 => x"642e2564",
         15138 => x"25640a00",
         15139 => x"536f4320",
         15140 => x"436f6e66",
         15141 => x"69677572",
         15142 => x"6174696f",
         15143 => x"6e000000",
         15144 => x"3a0a4465",
         15145 => x"76696365",
         15146 => x"7320696d",
         15147 => x"706c656d",
         15148 => x"656e7465",
         15149 => x"643a0000",
         15150 => x"41646472",
         15151 => x"65737365",
         15152 => x"733a0000",
         15153 => x"20202020",
         15154 => x"43505520",
         15155 => x"52657365",
         15156 => x"74205665",
         15157 => x"63746f72",
         15158 => x"20416464",
         15159 => x"72657373",
         15160 => x"203d2025",
         15161 => x"3038580a",
         15162 => x"00000000",
         15163 => x"20202020",
         15164 => x"43505520",
         15165 => x"4d656d6f",
         15166 => x"72792053",
         15167 => x"74617274",
         15168 => x"20416464",
         15169 => x"72657373",
         15170 => x"203d2025",
         15171 => x"3038580a",
         15172 => x"00000000",
         15173 => x"20202020",
         15174 => x"53746163",
         15175 => x"6b205374",
         15176 => x"61727420",
         15177 => x"41646472",
         15178 => x"65737320",
         15179 => x"20202020",
         15180 => x"203d2025",
         15181 => x"3038580a",
         15182 => x"00000000",
         15183 => x"4d697363",
         15184 => x"3a000000",
         15185 => x"20202020",
         15186 => x"5a505520",
         15187 => x"49642020",
         15188 => x"20202020",
         15189 => x"20202020",
         15190 => x"20202020",
         15191 => x"20202020",
         15192 => x"203d2025",
         15193 => x"3034580a",
         15194 => x"00000000",
         15195 => x"20202020",
         15196 => x"53797374",
         15197 => x"656d2043",
         15198 => x"6c6f636b",
         15199 => x"20467265",
         15200 => x"71202020",
         15201 => x"20202020",
         15202 => x"203d2025",
         15203 => x"642e2530",
         15204 => x"34644d48",
         15205 => x"7a0a0000",
         15206 => x"20202020",
         15207 => x"57697368",
         15208 => x"626f6e65",
         15209 => x"20534452",
         15210 => x"414d2043",
         15211 => x"6c6f636b",
         15212 => x"20467265",
         15213 => x"713d2025",
         15214 => x"642e2530",
         15215 => x"34644d48",
         15216 => x"7a0a0000",
         15217 => x"20202020",
         15218 => x"53445241",
         15219 => x"4d20436c",
         15220 => x"6f636b20",
         15221 => x"46726571",
         15222 => x"20202020",
         15223 => x"20202020",
         15224 => x"203d2025",
         15225 => x"642e2530",
         15226 => x"34644d48",
         15227 => x"7a0a0000",
         15228 => x"20202020",
         15229 => x"53504900",
         15230 => x"20202020",
         15231 => x"50533200",
         15232 => x"20202020",
         15233 => x"494f4354",
         15234 => x"4c000000",
         15235 => x"20202020",
         15236 => x"57422049",
         15237 => x"32430000",
         15238 => x"20202020",
         15239 => x"57495348",
         15240 => x"424f4e45",
         15241 => x"20425553",
         15242 => x"00000000",
         15243 => x"20202020",
         15244 => x"494e5452",
         15245 => x"20435452",
         15246 => x"4c202843",
         15247 => x"68616e6e",
         15248 => x"656c733d",
         15249 => x"25303264",
         15250 => x"292e0a00",
         15251 => x"20202020",
         15252 => x"54494d45",
         15253 => x"52312020",
         15254 => x"20202854",
         15255 => x"696d6572",
         15256 => x"7320203d",
         15257 => x"25303264",
         15258 => x"292e0a00",
         15259 => x"20202020",
         15260 => x"53442043",
         15261 => x"41524420",
         15262 => x"20202844",
         15263 => x"65766963",
         15264 => x"6573203d",
         15265 => x"25303264",
         15266 => x"292e0a00",
         15267 => x"20202020",
         15268 => x"52414d20",
         15269 => x"20202020",
         15270 => x"20202825",
         15271 => x"3038583a",
         15272 => x"25303858",
         15273 => x"292e0a00",
         15274 => x"20202020",
         15275 => x"4252414d",
         15276 => x"20202020",
         15277 => x"20202825",
         15278 => x"3038583a",
         15279 => x"25303858",
         15280 => x"292e0a00",
         15281 => x"20202020",
         15282 => x"494e534e",
         15283 => x"20425241",
         15284 => x"4d202825",
         15285 => x"3038583a",
         15286 => x"25303858",
         15287 => x"292e0a00",
         15288 => x"20202020",
         15289 => x"53445241",
         15290 => x"4d202020",
         15291 => x"20202825",
         15292 => x"3038583a",
         15293 => x"25303858",
         15294 => x"292e0a00",
         15295 => x"20202020",
         15296 => x"57422053",
         15297 => x"4452414d",
         15298 => x"20202825",
         15299 => x"3038583a",
         15300 => x"25303858",
         15301 => x"292e0a00",
         15302 => x"20286672",
         15303 => x"6f6d2053",
         15304 => x"6f432063",
         15305 => x"6f6e6669",
         15306 => x"67290000",
         15307 => x"556e6b6e",
         15308 => x"6f776e00",
         15309 => x"45564f6d",
         15310 => x"00000000",
         15311 => x"536d616c",
         15312 => x"6c000000",
         15313 => x"4d656469",
         15314 => x"756d0000",
         15315 => x"466c6578",
         15316 => x"00000000",
         15317 => x"45564f00",
         15318 => x"0000f0b4",
         15319 => x"01000000",
         15320 => x"00000002",
         15321 => x"0000f0b0",
         15322 => x"01000000",
         15323 => x"00000003",
         15324 => x"0000f0ac",
         15325 => x"01000000",
         15326 => x"00000004",
         15327 => x"0000f0a8",
         15328 => x"01000000",
         15329 => x"00000005",
         15330 => x"0000f0a4",
         15331 => x"01000000",
         15332 => x"00000006",
         15333 => x"0000f0a0",
         15334 => x"01000000",
         15335 => x"00000007",
         15336 => x"0000f09c",
         15337 => x"01000000",
         15338 => x"00000001",
         15339 => x"0000f098",
         15340 => x"01000000",
         15341 => x"00000008",
         15342 => x"0000f094",
         15343 => x"01000000",
         15344 => x"0000000b",
         15345 => x"0000f090",
         15346 => x"01000000",
         15347 => x"00000009",
         15348 => x"0000f08c",
         15349 => x"01000000",
         15350 => x"0000000a",
         15351 => x"0000f088",
         15352 => x"04000000",
         15353 => x"0000000d",
         15354 => x"0000f084",
         15355 => x"04000000",
         15356 => x"0000000c",
         15357 => x"0000f080",
         15358 => x"04000000",
         15359 => x"0000000e",
         15360 => x"0000f07c",
         15361 => x"03000000",
         15362 => x"0000000f",
         15363 => x"0000f078",
         15364 => x"04000000",
         15365 => x"0000000f",
         15366 => x"0000f074",
         15367 => x"04000000",
         15368 => x"00000010",
         15369 => x"0000f070",
         15370 => x"04000000",
         15371 => x"00000011",
         15372 => x"0000f06c",
         15373 => x"03000000",
         15374 => x"00000012",
         15375 => x"0000f068",
         15376 => x"03000000",
         15377 => x"00000013",
         15378 => x"0000f064",
         15379 => x"03000000",
         15380 => x"00000014",
         15381 => x"0000f060",
         15382 => x"03000000",
         15383 => x"00000015",
         15384 => x"1b5b4400",
         15385 => x"1b5b4300",
         15386 => x"1b5b4200",
         15387 => x"1b5b4100",
         15388 => x"1b5b367e",
         15389 => x"1b5b357e",
         15390 => x"1b5b347e",
         15391 => x"1b304600",
         15392 => x"1b5b337e",
         15393 => x"1b5b327e",
         15394 => x"1b5b317e",
         15395 => x"10000000",
         15396 => x"0e000000",
         15397 => x"0d000000",
         15398 => x"0b000000",
         15399 => x"08000000",
         15400 => x"06000000",
         15401 => x"05000000",
         15402 => x"04000000",
         15403 => x"03000000",
         15404 => x"02000000",
         15405 => x"01000000",
         15406 => x"43616e6e",
         15407 => x"6f74206f",
         15408 => x"70656e2f",
         15409 => x"63726561",
         15410 => x"74652068",
         15411 => x"6973746f",
         15412 => x"72792066",
         15413 => x"696c652c",
         15414 => x"20646973",
         15415 => x"61626c69",
         15416 => x"6e672e00",
         15417 => x"68697374",
         15418 => x"6f727900",
         15419 => x"68697374",
         15420 => x"00000000",
         15421 => x"21000000",
         15422 => x"2530366c",
         15423 => x"75202025",
         15424 => x"730a0000",
         15425 => x"4661696c",
         15426 => x"65642074",
         15427 => x"6f207265",
         15428 => x"73657420",
         15429 => x"74686520",
         15430 => x"68697374",
         15431 => x"6f727920",
         15432 => x"66696c65",
         15433 => x"20746f20",
         15434 => x"454f462e",
         15435 => x"00000000",
         15436 => x"3e25730a",
         15437 => x"00000000",
         15438 => x"1b5b317e",
         15439 => x"00000000",
         15440 => x"1b5b4100",
         15441 => x"1b5b4200",
         15442 => x"1b5b4300",
         15443 => x"1b5b4400",
         15444 => x"1b5b3130",
         15445 => x"7e000000",
         15446 => x"1b5b3131",
         15447 => x"7e000000",
         15448 => x"1b5b3132",
         15449 => x"7e000000",
         15450 => x"1b5b3133",
         15451 => x"7e000000",
         15452 => x"1b5b3134",
         15453 => x"7e000000",
         15454 => x"1b5b3135",
         15455 => x"7e000000",
         15456 => x"1b5b3137",
         15457 => x"7e000000",
         15458 => x"1b5b3138",
         15459 => x"7e000000",
         15460 => x"1b5b3139",
         15461 => x"7e000000",
         15462 => x"1b5b3230",
         15463 => x"7e000000",
         15464 => x"1b5b327e",
         15465 => x"00000000",
         15466 => x"1b5b337e",
         15467 => x"00000000",
         15468 => x"1b5b4600",
         15469 => x"1b5b357e",
         15470 => x"00000000",
         15471 => x"1b5b367e",
         15472 => x"00000000",
         15473 => x"583a2564",
         15474 => x"2c25642c",
         15475 => x"25642c25",
         15476 => x"642c2564",
         15477 => x"2c25643a",
         15478 => x"25303278",
         15479 => x"00000000",
         15480 => x"443a2564",
         15481 => x"2d25642d",
         15482 => x"25643a25",
         15483 => x"633a2564",
         15484 => x"2c25642c",
         15485 => x"25643a00",
         15486 => x"25642c00",
         15487 => x"4b3a2564",
         15488 => x"3a000000",
         15489 => x"25303278",
         15490 => x"2c000000",
         15491 => x"25635b25",
         15492 => x"643b2564",
         15493 => x"52000000",
         15494 => x"5265706f",
         15495 => x"72742043",
         15496 => x"7572736f",
         15497 => x"723a0000",
         15498 => x"55703a25",
         15499 => x"30327820",
         15500 => x"25303278",
         15501 => x"00000000",
         15502 => x"44773a25",
         15503 => x"30327820",
         15504 => x"25303278",
         15505 => x"00000000",
         15506 => x"48643a25",
         15507 => x"30327820",
         15508 => x"00000000",
         15509 => x"42616420",
         15510 => x"65786974",
         15511 => x"2c205344",
         15512 => x"20496e69",
         15513 => x"74000000",
         15514 => x"42616420",
         15515 => x"65786974",
         15516 => x"2c205344",
         15517 => x"20526561",
         15518 => x"64000000",
         15519 => x"42616420",
         15520 => x"65786974",
         15521 => x"2c205344",
         15522 => x"20577269",
         15523 => x"74650000",
         15524 => x"4e6f2074",
         15525 => x"65737420",
         15526 => x"64656669",
         15527 => x"6e65642e",
         15528 => x"00000000",
         15529 => x"53440000",
         15530 => x"222a3a3c",
         15531 => x"3e3f7c7f",
         15532 => x"00000000",
         15533 => x"2b2c3b3d",
         15534 => x"5b5d0000",
         15535 => x"46415400",
         15536 => x"46415433",
         15537 => x"32000000",
         15538 => x"ebfe904d",
         15539 => x"53444f53",
         15540 => x"352e3000",
         15541 => x"4e4f204e",
         15542 => x"414d4520",
         15543 => x"20202046",
         15544 => x"41542020",
         15545 => x"20202000",
         15546 => x"4e4f204e",
         15547 => x"414d4520",
         15548 => x"20202046",
         15549 => x"41543332",
         15550 => x"20202000",
         15551 => x"0000f2a4",
         15552 => x"00000000",
         15553 => x"00000000",
         15554 => x"00000000",
         15555 => x"01030507",
         15556 => x"090e1012",
         15557 => x"1416181c",
         15558 => x"1e000000",
         15559 => x"809a4541",
         15560 => x"8e418f80",
         15561 => x"45454549",
         15562 => x"49498e8f",
         15563 => x"9092924f",
         15564 => x"994f5555",
         15565 => x"59999a9b",
         15566 => x"9c9d9e9f",
         15567 => x"41494f55",
         15568 => x"a5a5a6a7",
         15569 => x"a8a9aaab",
         15570 => x"acadaeaf",
         15571 => x"b0b1b2b3",
         15572 => x"b4b5b6b7",
         15573 => x"b8b9babb",
         15574 => x"bcbdbebf",
         15575 => x"c0c1c2c3",
         15576 => x"c4c5c6c7",
         15577 => x"c8c9cacb",
         15578 => x"cccdcecf",
         15579 => x"d0d1d2d3",
         15580 => x"d4d5d6d7",
         15581 => x"d8d9dadb",
         15582 => x"dcdddedf",
         15583 => x"e0e1e2e3",
         15584 => x"e4e5e6e7",
         15585 => x"e8e9eaeb",
         15586 => x"ecedeeef",
         15587 => x"f0f1f2f3",
         15588 => x"f4f5f6f7",
         15589 => x"f8f9fafb",
         15590 => x"fcfdfeff",
         15591 => x"2b2e2c3b",
         15592 => x"3d5b5d2f",
         15593 => x"5c222a3a",
         15594 => x"3c3e3f7c",
         15595 => x"7f000000",
         15596 => x"00010004",
         15597 => x"00100040",
         15598 => x"01000200",
         15599 => x"00000000",
         15600 => x"00010002",
         15601 => x"00040008",
         15602 => x"00100020",
         15603 => x"00000000",
         15604 => x"00c700fc",
         15605 => x"00e900e2",
         15606 => x"00e400e0",
         15607 => x"00e500e7",
         15608 => x"00ea00eb",
         15609 => x"00e800ef",
         15610 => x"00ee00ec",
         15611 => x"00c400c5",
         15612 => x"00c900e6",
         15613 => x"00c600f4",
         15614 => x"00f600f2",
         15615 => x"00fb00f9",
         15616 => x"00ff00d6",
         15617 => x"00dc00a2",
         15618 => x"00a300a5",
         15619 => x"20a70192",
         15620 => x"00e100ed",
         15621 => x"00f300fa",
         15622 => x"00f100d1",
         15623 => x"00aa00ba",
         15624 => x"00bf2310",
         15625 => x"00ac00bd",
         15626 => x"00bc00a1",
         15627 => x"00ab00bb",
         15628 => x"25912592",
         15629 => x"25932502",
         15630 => x"25242561",
         15631 => x"25622556",
         15632 => x"25552563",
         15633 => x"25512557",
         15634 => x"255d255c",
         15635 => x"255b2510",
         15636 => x"25142534",
         15637 => x"252c251c",
         15638 => x"2500253c",
         15639 => x"255e255f",
         15640 => x"255a2554",
         15641 => x"25692566",
         15642 => x"25602550",
         15643 => x"256c2567",
         15644 => x"25682564",
         15645 => x"25652559",
         15646 => x"25582552",
         15647 => x"2553256b",
         15648 => x"256a2518",
         15649 => x"250c2588",
         15650 => x"2584258c",
         15651 => x"25902580",
         15652 => x"03b100df",
         15653 => x"039303c0",
         15654 => x"03a303c3",
         15655 => x"00b503c4",
         15656 => x"03a60398",
         15657 => x"03a903b4",
         15658 => x"221e03c6",
         15659 => x"03b52229",
         15660 => x"226100b1",
         15661 => x"22652264",
         15662 => x"23202321",
         15663 => x"00f72248",
         15664 => x"00b02219",
         15665 => x"00b7221a",
         15666 => x"207f00b2",
         15667 => x"25a000a0",
         15668 => x"0061031a",
         15669 => x"00e00317",
         15670 => x"00f80307",
         15671 => x"00ff0001",
         15672 => x"01780100",
         15673 => x"01300132",
         15674 => x"01060139",
         15675 => x"0110014a",
         15676 => x"012e0179",
         15677 => x"01060180",
         15678 => x"004d0243",
         15679 => x"01810182",
         15680 => x"01820184",
         15681 => x"01840186",
         15682 => x"01870187",
         15683 => x"0189018a",
         15684 => x"018b018b",
         15685 => x"018d018e",
         15686 => x"018f0190",
         15687 => x"01910191",
         15688 => x"01930194",
         15689 => x"01f60196",
         15690 => x"01970198",
         15691 => x"0198023d",
         15692 => x"019b019c",
         15693 => x"019d0220",
         15694 => x"019f01a0",
         15695 => x"01a001a2",
         15696 => x"01a201a4",
         15697 => x"01a401a6",
         15698 => x"01a701a7",
         15699 => x"01a901aa",
         15700 => x"01ab01ac",
         15701 => x"01ac01ae",
         15702 => x"01af01af",
         15703 => x"01b101b2",
         15704 => x"01b301b3",
         15705 => x"01b501b5",
         15706 => x"01b701b8",
         15707 => x"01b801ba",
         15708 => x"01bb01bc",
         15709 => x"01bc01be",
         15710 => x"01f701c0",
         15711 => x"01c101c2",
         15712 => x"01c301c4",
         15713 => x"01c501c4",
         15714 => x"01c701c8",
         15715 => x"01c701ca",
         15716 => x"01cb01ca",
         15717 => x"01cd0110",
         15718 => x"01dd0001",
         15719 => x"018e01de",
         15720 => x"011201f3",
         15721 => x"000301f1",
         15722 => x"01f401f4",
         15723 => x"01f80128",
         15724 => x"02220112",
         15725 => x"023a0009",
         15726 => x"2c65023b",
         15727 => x"023b023d",
         15728 => x"2c66023f",
         15729 => x"02400241",
         15730 => x"02410246",
         15731 => x"010a0253",
         15732 => x"00400181",
         15733 => x"01860255",
         15734 => x"0189018a",
         15735 => x"0258018f",
         15736 => x"025a0190",
         15737 => x"025c025d",
         15738 => x"025e025f",
         15739 => x"01930261",
         15740 => x"02620194",
         15741 => x"02640265",
         15742 => x"02660267",
         15743 => x"01970196",
         15744 => x"026a2c62",
         15745 => x"026c026d",
         15746 => x"026e019c",
         15747 => x"02700271",
         15748 => x"019d0273",
         15749 => x"0274019f",
         15750 => x"02760277",
         15751 => x"02780279",
         15752 => x"027a027b",
         15753 => x"027c2c64",
         15754 => x"027e027f",
         15755 => x"01a60281",
         15756 => x"028201a9",
         15757 => x"02840285",
         15758 => x"02860287",
         15759 => x"01ae0244",
         15760 => x"01b101b2",
         15761 => x"0245028d",
         15762 => x"028e028f",
         15763 => x"02900291",
         15764 => x"01b7037b",
         15765 => x"000303fd",
         15766 => x"03fe03ff",
         15767 => x"03ac0004",
         15768 => x"03860388",
         15769 => x"0389038a",
         15770 => x"03b10311",
         15771 => x"03c20002",
         15772 => x"03a303a3",
         15773 => x"03c40308",
         15774 => x"03cc0003",
         15775 => x"038c038e",
         15776 => x"038f03d8",
         15777 => x"011803f2",
         15778 => x"000a03f9",
         15779 => x"03f303f4",
         15780 => x"03f503f6",
         15781 => x"03f703f7",
         15782 => x"03f903fa",
         15783 => x"03fa0430",
         15784 => x"03200450",
         15785 => x"07100460",
         15786 => x"0122048a",
         15787 => x"013604c1",
         15788 => x"010e04cf",
         15789 => x"000104c0",
         15790 => x"04d00144",
         15791 => x"05610426",
         15792 => x"00000000",
         15793 => x"1d7d0001",
         15794 => x"2c631e00",
         15795 => x"01961ea0",
         15796 => x"015a1f00",
         15797 => x"06081f10",
         15798 => x"06061f20",
         15799 => x"06081f30",
         15800 => x"06081f40",
         15801 => x"06061f51",
         15802 => x"00071f59",
         15803 => x"1f521f5b",
         15804 => x"1f541f5d",
         15805 => x"1f561f5f",
         15806 => x"1f600608",
         15807 => x"1f70000e",
         15808 => x"1fba1fbb",
         15809 => x"1fc81fc9",
         15810 => x"1fca1fcb",
         15811 => x"1fda1fdb",
         15812 => x"1ff81ff9",
         15813 => x"1fea1feb",
         15814 => x"1ffa1ffb",
         15815 => x"1f800608",
         15816 => x"1f900608",
         15817 => x"1fa00608",
         15818 => x"1fb00004",
         15819 => x"1fb81fb9",
         15820 => x"1fb21fbc",
         15821 => x"1fcc0001",
         15822 => x"1fc31fd0",
         15823 => x"06021fe0",
         15824 => x"06021fe5",
         15825 => x"00011fec",
         15826 => x"1ff30001",
         15827 => x"1ffc214e",
         15828 => x"00012132",
         15829 => x"21700210",
         15830 => x"21840001",
         15831 => x"218324d0",
         15832 => x"051a2c30",
         15833 => x"042f2c60",
         15834 => x"01022c67",
         15835 => x"01062c75",
         15836 => x"01022c80",
         15837 => x"01642d00",
         15838 => x"0826ff41",
         15839 => x"031a0000",
         15840 => x"00000000",
         15841 => x"0000e6b0",
         15842 => x"01020100",
         15843 => x"00000000",
         15844 => x"00000000",
         15845 => x"0000e6b8",
         15846 => x"01040100",
         15847 => x"00000000",
         15848 => x"00000000",
         15849 => x"0000e6c0",
         15850 => x"01140300",
         15851 => x"00000000",
         15852 => x"00000000",
         15853 => x"0000e6c8",
         15854 => x"012b0300",
         15855 => x"00000000",
         15856 => x"00000000",
         15857 => x"0000e6d0",
         15858 => x"01300300",
         15859 => x"00000000",
         15860 => x"00000000",
         15861 => x"0000e6d8",
         15862 => x"013c0400",
         15863 => x"00000000",
         15864 => x"00000000",
         15865 => x"0000e6e0",
         15866 => x"013d0400",
         15867 => x"00000000",
         15868 => x"00000000",
         15869 => x"0000e6e8",
         15870 => x"013f0400",
         15871 => x"00000000",
         15872 => x"00000000",
         15873 => x"0000e6f0",
         15874 => x"01400400",
         15875 => x"00000000",
         15876 => x"00000000",
         15877 => x"0000e6f8",
         15878 => x"01410400",
         15879 => x"00000000",
         15880 => x"00000000",
         15881 => x"0000e6fc",
         15882 => x"01420400",
         15883 => x"00000000",
         15884 => x"00000000",
         15885 => x"0000e700",
         15886 => x"01430400",
         15887 => x"00000000",
         15888 => x"00000000",
         15889 => x"0000e704",
         15890 => x"01500500",
         15891 => x"00000000",
         15892 => x"00000000",
         15893 => x"0000e708",
         15894 => x"01510500",
         15895 => x"00000000",
         15896 => x"00000000",
         15897 => x"0000e70c",
         15898 => x"01540500",
         15899 => x"00000000",
         15900 => x"00000000",
         15901 => x"0000e710",
         15902 => x"01550500",
         15903 => x"00000000",
         15904 => x"00000000",
         15905 => x"0000e714",
         15906 => x"01790700",
         15907 => x"00000000",
         15908 => x"00000000",
         15909 => x"0000e71c",
         15910 => x"01780700",
         15911 => x"00000000",
         15912 => x"00000000",
         15913 => x"0000e720",
         15914 => x"01820800",
         15915 => x"00000000",
         15916 => x"00000000",
         15917 => x"0000e728",
         15918 => x"01830800",
         15919 => x"00000000",
         15920 => x"00000000",
         15921 => x"0000e730",
         15922 => x"01850800",
         15923 => x"00000000",
         15924 => x"00000000",
         15925 => x"0000e738",
         15926 => x"01870800",
         15927 => x"00000000",
         15928 => x"00000000",
         15929 => x"0000e740",
         15930 => x"01880800",
         15931 => x"00000000",
         15932 => x"00000000",
         15933 => x"0000e744",
         15934 => x"01890800",
         15935 => x"00000000",
         15936 => x"00000000",
         15937 => x"0000e748",
         15938 => x"018c0900",
         15939 => x"00000000",
         15940 => x"00000000",
         15941 => x"0000e750",
         15942 => x"018d0900",
         15943 => x"00000000",
         15944 => x"00000000",
         15945 => x"0000e758",
         15946 => x"018e0900",
         15947 => x"00000000",
         15948 => x"00000000",
         15949 => x"0000e760",
         15950 => x"018f0900",
         15951 => x"00000000",
         15952 => x"00000000",
         15953 => x"00000000",
         15954 => x"00000000",
         15955 => x"00007fff",
         15956 => x"00000000",
         15957 => x"00007fff",
         15958 => x"00010000",
         15959 => x"00007fff",
         15960 => x"00010000",
         15961 => x"00810000",
         15962 => x"01000000",
         15963 => x"017fffff",
         15964 => x"00000000",
         15965 => x"00000000",
         15966 => x"00007800",
         15967 => x"00000000",
         15968 => x"05f5e100",
         15969 => x"05f5e100",
         15970 => x"05f5e100",
         15971 => x"00000000",
         15972 => x"01010101",
         15973 => x"01010101",
         15974 => x"01011001",
         15975 => x"01000000",
         15976 => x"00000000",
         15977 => x"00000000",
         15978 => x"00000000",
         15979 => x"00000000",
         15980 => x"00000000",
         15981 => x"00000000",
         15982 => x"00000000",
         15983 => x"00000000",
         15984 => x"00000000",
         15985 => x"00000000",
         15986 => x"00000000",
         15987 => x"00000000",
         15988 => x"00000000",
         15989 => x"00000000",
         15990 => x"00000000",
         15991 => x"00000000",
         15992 => x"00000000",
         15993 => x"00000000",
         15994 => x"00000000",
         15995 => x"00000000",
         15996 => x"00000000",
         15997 => x"00000000",
         15998 => x"00000000",
         15999 => x"00000000",
         16000 => x"0000f0e4",
         16001 => x"01000000",
         16002 => x"0000f0ec",
         16003 => x"01000000",
         16004 => x"0000f0f4",
         16005 => x"02000000",
         16006 => x"0001fd80",
         16007 => x"1bfc5ffd",
         16008 => x"f03b3a0d",
         16009 => x"797a405b",
         16010 => x"5df0f0f0",
         16011 => x"71727374",
         16012 => x"75767778",
         16013 => x"696a6b6c",
         16014 => x"6d6e6f70",
         16015 => x"61626364",
         16016 => x"65666768",
         16017 => x"31323334",
         16018 => x"35363738",
         16019 => x"5cf32d20",
         16020 => x"30392c2e",
         16021 => x"f67ff3f4",
         16022 => x"f1f23f2f",
         16023 => x"08f0f0f0",
         16024 => x"f0f0f0f0",
         16025 => x"80818283",
         16026 => x"84f0f0f0",
         16027 => x"1bfc58fd",
         16028 => x"f03a3b0d",
         16029 => x"595a405b",
         16030 => x"5df0f0f0",
         16031 => x"51525354",
         16032 => x"55565758",
         16033 => x"494a4b4c",
         16034 => x"4d4e4f50",
         16035 => x"41424344",
         16036 => x"45464748",
         16037 => x"31323334",
         16038 => x"35363738",
         16039 => x"5cf32d20",
         16040 => x"30392c2e",
         16041 => x"f67ff3f4",
         16042 => x"f1f23f2f",
         16043 => x"08f0f0f0",
         16044 => x"f0f0f0f0",
         16045 => x"80818283",
         16046 => x"84f0f0f0",
         16047 => x"1bfc58fd",
         16048 => x"f02b2a0d",
         16049 => x"595a607b",
         16050 => x"7df0f0f0",
         16051 => x"51525354",
         16052 => x"55565758",
         16053 => x"494a4b4c",
         16054 => x"4d4e4f50",
         16055 => x"41424344",
         16056 => x"45464748",
         16057 => x"21222324",
         16058 => x"25262728",
         16059 => x"7c7e3d20",
         16060 => x"20293c3e",
         16061 => x"f7e2e0e1",
         16062 => x"f9f83f2f",
         16063 => x"fbf0f0f0",
         16064 => x"f0f0f0f0",
         16065 => x"85868788",
         16066 => x"89f0f0f0",
         16067 => x"1bfe1efa",
         16068 => x"f0f0f0f0",
         16069 => x"191a001b",
         16070 => x"1df0f0f0",
         16071 => x"11121314",
         16072 => x"15161718",
         16073 => x"090a0b0c",
         16074 => x"0d0e0f10",
         16075 => x"01020304",
         16076 => x"05060708",
         16077 => x"f0f0f0f0",
         16078 => x"f0f0f0f0",
         16079 => x"f01ef0f0",
         16080 => x"f01ff0f0",
         16081 => x"f0f0f0f0",
         16082 => x"f0f0f01c",
         16083 => x"f0f0f0f0",
         16084 => x"f0f0f0f0",
         16085 => x"80818283",
         16086 => x"84f0f0f0",
         16087 => x"bff0cfc9",
         16088 => x"f0b54dcd",
         16089 => x"3577d7b3",
         16090 => x"b7f0f0f0",
         16091 => x"7c704131",
         16092 => x"39a678dd",
         16093 => x"3d5d6c56",
         16094 => x"1d33d5b1",
         16095 => x"466ed948",
         16096 => x"74434c73",
         16097 => x"3f367e3b",
         16098 => x"7a1e5fa2",
         16099 => x"d39fd100",
         16100 => x"9da3d0b9",
         16101 => x"c6c5c2c1",
         16102 => x"c3c4bbbe",
         16103 => x"f0f0f0f0",
         16104 => x"f0f0f0f0",
         16105 => x"80818283",
         16106 => x"84f0f0f0",
         16107 => x"00000000",
         16108 => x"00000000",
         16109 => x"00000000",
         16110 => x"00000000",
         16111 => x"00000000",
         16112 => x"00000000",
         16113 => x"00000000",
         16114 => x"00000000",
         16115 => x"00000000",
         16116 => x"00000000",
         16117 => x"00000000",
         16118 => x"00000000",
         16119 => x"00000000",
         16120 => x"00000000",
         16121 => x"00000000",
         16122 => x"00000000",
         16123 => x"00000000",
         16124 => x"00000000",
         16125 => x"00000000",
         16126 => x"00000000",
         16127 => x"00000000",
         16128 => x"00000000",
         16129 => x"00000000",
         16130 => x"00000000",
         16131 => x"00000000",
         16132 => x"00010000",
         16133 => x"00000000",
         16134 => x"f8000000",
         16135 => x"0000f138",
         16136 => x"f3000000",
         16137 => x"0000f140",
         16138 => x"f4000000",
         16139 => x"0000f144",
         16140 => x"f1000000",
         16141 => x"0000f148",
         16142 => x"f2000000",
         16143 => x"0000f14c",
         16144 => x"80000000",
         16145 => x"0000f150",
         16146 => x"81000000",
         16147 => x"0000f158",
         16148 => x"82000000",
         16149 => x"0000f160",
         16150 => x"83000000",
         16151 => x"0000f168",
         16152 => x"84000000",
         16153 => x"0000f170",
         16154 => x"85000000",
         16155 => x"0000f178",
         16156 => x"86000000",
         16157 => x"0000f180",
         16158 => x"87000000",
         16159 => x"0000f188",
         16160 => x"88000000",
         16161 => x"0000f190",
         16162 => x"89000000",
         16163 => x"0000f198",
         16164 => x"f6000000",
         16165 => x"0000f1a0",
         16166 => x"7f000000",
         16167 => x"0000f1a8",
         16168 => x"f9000000",
         16169 => x"0000f1b0",
         16170 => x"e0000000",
         16171 => x"0000f1b4",
         16172 => x"e1000000",
         16173 => x"0000f1bc",
         16174 => x"71000000",
         16175 => x"00000000",
         16176 => x"00000000",
         16177 => x"00000000",
         16178 => x"00000000",
         16179 => x"00000000",
         16180 => x"00000000",
         16181 => x"00000000",
         16182 => x"00000000",
         16183 => x"00000000",
         16184 => x"00000000",
         16185 => x"00000000",
         16186 => x"00000000",
         16187 => x"00000000",
         16188 => x"00000000",
         16189 => x"00000000",
         16190 => x"00000000",
         16191 => x"00000000",
         16192 => x"00000000",
         16193 => x"00000000",
         16194 => x"00000000",
         16195 => x"00000000",
         16196 => x"00000000",
         16197 => x"00000000",
         16198 => x"00000000",
         16199 => x"00000000",
         16200 => x"00000000",
         16201 => x"00000000",
         16202 => x"00000000",
         16203 => x"00000000",
         16204 => x"00000000",
         16205 => x"00000000",
         16206 => x"00000000",
         16207 => x"00000000",
         16208 => x"00000000",
         16209 => x"00000000",
         16210 => x"00000000",
         16211 => x"00000000",
         16212 => x"00000000",
         16213 => x"00000000",
         16214 => x"00000000",
         16215 => x"00000000",
         16216 => x"00000000",
         16217 => x"00000000",
         16218 => x"00000000",
         16219 => x"00000000",
         16220 => x"00000000",
         16221 => x"00000000",
         16222 => x"00000000",
         16223 => x"00000000",
         16224 => x"00000000",
         16225 => x"00000000",
         16226 => x"00000000",
         16227 => x"00000000",
         16228 => x"00000000",
         16229 => x"00000000",
         16230 => x"00000000",
         16231 => x"00000000",
         16232 => x"00000000",
         16233 => x"00000000",
         16234 => x"00000000",
         16235 => x"00000000",
         16236 => x"00000000",
         16237 => x"00000000",
         16238 => x"00000000",
         16239 => x"00000000",
         16240 => x"00000000",
         16241 => x"00000000",
         16242 => x"00000000",
         16243 => x"00000000",
         16244 => x"00000000",
         16245 => x"00000000",
         16246 => x"00000000",
         16247 => x"00000000",
         16248 => x"00000000",
         16249 => x"00000000",
         16250 => x"00000000",
         16251 => x"00000000",
         16252 => x"00000000",
         16253 => x"00000000",
         16254 => x"00000000",
         16255 => x"00000000",
         16256 => x"00000000",
         16257 => x"00000000",
         16258 => x"00000000",
         16259 => x"00000000",
         16260 => x"00000000",
         16261 => x"00000000",
         16262 => x"00000000",
         16263 => x"00000000",
         16264 => x"00000000",
         16265 => x"00000000",
         16266 => x"00000000",
         16267 => x"00000000",
         16268 => x"00000000",
         16269 => x"00000000",
         16270 => x"00000000",
         16271 => x"00000000",
         16272 => x"00000000",
         16273 => x"00000000",
         16274 => x"00000000",
         16275 => x"00000000",
         16276 => x"00000000",
         16277 => x"00000000",
         16278 => x"00000000",
         16279 => x"00000000",
         16280 => x"00000000",
         16281 => x"00000000",
         16282 => x"00000000",
         16283 => x"00000000",
         16284 => x"00000000",
         16285 => x"00000000",
         16286 => x"00000000",
         16287 => x"00000000",
         16288 => x"00000000",
         16289 => x"00000000",
         16290 => x"00000000",
         16291 => x"00000000",
         16292 => x"00000000",
         16293 => x"00000000",
         16294 => x"00000000",
         16295 => x"00000000",
         16296 => x"00000000",
         16297 => x"00000000",
         16298 => x"00000000",
         16299 => x"00000000",
         16300 => x"00000000",
         16301 => x"00000000",
         16302 => x"00000000",
         16303 => x"00000000",
         16304 => x"00000000",
         16305 => x"00000000",
         16306 => x"00000000",
         16307 => x"00000000",
         16308 => x"00000000",
         16309 => x"00000000",
         16310 => x"00000000",
         16311 => x"00000000",
         16312 => x"00000000",
         16313 => x"00000000",
         16314 => x"00000000",
         16315 => x"00000000",
         16316 => x"00000000",
         16317 => x"00000000",
         16318 => x"00000000",
         16319 => x"00000000",
         16320 => x"00000000",
         16321 => x"00000000",
         16322 => x"00000000",
         16323 => x"00000000",
         16324 => x"00000000",
         16325 => x"00000000",
         16326 => x"00000000",
         16327 => x"00000000",
         16328 => x"00000000",
         16329 => x"00000000",
         16330 => x"00000000",
         16331 => x"00000000",
         16332 => x"00000000",
         16333 => x"00000000",
         16334 => x"00000000",
         16335 => x"00000000",
         16336 => x"00000000",
         16337 => x"00000000",
         16338 => x"00000000",
         16339 => x"00000000",
         16340 => x"00000000",
         16341 => x"00000000",
         16342 => x"00000000",
         16343 => x"00000000",
         16344 => x"00000000",
         16345 => x"00000000",
         16346 => x"00000000",
         16347 => x"00000000",
         16348 => x"00000000",
         16349 => x"00000000",
         16350 => x"00000000",
         16351 => x"00000000",
         16352 => x"00000000",
         16353 => x"00000000",
         16354 => x"00000000",
         16355 => x"00000000",
         16356 => x"00000000",
         16357 => x"00000000",
         16358 => x"00000000",
         16359 => x"00000000",
         16360 => x"00000000",
         16361 => x"00000000",
         16362 => x"00000000",
         16363 => x"00000000",
         16364 => x"00000000",
         16365 => x"00000000",
         16366 => x"00000000",
         16367 => x"00000000",
         16368 => x"00000000",
         16369 => x"00000000",
         16370 => x"00000000",
         16371 => x"00000000",
         16372 => x"00000000",
         16373 => x"00000000",
         16374 => x"00000000",
         16375 => x"00000000",
         16376 => x"00000000",
         16377 => x"00000000",
         16378 => x"00000000",
         16379 => x"00000000",
         16380 => x"00000000",
         16381 => x"00000000",
         16382 => x"00000000",
         16383 => x"00000000",
         16384 => x"00000000",
         16385 => x"00000000",
         16386 => x"00000000",
         16387 => x"00000000",
         16388 => x"00000000",
         16389 => x"00000000",
         16390 => x"00000000",
         16391 => x"00000000",
         16392 => x"00000000",
         16393 => x"00000000",
         16394 => x"00000000",
         16395 => x"00000000",
         16396 => x"00000000",
         16397 => x"00000000",
         16398 => x"00000000",
         16399 => x"00000000",
         16400 => x"00000000",
         16401 => x"00000000",
         16402 => x"00000000",
         16403 => x"00000000",
         16404 => x"00000000",
         16405 => x"00000000",
         16406 => x"00000000",
         16407 => x"00000000",
         16408 => x"00000000",
         16409 => x"00000000",
         16410 => x"00000000",
         16411 => x"00000000",
         16412 => x"00000000",
         16413 => x"00000000",
         16414 => x"00000000",
         16415 => x"00000000",
         16416 => x"00000000",
         16417 => x"00000000",
         16418 => x"00000000",
         16419 => x"00000000",
         16420 => x"00000000",
         16421 => x"00000000",
         16422 => x"00000000",
         16423 => x"00000000",
         16424 => x"00000000",
         16425 => x"00000000",
         16426 => x"00000000",
         16427 => x"00000000",
         16428 => x"00000000",
         16429 => x"00000000",
         16430 => x"00000000",
         16431 => x"00000000",
         16432 => x"00000000",
         16433 => x"00000000",
         16434 => x"00000000",
         16435 => x"00000000",
         16436 => x"00000000",
         16437 => x"00000000",
         16438 => x"00000000",
         16439 => x"00000000",
         16440 => x"00000000",
         16441 => x"00000000",
         16442 => x"00000000",
         16443 => x"00000000",
         16444 => x"00000000",
         16445 => x"00000000",
         16446 => x"00000000",
         16447 => x"00000000",
         16448 => x"00000000",
         16449 => x"00000000",
         16450 => x"00000000",
         16451 => x"00000000",
         16452 => x"00000000",
         16453 => x"00000000",
         16454 => x"00000000",
         16455 => x"00000000",
         16456 => x"00000000",
         16457 => x"00000000",
         16458 => x"00000000",
         16459 => x"00000000",
         16460 => x"00000000",
         16461 => x"00000000",
         16462 => x"00000000",
         16463 => x"00000000",
         16464 => x"00000000",
         16465 => x"00000000",
         16466 => x"00000000",
         16467 => x"00000000",
         16468 => x"00000000",
         16469 => x"00000000",
         16470 => x"00000000",
         16471 => x"00000000",
         16472 => x"00000000",
         16473 => x"00000000",
         16474 => x"00000000",
         16475 => x"00000000",
         16476 => x"00000000",
         16477 => x"00000000",
         16478 => x"00000000",
         16479 => x"00000000",
         16480 => x"00000000",
         16481 => x"00000000",
         16482 => x"00000000",
         16483 => x"00000000",
         16484 => x"00000000",
         16485 => x"00000000",
         16486 => x"00000000",
         16487 => x"00000000",
         16488 => x"00000000",
         16489 => x"00000000",
         16490 => x"00000000",
         16491 => x"00000000",
         16492 => x"00000000",
         16493 => x"00000000",
         16494 => x"00000000",
         16495 => x"00000000",
         16496 => x"00000000",
         16497 => x"00000000",
         16498 => x"00000000",
         16499 => x"00000000",
         16500 => x"00000000",
         16501 => x"00000000",
         16502 => x"00000000",
         16503 => x"00000000",
         16504 => x"00000000",
         16505 => x"00000000",
         16506 => x"00000000",
         16507 => x"00000000",
         16508 => x"00000000",
         16509 => x"00000000",
         16510 => x"00000000",
         16511 => x"00000000",
         16512 => x"00000000",
         16513 => x"00000000",
         16514 => x"00000000",
         16515 => x"00000000",
         16516 => x"00000000",
         16517 => x"00000000",
         16518 => x"00000000",
         16519 => x"00000000",
         16520 => x"00000000",
         16521 => x"00000000",
         16522 => x"00000000",
         16523 => x"00000000",
         16524 => x"00000000",
         16525 => x"00000000",
         16526 => x"00000000",
         16527 => x"00000000",
         16528 => x"00000000",
         16529 => x"00000000",
         16530 => x"00000000",
         16531 => x"00000000",
         16532 => x"00000000",
         16533 => x"00000000",
         16534 => x"00000000",
         16535 => x"00000000",
         16536 => x"00000000",
         16537 => x"00000000",
         16538 => x"00000000",
         16539 => x"00000000",
         16540 => x"00000000",
         16541 => x"00000000",
         16542 => x"00000000",
         16543 => x"00000000",
         16544 => x"00000000",
         16545 => x"00000000",
         16546 => x"00000000",
         16547 => x"00000000",
         16548 => x"00000000",
         16549 => x"00000000",
         16550 => x"00000000",
         16551 => x"00000000",
         16552 => x"00000000",
         16553 => x"00000000",
         16554 => x"00000000",
         16555 => x"00000000",
         16556 => x"00000000",
         16557 => x"00000000",
         16558 => x"00000000",
         16559 => x"00000000",
         16560 => x"00000000",
         16561 => x"00000000",
         16562 => x"00000000",
         16563 => x"00000000",
         16564 => x"00000000",
         16565 => x"00000000",
         16566 => x"00000000",
         16567 => x"00000000",
         16568 => x"00000000",
         16569 => x"00000000",
         16570 => x"00000000",
         16571 => x"00000000",
         16572 => x"00000000",
         16573 => x"00000000",
         16574 => x"00000000",
         16575 => x"00000000",
         16576 => x"00000000",
         16577 => x"00000000",
         16578 => x"00000000",
         16579 => x"00000000",
         16580 => x"00000000",
         16581 => x"00000000",
         16582 => x"00000000",
         16583 => x"00000000",
         16584 => x"00000000",
         16585 => x"00000000",
         16586 => x"00000000",
         16587 => x"00000000",
         16588 => x"00000000",
         16589 => x"00000000",
         16590 => x"00000000",
         16591 => x"00000000",
         16592 => x"00000000",
         16593 => x"00000000",
         16594 => x"00000000",
         16595 => x"00000000",
         16596 => x"00000000",
         16597 => x"00000000",
         16598 => x"00000000",
         16599 => x"00000000",
         16600 => x"00000000",
         16601 => x"00000000",
         16602 => x"00000000",
         16603 => x"00000000",
         16604 => x"00000000",
         16605 => x"00000000",
         16606 => x"00000000",
         16607 => x"00000000",
         16608 => x"00000000",
         16609 => x"00000000",
         16610 => x"00000000",
         16611 => x"00000000",
         16612 => x"00000000",
         16613 => x"00000000",
         16614 => x"00000000",
         16615 => x"00000000",
         16616 => x"00000000",
         16617 => x"00000000",
         16618 => x"00000000",
         16619 => x"00000000",
         16620 => x"00000000",
         16621 => x"00000000",
         16622 => x"00000000",
         16623 => x"00000000",
         16624 => x"00000000",
         16625 => x"00000000",
         16626 => x"00000000",
         16627 => x"00000000",
         16628 => x"00000000",
         16629 => x"00000000",
         16630 => x"00000000",
         16631 => x"00000000",
         16632 => x"00000000",
         16633 => x"00000000",
         16634 => x"00000000",
         16635 => x"00000000",
         16636 => x"00000000",
         16637 => x"00000000",
         16638 => x"00000000",
         16639 => x"00000000",
         16640 => x"00000000",
         16641 => x"00000000",
         16642 => x"00000000",
         16643 => x"00000000",
         16644 => x"00000000",
         16645 => x"00000000",
         16646 => x"00000000",
         16647 => x"00000000",
         16648 => x"00000000",
         16649 => x"00000000",
         16650 => x"00000000",
         16651 => x"00000000",
         16652 => x"00000000",
         16653 => x"00000000",
         16654 => x"00000000",
         16655 => x"00000000",
         16656 => x"00000000",
         16657 => x"00000000",
         16658 => x"00000000",
         16659 => x"00000000",
         16660 => x"00000000",
         16661 => x"00000000",
         16662 => x"00000000",
         16663 => x"00000000",
         16664 => x"00000000",
         16665 => x"00000000",
         16666 => x"00000000",
         16667 => x"00000000",
         16668 => x"00000000",
         16669 => x"00000000",
         16670 => x"00000000",
         16671 => x"00000000",
         16672 => x"00000000",
         16673 => x"00000000",
         16674 => x"00000000",
         16675 => x"00000000",
         16676 => x"00000000",
         16677 => x"00000000",
         16678 => x"00000000",
         16679 => x"00000000",
         16680 => x"00000000",
         16681 => x"00000000",
         16682 => x"00000000",
         16683 => x"00000000",
         16684 => x"00000000",
         16685 => x"00000000",
         16686 => x"00000000",
         16687 => x"00000000",
         16688 => x"00000000",
         16689 => x"00000000",
         16690 => x"00000000",
         16691 => x"00000000",
         16692 => x"00000000",
         16693 => x"00000000",
         16694 => x"00000000",
         16695 => x"00000000",
         16696 => x"00000000",
         16697 => x"00000000",
         16698 => x"00000000",
         16699 => x"00000000",
         16700 => x"00000000",
         16701 => x"00000000",
         16702 => x"00000000",
         16703 => x"00000000",
         16704 => x"00000000",
         16705 => x"00000000",
         16706 => x"00000000",
         16707 => x"00000000",
         16708 => x"00000000",
         16709 => x"00000000",
         16710 => x"00000000",
         16711 => x"00000000",
         16712 => x"00000000",
         16713 => x"00000000",
         16714 => x"00000000",
         16715 => x"00000000",
         16716 => x"00000000",
         16717 => x"00000000",
         16718 => x"00000000",
         16719 => x"00000000",
         16720 => x"00000000",
         16721 => x"00000000",
         16722 => x"00000000",
         16723 => x"00000000",
         16724 => x"00000000",
         16725 => x"00000000",
         16726 => x"00000000",
         16727 => x"00000000",
         16728 => x"00000000",
         16729 => x"00000000",
         16730 => x"00000000",
         16731 => x"00000000",
         16732 => x"00000000",
         16733 => x"00000000",
         16734 => x"00000000",
         16735 => x"00000000",
         16736 => x"00000000",
         16737 => x"00000000",
         16738 => x"00000000",
         16739 => x"00000000",
         16740 => x"00000000",
         16741 => x"00000000",
         16742 => x"00000000",
         16743 => x"00000000",
         16744 => x"00000000",
         16745 => x"00000000",
         16746 => x"00000000",
         16747 => x"00000000",
         16748 => x"00000000",
         16749 => x"00000000",
         16750 => x"00000000",
         16751 => x"00000000",
         16752 => x"00000000",
         16753 => x"00000000",
         16754 => x"00000000",
         16755 => x"00000000",
         16756 => x"00000000",
         16757 => x"00000000",
         16758 => x"00000000",
         16759 => x"00000000",
         16760 => x"00000000",
         16761 => x"00000000",
         16762 => x"00000000",
         16763 => x"00000000",
         16764 => x"00000000",
         16765 => x"00000000",
         16766 => x"00000000",
         16767 => x"00000000",
         16768 => x"00000000",
         16769 => x"00000000",
         16770 => x"00000000",
         16771 => x"00000000",
         16772 => x"00000000",
         16773 => x"00000000",
         16774 => x"00000000",
         16775 => x"00000000",
         16776 => x"00000000",
         16777 => x"00000000",
         16778 => x"00000000",
         16779 => x"00000000",
         16780 => x"00000000",
         16781 => x"00000000",
         16782 => x"00000000",
         16783 => x"00000000",
         16784 => x"00000000",
         16785 => x"00000000",
         16786 => x"00000000",
         16787 => x"00000000",
         16788 => x"00000000",
         16789 => x"00000000",
         16790 => x"00000000",
         16791 => x"00000000",
         16792 => x"00000000",
         16793 => x"00000000",
         16794 => x"00000000",
         16795 => x"00000000",
         16796 => x"00000000",
         16797 => x"00000000",
         16798 => x"00000000",
         16799 => x"00000000",
         16800 => x"00000000",
         16801 => x"00000000",
         16802 => x"00000000",
         16803 => x"00000000",
         16804 => x"00000000",
         16805 => x"00000000",
         16806 => x"00000000",
         16807 => x"00000000",
         16808 => x"00000000",
         16809 => x"00000000",
         16810 => x"00000000",
         16811 => x"00000000",
         16812 => x"00000000",
         16813 => x"00000000",
         16814 => x"00000000",
         16815 => x"00000000",
         16816 => x"00000000",
         16817 => x"00000000",
         16818 => x"00000000",
         16819 => x"00000000",
         16820 => x"00000000",
         16821 => x"00000000",
         16822 => x"00000000",
         16823 => x"00000000",
         16824 => x"00000000",
         16825 => x"00000000",
         16826 => x"00000000",
         16827 => x"00000000",
         16828 => x"00000000",
         16829 => x"00000000",
         16830 => x"00000000",
         16831 => x"00000000",
         16832 => x"00000000",
         16833 => x"00000000",
         16834 => x"00000000",
         16835 => x"00000000",
         16836 => x"00000000",
         16837 => x"00000000",
         16838 => x"00000000",
         16839 => x"00000000",
         16840 => x"00000000",
         16841 => x"00000000",
         16842 => x"00000000",
         16843 => x"00000000",
         16844 => x"00000000",
         16845 => x"00000000",
         16846 => x"00000000",
         16847 => x"00000000",
         16848 => x"00000000",
         16849 => x"00000000",
         16850 => x"00000000",
         16851 => x"00000000",
         16852 => x"00000000",
         16853 => x"00000000",
         16854 => x"00000000",
         16855 => x"00000000",
         16856 => x"00000000",
         16857 => x"00000000",
         16858 => x"00000000",
         16859 => x"00000000",
         16860 => x"00000000",
         16861 => x"00000000",
         16862 => x"00000000",
         16863 => x"00000000",
         16864 => x"00000000",
         16865 => x"00000000",
         16866 => x"00000000",
         16867 => x"00000000",
         16868 => x"00000000",
         16869 => x"00000000",
         16870 => x"00000000",
         16871 => x"00000000",
         16872 => x"00000000",
         16873 => x"00000000",
         16874 => x"00000000",
         16875 => x"00000000",
         16876 => x"00000000",
         16877 => x"00000000",
         16878 => x"00000000",
         16879 => x"00000000",
         16880 => x"00000000",
         16881 => x"00000000",
         16882 => x"00000000",
         16883 => x"00000000",
         16884 => x"00000000",
         16885 => x"00000000",
         16886 => x"00000000",
         16887 => x"00000000",
         16888 => x"00000000",
         16889 => x"00000000",
         16890 => x"00000000",
         16891 => x"00000000",
         16892 => x"00000000",
         16893 => x"00000000",
         16894 => x"00000000",
         16895 => x"00000000",
         16896 => x"00000000",
         16897 => x"00000000",
         16898 => x"00000000",
         16899 => x"00000000",
         16900 => x"00000000",
         16901 => x"00000000",
         16902 => x"00000000",
         16903 => x"00000000",
         16904 => x"00000000",
         16905 => x"00000000",
         16906 => x"00000000",
         16907 => x"00000000",
         16908 => x"00000000",
         16909 => x"00000000",
         16910 => x"00000000",
         16911 => x"00000000",
         16912 => x"00000000",
         16913 => x"00000000",
         16914 => x"00000000",
         16915 => x"00000000",
         16916 => x"00000000",
         16917 => x"00000000",
         16918 => x"00000000",
         16919 => x"00000000",
         16920 => x"00000000",
         16921 => x"00000000",
         16922 => x"00000000",
         16923 => x"00000000",
         16924 => x"00000000",
         16925 => x"00000000",
         16926 => x"00000000",
         16927 => x"00000000",
         16928 => x"00000000",
         16929 => x"00000000",
         16930 => x"00000000",
         16931 => x"00000000",
         16932 => x"00000000",
         16933 => x"00000000",
         16934 => x"00000000",
         16935 => x"00000000",
         16936 => x"00000000",
         16937 => x"00000000",
         16938 => x"00000000",
         16939 => x"00000000",
         16940 => x"00000000",
         16941 => x"00000000",
         16942 => x"00000000",
         16943 => x"00000000",
         16944 => x"00000000",
         16945 => x"00000000",
         16946 => x"00000000",
         16947 => x"00000000",
         16948 => x"00000000",
         16949 => x"00000000",
         16950 => x"00000000",
         16951 => x"00000000",
         16952 => x"00000000",
         16953 => x"00000000",
         16954 => x"00000000",
         16955 => x"00000000",
         16956 => x"00000000",
         16957 => x"00000000",
         16958 => x"00000000",
         16959 => x"00000000",
         16960 => x"00000000",
         16961 => x"00000000",
         16962 => x"00000000",
         16963 => x"00000000",
         16964 => x"00000000",
         16965 => x"00000000",
         16966 => x"00000000",
         16967 => x"00000000",
         16968 => x"00000000",
         16969 => x"00000000",
         16970 => x"00000000",
         16971 => x"00000000",
         16972 => x"00000000",
         16973 => x"00000000",
         16974 => x"00000000",
         16975 => x"00000000",
         16976 => x"00000000",
         16977 => x"00000000",
         16978 => x"00000000",
         16979 => x"00000000",
         16980 => x"00000000",
         16981 => x"00000000",
         16982 => x"00000000",
         16983 => x"00000000",
         16984 => x"00000000",
         16985 => x"00000000",
         16986 => x"00000000",
         16987 => x"00000000",
         16988 => x"00000000",
         16989 => x"00000000",
         16990 => x"00000000",
         16991 => x"00000000",
         16992 => x"00000000",
         16993 => x"00000000",
         16994 => x"00000000",
         16995 => x"00000000",
         16996 => x"00000000",
         16997 => x"00000000",
         16998 => x"00000000",
         16999 => x"00000000",
         17000 => x"00000000",
         17001 => x"00000000",
         17002 => x"00000000",
         17003 => x"00000000",
         17004 => x"00000000",
         17005 => x"00000000",
         17006 => x"00000000",
         17007 => x"00000000",
         17008 => x"00000000",
         17009 => x"00000000",
         17010 => x"00000000",
         17011 => x"00000000",
         17012 => x"00000000",
         17013 => x"00000000",
         17014 => x"00000000",
         17015 => x"00000000",
         17016 => x"00000000",
         17017 => x"00000000",
         17018 => x"00000000",
         17019 => x"00000000",
         17020 => x"00000000",
         17021 => x"00000000",
         17022 => x"00000000",
         17023 => x"00000000",
         17024 => x"00000000",
         17025 => x"00000000",
         17026 => x"00000000",
         17027 => x"00000000",
         17028 => x"00000000",
         17029 => x"00000000",
         17030 => x"00000000",
         17031 => x"00000000",
         17032 => x"00000000",
         17033 => x"00000000",
         17034 => x"00000000",
         17035 => x"00000000",
         17036 => x"00000000",
         17037 => x"00000000",
         17038 => x"00000000",
         17039 => x"00000000",
         17040 => x"00000000",
         17041 => x"00000000",
         17042 => x"00000000",
         17043 => x"00000000",
         17044 => x"00000000",
         17045 => x"00000000",
         17046 => x"00000000",
         17047 => x"00000000",
         17048 => x"00000000",
         17049 => x"00000000",
         17050 => x"00000000",
         17051 => x"00000000",
         17052 => x"00000000",
         17053 => x"00000000",
         17054 => x"00000000",
         17055 => x"00000000",
         17056 => x"00000000",
         17057 => x"00000000",
         17058 => x"00000000",
         17059 => x"00000000",
         17060 => x"00000000",
         17061 => x"00000000",
         17062 => x"00000000",
         17063 => x"00000000",
         17064 => x"00000000",
         17065 => x"00000000",
         17066 => x"00000000",
         17067 => x"00000000",
         17068 => x"00000000",
         17069 => x"00000000",
         17070 => x"00000000",
         17071 => x"00000000",
         17072 => x"00000000",
         17073 => x"00000000",
         17074 => x"00000000",
         17075 => x"00000000",
         17076 => x"00000000",
         17077 => x"00000000",
         17078 => x"00000000",
         17079 => x"00000000",
         17080 => x"00000000",
         17081 => x"00000000",
         17082 => x"00000000",
         17083 => x"00000000",
         17084 => x"00000000",
         17085 => x"00000000",
         17086 => x"00000000",
         17087 => x"00000000",
         17088 => x"00000000",
         17089 => x"00000000",
         17090 => x"00000000",
         17091 => x"00000000",
         17092 => x"00000000",
         17093 => x"00000000",
         17094 => x"00000000",
         17095 => x"00000000",
         17096 => x"00000000",
         17097 => x"00000000",
         17098 => x"00000000",
         17099 => x"00000000",
         17100 => x"00000000",
         17101 => x"00000000",
         17102 => x"00000000",
         17103 => x"00000000",
         17104 => x"00000000",
         17105 => x"00000000",
         17106 => x"00000000",
         17107 => x"00000000",
         17108 => x"00000000",
         17109 => x"00000000",
         17110 => x"00000000",
         17111 => x"00000000",
         17112 => x"00000000",
         17113 => x"00000000",
         17114 => x"00000000",
         17115 => x"00000000",
         17116 => x"00000000",
         17117 => x"00000000",
         17118 => x"00000000",
         17119 => x"00000000",
         17120 => x"00000000",
         17121 => x"00000000",
         17122 => x"00000000",
         17123 => x"00000000",
         17124 => x"00000000",
         17125 => x"00000000",
         17126 => x"00000000",
         17127 => x"00000000",
         17128 => x"00000000",
         17129 => x"00000000",
         17130 => x"00000000",
         17131 => x"00000000",
         17132 => x"00000000",
         17133 => x"00000000",
         17134 => x"00000000",
         17135 => x"00000000",
         17136 => x"00000000",
         17137 => x"00000000",
         17138 => x"00000000",
         17139 => x"00000000",
         17140 => x"00000000",
         17141 => x"00000000",
         17142 => x"00000000",
         17143 => x"00000000",
         17144 => x"00000000",
         17145 => x"00000000",
         17146 => x"00000000",
         17147 => x"00000000",
         17148 => x"00000000",
         17149 => x"00000000",
         17150 => x"00000000",
         17151 => x"00000000",
         17152 => x"00000000",
         17153 => x"00000000",
         17154 => x"00000000",
         17155 => x"00000000",
         17156 => x"00000000",
         17157 => x"00000000",
         17158 => x"00000000",
         17159 => x"00000000",
         17160 => x"00000000",
         17161 => x"00000000",
         17162 => x"00000000",
         17163 => x"00000000",
         17164 => x"00000000",
         17165 => x"00000000",
         17166 => x"00000000",
         17167 => x"00000000",
         17168 => x"00000000",
         17169 => x"00000000",
         17170 => x"00000000",
         17171 => x"00000000",
         17172 => x"00000000",
         17173 => x"00000000",
         17174 => x"00000000",
         17175 => x"00000000",
         17176 => x"00000000",
         17177 => x"00000000",
         17178 => x"00000000",
         17179 => x"00000000",
         17180 => x"00000000",
         17181 => x"00000000",
         17182 => x"00000000",
         17183 => x"00000000",
         17184 => x"00000000",
         17185 => x"00000000",
         17186 => x"00000000",
         17187 => x"00000000",
         17188 => x"00000000",
         17189 => x"00000000",
         17190 => x"00000000",
         17191 => x"00000000",
         17192 => x"00000000",
         17193 => x"00000000",
         17194 => x"00000000",
         17195 => x"00000000",
         17196 => x"00000000",
         17197 => x"00000000",
         17198 => x"00000000",
         17199 => x"00000000",
         17200 => x"00000000",
         17201 => x"00000000",
         17202 => x"00000000",
         17203 => x"00000000",
         17204 => x"00000000",
         17205 => x"00000000",
         17206 => x"00000000",
         17207 => x"00000000",
         17208 => x"00000000",
         17209 => x"00000000",
         17210 => x"00000000",
         17211 => x"00000000",
         17212 => x"00000000",
         17213 => x"00000000",
         17214 => x"00000000",
         17215 => x"00000000",
         17216 => x"00000000",
         17217 => x"00000000",
         17218 => x"00000000",
         17219 => x"00000000",
         17220 => x"00000000",
         17221 => x"00000000",
         17222 => x"00000000",
         17223 => x"00000000",
         17224 => x"00000000",
         17225 => x"00000000",
         17226 => x"00000000",
         17227 => x"00000000",
         17228 => x"00000000",
         17229 => x"00000000",
         17230 => x"00000000",
         17231 => x"00000000",
         17232 => x"00000000",
         17233 => x"00000000",
         17234 => x"00000000",
         17235 => x"00000000",
         17236 => x"00000000",
         17237 => x"00000000",
         17238 => x"00000000",
         17239 => x"00000000",
         17240 => x"00000000",
         17241 => x"00000000",
         17242 => x"00000000",
         17243 => x"00000000",
         17244 => x"00000000",
         17245 => x"00000000",
         17246 => x"00000000",
         17247 => x"00000000",
         17248 => x"00000000",
         17249 => x"00000000",
         17250 => x"00000000",
         17251 => x"00000000",
         17252 => x"00000000",
         17253 => x"00000000",
         17254 => x"00000000",
         17255 => x"00000000",
         17256 => x"00000000",
         17257 => x"00000000",
         17258 => x"00000000",
         17259 => x"00000000",
         17260 => x"00000000",
         17261 => x"00000000",
         17262 => x"00000000",
         17263 => x"00000000",
         17264 => x"00000000",
         17265 => x"00000000",
         17266 => x"00000000",
         17267 => x"00000000",
         17268 => x"00000000",
         17269 => x"00000000",
         17270 => x"00000000",
         17271 => x"00000000",
         17272 => x"00000000",
         17273 => x"00000000",
         17274 => x"00000000",
         17275 => x"00000000",
         17276 => x"00000000",
         17277 => x"00000000",
         17278 => x"00000000",
         17279 => x"00000000",
         17280 => x"00000000",
         17281 => x"00000000",
         17282 => x"00000000",
         17283 => x"00000000",
         17284 => x"00000000",
         17285 => x"00000000",
         17286 => x"00000000",
         17287 => x"00000000",
         17288 => x"00000000",
         17289 => x"00000000",
         17290 => x"00000000",
         17291 => x"00000000",
         17292 => x"00000000",
         17293 => x"00000000",
         17294 => x"00000000",
         17295 => x"00000000",
         17296 => x"00000000",
         17297 => x"00000000",
         17298 => x"00000000",
         17299 => x"00000000",
         17300 => x"00000000",
         17301 => x"00000000",
         17302 => x"00000000",
         17303 => x"00000000",
         17304 => x"00000000",
         17305 => x"00000000",
         17306 => x"00000000",
         17307 => x"00000000",
         17308 => x"00000000",
         17309 => x"00000000",
         17310 => x"00000000",
         17311 => x"00000000",
         17312 => x"00000000",
         17313 => x"00000000",
         17314 => x"00000000",
         17315 => x"00000000",
         17316 => x"00000000",
         17317 => x"00000000",
         17318 => x"00000000",
         17319 => x"00000000",
         17320 => x"00000000",
         17321 => x"00000000",
         17322 => x"00000000",
         17323 => x"00000000",
         17324 => x"00000000",
         17325 => x"00000000",
         17326 => x"00000000",
         17327 => x"00000000",
         17328 => x"00000000",
         17329 => x"00000000",
         17330 => x"00000000",
         17331 => x"00000000",
         17332 => x"00000000",
         17333 => x"00000000",
         17334 => x"00000000",
         17335 => x"00000000",
         17336 => x"00000000",
         17337 => x"00000000",
         17338 => x"00000000",
         17339 => x"00000000",
         17340 => x"00000000",
         17341 => x"00000000",
         17342 => x"00000000",
         17343 => x"00000000",
         17344 => x"00000000",
         17345 => x"00000000",
         17346 => x"00000000",
         17347 => x"00000000",
         17348 => x"00000000",
         17349 => x"00000000",
         17350 => x"00000000",
         17351 => x"00000000",
         17352 => x"00000000",
         17353 => x"00000000",
         17354 => x"00000000",
         17355 => x"00000000",
         17356 => x"00000000",
         17357 => x"00000000",
         17358 => x"00000000",
         17359 => x"00000000",
         17360 => x"00000000",
         17361 => x"00000000",
         17362 => x"00000000",
         17363 => x"00000000",
         17364 => x"00000000",
         17365 => x"00000000",
         17366 => x"00000000",
         17367 => x"00000000",
         17368 => x"00000000",
         17369 => x"00000000",
         17370 => x"00000000",
         17371 => x"00000000",
         17372 => x"00000000",
         17373 => x"00000000",
         17374 => x"00000000",
         17375 => x"00000000",
         17376 => x"00000000",
         17377 => x"00000000",
         17378 => x"00000000",
         17379 => x"00000000",
         17380 => x"00000000",
         17381 => x"00000000",
         17382 => x"00000000",
         17383 => x"00000000",
         17384 => x"00000000",
         17385 => x"00000000",
         17386 => x"00000000",
         17387 => x"00000000",
         17388 => x"00000000",
         17389 => x"00000000",
         17390 => x"00000000",
         17391 => x"00000000",
         17392 => x"00000000",
         17393 => x"00000000",
         17394 => x"00000000",
         17395 => x"00000000",
         17396 => x"00000000",
         17397 => x"00000000",
         17398 => x"00000000",
         17399 => x"00000000",
         17400 => x"00000000",
         17401 => x"00000000",
         17402 => x"00000000",
         17403 => x"00000000",
         17404 => x"00000000",
         17405 => x"00000000",
         17406 => x"00000000",
         17407 => x"00000000",
         17408 => x"00000000",
         17409 => x"00000000",
         17410 => x"00000000",
         17411 => x"00000000",
         17412 => x"00000000",
         17413 => x"00000000",
         17414 => x"00000000",
         17415 => x"00000000",
         17416 => x"00000000",
         17417 => x"00000000",
         17418 => x"00000000",
         17419 => x"00000000",
         17420 => x"00000000",
         17421 => x"00000000",
         17422 => x"00000000",
         17423 => x"00000000",
         17424 => x"00000000",
         17425 => x"00000000",
         17426 => x"00000000",
         17427 => x"00000000",
         17428 => x"00000000",
         17429 => x"00000000",
         17430 => x"00000000",
         17431 => x"00000000",
         17432 => x"00000000",
         17433 => x"00000000",
         17434 => x"00000000",
         17435 => x"00000000",
         17436 => x"00000000",
         17437 => x"00000000",
         17438 => x"00000000",
         17439 => x"00000000",
         17440 => x"00000000",
         17441 => x"00000000",
         17442 => x"00000000",
         17443 => x"00000000",
         17444 => x"00000000",
         17445 => x"00000000",
         17446 => x"00000000",
         17447 => x"00000000",
         17448 => x"00000000",
         17449 => x"00000000",
         17450 => x"00000000",
         17451 => x"00000000",
         17452 => x"00000000",
         17453 => x"00000000",
         17454 => x"00000000",
         17455 => x"00000000",
         17456 => x"00000000",
         17457 => x"00000000",
         17458 => x"00000000",
         17459 => x"00000000",
         17460 => x"00000000",
         17461 => x"00000000",
         17462 => x"00000000",
         17463 => x"00000000",
         17464 => x"00000000",
         17465 => x"00000000",
         17466 => x"00000000",
         17467 => x"00000000",
         17468 => x"00000000",
         17469 => x"00000000",
         17470 => x"00000000",
         17471 => x"00000000",
         17472 => x"00000000",
         17473 => x"00000000",
         17474 => x"00000000",
         17475 => x"00000000",
         17476 => x"00000000",
         17477 => x"00000000",
         17478 => x"00000000",
         17479 => x"00000000",
         17480 => x"00000000",
         17481 => x"00000000",
         17482 => x"00000000",
         17483 => x"00000000",
         17484 => x"00000000",
         17485 => x"00000000",
         17486 => x"00000000",
         17487 => x"00000000",
         17488 => x"00000000",
         17489 => x"00000000",
         17490 => x"00000000",
         17491 => x"00000000",
         17492 => x"00000000",
         17493 => x"00000000",
         17494 => x"00000000",
         17495 => x"00000000",
         17496 => x"00000000",
         17497 => x"00000000",
         17498 => x"00000000",
         17499 => x"00000000",
         17500 => x"00000000",
         17501 => x"00000000",
         17502 => x"00000000",
         17503 => x"00000000",
         17504 => x"00000000",
         17505 => x"00000000",
         17506 => x"00000000",
         17507 => x"00000000",
         17508 => x"00000000",
         17509 => x"00000000",
         17510 => x"00000000",
         17511 => x"00000000",
         17512 => x"00000000",
         17513 => x"00000000",
         17514 => x"00000000",
         17515 => x"00000000",
         17516 => x"00000000",
         17517 => x"00000000",
         17518 => x"00000000",
         17519 => x"00000000",
         17520 => x"00000000",
         17521 => x"00000000",
         17522 => x"00000000",
         17523 => x"00000000",
         17524 => x"00000000",
         17525 => x"00000000",
         17526 => x"00000000",
         17527 => x"00000000",
         17528 => x"00000000",
         17529 => x"00000000",
         17530 => x"00000000",
         17531 => x"00000000",
         17532 => x"00000000",
         17533 => x"00000000",
         17534 => x"00000000",
         17535 => x"00000000",
         17536 => x"00000000",
         17537 => x"00000000",
         17538 => x"00000000",
         17539 => x"00000000",
         17540 => x"00000000",
         17541 => x"00000000",
         17542 => x"00000000",
         17543 => x"00000000",
         17544 => x"00000000",
         17545 => x"00000000",
         17546 => x"00000000",
         17547 => x"00000000",
         17548 => x"00000000",
         17549 => x"00000000",
         17550 => x"00000000",
         17551 => x"00000000",
         17552 => x"00000000",
         17553 => x"00000000",
         17554 => x"00000000",
         17555 => x"00000000",
         17556 => x"00000000",
         17557 => x"00000000",
         17558 => x"00000000",
         17559 => x"00000000",
         17560 => x"00000000",
         17561 => x"00000000",
         17562 => x"00000000",
         17563 => x"00000000",
         17564 => x"00000000",
         17565 => x"00000000",
         17566 => x"00000000",
         17567 => x"00000000",
         17568 => x"00000000",
         17569 => x"00000000",
         17570 => x"00000000",
         17571 => x"00000000",
         17572 => x"00000000",
         17573 => x"00000000",
         17574 => x"00000000",
         17575 => x"00000000",
         17576 => x"00000000",
         17577 => x"00000000",
         17578 => x"00000000",
         17579 => x"00000000",
         17580 => x"00000000",
         17581 => x"00000000",
         17582 => x"00000000",
         17583 => x"00000000",
         17584 => x"00000000",
         17585 => x"00000000",
         17586 => x"00000000",
         17587 => x"00000000",
         17588 => x"00000000",
         17589 => x"00000000",
         17590 => x"00000000",
         17591 => x"00000000",
         17592 => x"00000000",
         17593 => x"00000000",
         17594 => x"00000000",
         17595 => x"00000000",
         17596 => x"00000000",
         17597 => x"00000000",
         17598 => x"00000000",
         17599 => x"00000000",
         17600 => x"00000000",
         17601 => x"00000000",
         17602 => x"00000000",
         17603 => x"00000000",
         17604 => x"00000000",
         17605 => x"00000000",
         17606 => x"00000000",
         17607 => x"00000000",
         17608 => x"00000000",
         17609 => x"00000000",
         17610 => x"00000000",
         17611 => x"00000000",
         17612 => x"00000000",
         17613 => x"00000000",
         17614 => x"00000000",
         17615 => x"00000000",
         17616 => x"00000000",
         17617 => x"00000000",
         17618 => x"00000000",
         17619 => x"00000000",
         17620 => x"00000000",
         17621 => x"00000000",
         17622 => x"00000000",
         17623 => x"00000000",
         17624 => x"00000000",
         17625 => x"00000000",
         17626 => x"00000000",
         17627 => x"00000000",
         17628 => x"00000000",
         17629 => x"00000000",
         17630 => x"00000000",
         17631 => x"00000000",
         17632 => x"00000000",
         17633 => x"00000000",
         17634 => x"00000000",
         17635 => x"00000000",
         17636 => x"00000000",
         17637 => x"00000000",
         17638 => x"00000000",
         17639 => x"00000000",
         17640 => x"00000000",
         17641 => x"00000000",
         17642 => x"00000000",
         17643 => x"00000000",
         17644 => x"00000000",
         17645 => x"00000000",
         17646 => x"00000000",
         17647 => x"00000000",
         17648 => x"00000000",
         17649 => x"00000000",
         17650 => x"00000000",
         17651 => x"00000000",
         17652 => x"00000000",
         17653 => x"00000000",
         17654 => x"00000000",
         17655 => x"00000000",
         17656 => x"00000000",
         17657 => x"00000000",
         17658 => x"00000000",
         17659 => x"00000000",
         17660 => x"00000000",
         17661 => x"00000000",
         17662 => x"00000000",
         17663 => x"00000000",
         17664 => x"00000000",
         17665 => x"00000000",
         17666 => x"00000000",
         17667 => x"00000000",
         17668 => x"00000000",
         17669 => x"00000000",
         17670 => x"00000000",
         17671 => x"00000000",
         17672 => x"00000000",
         17673 => x"00000000",
         17674 => x"00000000",
         17675 => x"00000000",
         17676 => x"00000000",
         17677 => x"00000000",
         17678 => x"00000000",
         17679 => x"00000000",
         17680 => x"00000000",
         17681 => x"00000000",
         17682 => x"00000000",
         17683 => x"00000000",
         17684 => x"00000000",
         17685 => x"00000000",
         17686 => x"00000000",
         17687 => x"00000000",
         17688 => x"00000000",
         17689 => x"00000000",
         17690 => x"00000000",
         17691 => x"00000000",
         17692 => x"00000000",
         17693 => x"00000000",
         17694 => x"00000000",
         17695 => x"00000000",
         17696 => x"00000000",
         17697 => x"00000000",
         17698 => x"00000000",
         17699 => x"00000000",
         17700 => x"00000000",
         17701 => x"00000000",
         17702 => x"00000000",
         17703 => x"00000000",
         17704 => x"00000000",
         17705 => x"00000000",
         17706 => x"00000000",
         17707 => x"00000000",
         17708 => x"00000000",
         17709 => x"00000000",
         17710 => x"00000000",
         17711 => x"00000000",
         17712 => x"00000000",
         17713 => x"00000000",
         17714 => x"00000000",
         17715 => x"00000000",
         17716 => x"00000000",
         17717 => x"00000000",
         17718 => x"00000000",
         17719 => x"00000000",
         17720 => x"00000000",
         17721 => x"00000000",
         17722 => x"00000000",
         17723 => x"00000000",
         17724 => x"00000000",
         17725 => x"00000000",
         17726 => x"00000000",
         17727 => x"00000000",
         17728 => x"00000000",
         17729 => x"00000000",
         17730 => x"00000000",
         17731 => x"00000000",
         17732 => x"00000000",
         17733 => x"00000000",
         17734 => x"00000000",
         17735 => x"00000000",
         17736 => x"00000000",
         17737 => x"00000000",
         17738 => x"00000000",
         17739 => x"00000000",
         17740 => x"00000000",
         17741 => x"00000000",
         17742 => x"00000000",
         17743 => x"00000000",
         17744 => x"00000000",
         17745 => x"00000000",
         17746 => x"00000000",
         17747 => x"00000000",
         17748 => x"00000000",
         17749 => x"00000000",
         17750 => x"00000000",
         17751 => x"00000000",
         17752 => x"00000000",
         17753 => x"00000000",
         17754 => x"00000000",
         17755 => x"00000000",
         17756 => x"00000000",
         17757 => x"00000000",
         17758 => x"00000000",
         17759 => x"00000000",
         17760 => x"00000000",
         17761 => x"00000000",
         17762 => x"00000000",
         17763 => x"00000000",
         17764 => x"00000000",
         17765 => x"00000000",
         17766 => x"00000000",
         17767 => x"00000000",
         17768 => x"00000000",
         17769 => x"00000000",
         17770 => x"00000000",
         17771 => x"00000000",
         17772 => x"00000000",
         17773 => x"00000000",
         17774 => x"00000000",
         17775 => x"00000000",
         17776 => x"00000000",
         17777 => x"00000000",
         17778 => x"00000000",
         17779 => x"00000000",
         17780 => x"00000000",
         17781 => x"00000000",
         17782 => x"00000000",
         17783 => x"00000000",
         17784 => x"00000000",
         17785 => x"00000000",
         17786 => x"00000000",
         17787 => x"00000000",
         17788 => x"00000000",
         17789 => x"00000000",
         17790 => x"00000000",
         17791 => x"00000000",
         17792 => x"00000000",
         17793 => x"00000000",
         17794 => x"00000000",
         17795 => x"00000000",
         17796 => x"00000000",
         17797 => x"00000000",
         17798 => x"00000000",
         17799 => x"00000000",
         17800 => x"00000000",
         17801 => x"00000000",
         17802 => x"00000000",
         17803 => x"00000000",
         17804 => x"00000000",
         17805 => x"00000000",
         17806 => x"00000000",
         17807 => x"00000000",
         17808 => x"00000000",
         17809 => x"00000000",
         17810 => x"00000000",
         17811 => x"00000000",
         17812 => x"00000000",
         17813 => x"00000000",
         17814 => x"00000000",
         17815 => x"00000000",
         17816 => x"00000000",
         17817 => x"00000000",
         17818 => x"00000000",
         17819 => x"00000000",
         17820 => x"00000000",
         17821 => x"00000000",
         17822 => x"00000000",
         17823 => x"00000000",
         17824 => x"00000000",
         17825 => x"00000000",
         17826 => x"00000000",
         17827 => x"00000000",
         17828 => x"00000000",
         17829 => x"00000000",
         17830 => x"00000000",
         17831 => x"00000000",
         17832 => x"00000000",
         17833 => x"00000000",
         17834 => x"00000000",
         17835 => x"00000000",
         17836 => x"00000000",
         17837 => x"00000000",
         17838 => x"00000000",
         17839 => x"00000000",
         17840 => x"00000000",
         17841 => x"00000000",
         17842 => x"00000000",
         17843 => x"00000000",
         17844 => x"00000000",
         17845 => x"00000000",
         17846 => x"00000000",
         17847 => x"00000000",
         17848 => x"00000000",
         17849 => x"00000000",
         17850 => x"00000000",
         17851 => x"00000000",
         17852 => x"00000000",
         17853 => x"00000000",
         17854 => x"00000000",
         17855 => x"00000000",
         17856 => x"00000000",
         17857 => x"00000000",
         17858 => x"00000000",
         17859 => x"00000000",
         17860 => x"00000000",
         17861 => x"00000000",
         17862 => x"00000000",
         17863 => x"00000000",
         17864 => x"00000000",
         17865 => x"00000000",
         17866 => x"00000000",
         17867 => x"00000000",
         17868 => x"00000000",
         17869 => x"00000000",
         17870 => x"00000000",
         17871 => x"00000000",
         17872 => x"00000000",
         17873 => x"00000000",
         17874 => x"00000000",
         17875 => x"00000000",
         17876 => x"00000000",
         17877 => x"00000000",
         17878 => x"00000000",
         17879 => x"00000000",
         17880 => x"00000000",
         17881 => x"00000000",
         17882 => x"00000000",
         17883 => x"00000000",
         17884 => x"00000000",
         17885 => x"00000000",
         17886 => x"00000000",
         17887 => x"00000000",
         17888 => x"00000000",
         17889 => x"00000000",
         17890 => x"00000000",
         17891 => x"00000000",
         17892 => x"00000000",
         17893 => x"00000000",
         17894 => x"00000000",
         17895 => x"00000000",
         17896 => x"00000000",
         17897 => x"00000000",
         17898 => x"00000000",
         17899 => x"00000000",
         17900 => x"00000000",
         17901 => x"00000000",
         17902 => x"00000000",
         17903 => x"00000000",
         17904 => x"00000000",
         17905 => x"00000000",
         17906 => x"00000000",
         17907 => x"00000000",
         17908 => x"00000000",
         17909 => x"00000000",
         17910 => x"00000000",
         17911 => x"00000000",
         17912 => x"00000000",
         17913 => x"00000000",
         17914 => x"00000000",
         17915 => x"00000000",
         17916 => x"00000000",
         17917 => x"00000000",
         17918 => x"00000000",
         17919 => x"00000000",
         17920 => x"00000000",
         17921 => x"00000000",
         17922 => x"00000000",
         17923 => x"00000000",
         17924 => x"00000000",
         17925 => x"00000000",
         17926 => x"00000000",
         17927 => x"00000000",
         17928 => x"00000000",
         17929 => x"00000000",
         17930 => x"00000000",
         17931 => x"00000000",
         17932 => x"00000000",
         17933 => x"00000000",
         17934 => x"00000000",
         17935 => x"00000000",
         17936 => x"00000000",
         17937 => x"00000000",
         17938 => x"00000000",
         17939 => x"00000000",
         17940 => x"00000000",
         17941 => x"00000000",
         17942 => x"00000000",
         17943 => x"00000000",
         17944 => x"00000000",
         17945 => x"00000000",
         17946 => x"00000000",
         17947 => x"00000000",
         17948 => x"00000000",
         17949 => x"00000000",
         17950 => x"00000000",
         17951 => x"00000000",
         17952 => x"00000000",
         17953 => x"00000000",
         17954 => x"00000000",
         17955 => x"00000000",
         17956 => x"00000000",
         17957 => x"00000000",
         17958 => x"00000000",
         17959 => x"00000000",
         17960 => x"00000000",
         17961 => x"00000000",
         17962 => x"00000000",
         17963 => x"00000000",
         17964 => x"00000000",
         17965 => x"00000000",
         17966 => x"00000000",
         17967 => x"00000000",
         17968 => x"00000000",
         17969 => x"00000000",
         17970 => x"00000000",
         17971 => x"00000000",
         17972 => x"00000000",
         17973 => x"00000000",
         17974 => x"00000000",
         17975 => x"00000000",
         17976 => x"00000000",
         17977 => x"00000000",
         17978 => x"00000000",
         17979 => x"00000000",
         17980 => x"00000000",
         17981 => x"00000000",
         17982 => x"00000000",
         17983 => x"00000000",
         17984 => x"00000000",
         17985 => x"00000000",
         17986 => x"00000000",
         17987 => x"00000000",
         17988 => x"00000000",
         17989 => x"00000000",
         17990 => x"00000000",
         17991 => x"00000000",
         17992 => x"00000000",
         17993 => x"00000000",
         17994 => x"00000000",
         17995 => x"00000000",
         17996 => x"00000000",
         17997 => x"00000000",
         17998 => x"00000000",
         17999 => x"00000000",
         18000 => x"00000000",
         18001 => x"00000000",
         18002 => x"00000000",
         18003 => x"00000000",
         18004 => x"00000000",
         18005 => x"00000000",
         18006 => x"00000000",
         18007 => x"00000000",
         18008 => x"00000000",
         18009 => x"00000000",
         18010 => x"00000000",
         18011 => x"00000000",
         18012 => x"00000000",
         18013 => x"00000000",
         18014 => x"00000000",
         18015 => x"00000000",
         18016 => x"00000000",
         18017 => x"00000000",
         18018 => x"00000000",
         18019 => x"00000000",
         18020 => x"00000000",
         18021 => x"00000000",
         18022 => x"00000000",
         18023 => x"00000000",
         18024 => x"00000000",
         18025 => x"00000000",
         18026 => x"00000000",
         18027 => x"00000000",
         18028 => x"00000000",
         18029 => x"00000000",
         18030 => x"00000000",
         18031 => x"00000000",
         18032 => x"00000000",
         18033 => x"00000000",
         18034 => x"00000000",
         18035 => x"00000000",
         18036 => x"00000000",
         18037 => x"00000000",
         18038 => x"00000000",
         18039 => x"00000000",
         18040 => x"00000000",
         18041 => x"00000000",
         18042 => x"00000000",
         18043 => x"00000000",
         18044 => x"00000000",
         18045 => x"00000000",
         18046 => x"00000000",
         18047 => x"00000000",
         18048 => x"00000000",
         18049 => x"00000000",
         18050 => x"00000000",
         18051 => x"00000000",
         18052 => x"00000000",
         18053 => x"00000000",
         18054 => x"00000000",
         18055 => x"00000000",
         18056 => x"00000000",
         18057 => x"00000000",
         18058 => x"00000000",
         18059 => x"00000000",
         18060 => x"00000000",
         18061 => x"00000000",
         18062 => x"00000000",
         18063 => x"00000000",
         18064 => x"00000000",
         18065 => x"00000000",
         18066 => x"00000000",
         18067 => x"00000000",
         18068 => x"00000000",
         18069 => x"00000000",
         18070 => x"00000000",
         18071 => x"00000000",
         18072 => x"00000000",
         18073 => x"00000000",
         18074 => x"00000000",
         18075 => x"00000000",
         18076 => x"00000000",
         18077 => x"00000000",
         18078 => x"00000000",
         18079 => x"00000000",
         18080 => x"00000000",
         18081 => x"00000000",
         18082 => x"00000000",
         18083 => x"00000000",
         18084 => x"00000000",
         18085 => x"00000000",
         18086 => x"00000000",
         18087 => x"00000000",
         18088 => x"00000000",
         18089 => x"00000000",
         18090 => x"00000000",
         18091 => x"00000000",
         18092 => x"00000000",
         18093 => x"00000000",
         18094 => x"00000000",
         18095 => x"00000000",
         18096 => x"00000000",
         18097 => x"00000000",
         18098 => x"00000000",
         18099 => x"00000000",
         18100 => x"00000000",
         18101 => x"00000000",
         18102 => x"00000000",
         18103 => x"00000000",
         18104 => x"00000000",
         18105 => x"00000000",
         18106 => x"00000000",
         18107 => x"00000000",
         18108 => x"00000000",
         18109 => x"00000000",
         18110 => x"00000000",
         18111 => x"00000000",
         18112 => x"00000000",
         18113 => x"00000000",
         18114 => x"00000000",
         18115 => x"00000000",
         18116 => x"00000000",
         18117 => x"00000000",
         18118 => x"00000000",
         18119 => x"00000000",
         18120 => x"00000000",
         18121 => x"00000000",
         18122 => x"00000000",
         18123 => x"00000000",
         18124 => x"00000000",
         18125 => x"00000000",
         18126 => x"00000000",
         18127 => x"00000000",
         18128 => x"00000000",
         18129 => x"00000000",
         18130 => x"00000000",
         18131 => x"00000000",
         18132 => x"00000000",
         18133 => x"00000000",
         18134 => x"00000000",
         18135 => x"00000000",
         18136 => x"00000000",
         18137 => x"00000000",
         18138 => x"00000000",
         18139 => x"00000000",
         18140 => x"00000000",
         18141 => x"00000000",
         18142 => x"00000000",
         18143 => x"00000000",
         18144 => x"00000000",
         18145 => x"00000000",
         18146 => x"00000000",
         18147 => x"00000000",
         18148 => x"00000000",
         18149 => x"00000000",
         18150 => x"00000000",
         18151 => x"00000000",
         18152 => x"00000000",
         18153 => x"00000000",
         18154 => x"00000000",
         18155 => x"00000000",
         18156 => x"00000000",
         18157 => x"00000000",
         18158 => x"00000000",
         18159 => x"00000000",
         18160 => x"00000000",
         18161 => x"00000000",
         18162 => x"00000000",
         18163 => x"00000000",
         18164 => x"00000000",
         18165 => x"00000000",
         18166 => x"00000000",
         18167 => x"00000000",
         18168 => x"00000000",
         18169 => x"00000000",
         18170 => x"00000000",
         18171 => x"00000000",
         18172 => x"00000000",
         18173 => x"00000000",
         18174 => x"00000000",
         18175 => x"00003219",
         18176 => x"50000101",
         18177 => x"00000000",
         18178 => x"cce0f2f3",
         18179 => x"cecff6f7",
         18180 => x"f8f9fafb",
         18181 => x"fcfdfeff",
         18182 => x"e1c1c2c3",
         18183 => x"c4c5c6e2",
         18184 => x"e3e4e5e6",
         18185 => x"ebeeeff4",
         18186 => x"00616263",
         18187 => x"64656667",
         18188 => x"68696b6a",
         18189 => x"2f2a2e2d",
         18190 => x"20212223",
         18191 => x"24252627",
         18192 => x"28294f2c",
         18193 => x"512b5749",
         18194 => x"55010203",
         18195 => x"04050607",
         18196 => x"08090a0b",
         18197 => x"0c0d0e0f",
         18198 => x"10111213",
         18199 => x"14151617",
         18200 => x"18191a52",
         18201 => x"5954be3c",
         18202 => x"c7818283",
         18203 => x"84858687",
         18204 => x"88898a8b",
         18205 => x"8c8d8e8f",
         18206 => x"90919293",
         18207 => x"94959697",
         18208 => x"98999abc",
         18209 => x"8040a5c0",
         18210 => x"00000000",
         18211 => x"00000000",
         18212 => x"00000000",
         18213 => x"00000000",
         18214 => x"00000000",
         18215 => x"00000000",
         18216 => x"00000000",
         18217 => x"00000000",
         18218 => x"00000000",
         18219 => x"00000000",
         18220 => x"00000000",
         18221 => x"00000000",
         18222 => x"00000000",
         18223 => x"00000000",
         18224 => x"00000000",
         18225 => x"00000000",
         18226 => x"00000000",
         18227 => x"00000000",
         18228 => x"00000000",
         18229 => x"00000000",
         18230 => x"00000000",
         18231 => x"00000000",
         18232 => x"00000000",
         18233 => x"00000000",
         18234 => x"00000000",
         18235 => x"00000000",
         18236 => x"00000000",
         18237 => x"00000000",
         18238 => x"00000000",
         18239 => x"00000000",
         18240 => x"00020003",
         18241 => x"00040101",
         18242 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

