-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"ff",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"80",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"95",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"c3",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"c5",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"d4",
           386 => x"da",
           387 => x"d4",
           388 => x"90",
           389 => x"d4",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"82",
           395 => x"82",
           396 => x"82",
           397 => x"af",
           398 => x"b5",
           399 => x"d0",
           400 => x"b5",
           401 => x"ad",
           402 => x"d4",
           403 => x"90",
           404 => x"d4",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"82",
           418 => x"82",
           419 => x"82",
           420 => x"96",
           421 => x"b5",
           422 => x"d0",
           423 => x"b5",
           424 => x"cd",
           425 => x"d4",
           426 => x"90",
           427 => x"d4",
           428 => x"84",
           429 => x"d4",
           430 => x"90",
           431 => x"d4",
           432 => x"e2",
           433 => x"d4",
           434 => x"90",
           435 => x"d4",
           436 => x"9f",
           437 => x"d4",
           438 => x"90",
           439 => x"d4",
           440 => x"96",
           441 => x"d4",
           442 => x"90",
           443 => x"d4",
           444 => x"c9",
           445 => x"d4",
           446 => x"90",
           447 => x"d4",
           448 => x"fc",
           449 => x"d4",
           450 => x"90",
           451 => x"d4",
           452 => x"ed",
           453 => x"d4",
           454 => x"90",
           455 => x"d4",
           456 => x"e1",
           457 => x"d4",
           458 => x"90",
           459 => x"d4",
           460 => x"de",
           461 => x"d4",
           462 => x"90",
           463 => x"d4",
           464 => x"fc",
           465 => x"d4",
           466 => x"90",
           467 => x"d4",
           468 => x"dc",
           469 => x"d4",
           470 => x"90",
           471 => x"d4",
           472 => x"cf",
           473 => x"d4",
           474 => x"90",
           475 => x"d4",
           476 => x"9b",
           477 => x"d4",
           478 => x"90",
           479 => x"d4",
           480 => x"ba",
           481 => x"d4",
           482 => x"90",
           483 => x"d4",
           484 => x"d9",
           485 => x"d4",
           486 => x"90",
           487 => x"d4",
           488 => x"c3",
           489 => x"d4",
           490 => x"90",
           491 => x"d4",
           492 => x"a9",
           493 => x"d4",
           494 => x"90",
           495 => x"d4",
           496 => x"97",
           497 => x"d4",
           498 => x"90",
           499 => x"d4",
           500 => x"dd",
           501 => x"d4",
           502 => x"90",
           503 => x"d4",
           504 => x"97",
           505 => x"d4",
           506 => x"90",
           507 => x"d4",
           508 => x"98",
           509 => x"d4",
           510 => x"90",
           511 => x"d4",
           512 => x"cd",
           513 => x"d4",
           514 => x"90",
           515 => x"d4",
           516 => x"a6",
           517 => x"d4",
           518 => x"90",
           519 => x"d4",
           520 => x"d1",
           521 => x"d4",
           522 => x"90",
           523 => x"d4",
           524 => x"b4",
           525 => x"d4",
           526 => x"90",
           527 => x"d4",
           528 => x"89",
           529 => x"d4",
           530 => x"90",
           531 => x"d4",
           532 => x"93",
           533 => x"d4",
           534 => x"90",
           535 => x"d4",
           536 => x"d5",
           537 => x"d4",
           538 => x"90",
           539 => x"d4",
           540 => x"9b",
           541 => x"d4",
           542 => x"90",
           543 => x"d4",
           544 => x"c1",
           545 => x"d4",
           546 => x"90",
           547 => x"d4",
           548 => x"f6",
           549 => x"d4",
           550 => x"90",
           551 => x"d4",
           552 => x"e2",
           553 => x"d4",
           554 => x"90",
           555 => x"d4",
           556 => x"d6",
           557 => x"d4",
           558 => x"90",
           559 => x"d4",
           560 => x"c0",
           561 => x"d4",
           562 => x"90",
           563 => x"d4",
           564 => x"a4",
           565 => x"d4",
           566 => x"90",
           567 => x"d4",
           568 => x"c8",
           569 => x"d4",
           570 => x"90",
           571 => x"d4",
           572 => x"ec",
           573 => x"d4",
           574 => x"90",
           575 => x"d4",
           576 => x"cf",
           577 => x"d4",
           578 => x"90",
           579 => x"d4",
           580 => x"98",
           581 => x"d4",
           582 => x"90",
           583 => x"d4",
           584 => x"ea",
           585 => x"d4",
           586 => x"90",
           587 => x"d4",
           588 => x"92",
           589 => x"d4",
           590 => x"90",
           591 => x"d4",
           592 => x"8a",
           593 => x"d4",
           594 => x"90",
           595 => x"d4",
           596 => x"d4",
           597 => x"d4",
           598 => x"90",
           599 => x"00",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"00",
           609 => x"ff",
           610 => x"06",
           611 => x"83",
           612 => x"10",
           613 => x"fc",
           614 => x"51",
           615 => x"80",
           616 => x"ff",
           617 => x"06",
           618 => x"52",
           619 => x"0a",
           620 => x"38",
           621 => x"51",
           622 => x"c8",
           623 => x"a4",
           624 => x"80",
           625 => x"05",
           626 => x"0b",
           627 => x"04",
           628 => x"80",
           629 => x"00",
           630 => x"08",
           631 => x"d4",
           632 => x"0d",
           633 => x"08",
           634 => x"82",
           635 => x"fc",
           636 => x"b5",
           637 => x"05",
           638 => x"b5",
           639 => x"05",
           640 => x"cd",
           641 => x"54",
           642 => x"82",
           643 => x"70",
           644 => x"08",
           645 => x"82",
           646 => x"f8",
           647 => x"82",
           648 => x"51",
           649 => x"0d",
           650 => x"0c",
           651 => x"d4",
           652 => x"b5",
           653 => x"3d",
           654 => x"d4",
           655 => x"08",
           656 => x"70",
           657 => x"81",
           658 => x"51",
           659 => x"38",
           660 => x"b5",
           661 => x"05",
           662 => x"38",
           663 => x"0b",
           664 => x"08",
           665 => x"81",
           666 => x"b5",
           667 => x"05",
           668 => x"82",
           669 => x"8c",
           670 => x"0b",
           671 => x"08",
           672 => x"82",
           673 => x"88",
           674 => x"b5",
           675 => x"05",
           676 => x"d4",
           677 => x"08",
           678 => x"f6",
           679 => x"82",
           680 => x"8c",
           681 => x"80",
           682 => x"b5",
           683 => x"05",
           684 => x"90",
           685 => x"c8",
           686 => x"b5",
           687 => x"05",
           688 => x"b5",
           689 => x"05",
           690 => x"09",
           691 => x"38",
           692 => x"b5",
           693 => x"05",
           694 => x"39",
           695 => x"08",
           696 => x"82",
           697 => x"f8",
           698 => x"53",
           699 => x"82",
           700 => x"8c",
           701 => x"05",
           702 => x"08",
           703 => x"82",
           704 => x"fc",
           705 => x"05",
           706 => x"08",
           707 => x"ff",
           708 => x"b5",
           709 => x"05",
           710 => x"72",
           711 => x"d4",
           712 => x"08",
           713 => x"d4",
           714 => x"0c",
           715 => x"d4",
           716 => x"08",
           717 => x"0c",
           718 => x"82",
           719 => x"04",
           720 => x"08",
           721 => x"d4",
           722 => x"0d",
           723 => x"b5",
           724 => x"05",
           725 => x"d4",
           726 => x"08",
           727 => x"08",
           728 => x"fe",
           729 => x"b5",
           730 => x"05",
           731 => x"d4",
           732 => x"70",
           733 => x"08",
           734 => x"82",
           735 => x"fc",
           736 => x"82",
           737 => x"8c",
           738 => x"82",
           739 => x"e0",
           740 => x"51",
           741 => x"3f",
           742 => x"08",
           743 => x"d4",
           744 => x"0c",
           745 => x"08",
           746 => x"82",
           747 => x"88",
           748 => x"51",
           749 => x"34",
           750 => x"08",
           751 => x"70",
           752 => x"0c",
           753 => x"0d",
           754 => x"0c",
           755 => x"d4",
           756 => x"b5",
           757 => x"3d",
           758 => x"d4",
           759 => x"70",
           760 => x"08",
           761 => x"82",
           762 => x"fc",
           763 => x"82",
           764 => x"8c",
           765 => x"82",
           766 => x"88",
           767 => x"54",
           768 => x"b5",
           769 => x"82",
           770 => x"f8",
           771 => x"b5",
           772 => x"05",
           773 => x"b5",
           774 => x"54",
           775 => x"82",
           776 => x"04",
           777 => x"08",
           778 => x"d4",
           779 => x"0d",
           780 => x"b5",
           781 => x"05",
           782 => x"d4",
           783 => x"08",
           784 => x"8c",
           785 => x"b5",
           786 => x"05",
           787 => x"33",
           788 => x"70",
           789 => x"81",
           790 => x"51",
           791 => x"80",
           792 => x"ff",
           793 => x"d4",
           794 => x"0c",
           795 => x"82",
           796 => x"8c",
           797 => x"72",
           798 => x"82",
           799 => x"f8",
           800 => x"81",
           801 => x"72",
           802 => x"fa",
           803 => x"d4",
           804 => x"08",
           805 => x"b5",
           806 => x"05",
           807 => x"d4",
           808 => x"22",
           809 => x"51",
           810 => x"2e",
           811 => x"82",
           812 => x"f8",
           813 => x"af",
           814 => x"fc",
           815 => x"d4",
           816 => x"33",
           817 => x"26",
           818 => x"82",
           819 => x"f8",
           820 => x"72",
           821 => x"81",
           822 => x"38",
           823 => x"08",
           824 => x"70",
           825 => x"98",
           826 => x"53",
           827 => x"82",
           828 => x"e4",
           829 => x"83",
           830 => x"32",
           831 => x"51",
           832 => x"72",
           833 => x"38",
           834 => x"08",
           835 => x"70",
           836 => x"51",
           837 => x"b5",
           838 => x"05",
           839 => x"39",
           840 => x"08",
           841 => x"70",
           842 => x"98",
           843 => x"83",
           844 => x"73",
           845 => x"51",
           846 => x"53",
           847 => x"d4",
           848 => x"34",
           849 => x"08",
           850 => x"54",
           851 => x"08",
           852 => x"70",
           853 => x"51",
           854 => x"82",
           855 => x"e8",
           856 => x"b5",
           857 => x"05",
           858 => x"2b",
           859 => x"51",
           860 => x"80",
           861 => x"80",
           862 => x"b5",
           863 => x"05",
           864 => x"d4",
           865 => x"22",
           866 => x"70",
           867 => x"51",
           868 => x"db",
           869 => x"d4",
           870 => x"33",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"b5",
           876 => x"05",
           877 => x"39",
           878 => x"08",
           879 => x"70",
           880 => x"81",
           881 => x"53",
           882 => x"9d",
           883 => x"d4",
           884 => x"33",
           885 => x"70",
           886 => x"51",
           887 => x"38",
           888 => x"b5",
           889 => x"05",
           890 => x"d4",
           891 => x"33",
           892 => x"b5",
           893 => x"05",
           894 => x"b5",
           895 => x"05",
           896 => x"26",
           897 => x"82",
           898 => x"c4",
           899 => x"82",
           900 => x"e4",
           901 => x"51",
           902 => x"72",
           903 => x"d4",
           904 => x"22",
           905 => x"51",
           906 => x"b5",
           907 => x"05",
           908 => x"d4",
           909 => x"22",
           910 => x"51",
           911 => x"b5",
           912 => x"05",
           913 => x"39",
           914 => x"08",
           915 => x"70",
           916 => x"51",
           917 => x"b5",
           918 => x"05",
           919 => x"39",
           920 => x"08",
           921 => x"70",
           922 => x"51",
           923 => x"b5",
           924 => x"05",
           925 => x"39",
           926 => x"08",
           927 => x"70",
           928 => x"53",
           929 => x"d4",
           930 => x"23",
           931 => x"b5",
           932 => x"05",
           933 => x"39",
           934 => x"08",
           935 => x"70",
           936 => x"53",
           937 => x"d4",
           938 => x"23",
           939 => x"bf",
           940 => x"d4",
           941 => x"34",
           942 => x"08",
           943 => x"ff",
           944 => x"72",
           945 => x"08",
           946 => x"80",
           947 => x"b5",
           948 => x"05",
           949 => x"39",
           950 => x"08",
           951 => x"82",
           952 => x"90",
           953 => x"05",
           954 => x"08",
           955 => x"70",
           956 => x"72",
           957 => x"08",
           958 => x"82",
           959 => x"ec",
           960 => x"11",
           961 => x"82",
           962 => x"ec",
           963 => x"ef",
           964 => x"d4",
           965 => x"08",
           966 => x"08",
           967 => x"84",
           968 => x"d4",
           969 => x"0c",
           970 => x"b5",
           971 => x"05",
           972 => x"d4",
           973 => x"22",
           974 => x"70",
           975 => x"51",
           976 => x"80",
           977 => x"82",
           978 => x"e8",
           979 => x"98",
           980 => x"98",
           981 => x"b5",
           982 => x"05",
           983 => x"a2",
           984 => x"b5",
           985 => x"72",
           986 => x"08",
           987 => x"99",
           988 => x"d4",
           989 => x"08",
           990 => x"3f",
           991 => x"08",
           992 => x"b5",
           993 => x"05",
           994 => x"d4",
           995 => x"22",
           996 => x"d4",
           997 => x"22",
           998 => x"54",
           999 => x"b5",
          1000 => x"05",
          1001 => x"39",
          1002 => x"08",
          1003 => x"82",
          1004 => x"90",
          1005 => x"05",
          1006 => x"08",
          1007 => x"70",
          1008 => x"d4",
          1009 => x"0c",
          1010 => x"08",
          1011 => x"70",
          1012 => x"81",
          1013 => x"51",
          1014 => x"2e",
          1015 => x"b5",
          1016 => x"05",
          1017 => x"2b",
          1018 => x"2c",
          1019 => x"d4",
          1020 => x"08",
          1021 => x"c1",
          1022 => x"c8",
          1023 => x"82",
          1024 => x"f4",
          1025 => x"39",
          1026 => x"08",
          1027 => x"51",
          1028 => x"82",
          1029 => x"53",
          1030 => x"d4",
          1031 => x"23",
          1032 => x"08",
          1033 => x"53",
          1034 => x"08",
          1035 => x"73",
          1036 => x"54",
          1037 => x"d4",
          1038 => x"23",
          1039 => x"82",
          1040 => x"e4",
          1041 => x"82",
          1042 => x"06",
          1043 => x"72",
          1044 => x"38",
          1045 => x"08",
          1046 => x"82",
          1047 => x"90",
          1048 => x"05",
          1049 => x"08",
          1050 => x"70",
          1051 => x"d4",
          1052 => x"0c",
          1053 => x"82",
          1054 => x"90",
          1055 => x"b5",
          1056 => x"05",
          1057 => x"82",
          1058 => x"90",
          1059 => x"08",
          1060 => x"08",
          1061 => x"53",
          1062 => x"08",
          1063 => x"82",
          1064 => x"fc",
          1065 => x"b5",
          1066 => x"05",
          1067 => x"a4",
          1068 => x"d4",
          1069 => x"22",
          1070 => x"51",
          1071 => x"b5",
          1072 => x"05",
          1073 => x"d4",
          1074 => x"08",
          1075 => x"d4",
          1076 => x"0c",
          1077 => x"08",
          1078 => x"70",
          1079 => x"51",
          1080 => x"b5",
          1081 => x"05",
          1082 => x"39",
          1083 => x"b5",
          1084 => x"05",
          1085 => x"82",
          1086 => x"e4",
          1087 => x"80",
          1088 => x"53",
          1089 => x"d4",
          1090 => x"23",
          1091 => x"82",
          1092 => x"f8",
          1093 => x"0b",
          1094 => x"08",
          1095 => x"82",
          1096 => x"e4",
          1097 => x"82",
          1098 => x"06",
          1099 => x"72",
          1100 => x"38",
          1101 => x"08",
          1102 => x"82",
          1103 => x"90",
          1104 => x"05",
          1105 => x"08",
          1106 => x"70",
          1107 => x"d4",
          1108 => x"0c",
          1109 => x"82",
          1110 => x"90",
          1111 => x"b5",
          1112 => x"05",
          1113 => x"82",
          1114 => x"90",
          1115 => x"08",
          1116 => x"08",
          1117 => x"53",
          1118 => x"08",
          1119 => x"82",
          1120 => x"fc",
          1121 => x"b5",
          1122 => x"05",
          1123 => x"06",
          1124 => x"82",
          1125 => x"e4",
          1126 => x"b5",
          1127 => x"b5",
          1128 => x"05",
          1129 => x"d4",
          1130 => x"08",
          1131 => x"08",
          1132 => x"82",
          1133 => x"fc",
          1134 => x"55",
          1135 => x"54",
          1136 => x"3f",
          1137 => x"08",
          1138 => x"34",
          1139 => x"08",
          1140 => x"82",
          1141 => x"d4",
          1142 => x"b5",
          1143 => x"05",
          1144 => x"51",
          1145 => x"27",
          1146 => x"b5",
          1147 => x"05",
          1148 => x"33",
          1149 => x"d4",
          1150 => x"33",
          1151 => x"11",
          1152 => x"72",
          1153 => x"08",
          1154 => x"97",
          1155 => x"d4",
          1156 => x"08",
          1157 => x"b0",
          1158 => x"72",
          1159 => x"08",
          1160 => x"82",
          1161 => x"d4",
          1162 => x"82",
          1163 => x"d0",
          1164 => x"34",
          1165 => x"08",
          1166 => x"81",
          1167 => x"d4",
          1168 => x"0c",
          1169 => x"08",
          1170 => x"70",
          1171 => x"d4",
          1172 => x"08",
          1173 => x"ab",
          1174 => x"c8",
          1175 => x"b5",
          1176 => x"05",
          1177 => x"b5",
          1178 => x"05",
          1179 => x"84",
          1180 => x"39",
          1181 => x"08",
          1182 => x"82",
          1183 => x"55",
          1184 => x"70",
          1185 => x"53",
          1186 => x"d4",
          1187 => x"34",
          1188 => x"08",
          1189 => x"70",
          1190 => x"53",
          1191 => x"94",
          1192 => x"d4",
          1193 => x"22",
          1194 => x"53",
          1195 => x"d4",
          1196 => x"23",
          1197 => x"08",
          1198 => x"70",
          1199 => x"81",
          1200 => x"53",
          1201 => x"80",
          1202 => x"b5",
          1203 => x"05",
          1204 => x"2b",
          1205 => x"08",
          1206 => x"82",
          1207 => x"cc",
          1208 => x"2c",
          1209 => x"08",
          1210 => x"82",
          1211 => x"f4",
          1212 => x"53",
          1213 => x"09",
          1214 => x"38",
          1215 => x"08",
          1216 => x"fe",
          1217 => x"82",
          1218 => x"c8",
          1219 => x"39",
          1220 => x"08",
          1221 => x"ff",
          1222 => x"82",
          1223 => x"c8",
          1224 => x"b5",
          1225 => x"05",
          1226 => x"d4",
          1227 => x"23",
          1228 => x"08",
          1229 => x"70",
          1230 => x"81",
          1231 => x"53",
          1232 => x"80",
          1233 => x"b5",
          1234 => x"05",
          1235 => x"2b",
          1236 => x"82",
          1237 => x"fc",
          1238 => x"51",
          1239 => x"74",
          1240 => x"82",
          1241 => x"e4",
          1242 => x"f7",
          1243 => x"72",
          1244 => x"08",
          1245 => x"9d",
          1246 => x"d4",
          1247 => x"33",
          1248 => x"d4",
          1249 => x"33",
          1250 => x"54",
          1251 => x"b5",
          1252 => x"05",
          1253 => x"d4",
          1254 => x"22",
          1255 => x"70",
          1256 => x"51",
          1257 => x"2e",
          1258 => x"b5",
          1259 => x"05",
          1260 => x"2b",
          1261 => x"70",
          1262 => x"88",
          1263 => x"51",
          1264 => x"54",
          1265 => x"08",
          1266 => x"70",
          1267 => x"53",
          1268 => x"d4",
          1269 => x"23",
          1270 => x"b5",
          1271 => x"05",
          1272 => x"2b",
          1273 => x"70",
          1274 => x"88",
          1275 => x"51",
          1276 => x"54",
          1277 => x"08",
          1278 => x"70",
          1279 => x"53",
          1280 => x"d4",
          1281 => x"23",
          1282 => x"08",
          1283 => x"70",
          1284 => x"51",
          1285 => x"38",
          1286 => x"08",
          1287 => x"ff",
          1288 => x"72",
          1289 => x"08",
          1290 => x"73",
          1291 => x"90",
          1292 => x"80",
          1293 => x"38",
          1294 => x"08",
          1295 => x"52",
          1296 => x"ee",
          1297 => x"82",
          1298 => x"e4",
          1299 => x"81",
          1300 => x"06",
          1301 => x"72",
          1302 => x"38",
          1303 => x"08",
          1304 => x"52",
          1305 => x"ca",
          1306 => x"39",
          1307 => x"08",
          1308 => x"70",
          1309 => x"81",
          1310 => x"53",
          1311 => x"90",
          1312 => x"d4",
          1313 => x"08",
          1314 => x"8a",
          1315 => x"39",
          1316 => x"08",
          1317 => x"70",
          1318 => x"81",
          1319 => x"53",
          1320 => x"8e",
          1321 => x"d4",
          1322 => x"08",
          1323 => x"8a",
          1324 => x"b5",
          1325 => x"05",
          1326 => x"2a",
          1327 => x"51",
          1328 => x"80",
          1329 => x"82",
          1330 => x"88",
          1331 => x"b0",
          1332 => x"3f",
          1333 => x"08",
          1334 => x"53",
          1335 => x"09",
          1336 => x"38",
          1337 => x"08",
          1338 => x"52",
          1339 => x"08",
          1340 => x"51",
          1341 => x"82",
          1342 => x"e4",
          1343 => x"88",
          1344 => x"06",
          1345 => x"72",
          1346 => x"38",
          1347 => x"08",
          1348 => x"ff",
          1349 => x"72",
          1350 => x"08",
          1351 => x"73",
          1352 => x"90",
          1353 => x"80",
          1354 => x"38",
          1355 => x"08",
          1356 => x"52",
          1357 => x"fa",
          1358 => x"82",
          1359 => x"e4",
          1360 => x"83",
          1361 => x"06",
          1362 => x"72",
          1363 => x"38",
          1364 => x"08",
          1365 => x"ff",
          1366 => x"72",
          1367 => x"08",
          1368 => x"73",
          1369 => x"98",
          1370 => x"80",
          1371 => x"38",
          1372 => x"08",
          1373 => x"52",
          1374 => x"b6",
          1375 => x"82",
          1376 => x"e4",
          1377 => x"87",
          1378 => x"06",
          1379 => x"72",
          1380 => x"b5",
          1381 => x"05",
          1382 => x"54",
          1383 => x"b5",
          1384 => x"05",
          1385 => x"2b",
          1386 => x"51",
          1387 => x"25",
          1388 => x"b5",
          1389 => x"05",
          1390 => x"51",
          1391 => x"d2",
          1392 => x"d4",
          1393 => x"33",
          1394 => x"e3",
          1395 => x"06",
          1396 => x"b5",
          1397 => x"05",
          1398 => x"b5",
          1399 => x"05",
          1400 => x"ce",
          1401 => x"39",
          1402 => x"08",
          1403 => x"53",
          1404 => x"2e",
          1405 => x"80",
          1406 => x"b5",
          1407 => x"05",
          1408 => x"51",
          1409 => x"b5",
          1410 => x"05",
          1411 => x"ff",
          1412 => x"72",
          1413 => x"2e",
          1414 => x"82",
          1415 => x"88",
          1416 => x"82",
          1417 => x"fc",
          1418 => x"33",
          1419 => x"d4",
          1420 => x"08",
          1421 => x"b5",
          1422 => x"05",
          1423 => x"f2",
          1424 => x"39",
          1425 => x"08",
          1426 => x"53",
          1427 => x"2e",
          1428 => x"80",
          1429 => x"b5",
          1430 => x"05",
          1431 => x"51",
          1432 => x"b5",
          1433 => x"05",
          1434 => x"ff",
          1435 => x"72",
          1436 => x"2e",
          1437 => x"82",
          1438 => x"88",
          1439 => x"82",
          1440 => x"fc",
          1441 => x"33",
          1442 => x"a6",
          1443 => x"d4",
          1444 => x"08",
          1445 => x"b5",
          1446 => x"05",
          1447 => x"39",
          1448 => x"08",
          1449 => x"82",
          1450 => x"a9",
          1451 => x"d4",
          1452 => x"08",
          1453 => x"d4",
          1454 => x"08",
          1455 => x"b5",
          1456 => x"05",
          1457 => x"d4",
          1458 => x"08",
          1459 => x"53",
          1460 => x"cc",
          1461 => x"d4",
          1462 => x"22",
          1463 => x"70",
          1464 => x"51",
          1465 => x"2e",
          1466 => x"82",
          1467 => x"ec",
          1468 => x"11",
          1469 => x"82",
          1470 => x"ec",
          1471 => x"90",
          1472 => x"2c",
          1473 => x"73",
          1474 => x"82",
          1475 => x"88",
          1476 => x"a0",
          1477 => x"3f",
          1478 => x"b5",
          1479 => x"05",
          1480 => x"b5",
          1481 => x"05",
          1482 => x"86",
          1483 => x"82",
          1484 => x"e4",
          1485 => x"b7",
          1486 => x"d4",
          1487 => x"33",
          1488 => x"2e",
          1489 => x"a8",
          1490 => x"82",
          1491 => x"e4",
          1492 => x"0b",
          1493 => x"08",
          1494 => x"80",
          1495 => x"d4",
          1496 => x"34",
          1497 => x"b5",
          1498 => x"05",
          1499 => x"39",
          1500 => x"08",
          1501 => x"52",
          1502 => x"08",
          1503 => x"51",
          1504 => x"e9",
          1505 => x"b5",
          1506 => x"05",
          1507 => x"08",
          1508 => x"d4",
          1509 => x"0c",
          1510 => x"b5",
          1511 => x"05",
          1512 => x"c8",
          1513 => x"0d",
          1514 => x"0c",
          1515 => x"d4",
          1516 => x"b5",
          1517 => x"3d",
          1518 => x"98",
          1519 => x"b5",
          1520 => x"05",
          1521 => x"b5",
          1522 => x"05",
          1523 => x"dd",
          1524 => x"c8",
          1525 => x"b5",
          1526 => x"85",
          1527 => x"b5",
          1528 => x"82",
          1529 => x"02",
          1530 => x"0c",
          1531 => x"80",
          1532 => x"d4",
          1533 => x"0c",
          1534 => x"08",
          1535 => x"70",
          1536 => x"81",
          1537 => x"06",
          1538 => x"51",
          1539 => x"2e",
          1540 => x"0b",
          1541 => x"08",
          1542 => x"81",
          1543 => x"b5",
          1544 => x"05",
          1545 => x"33",
          1546 => x"08",
          1547 => x"81",
          1548 => x"d4",
          1549 => x"0c",
          1550 => x"b5",
          1551 => x"05",
          1552 => x"ff",
          1553 => x"80",
          1554 => x"82",
          1555 => x"82",
          1556 => x"53",
          1557 => x"08",
          1558 => x"52",
          1559 => x"51",
          1560 => x"82",
          1561 => x"53",
          1562 => x"ff",
          1563 => x"0b",
          1564 => x"08",
          1565 => x"ff",
          1566 => x"cd",
          1567 => x"cd",
          1568 => x"53",
          1569 => x"13",
          1570 => x"2d",
          1571 => x"08",
          1572 => x"2e",
          1573 => x"0b",
          1574 => x"08",
          1575 => x"82",
          1576 => x"f8",
          1577 => x"82",
          1578 => x"f4",
          1579 => x"82",
          1580 => x"f4",
          1581 => x"b5",
          1582 => x"3d",
          1583 => x"d4",
          1584 => x"b5",
          1585 => x"82",
          1586 => x"fb",
          1587 => x"0b",
          1588 => x"08",
          1589 => x"82",
          1590 => x"8c",
          1591 => x"11",
          1592 => x"2a",
          1593 => x"70",
          1594 => x"51",
          1595 => x"72",
          1596 => x"38",
          1597 => x"b5",
          1598 => x"05",
          1599 => x"39",
          1600 => x"08",
          1601 => x"53",
          1602 => x"b5",
          1603 => x"05",
          1604 => x"82",
          1605 => x"88",
          1606 => x"72",
          1607 => x"08",
          1608 => x"72",
          1609 => x"53",
          1610 => x"b6",
          1611 => x"d4",
          1612 => x"08",
          1613 => x"08",
          1614 => x"53",
          1615 => x"08",
          1616 => x"52",
          1617 => x"51",
          1618 => x"82",
          1619 => x"53",
          1620 => x"ff",
          1621 => x"0b",
          1622 => x"08",
          1623 => x"ff",
          1624 => x"b5",
          1625 => x"05",
          1626 => x"b5",
          1627 => x"05",
          1628 => x"b5",
          1629 => x"05",
          1630 => x"c8",
          1631 => x"0d",
          1632 => x"0c",
          1633 => x"d4",
          1634 => x"b5",
          1635 => x"3d",
          1636 => x"9c",
          1637 => x"b5",
          1638 => x"05",
          1639 => x"3f",
          1640 => x"08",
          1641 => x"c8",
          1642 => x"3d",
          1643 => x"d4",
          1644 => x"b5",
          1645 => x"82",
          1646 => x"fb",
          1647 => x"b5",
          1648 => x"05",
          1649 => x"33",
          1650 => x"70",
          1651 => x"81",
          1652 => x"51",
          1653 => x"80",
          1654 => x"ff",
          1655 => x"d4",
          1656 => x"0c",
          1657 => x"82",
          1658 => x"8c",
          1659 => x"11",
          1660 => x"2a",
          1661 => x"51",
          1662 => x"72",
          1663 => x"db",
          1664 => x"d4",
          1665 => x"08",
          1666 => x"08",
          1667 => x"54",
          1668 => x"08",
          1669 => x"25",
          1670 => x"b5",
          1671 => x"05",
          1672 => x"70",
          1673 => x"08",
          1674 => x"52",
          1675 => x"72",
          1676 => x"08",
          1677 => x"0c",
          1678 => x"08",
          1679 => x"8c",
          1680 => x"05",
          1681 => x"82",
          1682 => x"88",
          1683 => x"82",
          1684 => x"fc",
          1685 => x"53",
          1686 => x"82",
          1687 => x"8c",
          1688 => x"b5",
          1689 => x"05",
          1690 => x"b5",
          1691 => x"05",
          1692 => x"ff",
          1693 => x"12",
          1694 => x"54",
          1695 => x"b5",
          1696 => x"72",
          1697 => x"b5",
          1698 => x"05",
          1699 => x"08",
          1700 => x"12",
          1701 => x"d4",
          1702 => x"08",
          1703 => x"d4",
          1704 => x"0c",
          1705 => x"39",
          1706 => x"b5",
          1707 => x"05",
          1708 => x"d4",
          1709 => x"08",
          1710 => x"0c",
          1711 => x"82",
          1712 => x"04",
          1713 => x"08",
          1714 => x"d4",
          1715 => x"0d",
          1716 => x"08",
          1717 => x"85",
          1718 => x"81",
          1719 => x"06",
          1720 => x"52",
          1721 => x"8d",
          1722 => x"82",
          1723 => x"f8",
          1724 => x"94",
          1725 => x"d4",
          1726 => x"08",
          1727 => x"70",
          1728 => x"81",
          1729 => x"51",
          1730 => x"2e",
          1731 => x"82",
          1732 => x"88",
          1733 => x"b5",
          1734 => x"05",
          1735 => x"85",
          1736 => x"ff",
          1737 => x"52",
          1738 => x"34",
          1739 => x"08",
          1740 => x"8c",
          1741 => x"05",
          1742 => x"82",
          1743 => x"88",
          1744 => x"11",
          1745 => x"b5",
          1746 => x"05",
          1747 => x"52",
          1748 => x"82",
          1749 => x"88",
          1750 => x"11",
          1751 => x"2a",
          1752 => x"51",
          1753 => x"71",
          1754 => x"d7",
          1755 => x"d4",
          1756 => x"08",
          1757 => x"33",
          1758 => x"08",
          1759 => x"51",
          1760 => x"d4",
          1761 => x"08",
          1762 => x"b5",
          1763 => x"05",
          1764 => x"d4",
          1765 => x"08",
          1766 => x"12",
          1767 => x"07",
          1768 => x"85",
          1769 => x"0b",
          1770 => x"08",
          1771 => x"81",
          1772 => x"b5",
          1773 => x"05",
          1774 => x"81",
          1775 => x"52",
          1776 => x"82",
          1777 => x"88",
          1778 => x"b5",
          1779 => x"05",
          1780 => x"11",
          1781 => x"71",
          1782 => x"c8",
          1783 => x"b5",
          1784 => x"05",
          1785 => x"b5",
          1786 => x"05",
          1787 => x"80",
          1788 => x"b5",
          1789 => x"05",
          1790 => x"d4",
          1791 => x"0c",
          1792 => x"08",
          1793 => x"85",
          1794 => x"b5",
          1795 => x"05",
          1796 => x"b5",
          1797 => x"05",
          1798 => x"09",
          1799 => x"38",
          1800 => x"08",
          1801 => x"90",
          1802 => x"82",
          1803 => x"ec",
          1804 => x"39",
          1805 => x"08",
          1806 => x"a0",
          1807 => x"82",
          1808 => x"ec",
          1809 => x"b5",
          1810 => x"05",
          1811 => x"b5",
          1812 => x"05",
          1813 => x"34",
          1814 => x"b5",
          1815 => x"05",
          1816 => x"82",
          1817 => x"88",
          1818 => x"11",
          1819 => x"8c",
          1820 => x"b5",
          1821 => x"05",
          1822 => x"ff",
          1823 => x"b5",
          1824 => x"05",
          1825 => x"52",
          1826 => x"08",
          1827 => x"82",
          1828 => x"89",
          1829 => x"b5",
          1830 => x"82",
          1831 => x"02",
          1832 => x"0c",
          1833 => x"82",
          1834 => x"88",
          1835 => x"b5",
          1836 => x"05",
          1837 => x"d4",
          1838 => x"08",
          1839 => x"08",
          1840 => x"82",
          1841 => x"90",
          1842 => x"2e",
          1843 => x"82",
          1844 => x"f8",
          1845 => x"b5",
          1846 => x"05",
          1847 => x"ac",
          1848 => x"d4",
          1849 => x"08",
          1850 => x"08",
          1851 => x"05",
          1852 => x"d4",
          1853 => x"08",
          1854 => x"90",
          1855 => x"d4",
          1856 => x"08",
          1857 => x"08",
          1858 => x"05",
          1859 => x"08",
          1860 => x"82",
          1861 => x"f8",
          1862 => x"b5",
          1863 => x"05",
          1864 => x"b5",
          1865 => x"05",
          1866 => x"d4",
          1867 => x"08",
          1868 => x"b5",
          1869 => x"05",
          1870 => x"d4",
          1871 => x"08",
          1872 => x"b5",
          1873 => x"05",
          1874 => x"d4",
          1875 => x"08",
          1876 => x"9c",
          1877 => x"d4",
          1878 => x"08",
          1879 => x"b5",
          1880 => x"05",
          1881 => x"d4",
          1882 => x"08",
          1883 => x"b5",
          1884 => x"05",
          1885 => x"d4",
          1886 => x"08",
          1887 => x"08",
          1888 => x"53",
          1889 => x"71",
          1890 => x"39",
          1891 => x"08",
          1892 => x"81",
          1893 => x"d4",
          1894 => x"0c",
          1895 => x"08",
          1896 => x"ff",
          1897 => x"d4",
          1898 => x"0c",
          1899 => x"08",
          1900 => x"80",
          1901 => x"82",
          1902 => x"f8",
          1903 => x"70",
          1904 => x"d4",
          1905 => x"08",
          1906 => x"b5",
          1907 => x"05",
          1908 => x"d4",
          1909 => x"08",
          1910 => x"71",
          1911 => x"d4",
          1912 => x"08",
          1913 => x"b5",
          1914 => x"05",
          1915 => x"39",
          1916 => x"08",
          1917 => x"70",
          1918 => x"0c",
          1919 => x"0d",
          1920 => x"0c",
          1921 => x"d4",
          1922 => x"b5",
          1923 => x"3d",
          1924 => x"d4",
          1925 => x"08",
          1926 => x"08",
          1927 => x"82",
          1928 => x"fc",
          1929 => x"71",
          1930 => x"d4",
          1931 => x"08",
          1932 => x"b5",
          1933 => x"05",
          1934 => x"ff",
          1935 => x"70",
          1936 => x"38",
          1937 => x"b5",
          1938 => x"05",
          1939 => x"82",
          1940 => x"fc",
          1941 => x"b5",
          1942 => x"05",
          1943 => x"d4",
          1944 => x"08",
          1945 => x"b5",
          1946 => x"84",
          1947 => x"b5",
          1948 => x"82",
          1949 => x"02",
          1950 => x"0c",
          1951 => x"82",
          1952 => x"88",
          1953 => x"b5",
          1954 => x"05",
          1955 => x"d4",
          1956 => x"08",
          1957 => x"82",
          1958 => x"8c",
          1959 => x"05",
          1960 => x"08",
          1961 => x"82",
          1962 => x"fc",
          1963 => x"51",
          1964 => x"82",
          1965 => x"fc",
          1966 => x"05",
          1967 => x"08",
          1968 => x"70",
          1969 => x"51",
          1970 => x"84",
          1971 => x"39",
          1972 => x"08",
          1973 => x"70",
          1974 => x"0c",
          1975 => x"0d",
          1976 => x"0c",
          1977 => x"d4",
          1978 => x"b5",
          1979 => x"3d",
          1980 => x"d4",
          1981 => x"08",
          1982 => x"08",
          1983 => x"82",
          1984 => x"8c",
          1985 => x"b5",
          1986 => x"05",
          1987 => x"d4",
          1988 => x"08",
          1989 => x"e5",
          1990 => x"d4",
          1991 => x"08",
          1992 => x"b5",
          1993 => x"05",
          1994 => x"d4",
          1995 => x"08",
          1996 => x"b5",
          1997 => x"05",
          1998 => x"d4",
          1999 => x"08",
          2000 => x"38",
          2001 => x"08",
          2002 => x"51",
          2003 => x"b5",
          2004 => x"05",
          2005 => x"82",
          2006 => x"f8",
          2007 => x"b5",
          2008 => x"05",
          2009 => x"71",
          2010 => x"b5",
          2011 => x"05",
          2012 => x"82",
          2013 => x"fc",
          2014 => x"ad",
          2015 => x"d4",
          2016 => x"08",
          2017 => x"c8",
          2018 => x"3d",
          2019 => x"d4",
          2020 => x"b5",
          2021 => x"82",
          2022 => x"fd",
          2023 => x"b5",
          2024 => x"05",
          2025 => x"81",
          2026 => x"b5",
          2027 => x"05",
          2028 => x"33",
          2029 => x"08",
          2030 => x"81",
          2031 => x"d4",
          2032 => x"0c",
          2033 => x"08",
          2034 => x"70",
          2035 => x"ff",
          2036 => x"54",
          2037 => x"2e",
          2038 => x"ce",
          2039 => x"d4",
          2040 => x"08",
          2041 => x"82",
          2042 => x"88",
          2043 => x"05",
          2044 => x"08",
          2045 => x"70",
          2046 => x"51",
          2047 => x"38",
          2048 => x"b5",
          2049 => x"05",
          2050 => x"39",
          2051 => x"08",
          2052 => x"ff",
          2053 => x"d4",
          2054 => x"0c",
          2055 => x"08",
          2056 => x"80",
          2057 => x"ff",
          2058 => x"b5",
          2059 => x"05",
          2060 => x"80",
          2061 => x"b5",
          2062 => x"05",
          2063 => x"52",
          2064 => x"38",
          2065 => x"b5",
          2066 => x"05",
          2067 => x"39",
          2068 => x"08",
          2069 => x"ff",
          2070 => x"d4",
          2071 => x"0c",
          2072 => x"08",
          2073 => x"70",
          2074 => x"70",
          2075 => x"0b",
          2076 => x"08",
          2077 => x"ae",
          2078 => x"d4",
          2079 => x"08",
          2080 => x"b5",
          2081 => x"05",
          2082 => x"72",
          2083 => x"82",
          2084 => x"fc",
          2085 => x"55",
          2086 => x"8a",
          2087 => x"82",
          2088 => x"fc",
          2089 => x"b5",
          2090 => x"05",
          2091 => x"c8",
          2092 => x"0d",
          2093 => x"0c",
          2094 => x"d4",
          2095 => x"b5",
          2096 => x"3d",
          2097 => x"d4",
          2098 => x"08",
          2099 => x"08",
          2100 => x"82",
          2101 => x"8c",
          2102 => x"38",
          2103 => x"b5",
          2104 => x"05",
          2105 => x"39",
          2106 => x"08",
          2107 => x"52",
          2108 => x"b5",
          2109 => x"05",
          2110 => x"82",
          2111 => x"f8",
          2112 => x"81",
          2113 => x"51",
          2114 => x"9f",
          2115 => x"d4",
          2116 => x"08",
          2117 => x"b5",
          2118 => x"05",
          2119 => x"d4",
          2120 => x"08",
          2121 => x"38",
          2122 => x"82",
          2123 => x"f8",
          2124 => x"05",
          2125 => x"08",
          2126 => x"82",
          2127 => x"f8",
          2128 => x"b5",
          2129 => x"05",
          2130 => x"82",
          2131 => x"fc",
          2132 => x"82",
          2133 => x"fc",
          2134 => x"b5",
          2135 => x"3d",
          2136 => x"d4",
          2137 => x"b5",
          2138 => x"82",
          2139 => x"fe",
          2140 => x"b5",
          2141 => x"05",
          2142 => x"d4",
          2143 => x"0c",
          2144 => x"08",
          2145 => x"80",
          2146 => x"38",
          2147 => x"08",
          2148 => x"81",
          2149 => x"d4",
          2150 => x"0c",
          2151 => x"08",
          2152 => x"ff",
          2153 => x"d4",
          2154 => x"0c",
          2155 => x"08",
          2156 => x"80",
          2157 => x"82",
          2158 => x"8c",
          2159 => x"70",
          2160 => x"08",
          2161 => x"52",
          2162 => x"34",
          2163 => x"08",
          2164 => x"81",
          2165 => x"d4",
          2166 => x"0c",
          2167 => x"82",
          2168 => x"88",
          2169 => x"82",
          2170 => x"51",
          2171 => x"82",
          2172 => x"04",
          2173 => x"08",
          2174 => x"d4",
          2175 => x"0d",
          2176 => x"b5",
          2177 => x"05",
          2178 => x"d4",
          2179 => x"08",
          2180 => x"38",
          2181 => x"08",
          2182 => x"30",
          2183 => x"08",
          2184 => x"80",
          2185 => x"d4",
          2186 => x"0c",
          2187 => x"08",
          2188 => x"8a",
          2189 => x"82",
          2190 => x"f4",
          2191 => x"b5",
          2192 => x"05",
          2193 => x"d4",
          2194 => x"0c",
          2195 => x"08",
          2196 => x"80",
          2197 => x"82",
          2198 => x"8c",
          2199 => x"82",
          2200 => x"8c",
          2201 => x"0b",
          2202 => x"08",
          2203 => x"82",
          2204 => x"fc",
          2205 => x"38",
          2206 => x"b5",
          2207 => x"05",
          2208 => x"d4",
          2209 => x"08",
          2210 => x"08",
          2211 => x"80",
          2212 => x"d4",
          2213 => x"08",
          2214 => x"d4",
          2215 => x"08",
          2216 => x"3f",
          2217 => x"08",
          2218 => x"d4",
          2219 => x"0c",
          2220 => x"d4",
          2221 => x"08",
          2222 => x"38",
          2223 => x"08",
          2224 => x"30",
          2225 => x"08",
          2226 => x"82",
          2227 => x"f8",
          2228 => x"82",
          2229 => x"54",
          2230 => x"82",
          2231 => x"04",
          2232 => x"08",
          2233 => x"d4",
          2234 => x"0d",
          2235 => x"b5",
          2236 => x"05",
          2237 => x"d4",
          2238 => x"08",
          2239 => x"38",
          2240 => x"08",
          2241 => x"30",
          2242 => x"08",
          2243 => x"81",
          2244 => x"d4",
          2245 => x"0c",
          2246 => x"08",
          2247 => x"80",
          2248 => x"82",
          2249 => x"8c",
          2250 => x"82",
          2251 => x"8c",
          2252 => x"53",
          2253 => x"08",
          2254 => x"52",
          2255 => x"08",
          2256 => x"51",
          2257 => x"82",
          2258 => x"70",
          2259 => x"08",
          2260 => x"54",
          2261 => x"08",
          2262 => x"80",
          2263 => x"82",
          2264 => x"f8",
          2265 => x"82",
          2266 => x"f8",
          2267 => x"b5",
          2268 => x"05",
          2269 => x"b5",
          2270 => x"87",
          2271 => x"b5",
          2272 => x"82",
          2273 => x"02",
          2274 => x"0c",
          2275 => x"80",
          2276 => x"d4",
          2277 => x"08",
          2278 => x"d4",
          2279 => x"08",
          2280 => x"3f",
          2281 => x"08",
          2282 => x"c8",
          2283 => x"3d",
          2284 => x"d4",
          2285 => x"b5",
          2286 => x"82",
          2287 => x"fd",
          2288 => x"53",
          2289 => x"08",
          2290 => x"52",
          2291 => x"08",
          2292 => x"51",
          2293 => x"b5",
          2294 => x"82",
          2295 => x"54",
          2296 => x"82",
          2297 => x"04",
          2298 => x"08",
          2299 => x"d4",
          2300 => x"0d",
          2301 => x"b5",
          2302 => x"05",
          2303 => x"82",
          2304 => x"f8",
          2305 => x"b5",
          2306 => x"05",
          2307 => x"d4",
          2308 => x"08",
          2309 => x"82",
          2310 => x"fc",
          2311 => x"2e",
          2312 => x"0b",
          2313 => x"08",
          2314 => x"24",
          2315 => x"b5",
          2316 => x"05",
          2317 => x"b5",
          2318 => x"05",
          2319 => x"d4",
          2320 => x"08",
          2321 => x"d4",
          2322 => x"0c",
          2323 => x"82",
          2324 => x"fc",
          2325 => x"2e",
          2326 => x"82",
          2327 => x"8c",
          2328 => x"b5",
          2329 => x"05",
          2330 => x"38",
          2331 => x"08",
          2332 => x"82",
          2333 => x"8c",
          2334 => x"82",
          2335 => x"88",
          2336 => x"b5",
          2337 => x"05",
          2338 => x"d4",
          2339 => x"08",
          2340 => x"d4",
          2341 => x"0c",
          2342 => x"08",
          2343 => x"81",
          2344 => x"d4",
          2345 => x"0c",
          2346 => x"08",
          2347 => x"81",
          2348 => x"d4",
          2349 => x"0c",
          2350 => x"82",
          2351 => x"90",
          2352 => x"2e",
          2353 => x"b5",
          2354 => x"05",
          2355 => x"b5",
          2356 => x"05",
          2357 => x"39",
          2358 => x"08",
          2359 => x"70",
          2360 => x"08",
          2361 => x"51",
          2362 => x"08",
          2363 => x"82",
          2364 => x"85",
          2365 => x"b5",
          2366 => x"82",
          2367 => x"02",
          2368 => x"0c",
          2369 => x"80",
          2370 => x"d4",
          2371 => x"34",
          2372 => x"08",
          2373 => x"53",
          2374 => x"82",
          2375 => x"88",
          2376 => x"08",
          2377 => x"33",
          2378 => x"b5",
          2379 => x"05",
          2380 => x"ff",
          2381 => x"a0",
          2382 => x"06",
          2383 => x"b5",
          2384 => x"05",
          2385 => x"81",
          2386 => x"53",
          2387 => x"b5",
          2388 => x"05",
          2389 => x"ad",
          2390 => x"06",
          2391 => x"0b",
          2392 => x"08",
          2393 => x"82",
          2394 => x"88",
          2395 => x"08",
          2396 => x"0c",
          2397 => x"53",
          2398 => x"b5",
          2399 => x"05",
          2400 => x"d4",
          2401 => x"33",
          2402 => x"2e",
          2403 => x"81",
          2404 => x"b5",
          2405 => x"05",
          2406 => x"81",
          2407 => x"70",
          2408 => x"72",
          2409 => x"d4",
          2410 => x"34",
          2411 => x"08",
          2412 => x"82",
          2413 => x"e8",
          2414 => x"b5",
          2415 => x"05",
          2416 => x"2e",
          2417 => x"b5",
          2418 => x"05",
          2419 => x"2e",
          2420 => x"cd",
          2421 => x"82",
          2422 => x"f4",
          2423 => x"b5",
          2424 => x"05",
          2425 => x"81",
          2426 => x"70",
          2427 => x"72",
          2428 => x"d4",
          2429 => x"34",
          2430 => x"82",
          2431 => x"d4",
          2432 => x"34",
          2433 => x"08",
          2434 => x"70",
          2435 => x"71",
          2436 => x"51",
          2437 => x"82",
          2438 => x"f8",
          2439 => x"fe",
          2440 => x"d4",
          2441 => x"33",
          2442 => x"26",
          2443 => x"0b",
          2444 => x"08",
          2445 => x"83",
          2446 => x"b5",
          2447 => x"05",
          2448 => x"73",
          2449 => x"82",
          2450 => x"f8",
          2451 => x"72",
          2452 => x"38",
          2453 => x"0b",
          2454 => x"08",
          2455 => x"82",
          2456 => x"0b",
          2457 => x"08",
          2458 => x"b2",
          2459 => x"d4",
          2460 => x"33",
          2461 => x"27",
          2462 => x"b5",
          2463 => x"05",
          2464 => x"b9",
          2465 => x"8d",
          2466 => x"82",
          2467 => x"ec",
          2468 => x"a5",
          2469 => x"82",
          2470 => x"f4",
          2471 => x"0b",
          2472 => x"08",
          2473 => x"82",
          2474 => x"f8",
          2475 => x"a0",
          2476 => x"cf",
          2477 => x"d4",
          2478 => x"33",
          2479 => x"73",
          2480 => x"82",
          2481 => x"f8",
          2482 => x"11",
          2483 => x"82",
          2484 => x"f8",
          2485 => x"b5",
          2486 => x"05",
          2487 => x"51",
          2488 => x"b5",
          2489 => x"05",
          2490 => x"d4",
          2491 => x"33",
          2492 => x"27",
          2493 => x"b5",
          2494 => x"05",
          2495 => x"51",
          2496 => x"b5",
          2497 => x"05",
          2498 => x"d4",
          2499 => x"33",
          2500 => x"26",
          2501 => x"0b",
          2502 => x"08",
          2503 => x"81",
          2504 => x"b5",
          2505 => x"05",
          2506 => x"d4",
          2507 => x"33",
          2508 => x"74",
          2509 => x"80",
          2510 => x"d4",
          2511 => x"0c",
          2512 => x"82",
          2513 => x"f4",
          2514 => x"82",
          2515 => x"fc",
          2516 => x"82",
          2517 => x"f8",
          2518 => x"12",
          2519 => x"08",
          2520 => x"82",
          2521 => x"88",
          2522 => x"08",
          2523 => x"0c",
          2524 => x"51",
          2525 => x"72",
          2526 => x"d4",
          2527 => x"34",
          2528 => x"82",
          2529 => x"f0",
          2530 => x"72",
          2531 => x"38",
          2532 => x"08",
          2533 => x"30",
          2534 => x"08",
          2535 => x"82",
          2536 => x"8c",
          2537 => x"b5",
          2538 => x"05",
          2539 => x"53",
          2540 => x"b5",
          2541 => x"05",
          2542 => x"d4",
          2543 => x"08",
          2544 => x"0c",
          2545 => x"82",
          2546 => x"04",
          2547 => x"08",
          2548 => x"d4",
          2549 => x"0d",
          2550 => x"b5",
          2551 => x"05",
          2552 => x"d4",
          2553 => x"08",
          2554 => x"0c",
          2555 => x"08",
          2556 => x"70",
          2557 => x"72",
          2558 => x"82",
          2559 => x"f8",
          2560 => x"81",
          2561 => x"72",
          2562 => x"81",
          2563 => x"82",
          2564 => x"88",
          2565 => x"08",
          2566 => x"0c",
          2567 => x"82",
          2568 => x"f8",
          2569 => x"72",
          2570 => x"81",
          2571 => x"81",
          2572 => x"d4",
          2573 => x"34",
          2574 => x"08",
          2575 => x"70",
          2576 => x"71",
          2577 => x"51",
          2578 => x"82",
          2579 => x"f8",
          2580 => x"b5",
          2581 => x"05",
          2582 => x"b0",
          2583 => x"06",
          2584 => x"82",
          2585 => x"88",
          2586 => x"08",
          2587 => x"0c",
          2588 => x"53",
          2589 => x"b5",
          2590 => x"05",
          2591 => x"d4",
          2592 => x"33",
          2593 => x"08",
          2594 => x"82",
          2595 => x"e8",
          2596 => x"e2",
          2597 => x"82",
          2598 => x"e8",
          2599 => x"f8",
          2600 => x"80",
          2601 => x"0b",
          2602 => x"08",
          2603 => x"82",
          2604 => x"88",
          2605 => x"08",
          2606 => x"0c",
          2607 => x"53",
          2608 => x"b5",
          2609 => x"05",
          2610 => x"39",
          2611 => x"b5",
          2612 => x"05",
          2613 => x"d4",
          2614 => x"08",
          2615 => x"05",
          2616 => x"08",
          2617 => x"33",
          2618 => x"08",
          2619 => x"80",
          2620 => x"b5",
          2621 => x"05",
          2622 => x"a0",
          2623 => x"81",
          2624 => x"d4",
          2625 => x"0c",
          2626 => x"82",
          2627 => x"f8",
          2628 => x"af",
          2629 => x"38",
          2630 => x"08",
          2631 => x"53",
          2632 => x"83",
          2633 => x"80",
          2634 => x"d4",
          2635 => x"0c",
          2636 => x"88",
          2637 => x"d4",
          2638 => x"34",
          2639 => x"b5",
          2640 => x"05",
          2641 => x"73",
          2642 => x"82",
          2643 => x"f8",
          2644 => x"72",
          2645 => x"38",
          2646 => x"0b",
          2647 => x"08",
          2648 => x"82",
          2649 => x"0b",
          2650 => x"08",
          2651 => x"80",
          2652 => x"d4",
          2653 => x"0c",
          2654 => x"08",
          2655 => x"53",
          2656 => x"81",
          2657 => x"b5",
          2658 => x"05",
          2659 => x"e0",
          2660 => x"38",
          2661 => x"08",
          2662 => x"e0",
          2663 => x"72",
          2664 => x"08",
          2665 => x"82",
          2666 => x"f8",
          2667 => x"11",
          2668 => x"82",
          2669 => x"f8",
          2670 => x"b5",
          2671 => x"05",
          2672 => x"73",
          2673 => x"82",
          2674 => x"f8",
          2675 => x"11",
          2676 => x"82",
          2677 => x"f8",
          2678 => x"b5",
          2679 => x"05",
          2680 => x"89",
          2681 => x"80",
          2682 => x"d4",
          2683 => x"0c",
          2684 => x"82",
          2685 => x"f8",
          2686 => x"b5",
          2687 => x"05",
          2688 => x"72",
          2689 => x"38",
          2690 => x"b5",
          2691 => x"05",
          2692 => x"39",
          2693 => x"08",
          2694 => x"70",
          2695 => x"08",
          2696 => x"29",
          2697 => x"08",
          2698 => x"70",
          2699 => x"d4",
          2700 => x"0c",
          2701 => x"08",
          2702 => x"70",
          2703 => x"71",
          2704 => x"51",
          2705 => x"53",
          2706 => x"b5",
          2707 => x"05",
          2708 => x"39",
          2709 => x"08",
          2710 => x"53",
          2711 => x"90",
          2712 => x"d4",
          2713 => x"08",
          2714 => x"d4",
          2715 => x"0c",
          2716 => x"08",
          2717 => x"82",
          2718 => x"fc",
          2719 => x"0c",
          2720 => x"82",
          2721 => x"ec",
          2722 => x"b5",
          2723 => x"05",
          2724 => x"c8",
          2725 => x"0d",
          2726 => x"0c",
          2727 => x"0d",
          2728 => x"70",
          2729 => x"74",
          2730 => x"e3",
          2731 => x"75",
          2732 => x"d1",
          2733 => x"c8",
          2734 => x"0c",
          2735 => x"54",
          2736 => x"74",
          2737 => x"a0",
          2738 => x"06",
          2739 => x"15",
          2740 => x"80",
          2741 => x"29",
          2742 => x"05",
          2743 => x"56",
          2744 => x"82",
          2745 => x"53",
          2746 => x"08",
          2747 => x"3f",
          2748 => x"08",
          2749 => x"16",
          2750 => x"81",
          2751 => x"38",
          2752 => x"81",
          2753 => x"54",
          2754 => x"c9",
          2755 => x"73",
          2756 => x"0c",
          2757 => x"04",
          2758 => x"73",
          2759 => x"26",
          2760 => x"71",
          2761 => x"95",
          2762 => x"71",
          2763 => x"9a",
          2764 => x"80",
          2765 => x"80",
          2766 => x"39",
          2767 => x"51",
          2768 => x"82",
          2769 => x"80",
          2770 => x"9b",
          2771 => x"e4",
          2772 => x"c0",
          2773 => x"39",
          2774 => x"51",
          2775 => x"82",
          2776 => x"80",
          2777 => x"9b",
          2778 => x"c8",
          2779 => x"94",
          2780 => x"39",
          2781 => x"51",
          2782 => x"9c",
          2783 => x"39",
          2784 => x"51",
          2785 => x"9d",
          2786 => x"39",
          2787 => x"51",
          2788 => x"9d",
          2789 => x"39",
          2790 => x"51",
          2791 => x"9d",
          2792 => x"39",
          2793 => x"51",
          2794 => x"9e",
          2795 => x"39",
          2796 => x"51",
          2797 => x"83",
          2798 => x"fb",
          2799 => x"79",
          2800 => x"87",
          2801 => x"38",
          2802 => x"87",
          2803 => x"90",
          2804 => x"52",
          2805 => x"ab",
          2806 => x"c8",
          2807 => x"51",
          2808 => x"82",
          2809 => x"54",
          2810 => x"52",
          2811 => x"51",
          2812 => x"3f",
          2813 => x"04",
          2814 => x"66",
          2815 => x"80",
          2816 => x"5b",
          2817 => x"78",
          2818 => x"07",
          2819 => x"57",
          2820 => x"56",
          2821 => x"26",
          2822 => x"56",
          2823 => x"70",
          2824 => x"51",
          2825 => x"74",
          2826 => x"81",
          2827 => x"8c",
          2828 => x"56",
          2829 => x"3f",
          2830 => x"08",
          2831 => x"c8",
          2832 => x"82",
          2833 => x"87",
          2834 => x"0c",
          2835 => x"08",
          2836 => x"d4",
          2837 => x"80",
          2838 => x"75",
          2839 => x"81",
          2840 => x"c8",
          2841 => x"b5",
          2842 => x"38",
          2843 => x"80",
          2844 => x"74",
          2845 => x"59",
          2846 => x"96",
          2847 => x"51",
          2848 => x"3f",
          2849 => x"78",
          2850 => x"7b",
          2851 => x"2a",
          2852 => x"57",
          2853 => x"80",
          2854 => x"82",
          2855 => x"87",
          2856 => x"08",
          2857 => x"fe",
          2858 => x"56",
          2859 => x"c8",
          2860 => x"0d",
          2861 => x"0d",
          2862 => x"05",
          2863 => x"58",
          2864 => x"80",
          2865 => x"7a",
          2866 => x"3f",
          2867 => x"08",
          2868 => x"80",
          2869 => x"76",
          2870 => x"38",
          2871 => x"cd",
          2872 => x"55",
          2873 => x"b5",
          2874 => x"52",
          2875 => x"2d",
          2876 => x"08",
          2877 => x"78",
          2878 => x"b5",
          2879 => x"3d",
          2880 => x"3d",
          2881 => x"63",
          2882 => x"80",
          2883 => x"73",
          2884 => x"41",
          2885 => x"5e",
          2886 => x"52",
          2887 => x"51",
          2888 => x"3f",
          2889 => x"51",
          2890 => x"3f",
          2891 => x"79",
          2892 => x"38",
          2893 => x"89",
          2894 => x"2e",
          2895 => x"c6",
          2896 => x"53",
          2897 => x"8e",
          2898 => x"52",
          2899 => x"51",
          2900 => x"3f",
          2901 => x"9e",
          2902 => x"b8",
          2903 => x"15",
          2904 => x"39",
          2905 => x"72",
          2906 => x"38",
          2907 => x"82",
          2908 => x"ff",
          2909 => x"89",
          2910 => x"e8",
          2911 => x"d8",
          2912 => x"55",
          2913 => x"18",
          2914 => x"27",
          2915 => x"33",
          2916 => x"f4",
          2917 => x"c0",
          2918 => x"82",
          2919 => x"ff",
          2920 => x"81",
          2921 => x"cd",
          2922 => x"a0",
          2923 => x"3f",
          2924 => x"82",
          2925 => x"ff",
          2926 => x"80",
          2927 => x"27",
          2928 => x"74",
          2929 => x"55",
          2930 => x"72",
          2931 => x"38",
          2932 => x"53",
          2933 => x"83",
          2934 => x"75",
          2935 => x"81",
          2936 => x"53",
          2937 => x"90",
          2938 => x"fe",
          2939 => x"82",
          2940 => x"52",
          2941 => x"39",
          2942 => x"08",
          2943 => x"d7",
          2944 => x"15",
          2945 => x"39",
          2946 => x"51",
          2947 => x"78",
          2948 => x"5c",
          2949 => x"3f",
          2950 => x"08",
          2951 => x"98",
          2952 => x"76",
          2953 => x"81",
          2954 => x"9c",
          2955 => x"b5",
          2956 => x"2b",
          2957 => x"70",
          2958 => x"30",
          2959 => x"70",
          2960 => x"07",
          2961 => x"06",
          2962 => x"59",
          2963 => x"80",
          2964 => x"38",
          2965 => x"09",
          2966 => x"38",
          2967 => x"39",
          2968 => x"72",
          2969 => x"b2",
          2970 => x"72",
          2971 => x"0c",
          2972 => x"04",
          2973 => x"02",
          2974 => x"82",
          2975 => x"82",
          2976 => x"55",
          2977 => x"3f",
          2978 => x"22",
          2979 => x"3f",
          2980 => x"54",
          2981 => x"53",
          2982 => x"33",
          2983 => x"ac",
          2984 => x"b4",
          2985 => x"2e",
          2986 => x"d8",
          2987 => x"0d",
          2988 => x"0d",
          2989 => x"80",
          2990 => x"c2",
          2991 => x"98",
          2992 => x"9f",
          2993 => x"a3",
          2994 => x"98",
          2995 => x"81",
          2996 => x"06",
          2997 => x"80",
          2998 => x"81",
          2999 => x"3f",
          3000 => x"51",
          3001 => x"80",
          3002 => x"3f",
          3003 => x"70",
          3004 => x"52",
          3005 => x"92",
          3006 => x"97",
          3007 => x"9f",
          3008 => x"e7",
          3009 => x"97",
          3010 => x"83",
          3011 => x"06",
          3012 => x"80",
          3013 => x"81",
          3014 => x"3f",
          3015 => x"51",
          3016 => x"80",
          3017 => x"3f",
          3018 => x"70",
          3019 => x"52",
          3020 => x"92",
          3021 => x"97",
          3022 => x"a0",
          3023 => x"ab",
          3024 => x"97",
          3025 => x"85",
          3026 => x"06",
          3027 => x"80",
          3028 => x"81",
          3029 => x"3f",
          3030 => x"51",
          3031 => x"80",
          3032 => x"3f",
          3033 => x"70",
          3034 => x"52",
          3035 => x"92",
          3036 => x"96",
          3037 => x"a0",
          3038 => x"ef",
          3039 => x"96",
          3040 => x"87",
          3041 => x"06",
          3042 => x"80",
          3043 => x"81",
          3044 => x"3f",
          3045 => x"51",
          3046 => x"80",
          3047 => x"3f",
          3048 => x"70",
          3049 => x"52",
          3050 => x"92",
          3051 => x"96",
          3052 => x"a0",
          3053 => x"b3",
          3054 => x"96",
          3055 => x"c6",
          3056 => x"0d",
          3057 => x"0d",
          3058 => x"05",
          3059 => x"70",
          3060 => x"80",
          3061 => x"e3",
          3062 => x"0b",
          3063 => x"33",
          3064 => x"38",
          3065 => x"a1",
          3066 => x"cc",
          3067 => x"f8",
          3068 => x"b5",
          3069 => x"70",
          3070 => x"08",
          3071 => x"82",
          3072 => x"51",
          3073 => x"0b",
          3074 => x"34",
          3075 => x"b0",
          3076 => x"73",
          3077 => x"81",
          3078 => x"82",
          3079 => x"74",
          3080 => x"81",
          3081 => x"82",
          3082 => x"80",
          3083 => x"82",
          3084 => x"51",
          3085 => x"91",
          3086 => x"c8",
          3087 => x"ad",
          3088 => x"0b",
          3089 => x"c4",
          3090 => x"82",
          3091 => x"54",
          3092 => x"09",
          3093 => x"38",
          3094 => x"53",
          3095 => x"51",
          3096 => x"80",
          3097 => x"c8",
          3098 => x"0d",
          3099 => x"0d",
          3100 => x"82",
          3101 => x"5f",
          3102 => x"7c",
          3103 => x"d7",
          3104 => x"c8",
          3105 => x"06",
          3106 => x"2e",
          3107 => x"a3",
          3108 => x"59",
          3109 => x"a1",
          3110 => x"51",
          3111 => x"7c",
          3112 => x"82",
          3113 => x"80",
          3114 => x"82",
          3115 => x"7d",
          3116 => x"82",
          3117 => x"8d",
          3118 => x"70",
          3119 => x"a1",
          3120 => x"b2",
          3121 => x"3d",
          3122 => x"80",
          3123 => x"51",
          3124 => x"b4",
          3125 => x"05",
          3126 => x"3f",
          3127 => x"08",
          3128 => x"90",
          3129 => x"78",
          3130 => x"87",
          3131 => x"80",
          3132 => x"38",
          3133 => x"81",
          3134 => x"bd",
          3135 => x"78",
          3136 => x"ba",
          3137 => x"2e",
          3138 => x"8a",
          3139 => x"80",
          3140 => x"99",
          3141 => x"c0",
          3142 => x"38",
          3143 => x"82",
          3144 => x"bd",
          3145 => x"f9",
          3146 => x"38",
          3147 => x"24",
          3148 => x"80",
          3149 => x"88",
          3150 => x"f8",
          3151 => x"38",
          3152 => x"78",
          3153 => x"8a",
          3154 => x"81",
          3155 => x"38",
          3156 => x"2e",
          3157 => x"8a",
          3158 => x"81",
          3159 => x"fb",
          3160 => x"39",
          3161 => x"80",
          3162 => x"84",
          3163 => x"dc",
          3164 => x"c8",
          3165 => x"fe",
          3166 => x"3d",
          3167 => x"53",
          3168 => x"51",
          3169 => x"82",
          3170 => x"80",
          3171 => x"38",
          3172 => x"f8",
          3173 => x"84",
          3174 => x"b0",
          3175 => x"c8",
          3176 => x"82",
          3177 => x"42",
          3178 => x"51",
          3179 => x"3f",
          3180 => x"5a",
          3181 => x"81",
          3182 => x"59",
          3183 => x"84",
          3184 => x"7a",
          3185 => x"38",
          3186 => x"b4",
          3187 => x"11",
          3188 => x"05",
          3189 => x"3f",
          3190 => x"08",
          3191 => x"de",
          3192 => x"fe",
          3193 => x"ff",
          3194 => x"eb",
          3195 => x"b5",
          3196 => x"2e",
          3197 => x"b4",
          3198 => x"11",
          3199 => x"05",
          3200 => x"3f",
          3201 => x"08",
          3202 => x"b2",
          3203 => x"88",
          3204 => x"c4",
          3205 => x"79",
          3206 => x"89",
          3207 => x"79",
          3208 => x"5b",
          3209 => x"61",
          3210 => x"eb",
          3211 => x"ff",
          3212 => x"ff",
          3213 => x"eb",
          3214 => x"b5",
          3215 => x"2e",
          3216 => x"b4",
          3217 => x"11",
          3218 => x"05",
          3219 => x"3f",
          3220 => x"08",
          3221 => x"e6",
          3222 => x"fe",
          3223 => x"ff",
          3224 => x"ea",
          3225 => x"b5",
          3226 => x"2e",
          3227 => x"82",
          3228 => x"ff",
          3229 => x"63",
          3230 => x"27",
          3231 => x"70",
          3232 => x"5e",
          3233 => x"7c",
          3234 => x"78",
          3235 => x"79",
          3236 => x"52",
          3237 => x"51",
          3238 => x"3f",
          3239 => x"81",
          3240 => x"d5",
          3241 => x"cd",
          3242 => x"92",
          3243 => x"ff",
          3244 => x"ff",
          3245 => x"ea",
          3246 => x"b5",
          3247 => x"df",
          3248 => x"b4",
          3249 => x"80",
          3250 => x"82",
          3251 => x"44",
          3252 => x"82",
          3253 => x"59",
          3254 => x"88",
          3255 => x"f4",
          3256 => x"39",
          3257 => x"33",
          3258 => x"2e",
          3259 => x"b3",
          3260 => x"ab",
          3261 => x"b7",
          3262 => x"80",
          3263 => x"82",
          3264 => x"44",
          3265 => x"b4",
          3266 => x"78",
          3267 => x"38",
          3268 => x"08",
          3269 => x"82",
          3270 => x"fc",
          3271 => x"b4",
          3272 => x"11",
          3273 => x"05",
          3274 => x"3f",
          3275 => x"08",
          3276 => x"82",
          3277 => x"59",
          3278 => x"89",
          3279 => x"f0",
          3280 => x"cc",
          3281 => x"b5",
          3282 => x"80",
          3283 => x"82",
          3284 => x"43",
          3285 => x"b4",
          3286 => x"78",
          3287 => x"38",
          3288 => x"08",
          3289 => x"82",
          3290 => x"59",
          3291 => x"88",
          3292 => x"88",
          3293 => x"39",
          3294 => x"33",
          3295 => x"2e",
          3296 => x"b4",
          3297 => x"88",
          3298 => x"9c",
          3299 => x"43",
          3300 => x"f8",
          3301 => x"84",
          3302 => x"b0",
          3303 => x"c8",
          3304 => x"a7",
          3305 => x"5c",
          3306 => x"2e",
          3307 => x"5c",
          3308 => x"70",
          3309 => x"07",
          3310 => x"7f",
          3311 => x"5a",
          3312 => x"2e",
          3313 => x"a0",
          3314 => x"88",
          3315 => x"c0",
          3316 => x"3f",
          3317 => x"54",
          3318 => x"52",
          3319 => x"a2",
          3320 => x"cc",
          3321 => x"39",
          3322 => x"80",
          3323 => x"84",
          3324 => x"d8",
          3325 => x"c8",
          3326 => x"f9",
          3327 => x"3d",
          3328 => x"53",
          3329 => x"51",
          3330 => x"82",
          3331 => x"80",
          3332 => x"63",
          3333 => x"cb",
          3334 => x"34",
          3335 => x"44",
          3336 => x"fc",
          3337 => x"84",
          3338 => x"a0",
          3339 => x"c8",
          3340 => x"f9",
          3341 => x"70",
          3342 => x"82",
          3343 => x"ff",
          3344 => x"82",
          3345 => x"53",
          3346 => x"79",
          3347 => x"dd",
          3348 => x"79",
          3349 => x"ae",
          3350 => x"38",
          3351 => x"9f",
          3352 => x"fe",
          3353 => x"ff",
          3354 => x"e6",
          3355 => x"b5",
          3356 => x"2e",
          3357 => x"59",
          3358 => x"05",
          3359 => x"63",
          3360 => x"ff",
          3361 => x"a2",
          3362 => x"d7",
          3363 => x"39",
          3364 => x"f4",
          3365 => x"84",
          3366 => x"df",
          3367 => x"c8",
          3368 => x"f8",
          3369 => x"3d",
          3370 => x"53",
          3371 => x"51",
          3372 => x"82",
          3373 => x"80",
          3374 => x"60",
          3375 => x"05",
          3376 => x"82",
          3377 => x"78",
          3378 => x"fe",
          3379 => x"ff",
          3380 => x"e0",
          3381 => x"b5",
          3382 => x"38",
          3383 => x"60",
          3384 => x"52",
          3385 => x"51",
          3386 => x"3f",
          3387 => x"08",
          3388 => x"52",
          3389 => x"aa",
          3390 => x"45",
          3391 => x"78",
          3392 => x"ba",
          3393 => x"26",
          3394 => x"82",
          3395 => x"39",
          3396 => x"f0",
          3397 => x"84",
          3398 => x"df",
          3399 => x"c8",
          3400 => x"92",
          3401 => x"02",
          3402 => x"79",
          3403 => x"5b",
          3404 => x"ff",
          3405 => x"a2",
          3406 => x"a7",
          3407 => x"39",
          3408 => x"f4",
          3409 => x"84",
          3410 => x"af",
          3411 => x"c8",
          3412 => x"f6",
          3413 => x"3d",
          3414 => x"53",
          3415 => x"51",
          3416 => x"82",
          3417 => x"80",
          3418 => x"60",
          3419 => x"59",
          3420 => x"41",
          3421 => x"f0",
          3422 => x"84",
          3423 => x"fb",
          3424 => x"c8",
          3425 => x"f6",
          3426 => x"70",
          3427 => x"82",
          3428 => x"ff",
          3429 => x"82",
          3430 => x"53",
          3431 => x"79",
          3432 => x"89",
          3433 => x"79",
          3434 => x"ae",
          3435 => x"38",
          3436 => x"9b",
          3437 => x"fe",
          3438 => x"ff",
          3439 => x"de",
          3440 => x"b5",
          3441 => x"2e",
          3442 => x"60",
          3443 => x"60",
          3444 => x"ff",
          3445 => x"a2",
          3446 => x"87",
          3447 => x"39",
          3448 => x"80",
          3449 => x"84",
          3450 => x"e0",
          3451 => x"c8",
          3452 => x"f5",
          3453 => x"52",
          3454 => x"51",
          3455 => x"3f",
          3456 => x"04",
          3457 => x"80",
          3458 => x"84",
          3459 => x"bc",
          3460 => x"c8",
          3461 => x"f5",
          3462 => x"52",
          3463 => x"51",
          3464 => x"3f",
          3465 => x"2d",
          3466 => x"08",
          3467 => x"8e",
          3468 => x"c8",
          3469 => x"a3",
          3470 => x"a7",
          3471 => x"fe",
          3472 => x"d8",
          3473 => x"3f",
          3474 => x"3f",
          3475 => x"82",
          3476 => x"c3",
          3477 => x"59",
          3478 => x"91",
          3479 => x"de",
          3480 => x"79",
          3481 => x"80",
          3482 => x"38",
          3483 => x"59",
          3484 => x"81",
          3485 => x"3d",
          3486 => x"51",
          3487 => x"82",
          3488 => x"5c",
          3489 => x"82",
          3490 => x"7a",
          3491 => x"38",
          3492 => x"8c",
          3493 => x"39",
          3494 => x"ad",
          3495 => x"39",
          3496 => x"56",
          3497 => x"a4",
          3498 => x"53",
          3499 => x"52",
          3500 => x"b0",
          3501 => x"a9",
          3502 => x"39",
          3503 => x"3d",
          3504 => x"51",
          3505 => x"ab",
          3506 => x"82",
          3507 => x"80",
          3508 => x"a0",
          3509 => x"ff",
          3510 => x"ff",
          3511 => x"93",
          3512 => x"80",
          3513 => x"ac",
          3514 => x"ff",
          3515 => x"ff",
          3516 => x"82",
          3517 => x"82",
          3518 => x"80",
          3519 => x"80",
          3520 => x"80",
          3521 => x"80",
          3522 => x"ff",
          3523 => x"eb",
          3524 => x"b5",
          3525 => x"b5",
          3526 => x"70",
          3527 => x"07",
          3528 => x"5b",
          3529 => x"5a",
          3530 => x"83",
          3531 => x"78",
          3532 => x"78",
          3533 => x"38",
          3534 => x"81",
          3535 => x"59",
          3536 => x"38",
          3537 => x"7d",
          3538 => x"59",
          3539 => x"7e",
          3540 => x"81",
          3541 => x"38",
          3542 => x"51",
          3543 => x"f2",
          3544 => x"3d",
          3545 => x"82",
          3546 => x"87",
          3547 => x"70",
          3548 => x"87",
          3549 => x"72",
          3550 => x"3f",
          3551 => x"08",
          3552 => x"08",
          3553 => x"84",
          3554 => x"51",
          3555 => x"72",
          3556 => x"08",
          3557 => x"87",
          3558 => x"70",
          3559 => x"87",
          3560 => x"72",
          3561 => x"3f",
          3562 => x"08",
          3563 => x"08",
          3564 => x"84",
          3565 => x"51",
          3566 => x"72",
          3567 => x"08",
          3568 => x"8c",
          3569 => x"87",
          3570 => x"0c",
          3571 => x"0b",
          3572 => x"94",
          3573 => x"e7",
          3574 => x"d3",
          3575 => x"84",
          3576 => x"34",
          3577 => x"cd",
          3578 => x"3d",
          3579 => x"0c",
          3580 => x"82",
          3581 => x"54",
          3582 => x"93",
          3583 => x"a4",
          3584 => x"bf",
          3585 => x"a4",
          3586 => x"bf",
          3587 => x"dd",
          3588 => x"e5",
          3589 => x"ec",
          3590 => x"d1",
          3591 => x"fe",
          3592 => x"52",
          3593 => x"88",
          3594 => x"d8",
          3595 => x"c8",
          3596 => x"06",
          3597 => x"14",
          3598 => x"80",
          3599 => x"71",
          3600 => x"0c",
          3601 => x"04",
          3602 => x"76",
          3603 => x"55",
          3604 => x"54",
          3605 => x"81",
          3606 => x"33",
          3607 => x"2e",
          3608 => x"86",
          3609 => x"53",
          3610 => x"33",
          3611 => x"2e",
          3612 => x"86",
          3613 => x"53",
          3614 => x"52",
          3615 => x"09",
          3616 => x"38",
          3617 => x"12",
          3618 => x"33",
          3619 => x"a2",
          3620 => x"81",
          3621 => x"2e",
          3622 => x"ea",
          3623 => x"81",
          3624 => x"72",
          3625 => x"70",
          3626 => x"38",
          3627 => x"80",
          3628 => x"73",
          3629 => x"72",
          3630 => x"70",
          3631 => x"81",
          3632 => x"81",
          3633 => x"32",
          3634 => x"80",
          3635 => x"51",
          3636 => x"80",
          3637 => x"80",
          3638 => x"05",
          3639 => x"75",
          3640 => x"70",
          3641 => x"0c",
          3642 => x"04",
          3643 => x"76",
          3644 => x"80",
          3645 => x"86",
          3646 => x"52",
          3647 => x"fb",
          3648 => x"c8",
          3649 => x"80",
          3650 => x"74",
          3651 => x"b5",
          3652 => x"3d",
          3653 => x"3d",
          3654 => x"11",
          3655 => x"52",
          3656 => x"70",
          3657 => x"98",
          3658 => x"33",
          3659 => x"82",
          3660 => x"26",
          3661 => x"84",
          3662 => x"83",
          3663 => x"26",
          3664 => x"85",
          3665 => x"84",
          3666 => x"26",
          3667 => x"86",
          3668 => x"85",
          3669 => x"26",
          3670 => x"88",
          3671 => x"86",
          3672 => x"e7",
          3673 => x"38",
          3674 => x"54",
          3675 => x"87",
          3676 => x"cc",
          3677 => x"87",
          3678 => x"0c",
          3679 => x"c0",
          3680 => x"82",
          3681 => x"c0",
          3682 => x"83",
          3683 => x"c0",
          3684 => x"84",
          3685 => x"c0",
          3686 => x"85",
          3687 => x"c0",
          3688 => x"86",
          3689 => x"c0",
          3690 => x"74",
          3691 => x"a4",
          3692 => x"c0",
          3693 => x"80",
          3694 => x"98",
          3695 => x"52",
          3696 => x"c8",
          3697 => x"0d",
          3698 => x"0d",
          3699 => x"c0",
          3700 => x"81",
          3701 => x"c0",
          3702 => x"5e",
          3703 => x"87",
          3704 => x"08",
          3705 => x"1c",
          3706 => x"98",
          3707 => x"79",
          3708 => x"87",
          3709 => x"08",
          3710 => x"1c",
          3711 => x"98",
          3712 => x"79",
          3713 => x"87",
          3714 => x"08",
          3715 => x"1c",
          3716 => x"98",
          3717 => x"7b",
          3718 => x"87",
          3719 => x"08",
          3720 => x"1c",
          3721 => x"0c",
          3722 => x"ff",
          3723 => x"83",
          3724 => x"58",
          3725 => x"57",
          3726 => x"56",
          3727 => x"55",
          3728 => x"54",
          3729 => x"53",
          3730 => x"ff",
          3731 => x"a4",
          3732 => x"9f",
          3733 => x"3d",
          3734 => x"3d",
          3735 => x"05",
          3736 => x"e8",
          3737 => x"ff",
          3738 => x"55",
          3739 => x"84",
          3740 => x"2e",
          3741 => x"c0",
          3742 => x"70",
          3743 => x"2a",
          3744 => x"53",
          3745 => x"80",
          3746 => x"71",
          3747 => x"81",
          3748 => x"70",
          3749 => x"81",
          3750 => x"06",
          3751 => x"80",
          3752 => x"71",
          3753 => x"81",
          3754 => x"70",
          3755 => x"73",
          3756 => x"51",
          3757 => x"80",
          3758 => x"2e",
          3759 => x"c0",
          3760 => x"74",
          3761 => x"82",
          3762 => x"87",
          3763 => x"ff",
          3764 => x"8f",
          3765 => x"30",
          3766 => x"51",
          3767 => x"82",
          3768 => x"83",
          3769 => x"f9",
          3770 => x"a7",
          3771 => x"77",
          3772 => x"81",
          3773 => x"7a",
          3774 => x"eb",
          3775 => x"e8",
          3776 => x"ff",
          3777 => x"87",
          3778 => x"53",
          3779 => x"86",
          3780 => x"94",
          3781 => x"08",
          3782 => x"70",
          3783 => x"56",
          3784 => x"2e",
          3785 => x"91",
          3786 => x"06",
          3787 => x"d7",
          3788 => x"32",
          3789 => x"51",
          3790 => x"2e",
          3791 => x"93",
          3792 => x"06",
          3793 => x"ff",
          3794 => x"81",
          3795 => x"87",
          3796 => x"54",
          3797 => x"86",
          3798 => x"94",
          3799 => x"74",
          3800 => x"82",
          3801 => x"89",
          3802 => x"f9",
          3803 => x"54",
          3804 => x"70",
          3805 => x"53",
          3806 => x"77",
          3807 => x"38",
          3808 => x"06",
          3809 => x"b3",
          3810 => x"81",
          3811 => x"57",
          3812 => x"c0",
          3813 => x"75",
          3814 => x"38",
          3815 => x"94",
          3816 => x"70",
          3817 => x"81",
          3818 => x"52",
          3819 => x"8c",
          3820 => x"2a",
          3821 => x"51",
          3822 => x"38",
          3823 => x"70",
          3824 => x"51",
          3825 => x"8d",
          3826 => x"2a",
          3827 => x"51",
          3828 => x"be",
          3829 => x"ff",
          3830 => x"c0",
          3831 => x"70",
          3832 => x"38",
          3833 => x"90",
          3834 => x"0c",
          3835 => x"33",
          3836 => x"06",
          3837 => x"70",
          3838 => x"76",
          3839 => x"0c",
          3840 => x"04",
          3841 => x"82",
          3842 => x"70",
          3843 => x"54",
          3844 => x"94",
          3845 => x"80",
          3846 => x"87",
          3847 => x"51",
          3848 => x"82",
          3849 => x"06",
          3850 => x"70",
          3851 => x"38",
          3852 => x"06",
          3853 => x"94",
          3854 => x"80",
          3855 => x"87",
          3856 => x"52",
          3857 => x"81",
          3858 => x"b5",
          3859 => x"84",
          3860 => x"ff",
          3861 => x"b5",
          3862 => x"ff",
          3863 => x"c8",
          3864 => x"3d",
          3865 => x"e8",
          3866 => x"ff",
          3867 => x"87",
          3868 => x"52",
          3869 => x"86",
          3870 => x"94",
          3871 => x"08",
          3872 => x"70",
          3873 => x"51",
          3874 => x"70",
          3875 => x"38",
          3876 => x"06",
          3877 => x"94",
          3878 => x"80",
          3879 => x"87",
          3880 => x"52",
          3881 => x"98",
          3882 => x"2c",
          3883 => x"71",
          3884 => x"0c",
          3885 => x"04",
          3886 => x"87",
          3887 => x"08",
          3888 => x"8a",
          3889 => x"70",
          3890 => x"b4",
          3891 => x"9e",
          3892 => x"b3",
          3893 => x"c0",
          3894 => x"82",
          3895 => x"87",
          3896 => x"08",
          3897 => x"0c",
          3898 => x"98",
          3899 => x"f8",
          3900 => x"9e",
          3901 => x"b3",
          3902 => x"c0",
          3903 => x"82",
          3904 => x"87",
          3905 => x"08",
          3906 => x"0c",
          3907 => x"b0",
          3908 => x"88",
          3909 => x"9e",
          3910 => x"b4",
          3911 => x"c0",
          3912 => x"82",
          3913 => x"87",
          3914 => x"08",
          3915 => x"0c",
          3916 => x"c0",
          3917 => x"98",
          3918 => x"9e",
          3919 => x"b4",
          3920 => x"c0",
          3921 => x"51",
          3922 => x"a0",
          3923 => x"9e",
          3924 => x"b4",
          3925 => x"c0",
          3926 => x"82",
          3927 => x"87",
          3928 => x"08",
          3929 => x"0c",
          3930 => x"b4",
          3931 => x"0b",
          3932 => x"90",
          3933 => x"80",
          3934 => x"52",
          3935 => x"2e",
          3936 => x"52",
          3937 => x"b1",
          3938 => x"87",
          3939 => x"08",
          3940 => x"0a",
          3941 => x"52",
          3942 => x"83",
          3943 => x"71",
          3944 => x"34",
          3945 => x"c0",
          3946 => x"70",
          3947 => x"06",
          3948 => x"70",
          3949 => x"38",
          3950 => x"82",
          3951 => x"80",
          3952 => x"9e",
          3953 => x"88",
          3954 => x"51",
          3955 => x"80",
          3956 => x"81",
          3957 => x"b4",
          3958 => x"0b",
          3959 => x"90",
          3960 => x"80",
          3961 => x"52",
          3962 => x"2e",
          3963 => x"52",
          3964 => x"b5",
          3965 => x"87",
          3966 => x"08",
          3967 => x"80",
          3968 => x"52",
          3969 => x"83",
          3970 => x"71",
          3971 => x"34",
          3972 => x"c0",
          3973 => x"70",
          3974 => x"06",
          3975 => x"70",
          3976 => x"38",
          3977 => x"82",
          3978 => x"80",
          3979 => x"9e",
          3980 => x"82",
          3981 => x"51",
          3982 => x"80",
          3983 => x"81",
          3984 => x"b4",
          3985 => x"0b",
          3986 => x"90",
          3987 => x"80",
          3988 => x"52",
          3989 => x"2e",
          3990 => x"52",
          3991 => x"b9",
          3992 => x"87",
          3993 => x"08",
          3994 => x"80",
          3995 => x"52",
          3996 => x"83",
          3997 => x"71",
          3998 => x"34",
          3999 => x"c0",
          4000 => x"70",
          4001 => x"51",
          4002 => x"80",
          4003 => x"81",
          4004 => x"b4",
          4005 => x"c0",
          4006 => x"70",
          4007 => x"70",
          4008 => x"51",
          4009 => x"b4",
          4010 => x"0b",
          4011 => x"90",
          4012 => x"80",
          4013 => x"52",
          4014 => x"83",
          4015 => x"71",
          4016 => x"34",
          4017 => x"90",
          4018 => x"f0",
          4019 => x"2a",
          4020 => x"70",
          4021 => x"34",
          4022 => x"c0",
          4023 => x"70",
          4024 => x"52",
          4025 => x"2e",
          4026 => x"52",
          4027 => x"bf",
          4028 => x"9e",
          4029 => x"87",
          4030 => x"70",
          4031 => x"34",
          4032 => x"04",
          4033 => x"82",
          4034 => x"ff",
          4035 => x"82",
          4036 => x"54",
          4037 => x"89",
          4038 => x"94",
          4039 => x"c3",
          4040 => x"a8",
          4041 => x"bb",
          4042 => x"b2",
          4043 => x"80",
          4044 => x"82",
          4045 => x"82",
          4046 => x"11",
          4047 => x"a5",
          4048 => x"95",
          4049 => x"b4",
          4050 => x"73",
          4051 => x"38",
          4052 => x"08",
          4053 => x"08",
          4054 => x"82",
          4055 => x"ff",
          4056 => x"82",
          4057 => x"54",
          4058 => x"94",
          4059 => x"ec",
          4060 => x"f0",
          4061 => x"52",
          4062 => x"51",
          4063 => x"3f",
          4064 => x"33",
          4065 => x"2e",
          4066 => x"b3",
          4067 => x"b3",
          4068 => x"54",
          4069 => x"94",
          4070 => x"bc",
          4071 => x"b6",
          4072 => x"80",
          4073 => x"82",
          4074 => x"82",
          4075 => x"11",
          4076 => x"a6",
          4077 => x"94",
          4078 => x"b4",
          4079 => x"73",
          4080 => x"38",
          4081 => x"33",
          4082 => x"cc",
          4083 => x"88",
          4084 => x"bf",
          4085 => x"80",
          4086 => x"82",
          4087 => x"52",
          4088 => x"51",
          4089 => x"3f",
          4090 => x"33",
          4091 => x"2e",
          4092 => x"b4",
          4093 => x"82",
          4094 => x"ff",
          4095 => x"82",
          4096 => x"54",
          4097 => x"89",
          4098 => x"ac",
          4099 => x"d3",
          4100 => x"b3",
          4101 => x"80",
          4102 => x"82",
          4103 => x"ff",
          4104 => x"82",
          4105 => x"54",
          4106 => x"89",
          4107 => x"cc",
          4108 => x"af",
          4109 => x"b9",
          4110 => x"80",
          4111 => x"82",
          4112 => x"ff",
          4113 => x"82",
          4114 => x"54",
          4115 => x"89",
          4116 => x"e4",
          4117 => x"8b",
          4118 => x"f0",
          4119 => x"83",
          4120 => x"94",
          4121 => x"a7",
          4122 => x"92",
          4123 => x"b4",
          4124 => x"82",
          4125 => x"ff",
          4126 => x"82",
          4127 => x"52",
          4128 => x"51",
          4129 => x"3f",
          4130 => x"51",
          4131 => x"3f",
          4132 => x"22",
          4133 => x"fc",
          4134 => x"bc",
          4135 => x"a4",
          4136 => x"84",
          4137 => x"51",
          4138 => x"82",
          4139 => x"bd",
          4140 => x"76",
          4141 => x"54",
          4142 => x"08",
          4143 => x"a4",
          4144 => x"94",
          4145 => x"b7",
          4146 => x"80",
          4147 => x"82",
          4148 => x"56",
          4149 => x"52",
          4150 => x"a7",
          4151 => x"c8",
          4152 => x"c0",
          4153 => x"31",
          4154 => x"b5",
          4155 => x"82",
          4156 => x"ff",
          4157 => x"82",
          4158 => x"54",
          4159 => x"a9",
          4160 => x"ac",
          4161 => x"84",
          4162 => x"51",
          4163 => x"82",
          4164 => x"bd",
          4165 => x"76",
          4166 => x"54",
          4167 => x"08",
          4168 => x"fc",
          4169 => x"b0",
          4170 => x"bc",
          4171 => x"b3",
          4172 => x"0d",
          4173 => x"0d",
          4174 => x"33",
          4175 => x"71",
          4176 => x"38",
          4177 => x"82",
          4178 => x"52",
          4179 => x"82",
          4180 => x"9d",
          4181 => x"b0",
          4182 => x"82",
          4183 => x"91",
          4184 => x"c0",
          4185 => x"82",
          4186 => x"85",
          4187 => x"cc",
          4188 => x"ef",
          4189 => x"0d",
          4190 => x"80",
          4191 => x"0b",
          4192 => x"84",
          4193 => x"b4",
          4194 => x"c0",
          4195 => x"04",
          4196 => x"76",
          4197 => x"98",
          4198 => x"2b",
          4199 => x"72",
          4200 => x"82",
          4201 => x"51",
          4202 => x"80",
          4203 => x"d8",
          4204 => x"53",
          4205 => x"9c",
          4206 => x"d4",
          4207 => x"02",
          4208 => x"05",
          4209 => x"52",
          4210 => x"72",
          4211 => x"06",
          4212 => x"53",
          4213 => x"c8",
          4214 => x"0d",
          4215 => x"0d",
          4216 => x"05",
          4217 => x"71",
          4218 => x"54",
          4219 => x"b1",
          4220 => x"9c",
          4221 => x"51",
          4222 => x"3f",
          4223 => x"08",
          4224 => x"ff",
          4225 => x"82",
          4226 => x"52",
          4227 => x"af",
          4228 => x"33",
          4229 => x"72",
          4230 => x"81",
          4231 => x"cc",
          4232 => x"ff",
          4233 => x"74",
          4234 => x"3d",
          4235 => x"3d",
          4236 => x"84",
          4237 => x"33",
          4238 => x"bb",
          4239 => x"b5",
          4240 => x"84",
          4241 => x"c8",
          4242 => x"51",
          4243 => x"58",
          4244 => x"2e",
          4245 => x"51",
          4246 => x"82",
          4247 => x"70",
          4248 => x"b4",
          4249 => x"19",
          4250 => x"56",
          4251 => x"3f",
          4252 => x"08",
          4253 => x"b5",
          4254 => x"84",
          4255 => x"c8",
          4256 => x"51",
          4257 => x"80",
          4258 => x"75",
          4259 => x"74",
          4260 => x"d1",
          4261 => x"a0",
          4262 => x"55",
          4263 => x"a0",
          4264 => x"ff",
          4265 => x"75",
          4266 => x"80",
          4267 => x"a0",
          4268 => x"2e",
          4269 => x"b5",
          4270 => x"75",
          4271 => x"38",
          4272 => x"33",
          4273 => x"38",
          4274 => x"05",
          4275 => x"78",
          4276 => x"80",
          4277 => x"82",
          4278 => x"52",
          4279 => x"8f",
          4280 => x"b5",
          4281 => x"80",
          4282 => x"8c",
          4283 => x"fd",
          4284 => x"b4",
          4285 => x"54",
          4286 => x"71",
          4287 => x"38",
          4288 => x"d0",
          4289 => x"0c",
          4290 => x"14",
          4291 => x"80",
          4292 => x"80",
          4293 => x"a0",
          4294 => x"9c",
          4295 => x"80",
          4296 => x"71",
          4297 => x"c5",
          4298 => x"9c",
          4299 => x"a4",
          4300 => x"82",
          4301 => x"85",
          4302 => x"dc",
          4303 => x"57",
          4304 => x"b5",
          4305 => x"80",
          4306 => x"82",
          4307 => x"80",
          4308 => x"b5",
          4309 => x"80",
          4310 => x"3d",
          4311 => x"81",
          4312 => x"82",
          4313 => x"80",
          4314 => x"75",
          4315 => x"95",
          4316 => x"c8",
          4317 => x"0b",
          4318 => x"08",
          4319 => x"82",
          4320 => x"ff",
          4321 => x"55",
          4322 => x"34",
          4323 => x"52",
          4324 => x"ad",
          4325 => x"ff",
          4326 => x"74",
          4327 => x"81",
          4328 => x"38",
          4329 => x"04",
          4330 => x"aa",
          4331 => x"3d",
          4332 => x"81",
          4333 => x"80",
          4334 => x"9c",
          4335 => x"e2",
          4336 => x"b5",
          4337 => x"95",
          4338 => x"82",
          4339 => x"54",
          4340 => x"52",
          4341 => x"52",
          4342 => x"86",
          4343 => x"c8",
          4344 => x"a5",
          4345 => x"ff",
          4346 => x"82",
          4347 => x"81",
          4348 => x"80",
          4349 => x"c8",
          4350 => x"38",
          4351 => x"08",
          4352 => x"17",
          4353 => x"74",
          4354 => x"70",
          4355 => x"07",
          4356 => x"55",
          4357 => x"2e",
          4358 => x"ff",
          4359 => x"b5",
          4360 => x"11",
          4361 => x"80",
          4362 => x"82",
          4363 => x"80",
          4364 => x"82",
          4365 => x"ff",
          4366 => x"78",
          4367 => x"81",
          4368 => x"75",
          4369 => x"ff",
          4370 => x"79",
          4371 => x"b5",
          4372 => x"08",
          4373 => x"c8",
          4374 => x"80",
          4375 => x"b5",
          4376 => x"3d",
          4377 => x"3d",
          4378 => x"71",
          4379 => x"33",
          4380 => x"58",
          4381 => x"09",
          4382 => x"38",
          4383 => x"05",
          4384 => x"27",
          4385 => x"17",
          4386 => x"71",
          4387 => x"55",
          4388 => x"09",
          4389 => x"38",
          4390 => x"ea",
          4391 => x"73",
          4392 => x"b5",
          4393 => x"08",
          4394 => x"b2",
          4395 => x"b5",
          4396 => x"79",
          4397 => x"51",
          4398 => x"3f",
          4399 => x"08",
          4400 => x"84",
          4401 => x"74",
          4402 => x"38",
          4403 => x"88",
          4404 => x"fc",
          4405 => x"39",
          4406 => x"8c",
          4407 => x"53",
          4408 => x"c5",
          4409 => x"b5",
          4410 => x"2e",
          4411 => x"1b",
          4412 => x"77",
          4413 => x"3f",
          4414 => x"08",
          4415 => x"55",
          4416 => x"74",
          4417 => x"81",
          4418 => x"ff",
          4419 => x"82",
          4420 => x"8b",
          4421 => x"73",
          4422 => x"0c",
          4423 => x"04",
          4424 => x"b0",
          4425 => x"3d",
          4426 => x"08",
          4427 => x"80",
          4428 => x"34",
          4429 => x"33",
          4430 => x"08",
          4431 => x"81",
          4432 => x"82",
          4433 => x"55",
          4434 => x"38",
          4435 => x"80",
          4436 => x"38",
          4437 => x"06",
          4438 => x"80",
          4439 => x"38",
          4440 => x"86",
          4441 => x"c8",
          4442 => x"9c",
          4443 => x"c8",
          4444 => x"81",
          4445 => x"53",
          4446 => x"b5",
          4447 => x"80",
          4448 => x"82",
          4449 => x"80",
          4450 => x"82",
          4451 => x"ff",
          4452 => x"80",
          4453 => x"b5",
          4454 => x"82",
          4455 => x"53",
          4456 => x"90",
          4457 => x"54",
          4458 => x"3f",
          4459 => x"08",
          4460 => x"c8",
          4461 => x"09",
          4462 => x"d0",
          4463 => x"c8",
          4464 => x"b0",
          4465 => x"b5",
          4466 => x"80",
          4467 => x"c8",
          4468 => x"38",
          4469 => x"08",
          4470 => x"17",
          4471 => x"74",
          4472 => x"74",
          4473 => x"52",
          4474 => x"c2",
          4475 => x"70",
          4476 => x"5c",
          4477 => x"27",
          4478 => x"5b",
          4479 => x"09",
          4480 => x"97",
          4481 => x"75",
          4482 => x"34",
          4483 => x"82",
          4484 => x"80",
          4485 => x"f9",
          4486 => x"3d",
          4487 => x"3f",
          4488 => x"08",
          4489 => x"98",
          4490 => x"78",
          4491 => x"38",
          4492 => x"06",
          4493 => x"33",
          4494 => x"70",
          4495 => x"cc",
          4496 => x"98",
          4497 => x"2c",
          4498 => x"05",
          4499 => x"82",
          4500 => x"70",
          4501 => x"33",
          4502 => x"51",
          4503 => x"59",
          4504 => x"56",
          4505 => x"80",
          4506 => x"74",
          4507 => x"74",
          4508 => x"29",
          4509 => x"05",
          4510 => x"51",
          4511 => x"24",
          4512 => x"76",
          4513 => x"77",
          4514 => x"3f",
          4515 => x"08",
          4516 => x"54",
          4517 => x"d7",
          4518 => x"cc",
          4519 => x"56",
          4520 => x"81",
          4521 => x"81",
          4522 => x"70",
          4523 => x"81",
          4524 => x"51",
          4525 => x"26",
          4526 => x"53",
          4527 => x"51",
          4528 => x"82",
          4529 => x"81",
          4530 => x"73",
          4531 => x"39",
          4532 => x"80",
          4533 => x"38",
          4534 => x"74",
          4535 => x"34",
          4536 => x"70",
          4537 => x"cc",
          4538 => x"98",
          4539 => x"2c",
          4540 => x"70",
          4541 => x"aa",
          4542 => x"5e",
          4543 => x"57",
          4544 => x"74",
          4545 => x"81",
          4546 => x"38",
          4547 => x"14",
          4548 => x"80",
          4549 => x"f4",
          4550 => x"82",
          4551 => x"92",
          4552 => x"cc",
          4553 => x"82",
          4554 => x"78",
          4555 => x"75",
          4556 => x"54",
          4557 => x"fd",
          4558 => x"84",
          4559 => x"8c",
          4560 => x"08",
          4561 => x"fc",
          4562 => x"7e",
          4563 => x"38",
          4564 => x"33",
          4565 => x"27",
          4566 => x"98",
          4567 => x"2c",
          4568 => x"75",
          4569 => x"74",
          4570 => x"33",
          4571 => x"74",
          4572 => x"29",
          4573 => x"05",
          4574 => x"82",
          4575 => x"56",
          4576 => x"39",
          4577 => x"33",
          4578 => x"54",
          4579 => x"fc",
          4580 => x"54",
          4581 => x"74",
          4582 => x"f8",
          4583 => x"7e",
          4584 => x"81",
          4585 => x"82",
          4586 => x"82",
          4587 => x"70",
          4588 => x"29",
          4589 => x"05",
          4590 => x"82",
          4591 => x"5a",
          4592 => x"74",
          4593 => x"38",
          4594 => x"08",
          4595 => x"70",
          4596 => x"ff",
          4597 => x"74",
          4598 => x"29",
          4599 => x"05",
          4600 => x"82",
          4601 => x"56",
          4602 => x"75",
          4603 => x"82",
          4604 => x"70",
          4605 => x"98",
          4606 => x"f8",
          4607 => x"56",
          4608 => x"25",
          4609 => x"82",
          4610 => x"52",
          4611 => x"a3",
          4612 => x"81",
          4613 => x"81",
          4614 => x"70",
          4615 => x"cc",
          4616 => x"51",
          4617 => x"24",
          4618 => x"ee",
          4619 => x"34",
          4620 => x"1b",
          4621 => x"fc",
          4622 => x"82",
          4623 => x"f3",
          4624 => x"fd",
          4625 => x"fc",
          4626 => x"ff",
          4627 => x"73",
          4628 => x"c6",
          4629 => x"f8",
          4630 => x"54",
          4631 => x"f8",
          4632 => x"54",
          4633 => x"fc",
          4634 => x"9c",
          4635 => x"51",
          4636 => x"3f",
          4637 => x"33",
          4638 => x"70",
          4639 => x"cc",
          4640 => x"51",
          4641 => x"74",
          4642 => x"74",
          4643 => x"14",
          4644 => x"82",
          4645 => x"52",
          4646 => x"ff",
          4647 => x"74",
          4648 => x"29",
          4649 => x"05",
          4650 => x"82",
          4651 => x"58",
          4652 => x"75",
          4653 => x"82",
          4654 => x"52",
          4655 => x"a1",
          4656 => x"cc",
          4657 => x"98",
          4658 => x"2c",
          4659 => x"33",
          4660 => x"57",
          4661 => x"fa",
          4662 => x"cd",
          4663 => x"88",
          4664 => x"ce",
          4665 => x"80",
          4666 => x"80",
          4667 => x"98",
          4668 => x"f8",
          4669 => x"55",
          4670 => x"de",
          4671 => x"39",
          4672 => x"33",
          4673 => x"80",
          4674 => x"cd",
          4675 => x"8a",
          4676 => x"9e",
          4677 => x"f8",
          4678 => x"f6",
          4679 => x"b5",
          4680 => x"ff",
          4681 => x"96",
          4682 => x"f8",
          4683 => x"80",
          4684 => x"81",
          4685 => x"79",
          4686 => x"3f",
          4687 => x"7a",
          4688 => x"82",
          4689 => x"80",
          4690 => x"f8",
          4691 => x"b5",
          4692 => x"3d",
          4693 => x"cc",
          4694 => x"73",
          4695 => x"ba",
          4696 => x"9c",
          4697 => x"51",
          4698 => x"3f",
          4699 => x"33",
          4700 => x"73",
          4701 => x"34",
          4702 => x"06",
          4703 => x"82",
          4704 => x"82",
          4705 => x"55",
          4706 => x"2e",
          4707 => x"ff",
          4708 => x"82",
          4709 => x"74",
          4710 => x"98",
          4711 => x"ff",
          4712 => x"55",
          4713 => x"ad",
          4714 => x"54",
          4715 => x"74",
          4716 => x"9c",
          4717 => x"33",
          4718 => x"f6",
          4719 => x"80",
          4720 => x"80",
          4721 => x"98",
          4722 => x"f8",
          4723 => x"55",
          4724 => x"d5",
          4725 => x"9c",
          4726 => x"51",
          4727 => x"3f",
          4728 => x"33",
          4729 => x"70",
          4730 => x"cc",
          4731 => x"51",
          4732 => x"74",
          4733 => x"38",
          4734 => x"08",
          4735 => x"ff",
          4736 => x"74",
          4737 => x"29",
          4738 => x"05",
          4739 => x"82",
          4740 => x"58",
          4741 => x"75",
          4742 => x"f7",
          4743 => x"cc",
          4744 => x"81",
          4745 => x"cc",
          4746 => x"56",
          4747 => x"27",
          4748 => x"82",
          4749 => x"52",
          4750 => x"73",
          4751 => x"34",
          4752 => x"33",
          4753 => x"9e",
          4754 => x"cc",
          4755 => x"81",
          4756 => x"cc",
          4757 => x"56",
          4758 => x"26",
          4759 => x"ba",
          4760 => x"fc",
          4761 => x"82",
          4762 => x"ee",
          4763 => x"0b",
          4764 => x"34",
          4765 => x"cc",
          4766 => x"9e",
          4767 => x"38",
          4768 => x"08",
          4769 => x"2e",
          4770 => x"51",
          4771 => x"3f",
          4772 => x"08",
          4773 => x"34",
          4774 => x"08",
          4775 => x"81",
          4776 => x"52",
          4777 => x"a8",
          4778 => x"5b",
          4779 => x"7a",
          4780 => x"b4",
          4781 => x"11",
          4782 => x"74",
          4783 => x"38",
          4784 => x"a6",
          4785 => x"b5",
          4786 => x"cc",
          4787 => x"b5",
          4788 => x"ff",
          4789 => x"53",
          4790 => x"51",
          4791 => x"3f",
          4792 => x"80",
          4793 => x"08",
          4794 => x"2e",
          4795 => x"74",
          4796 => x"91",
          4797 => x"7a",
          4798 => x"81",
          4799 => x"82",
          4800 => x"55",
          4801 => x"a4",
          4802 => x"ff",
          4803 => x"82",
          4804 => x"82",
          4805 => x"82",
          4806 => x"81",
          4807 => x"05",
          4808 => x"79",
          4809 => x"bd",
          4810 => x"39",
          4811 => x"82",
          4812 => x"70",
          4813 => x"74",
          4814 => x"38",
          4815 => x"a5",
          4816 => x"b5",
          4817 => x"cc",
          4818 => x"b5",
          4819 => x"ff",
          4820 => x"53",
          4821 => x"51",
          4822 => x"3f",
          4823 => x"73",
          4824 => x"5b",
          4825 => x"82",
          4826 => x"74",
          4827 => x"cc",
          4828 => x"cc",
          4829 => x"79",
          4830 => x"3f",
          4831 => x"82",
          4832 => x"70",
          4833 => x"82",
          4834 => x"59",
          4835 => x"77",
          4836 => x"38",
          4837 => x"08",
          4838 => x"54",
          4839 => x"fc",
          4840 => x"70",
          4841 => x"ff",
          4842 => x"f4",
          4843 => x"cc",
          4844 => x"73",
          4845 => x"e2",
          4846 => x"9c",
          4847 => x"51",
          4848 => x"3f",
          4849 => x"33",
          4850 => x"73",
          4851 => x"34",
          4852 => x"f9",
          4853 => x"bf",
          4854 => x"b5",
          4855 => x"80",
          4856 => x"bc",
          4857 => x"53",
          4858 => x"bf",
          4859 => x"aa",
          4860 => x"b5",
          4861 => x"80",
          4862 => x"34",
          4863 => x"81",
          4864 => x"b5",
          4865 => x"77",
          4866 => x"76",
          4867 => x"82",
          4868 => x"54",
          4869 => x"34",
          4870 => x"34",
          4871 => x"08",
          4872 => x"22",
          4873 => x"80",
          4874 => x"83",
          4875 => x"70",
          4876 => x"51",
          4877 => x"88",
          4878 => x"89",
          4879 => x"b5",
          4880 => x"88",
          4881 => x"c0",
          4882 => x"11",
          4883 => x"77",
          4884 => x"76",
          4885 => x"89",
          4886 => x"ff",
          4887 => x"52",
          4888 => x"72",
          4889 => x"fb",
          4890 => x"82",
          4891 => x"ff",
          4892 => x"51",
          4893 => x"b5",
          4894 => x"3d",
          4895 => x"3d",
          4896 => x"05",
          4897 => x"05",
          4898 => x"71",
          4899 => x"c0",
          4900 => x"2b",
          4901 => x"83",
          4902 => x"70",
          4903 => x"33",
          4904 => x"07",
          4905 => x"ae",
          4906 => x"81",
          4907 => x"07",
          4908 => x"53",
          4909 => x"54",
          4910 => x"53",
          4911 => x"77",
          4912 => x"18",
          4913 => x"c0",
          4914 => x"88",
          4915 => x"70",
          4916 => x"74",
          4917 => x"82",
          4918 => x"70",
          4919 => x"81",
          4920 => x"88",
          4921 => x"83",
          4922 => x"f8",
          4923 => x"56",
          4924 => x"73",
          4925 => x"06",
          4926 => x"54",
          4927 => x"82",
          4928 => x"81",
          4929 => x"72",
          4930 => x"82",
          4931 => x"16",
          4932 => x"34",
          4933 => x"34",
          4934 => x"04",
          4935 => x"82",
          4936 => x"02",
          4937 => x"05",
          4938 => x"2b",
          4939 => x"11",
          4940 => x"33",
          4941 => x"71",
          4942 => x"58",
          4943 => x"55",
          4944 => x"84",
          4945 => x"13",
          4946 => x"2b",
          4947 => x"2a",
          4948 => x"52",
          4949 => x"34",
          4950 => x"34",
          4951 => x"08",
          4952 => x"11",
          4953 => x"33",
          4954 => x"71",
          4955 => x"56",
          4956 => x"72",
          4957 => x"33",
          4958 => x"71",
          4959 => x"70",
          4960 => x"56",
          4961 => x"86",
          4962 => x"87",
          4963 => x"b5",
          4964 => x"70",
          4965 => x"33",
          4966 => x"07",
          4967 => x"ff",
          4968 => x"2a",
          4969 => x"53",
          4970 => x"34",
          4971 => x"34",
          4972 => x"04",
          4973 => x"02",
          4974 => x"82",
          4975 => x"71",
          4976 => x"11",
          4977 => x"12",
          4978 => x"2b",
          4979 => x"29",
          4980 => x"81",
          4981 => x"98",
          4982 => x"2b",
          4983 => x"53",
          4984 => x"56",
          4985 => x"71",
          4986 => x"f6",
          4987 => x"fe",
          4988 => x"b5",
          4989 => x"16",
          4990 => x"12",
          4991 => x"2b",
          4992 => x"07",
          4993 => x"33",
          4994 => x"71",
          4995 => x"70",
          4996 => x"ff",
          4997 => x"52",
          4998 => x"5a",
          4999 => x"05",
          5000 => x"54",
          5001 => x"13",
          5002 => x"13",
          5003 => x"c0",
          5004 => x"70",
          5005 => x"33",
          5006 => x"71",
          5007 => x"56",
          5008 => x"72",
          5009 => x"81",
          5010 => x"88",
          5011 => x"81",
          5012 => x"70",
          5013 => x"51",
          5014 => x"72",
          5015 => x"81",
          5016 => x"3d",
          5017 => x"3d",
          5018 => x"c0",
          5019 => x"05",
          5020 => x"70",
          5021 => x"11",
          5022 => x"83",
          5023 => x"8b",
          5024 => x"2b",
          5025 => x"59",
          5026 => x"73",
          5027 => x"81",
          5028 => x"88",
          5029 => x"8c",
          5030 => x"22",
          5031 => x"88",
          5032 => x"53",
          5033 => x"73",
          5034 => x"14",
          5035 => x"c0",
          5036 => x"70",
          5037 => x"33",
          5038 => x"71",
          5039 => x"56",
          5040 => x"72",
          5041 => x"33",
          5042 => x"71",
          5043 => x"70",
          5044 => x"55",
          5045 => x"82",
          5046 => x"83",
          5047 => x"b5",
          5048 => x"82",
          5049 => x"12",
          5050 => x"2b",
          5051 => x"c8",
          5052 => x"87",
          5053 => x"f7",
          5054 => x"82",
          5055 => x"31",
          5056 => x"83",
          5057 => x"70",
          5058 => x"fd",
          5059 => x"b5",
          5060 => x"83",
          5061 => x"82",
          5062 => x"12",
          5063 => x"2b",
          5064 => x"07",
          5065 => x"33",
          5066 => x"71",
          5067 => x"90",
          5068 => x"42",
          5069 => x"5b",
          5070 => x"54",
          5071 => x"8d",
          5072 => x"80",
          5073 => x"fe",
          5074 => x"84",
          5075 => x"33",
          5076 => x"71",
          5077 => x"83",
          5078 => x"11",
          5079 => x"53",
          5080 => x"55",
          5081 => x"34",
          5082 => x"06",
          5083 => x"14",
          5084 => x"c0",
          5085 => x"84",
          5086 => x"13",
          5087 => x"2b",
          5088 => x"2a",
          5089 => x"56",
          5090 => x"16",
          5091 => x"16",
          5092 => x"c0",
          5093 => x"80",
          5094 => x"34",
          5095 => x"14",
          5096 => x"c0",
          5097 => x"84",
          5098 => x"85",
          5099 => x"b5",
          5100 => x"70",
          5101 => x"33",
          5102 => x"07",
          5103 => x"80",
          5104 => x"2a",
          5105 => x"56",
          5106 => x"34",
          5107 => x"34",
          5108 => x"04",
          5109 => x"73",
          5110 => x"c0",
          5111 => x"f7",
          5112 => x"80",
          5113 => x"71",
          5114 => x"3f",
          5115 => x"04",
          5116 => x"80",
          5117 => x"f8",
          5118 => x"b5",
          5119 => x"ff",
          5120 => x"b5",
          5121 => x"11",
          5122 => x"33",
          5123 => x"07",
          5124 => x"56",
          5125 => x"ff",
          5126 => x"78",
          5127 => x"38",
          5128 => x"17",
          5129 => x"12",
          5130 => x"2b",
          5131 => x"ff",
          5132 => x"31",
          5133 => x"ff",
          5134 => x"27",
          5135 => x"56",
          5136 => x"79",
          5137 => x"73",
          5138 => x"38",
          5139 => x"5b",
          5140 => x"85",
          5141 => x"88",
          5142 => x"54",
          5143 => x"78",
          5144 => x"2e",
          5145 => x"79",
          5146 => x"76",
          5147 => x"b5",
          5148 => x"70",
          5149 => x"33",
          5150 => x"07",
          5151 => x"ff",
          5152 => x"5a",
          5153 => x"73",
          5154 => x"38",
          5155 => x"54",
          5156 => x"81",
          5157 => x"54",
          5158 => x"81",
          5159 => x"7a",
          5160 => x"06",
          5161 => x"51",
          5162 => x"81",
          5163 => x"80",
          5164 => x"52",
          5165 => x"c6",
          5166 => x"c0",
          5167 => x"86",
          5168 => x"12",
          5169 => x"2b",
          5170 => x"07",
          5171 => x"55",
          5172 => x"17",
          5173 => x"ff",
          5174 => x"2a",
          5175 => x"54",
          5176 => x"34",
          5177 => x"06",
          5178 => x"15",
          5179 => x"c0",
          5180 => x"2b",
          5181 => x"1e",
          5182 => x"87",
          5183 => x"88",
          5184 => x"88",
          5185 => x"5e",
          5186 => x"54",
          5187 => x"34",
          5188 => x"34",
          5189 => x"08",
          5190 => x"11",
          5191 => x"33",
          5192 => x"71",
          5193 => x"53",
          5194 => x"74",
          5195 => x"86",
          5196 => x"87",
          5197 => x"b5",
          5198 => x"16",
          5199 => x"11",
          5200 => x"33",
          5201 => x"07",
          5202 => x"53",
          5203 => x"56",
          5204 => x"16",
          5205 => x"16",
          5206 => x"c0",
          5207 => x"05",
          5208 => x"b5",
          5209 => x"3d",
          5210 => x"3d",
          5211 => x"82",
          5212 => x"84",
          5213 => x"3f",
          5214 => x"80",
          5215 => x"71",
          5216 => x"3f",
          5217 => x"08",
          5218 => x"b5",
          5219 => x"3d",
          5220 => x"3d",
          5221 => x"40",
          5222 => x"42",
          5223 => x"c0",
          5224 => x"09",
          5225 => x"38",
          5226 => x"7b",
          5227 => x"51",
          5228 => x"82",
          5229 => x"54",
          5230 => x"7e",
          5231 => x"51",
          5232 => x"7e",
          5233 => x"39",
          5234 => x"8f",
          5235 => x"c8",
          5236 => x"ff",
          5237 => x"c0",
          5238 => x"31",
          5239 => x"83",
          5240 => x"70",
          5241 => x"11",
          5242 => x"12",
          5243 => x"2b",
          5244 => x"31",
          5245 => x"ff",
          5246 => x"29",
          5247 => x"88",
          5248 => x"33",
          5249 => x"71",
          5250 => x"70",
          5251 => x"44",
          5252 => x"41",
          5253 => x"5b",
          5254 => x"5b",
          5255 => x"25",
          5256 => x"81",
          5257 => x"75",
          5258 => x"ff",
          5259 => x"54",
          5260 => x"83",
          5261 => x"88",
          5262 => x"88",
          5263 => x"33",
          5264 => x"71",
          5265 => x"90",
          5266 => x"47",
          5267 => x"54",
          5268 => x"8b",
          5269 => x"31",
          5270 => x"ff",
          5271 => x"77",
          5272 => x"fe",
          5273 => x"54",
          5274 => x"09",
          5275 => x"38",
          5276 => x"c0",
          5277 => x"ff",
          5278 => x"81",
          5279 => x"8e",
          5280 => x"24",
          5281 => x"51",
          5282 => x"81",
          5283 => x"18",
          5284 => x"24",
          5285 => x"79",
          5286 => x"33",
          5287 => x"71",
          5288 => x"53",
          5289 => x"f4",
          5290 => x"78",
          5291 => x"3f",
          5292 => x"08",
          5293 => x"06",
          5294 => x"53",
          5295 => x"82",
          5296 => x"11",
          5297 => x"55",
          5298 => x"cf",
          5299 => x"c0",
          5300 => x"05",
          5301 => x"ff",
          5302 => x"81",
          5303 => x"15",
          5304 => x"24",
          5305 => x"78",
          5306 => x"3f",
          5307 => x"08",
          5308 => x"33",
          5309 => x"71",
          5310 => x"53",
          5311 => x"9c",
          5312 => x"78",
          5313 => x"3f",
          5314 => x"08",
          5315 => x"06",
          5316 => x"53",
          5317 => x"82",
          5318 => x"11",
          5319 => x"55",
          5320 => x"f7",
          5321 => x"c0",
          5322 => x"05",
          5323 => x"19",
          5324 => x"83",
          5325 => x"58",
          5326 => x"7f",
          5327 => x"b0",
          5328 => x"c8",
          5329 => x"b5",
          5330 => x"2e",
          5331 => x"53",
          5332 => x"b5",
          5333 => x"ff",
          5334 => x"73",
          5335 => x"3f",
          5336 => x"78",
          5337 => x"80",
          5338 => x"78",
          5339 => x"3f",
          5340 => x"2b",
          5341 => x"08",
          5342 => x"51",
          5343 => x"7b",
          5344 => x"b5",
          5345 => x"3d",
          5346 => x"3d",
          5347 => x"29",
          5348 => x"fb",
          5349 => x"b5",
          5350 => x"82",
          5351 => x"80",
          5352 => x"73",
          5353 => x"82",
          5354 => x"51",
          5355 => x"3f",
          5356 => x"c8",
          5357 => x"0d",
          5358 => x"0d",
          5359 => x"33",
          5360 => x"70",
          5361 => x"38",
          5362 => x"11",
          5363 => x"82",
          5364 => x"83",
          5365 => x"fc",
          5366 => x"9b",
          5367 => x"84",
          5368 => x"33",
          5369 => x"51",
          5370 => x"80",
          5371 => x"84",
          5372 => x"92",
          5373 => x"51",
          5374 => x"80",
          5375 => x"81",
          5376 => x"72",
          5377 => x"92",
          5378 => x"81",
          5379 => x"0b",
          5380 => x"8c",
          5381 => x"71",
          5382 => x"06",
          5383 => x"80",
          5384 => x"87",
          5385 => x"08",
          5386 => x"38",
          5387 => x"80",
          5388 => x"71",
          5389 => x"c0",
          5390 => x"51",
          5391 => x"87",
          5392 => x"b5",
          5393 => x"82",
          5394 => x"33",
          5395 => x"b5",
          5396 => x"3d",
          5397 => x"3d",
          5398 => x"64",
          5399 => x"bf",
          5400 => x"40",
          5401 => x"74",
          5402 => x"cd",
          5403 => x"c8",
          5404 => x"7a",
          5405 => x"81",
          5406 => x"72",
          5407 => x"87",
          5408 => x"11",
          5409 => x"8c",
          5410 => x"92",
          5411 => x"5a",
          5412 => x"58",
          5413 => x"c0",
          5414 => x"76",
          5415 => x"76",
          5416 => x"70",
          5417 => x"81",
          5418 => x"54",
          5419 => x"8e",
          5420 => x"52",
          5421 => x"81",
          5422 => x"81",
          5423 => x"74",
          5424 => x"53",
          5425 => x"83",
          5426 => x"78",
          5427 => x"8f",
          5428 => x"2e",
          5429 => x"c0",
          5430 => x"52",
          5431 => x"87",
          5432 => x"08",
          5433 => x"2e",
          5434 => x"84",
          5435 => x"38",
          5436 => x"87",
          5437 => x"15",
          5438 => x"70",
          5439 => x"52",
          5440 => x"ff",
          5441 => x"39",
          5442 => x"81",
          5443 => x"ff",
          5444 => x"57",
          5445 => x"90",
          5446 => x"80",
          5447 => x"71",
          5448 => x"78",
          5449 => x"38",
          5450 => x"80",
          5451 => x"80",
          5452 => x"81",
          5453 => x"72",
          5454 => x"0c",
          5455 => x"04",
          5456 => x"60",
          5457 => x"8c",
          5458 => x"33",
          5459 => x"5b",
          5460 => x"74",
          5461 => x"e1",
          5462 => x"c8",
          5463 => x"79",
          5464 => x"78",
          5465 => x"06",
          5466 => x"77",
          5467 => x"87",
          5468 => x"11",
          5469 => x"8c",
          5470 => x"92",
          5471 => x"59",
          5472 => x"85",
          5473 => x"98",
          5474 => x"7d",
          5475 => x"0c",
          5476 => x"08",
          5477 => x"70",
          5478 => x"53",
          5479 => x"2e",
          5480 => x"70",
          5481 => x"33",
          5482 => x"18",
          5483 => x"2a",
          5484 => x"51",
          5485 => x"2e",
          5486 => x"c0",
          5487 => x"52",
          5488 => x"87",
          5489 => x"08",
          5490 => x"2e",
          5491 => x"84",
          5492 => x"38",
          5493 => x"87",
          5494 => x"15",
          5495 => x"70",
          5496 => x"52",
          5497 => x"ff",
          5498 => x"39",
          5499 => x"81",
          5500 => x"80",
          5501 => x"52",
          5502 => x"90",
          5503 => x"80",
          5504 => x"71",
          5505 => x"7a",
          5506 => x"38",
          5507 => x"80",
          5508 => x"80",
          5509 => x"81",
          5510 => x"72",
          5511 => x"0c",
          5512 => x"04",
          5513 => x"7a",
          5514 => x"a3",
          5515 => x"88",
          5516 => x"33",
          5517 => x"56",
          5518 => x"3f",
          5519 => x"08",
          5520 => x"83",
          5521 => x"fe",
          5522 => x"87",
          5523 => x"0c",
          5524 => x"76",
          5525 => x"38",
          5526 => x"93",
          5527 => x"2b",
          5528 => x"8c",
          5529 => x"71",
          5530 => x"38",
          5531 => x"71",
          5532 => x"c6",
          5533 => x"39",
          5534 => x"81",
          5535 => x"06",
          5536 => x"71",
          5537 => x"38",
          5538 => x"8c",
          5539 => x"e8",
          5540 => x"98",
          5541 => x"71",
          5542 => x"73",
          5543 => x"92",
          5544 => x"72",
          5545 => x"06",
          5546 => x"f7",
          5547 => x"80",
          5548 => x"88",
          5549 => x"0c",
          5550 => x"80",
          5551 => x"56",
          5552 => x"56",
          5553 => x"82",
          5554 => x"88",
          5555 => x"fe",
          5556 => x"81",
          5557 => x"33",
          5558 => x"07",
          5559 => x"0c",
          5560 => x"3d",
          5561 => x"3d",
          5562 => x"11",
          5563 => x"33",
          5564 => x"71",
          5565 => x"81",
          5566 => x"72",
          5567 => x"75",
          5568 => x"82",
          5569 => x"52",
          5570 => x"54",
          5571 => x"0d",
          5572 => x"0d",
          5573 => x"05",
          5574 => x"52",
          5575 => x"70",
          5576 => x"34",
          5577 => x"51",
          5578 => x"83",
          5579 => x"ff",
          5580 => x"75",
          5581 => x"72",
          5582 => x"54",
          5583 => x"2a",
          5584 => x"70",
          5585 => x"34",
          5586 => x"51",
          5587 => x"81",
          5588 => x"70",
          5589 => x"70",
          5590 => x"3d",
          5591 => x"3d",
          5592 => x"77",
          5593 => x"70",
          5594 => x"38",
          5595 => x"05",
          5596 => x"70",
          5597 => x"34",
          5598 => x"eb",
          5599 => x"0d",
          5600 => x"0d",
          5601 => x"54",
          5602 => x"72",
          5603 => x"54",
          5604 => x"51",
          5605 => x"84",
          5606 => x"fc",
          5607 => x"77",
          5608 => x"53",
          5609 => x"05",
          5610 => x"70",
          5611 => x"33",
          5612 => x"ff",
          5613 => x"52",
          5614 => x"2e",
          5615 => x"80",
          5616 => x"71",
          5617 => x"0c",
          5618 => x"04",
          5619 => x"74",
          5620 => x"89",
          5621 => x"2e",
          5622 => x"11",
          5623 => x"52",
          5624 => x"70",
          5625 => x"c8",
          5626 => x"0d",
          5627 => x"82",
          5628 => x"04",
          5629 => x"b5",
          5630 => x"f7",
          5631 => x"56",
          5632 => x"17",
          5633 => x"74",
          5634 => x"d6",
          5635 => x"b0",
          5636 => x"b4",
          5637 => x"81",
          5638 => x"59",
          5639 => x"82",
          5640 => x"7a",
          5641 => x"06",
          5642 => x"b5",
          5643 => x"17",
          5644 => x"08",
          5645 => x"08",
          5646 => x"08",
          5647 => x"74",
          5648 => x"38",
          5649 => x"55",
          5650 => x"09",
          5651 => x"38",
          5652 => x"18",
          5653 => x"81",
          5654 => x"f9",
          5655 => x"39",
          5656 => x"82",
          5657 => x"8b",
          5658 => x"fa",
          5659 => x"7a",
          5660 => x"57",
          5661 => x"08",
          5662 => x"75",
          5663 => x"3f",
          5664 => x"08",
          5665 => x"c8",
          5666 => x"81",
          5667 => x"b4",
          5668 => x"16",
          5669 => x"be",
          5670 => x"c8",
          5671 => x"85",
          5672 => x"81",
          5673 => x"17",
          5674 => x"b5",
          5675 => x"3d",
          5676 => x"3d",
          5677 => x"52",
          5678 => x"3f",
          5679 => x"08",
          5680 => x"c8",
          5681 => x"38",
          5682 => x"74",
          5683 => x"81",
          5684 => x"38",
          5685 => x"59",
          5686 => x"09",
          5687 => x"e3",
          5688 => x"53",
          5689 => x"08",
          5690 => x"70",
          5691 => x"91",
          5692 => x"d5",
          5693 => x"17",
          5694 => x"3f",
          5695 => x"a4",
          5696 => x"51",
          5697 => x"86",
          5698 => x"f2",
          5699 => x"17",
          5700 => x"3f",
          5701 => x"52",
          5702 => x"51",
          5703 => x"8c",
          5704 => x"84",
          5705 => x"fc",
          5706 => x"17",
          5707 => x"70",
          5708 => x"79",
          5709 => x"52",
          5710 => x"51",
          5711 => x"77",
          5712 => x"80",
          5713 => x"81",
          5714 => x"f9",
          5715 => x"b5",
          5716 => x"2e",
          5717 => x"58",
          5718 => x"c8",
          5719 => x"0d",
          5720 => x"0d",
          5721 => x"98",
          5722 => x"05",
          5723 => x"80",
          5724 => x"27",
          5725 => x"14",
          5726 => x"29",
          5727 => x"05",
          5728 => x"82",
          5729 => x"87",
          5730 => x"f9",
          5731 => x"7a",
          5732 => x"54",
          5733 => x"27",
          5734 => x"76",
          5735 => x"27",
          5736 => x"ff",
          5737 => x"58",
          5738 => x"80",
          5739 => x"82",
          5740 => x"72",
          5741 => x"38",
          5742 => x"72",
          5743 => x"8e",
          5744 => x"39",
          5745 => x"17",
          5746 => x"a4",
          5747 => x"53",
          5748 => x"fd",
          5749 => x"b5",
          5750 => x"9f",
          5751 => x"ff",
          5752 => x"11",
          5753 => x"70",
          5754 => x"18",
          5755 => x"76",
          5756 => x"53",
          5757 => x"82",
          5758 => x"80",
          5759 => x"83",
          5760 => x"b4",
          5761 => x"88",
          5762 => x"79",
          5763 => x"84",
          5764 => x"58",
          5765 => x"80",
          5766 => x"9f",
          5767 => x"80",
          5768 => x"88",
          5769 => x"08",
          5770 => x"51",
          5771 => x"82",
          5772 => x"80",
          5773 => x"10",
          5774 => x"74",
          5775 => x"51",
          5776 => x"82",
          5777 => x"83",
          5778 => x"58",
          5779 => x"87",
          5780 => x"08",
          5781 => x"51",
          5782 => x"82",
          5783 => x"9b",
          5784 => x"2b",
          5785 => x"74",
          5786 => x"51",
          5787 => x"82",
          5788 => x"f0",
          5789 => x"83",
          5790 => x"77",
          5791 => x"0c",
          5792 => x"04",
          5793 => x"7a",
          5794 => x"58",
          5795 => x"81",
          5796 => x"9e",
          5797 => x"17",
          5798 => x"96",
          5799 => x"53",
          5800 => x"81",
          5801 => x"79",
          5802 => x"72",
          5803 => x"38",
          5804 => x"72",
          5805 => x"b8",
          5806 => x"39",
          5807 => x"17",
          5808 => x"a4",
          5809 => x"53",
          5810 => x"fb",
          5811 => x"b5",
          5812 => x"82",
          5813 => x"81",
          5814 => x"83",
          5815 => x"b4",
          5816 => x"78",
          5817 => x"56",
          5818 => x"76",
          5819 => x"38",
          5820 => x"9f",
          5821 => x"33",
          5822 => x"07",
          5823 => x"74",
          5824 => x"83",
          5825 => x"89",
          5826 => x"08",
          5827 => x"51",
          5828 => x"82",
          5829 => x"59",
          5830 => x"08",
          5831 => x"74",
          5832 => x"16",
          5833 => x"84",
          5834 => x"76",
          5835 => x"88",
          5836 => x"81",
          5837 => x"8f",
          5838 => x"53",
          5839 => x"80",
          5840 => x"88",
          5841 => x"08",
          5842 => x"51",
          5843 => x"82",
          5844 => x"59",
          5845 => x"08",
          5846 => x"77",
          5847 => x"06",
          5848 => x"83",
          5849 => x"05",
          5850 => x"f7",
          5851 => x"39",
          5852 => x"a4",
          5853 => x"52",
          5854 => x"ef",
          5855 => x"c8",
          5856 => x"b5",
          5857 => x"38",
          5858 => x"06",
          5859 => x"83",
          5860 => x"18",
          5861 => x"54",
          5862 => x"f6",
          5863 => x"b5",
          5864 => x"0a",
          5865 => x"52",
          5866 => x"83",
          5867 => x"83",
          5868 => x"82",
          5869 => x"8a",
          5870 => x"f8",
          5871 => x"7c",
          5872 => x"59",
          5873 => x"81",
          5874 => x"38",
          5875 => x"08",
          5876 => x"73",
          5877 => x"38",
          5878 => x"52",
          5879 => x"a4",
          5880 => x"c8",
          5881 => x"b5",
          5882 => x"f2",
          5883 => x"82",
          5884 => x"39",
          5885 => x"e6",
          5886 => x"c8",
          5887 => x"de",
          5888 => x"78",
          5889 => x"3f",
          5890 => x"08",
          5891 => x"c8",
          5892 => x"80",
          5893 => x"b5",
          5894 => x"2e",
          5895 => x"b5",
          5896 => x"2e",
          5897 => x"53",
          5898 => x"51",
          5899 => x"82",
          5900 => x"c5",
          5901 => x"08",
          5902 => x"18",
          5903 => x"57",
          5904 => x"90",
          5905 => x"90",
          5906 => x"16",
          5907 => x"54",
          5908 => x"34",
          5909 => x"78",
          5910 => x"38",
          5911 => x"82",
          5912 => x"8a",
          5913 => x"f6",
          5914 => x"7e",
          5915 => x"5b",
          5916 => x"38",
          5917 => x"58",
          5918 => x"88",
          5919 => x"08",
          5920 => x"38",
          5921 => x"39",
          5922 => x"51",
          5923 => x"81",
          5924 => x"b5",
          5925 => x"82",
          5926 => x"b5",
          5927 => x"82",
          5928 => x"ff",
          5929 => x"38",
          5930 => x"82",
          5931 => x"26",
          5932 => x"79",
          5933 => x"08",
          5934 => x"73",
          5935 => x"b9",
          5936 => x"2e",
          5937 => x"80",
          5938 => x"1a",
          5939 => x"08",
          5940 => x"38",
          5941 => x"52",
          5942 => x"af",
          5943 => x"82",
          5944 => x"81",
          5945 => x"06",
          5946 => x"b5",
          5947 => x"82",
          5948 => x"09",
          5949 => x"72",
          5950 => x"70",
          5951 => x"b5",
          5952 => x"51",
          5953 => x"73",
          5954 => x"82",
          5955 => x"80",
          5956 => x"8c",
          5957 => x"81",
          5958 => x"38",
          5959 => x"08",
          5960 => x"73",
          5961 => x"75",
          5962 => x"77",
          5963 => x"56",
          5964 => x"76",
          5965 => x"82",
          5966 => x"26",
          5967 => x"75",
          5968 => x"f8",
          5969 => x"b5",
          5970 => x"2e",
          5971 => x"59",
          5972 => x"08",
          5973 => x"81",
          5974 => x"82",
          5975 => x"59",
          5976 => x"08",
          5977 => x"70",
          5978 => x"25",
          5979 => x"51",
          5980 => x"73",
          5981 => x"75",
          5982 => x"81",
          5983 => x"38",
          5984 => x"f5",
          5985 => x"75",
          5986 => x"f9",
          5987 => x"b5",
          5988 => x"b5",
          5989 => x"70",
          5990 => x"08",
          5991 => x"51",
          5992 => x"80",
          5993 => x"73",
          5994 => x"38",
          5995 => x"52",
          5996 => x"d0",
          5997 => x"c8",
          5998 => x"a5",
          5999 => x"18",
          6000 => x"08",
          6001 => x"18",
          6002 => x"74",
          6003 => x"38",
          6004 => x"18",
          6005 => x"33",
          6006 => x"73",
          6007 => x"97",
          6008 => x"74",
          6009 => x"38",
          6010 => x"55",
          6011 => x"b5",
          6012 => x"85",
          6013 => x"75",
          6014 => x"b5",
          6015 => x"3d",
          6016 => x"3d",
          6017 => x"52",
          6018 => x"3f",
          6019 => x"08",
          6020 => x"82",
          6021 => x"80",
          6022 => x"52",
          6023 => x"c1",
          6024 => x"c8",
          6025 => x"c8",
          6026 => x"0c",
          6027 => x"53",
          6028 => x"15",
          6029 => x"f2",
          6030 => x"56",
          6031 => x"16",
          6032 => x"22",
          6033 => x"27",
          6034 => x"54",
          6035 => x"76",
          6036 => x"33",
          6037 => x"3f",
          6038 => x"08",
          6039 => x"38",
          6040 => x"76",
          6041 => x"70",
          6042 => x"9f",
          6043 => x"56",
          6044 => x"b5",
          6045 => x"3d",
          6046 => x"3d",
          6047 => x"71",
          6048 => x"57",
          6049 => x"0a",
          6050 => x"38",
          6051 => x"53",
          6052 => x"38",
          6053 => x"0c",
          6054 => x"54",
          6055 => x"75",
          6056 => x"73",
          6057 => x"a8",
          6058 => x"73",
          6059 => x"85",
          6060 => x"0b",
          6061 => x"5a",
          6062 => x"27",
          6063 => x"a8",
          6064 => x"18",
          6065 => x"39",
          6066 => x"70",
          6067 => x"58",
          6068 => x"b2",
          6069 => x"76",
          6070 => x"3f",
          6071 => x"08",
          6072 => x"c8",
          6073 => x"bd",
          6074 => x"82",
          6075 => x"27",
          6076 => x"16",
          6077 => x"c8",
          6078 => x"38",
          6079 => x"39",
          6080 => x"55",
          6081 => x"52",
          6082 => x"d5",
          6083 => x"c8",
          6084 => x"0c",
          6085 => x"0c",
          6086 => x"53",
          6087 => x"80",
          6088 => x"85",
          6089 => x"94",
          6090 => x"2a",
          6091 => x"0c",
          6092 => x"06",
          6093 => x"9c",
          6094 => x"58",
          6095 => x"c8",
          6096 => x"0d",
          6097 => x"0d",
          6098 => x"90",
          6099 => x"05",
          6100 => x"f0",
          6101 => x"27",
          6102 => x"0b",
          6103 => x"98",
          6104 => x"84",
          6105 => x"2e",
          6106 => x"76",
          6107 => x"58",
          6108 => x"38",
          6109 => x"15",
          6110 => x"08",
          6111 => x"38",
          6112 => x"88",
          6113 => x"53",
          6114 => x"81",
          6115 => x"c0",
          6116 => x"22",
          6117 => x"89",
          6118 => x"72",
          6119 => x"74",
          6120 => x"f3",
          6121 => x"b5",
          6122 => x"82",
          6123 => x"82",
          6124 => x"27",
          6125 => x"81",
          6126 => x"c8",
          6127 => x"80",
          6128 => x"16",
          6129 => x"c8",
          6130 => x"ca",
          6131 => x"38",
          6132 => x"0c",
          6133 => x"dd",
          6134 => x"08",
          6135 => x"f9",
          6136 => x"b5",
          6137 => x"87",
          6138 => x"c8",
          6139 => x"80",
          6140 => x"55",
          6141 => x"08",
          6142 => x"38",
          6143 => x"b5",
          6144 => x"2e",
          6145 => x"b5",
          6146 => x"75",
          6147 => x"3f",
          6148 => x"08",
          6149 => x"94",
          6150 => x"52",
          6151 => x"c1",
          6152 => x"c8",
          6153 => x"0c",
          6154 => x"0c",
          6155 => x"05",
          6156 => x"80",
          6157 => x"b5",
          6158 => x"3d",
          6159 => x"3d",
          6160 => x"71",
          6161 => x"57",
          6162 => x"51",
          6163 => x"82",
          6164 => x"54",
          6165 => x"08",
          6166 => x"82",
          6167 => x"56",
          6168 => x"52",
          6169 => x"83",
          6170 => x"c8",
          6171 => x"b5",
          6172 => x"d2",
          6173 => x"c8",
          6174 => x"08",
          6175 => x"54",
          6176 => x"e5",
          6177 => x"06",
          6178 => x"58",
          6179 => x"08",
          6180 => x"38",
          6181 => x"75",
          6182 => x"80",
          6183 => x"81",
          6184 => x"7a",
          6185 => x"06",
          6186 => x"39",
          6187 => x"08",
          6188 => x"76",
          6189 => x"3f",
          6190 => x"08",
          6191 => x"c8",
          6192 => x"ff",
          6193 => x"84",
          6194 => x"06",
          6195 => x"54",
          6196 => x"c8",
          6197 => x"0d",
          6198 => x"0d",
          6199 => x"52",
          6200 => x"3f",
          6201 => x"08",
          6202 => x"06",
          6203 => x"51",
          6204 => x"83",
          6205 => x"06",
          6206 => x"14",
          6207 => x"3f",
          6208 => x"08",
          6209 => x"07",
          6210 => x"b5",
          6211 => x"3d",
          6212 => x"3d",
          6213 => x"70",
          6214 => x"06",
          6215 => x"53",
          6216 => x"ed",
          6217 => x"33",
          6218 => x"83",
          6219 => x"06",
          6220 => x"90",
          6221 => x"15",
          6222 => x"3f",
          6223 => x"04",
          6224 => x"7b",
          6225 => x"84",
          6226 => x"58",
          6227 => x"80",
          6228 => x"38",
          6229 => x"52",
          6230 => x"8f",
          6231 => x"c8",
          6232 => x"b5",
          6233 => x"f5",
          6234 => x"08",
          6235 => x"53",
          6236 => x"84",
          6237 => x"39",
          6238 => x"70",
          6239 => x"81",
          6240 => x"51",
          6241 => x"16",
          6242 => x"c8",
          6243 => x"81",
          6244 => x"38",
          6245 => x"ae",
          6246 => x"81",
          6247 => x"54",
          6248 => x"2e",
          6249 => x"8f",
          6250 => x"82",
          6251 => x"76",
          6252 => x"54",
          6253 => x"09",
          6254 => x"38",
          6255 => x"7a",
          6256 => x"80",
          6257 => x"fa",
          6258 => x"b5",
          6259 => x"82",
          6260 => x"89",
          6261 => x"08",
          6262 => x"86",
          6263 => x"98",
          6264 => x"82",
          6265 => x"8b",
          6266 => x"fb",
          6267 => x"70",
          6268 => x"81",
          6269 => x"fc",
          6270 => x"b5",
          6271 => x"82",
          6272 => x"b4",
          6273 => x"08",
          6274 => x"ec",
          6275 => x"b5",
          6276 => x"82",
          6277 => x"a0",
          6278 => x"82",
          6279 => x"52",
          6280 => x"51",
          6281 => x"8b",
          6282 => x"52",
          6283 => x"51",
          6284 => x"81",
          6285 => x"34",
          6286 => x"c8",
          6287 => x"0d",
          6288 => x"0d",
          6289 => x"98",
          6290 => x"70",
          6291 => x"ec",
          6292 => x"b5",
          6293 => x"38",
          6294 => x"53",
          6295 => x"81",
          6296 => x"34",
          6297 => x"04",
          6298 => x"78",
          6299 => x"80",
          6300 => x"34",
          6301 => x"80",
          6302 => x"38",
          6303 => x"18",
          6304 => x"9c",
          6305 => x"70",
          6306 => x"56",
          6307 => x"a0",
          6308 => x"71",
          6309 => x"81",
          6310 => x"81",
          6311 => x"89",
          6312 => x"06",
          6313 => x"73",
          6314 => x"55",
          6315 => x"55",
          6316 => x"81",
          6317 => x"81",
          6318 => x"74",
          6319 => x"75",
          6320 => x"52",
          6321 => x"13",
          6322 => x"08",
          6323 => x"33",
          6324 => x"9c",
          6325 => x"11",
          6326 => x"8a",
          6327 => x"c8",
          6328 => x"96",
          6329 => x"e7",
          6330 => x"c8",
          6331 => x"23",
          6332 => x"e7",
          6333 => x"b5",
          6334 => x"17",
          6335 => x"0d",
          6336 => x"0d",
          6337 => x"5e",
          6338 => x"70",
          6339 => x"55",
          6340 => x"83",
          6341 => x"73",
          6342 => x"91",
          6343 => x"2e",
          6344 => x"1d",
          6345 => x"0c",
          6346 => x"15",
          6347 => x"70",
          6348 => x"56",
          6349 => x"09",
          6350 => x"38",
          6351 => x"80",
          6352 => x"30",
          6353 => x"78",
          6354 => x"54",
          6355 => x"73",
          6356 => x"60",
          6357 => x"54",
          6358 => x"96",
          6359 => x"0b",
          6360 => x"80",
          6361 => x"f6",
          6362 => x"b5",
          6363 => x"85",
          6364 => x"3d",
          6365 => x"5c",
          6366 => x"53",
          6367 => x"51",
          6368 => x"80",
          6369 => x"88",
          6370 => x"5c",
          6371 => x"09",
          6372 => x"d4",
          6373 => x"70",
          6374 => x"71",
          6375 => x"30",
          6376 => x"73",
          6377 => x"51",
          6378 => x"57",
          6379 => x"38",
          6380 => x"75",
          6381 => x"17",
          6382 => x"75",
          6383 => x"30",
          6384 => x"51",
          6385 => x"80",
          6386 => x"38",
          6387 => x"87",
          6388 => x"26",
          6389 => x"77",
          6390 => x"a4",
          6391 => x"27",
          6392 => x"a0",
          6393 => x"39",
          6394 => x"33",
          6395 => x"57",
          6396 => x"27",
          6397 => x"75",
          6398 => x"30",
          6399 => x"32",
          6400 => x"80",
          6401 => x"25",
          6402 => x"56",
          6403 => x"80",
          6404 => x"84",
          6405 => x"58",
          6406 => x"70",
          6407 => x"55",
          6408 => x"09",
          6409 => x"38",
          6410 => x"80",
          6411 => x"30",
          6412 => x"77",
          6413 => x"54",
          6414 => x"81",
          6415 => x"ae",
          6416 => x"06",
          6417 => x"54",
          6418 => x"74",
          6419 => x"80",
          6420 => x"7b",
          6421 => x"30",
          6422 => x"70",
          6423 => x"25",
          6424 => x"07",
          6425 => x"51",
          6426 => x"a7",
          6427 => x"8b",
          6428 => x"39",
          6429 => x"54",
          6430 => x"8c",
          6431 => x"ff",
          6432 => x"90",
          6433 => x"54",
          6434 => x"e1",
          6435 => x"c8",
          6436 => x"b2",
          6437 => x"70",
          6438 => x"71",
          6439 => x"54",
          6440 => x"82",
          6441 => x"80",
          6442 => x"38",
          6443 => x"76",
          6444 => x"df",
          6445 => x"54",
          6446 => x"81",
          6447 => x"55",
          6448 => x"34",
          6449 => x"52",
          6450 => x"51",
          6451 => x"82",
          6452 => x"bf",
          6453 => x"16",
          6454 => x"26",
          6455 => x"16",
          6456 => x"06",
          6457 => x"17",
          6458 => x"34",
          6459 => x"fd",
          6460 => x"19",
          6461 => x"80",
          6462 => x"79",
          6463 => x"81",
          6464 => x"81",
          6465 => x"85",
          6466 => x"54",
          6467 => x"8f",
          6468 => x"86",
          6469 => x"39",
          6470 => x"f3",
          6471 => x"73",
          6472 => x"80",
          6473 => x"52",
          6474 => x"ce",
          6475 => x"c8",
          6476 => x"b5",
          6477 => x"d7",
          6478 => x"08",
          6479 => x"e6",
          6480 => x"b5",
          6481 => x"82",
          6482 => x"80",
          6483 => x"1b",
          6484 => x"55",
          6485 => x"2e",
          6486 => x"8b",
          6487 => x"06",
          6488 => x"1c",
          6489 => x"33",
          6490 => x"70",
          6491 => x"55",
          6492 => x"38",
          6493 => x"52",
          6494 => x"9f",
          6495 => x"c8",
          6496 => x"8b",
          6497 => x"7a",
          6498 => x"3f",
          6499 => x"75",
          6500 => x"57",
          6501 => x"2e",
          6502 => x"84",
          6503 => x"06",
          6504 => x"75",
          6505 => x"81",
          6506 => x"2a",
          6507 => x"73",
          6508 => x"38",
          6509 => x"54",
          6510 => x"fb",
          6511 => x"80",
          6512 => x"34",
          6513 => x"c1",
          6514 => x"06",
          6515 => x"38",
          6516 => x"39",
          6517 => x"70",
          6518 => x"54",
          6519 => x"86",
          6520 => x"84",
          6521 => x"06",
          6522 => x"73",
          6523 => x"38",
          6524 => x"83",
          6525 => x"b4",
          6526 => x"51",
          6527 => x"82",
          6528 => x"88",
          6529 => x"ea",
          6530 => x"b5",
          6531 => x"3d",
          6532 => x"3d",
          6533 => x"ff",
          6534 => x"71",
          6535 => x"5c",
          6536 => x"80",
          6537 => x"38",
          6538 => x"05",
          6539 => x"a0",
          6540 => x"71",
          6541 => x"38",
          6542 => x"71",
          6543 => x"81",
          6544 => x"38",
          6545 => x"11",
          6546 => x"06",
          6547 => x"70",
          6548 => x"38",
          6549 => x"81",
          6550 => x"05",
          6551 => x"76",
          6552 => x"38",
          6553 => x"af",
          6554 => x"77",
          6555 => x"57",
          6556 => x"05",
          6557 => x"70",
          6558 => x"33",
          6559 => x"53",
          6560 => x"99",
          6561 => x"e0",
          6562 => x"ff",
          6563 => x"ff",
          6564 => x"70",
          6565 => x"38",
          6566 => x"81",
          6567 => x"51",
          6568 => x"9f",
          6569 => x"72",
          6570 => x"81",
          6571 => x"70",
          6572 => x"72",
          6573 => x"32",
          6574 => x"72",
          6575 => x"73",
          6576 => x"53",
          6577 => x"70",
          6578 => x"38",
          6579 => x"19",
          6580 => x"75",
          6581 => x"38",
          6582 => x"83",
          6583 => x"74",
          6584 => x"59",
          6585 => x"39",
          6586 => x"33",
          6587 => x"b5",
          6588 => x"3d",
          6589 => x"3d",
          6590 => x"80",
          6591 => x"34",
          6592 => x"17",
          6593 => x"75",
          6594 => x"3f",
          6595 => x"b5",
          6596 => x"80",
          6597 => x"16",
          6598 => x"3f",
          6599 => x"08",
          6600 => x"06",
          6601 => x"73",
          6602 => x"2e",
          6603 => x"80",
          6604 => x"0b",
          6605 => x"56",
          6606 => x"e9",
          6607 => x"06",
          6608 => x"57",
          6609 => x"32",
          6610 => x"80",
          6611 => x"51",
          6612 => x"8a",
          6613 => x"e8",
          6614 => x"06",
          6615 => x"53",
          6616 => x"52",
          6617 => x"51",
          6618 => x"82",
          6619 => x"55",
          6620 => x"08",
          6621 => x"38",
          6622 => x"ae",
          6623 => x"86",
          6624 => x"97",
          6625 => x"c8",
          6626 => x"b5",
          6627 => x"2e",
          6628 => x"55",
          6629 => x"c8",
          6630 => x"0d",
          6631 => x"0d",
          6632 => x"05",
          6633 => x"33",
          6634 => x"75",
          6635 => x"fc",
          6636 => x"b5",
          6637 => x"8b",
          6638 => x"82",
          6639 => x"24",
          6640 => x"82",
          6641 => x"84",
          6642 => x"80",
          6643 => x"55",
          6644 => x"73",
          6645 => x"e6",
          6646 => x"0c",
          6647 => x"06",
          6648 => x"57",
          6649 => x"ae",
          6650 => x"33",
          6651 => x"3f",
          6652 => x"08",
          6653 => x"70",
          6654 => x"55",
          6655 => x"76",
          6656 => x"b8",
          6657 => x"2a",
          6658 => x"51",
          6659 => x"72",
          6660 => x"86",
          6661 => x"74",
          6662 => x"15",
          6663 => x"81",
          6664 => x"d7",
          6665 => x"b5",
          6666 => x"ff",
          6667 => x"06",
          6668 => x"56",
          6669 => x"38",
          6670 => x"8f",
          6671 => x"2a",
          6672 => x"51",
          6673 => x"72",
          6674 => x"80",
          6675 => x"52",
          6676 => x"3f",
          6677 => x"08",
          6678 => x"57",
          6679 => x"09",
          6680 => x"e2",
          6681 => x"74",
          6682 => x"56",
          6683 => x"33",
          6684 => x"72",
          6685 => x"38",
          6686 => x"51",
          6687 => x"82",
          6688 => x"57",
          6689 => x"84",
          6690 => x"ff",
          6691 => x"56",
          6692 => x"25",
          6693 => x"0b",
          6694 => x"56",
          6695 => x"05",
          6696 => x"83",
          6697 => x"2e",
          6698 => x"52",
          6699 => x"c6",
          6700 => x"c8",
          6701 => x"06",
          6702 => x"27",
          6703 => x"16",
          6704 => x"27",
          6705 => x"56",
          6706 => x"84",
          6707 => x"56",
          6708 => x"84",
          6709 => x"14",
          6710 => x"3f",
          6711 => x"08",
          6712 => x"06",
          6713 => x"80",
          6714 => x"06",
          6715 => x"80",
          6716 => x"db",
          6717 => x"b5",
          6718 => x"ff",
          6719 => x"77",
          6720 => x"d8",
          6721 => x"de",
          6722 => x"c8",
          6723 => x"9c",
          6724 => x"c4",
          6725 => x"15",
          6726 => x"14",
          6727 => x"70",
          6728 => x"51",
          6729 => x"56",
          6730 => x"84",
          6731 => x"81",
          6732 => x"71",
          6733 => x"16",
          6734 => x"53",
          6735 => x"23",
          6736 => x"8b",
          6737 => x"73",
          6738 => x"80",
          6739 => x"8d",
          6740 => x"39",
          6741 => x"51",
          6742 => x"82",
          6743 => x"53",
          6744 => x"08",
          6745 => x"72",
          6746 => x"8d",
          6747 => x"ce",
          6748 => x"14",
          6749 => x"3f",
          6750 => x"08",
          6751 => x"06",
          6752 => x"38",
          6753 => x"51",
          6754 => x"82",
          6755 => x"55",
          6756 => x"51",
          6757 => x"82",
          6758 => x"83",
          6759 => x"53",
          6760 => x"80",
          6761 => x"38",
          6762 => x"78",
          6763 => x"2a",
          6764 => x"78",
          6765 => x"86",
          6766 => x"22",
          6767 => x"31",
          6768 => x"bf",
          6769 => x"c8",
          6770 => x"b5",
          6771 => x"2e",
          6772 => x"82",
          6773 => x"80",
          6774 => x"f5",
          6775 => x"83",
          6776 => x"ff",
          6777 => x"38",
          6778 => x"9f",
          6779 => x"38",
          6780 => x"39",
          6781 => x"80",
          6782 => x"38",
          6783 => x"98",
          6784 => x"a0",
          6785 => x"1c",
          6786 => x"0c",
          6787 => x"17",
          6788 => x"76",
          6789 => x"81",
          6790 => x"80",
          6791 => x"d9",
          6792 => x"b5",
          6793 => x"ff",
          6794 => x"8d",
          6795 => x"8e",
          6796 => x"8a",
          6797 => x"14",
          6798 => x"3f",
          6799 => x"08",
          6800 => x"74",
          6801 => x"a2",
          6802 => x"79",
          6803 => x"ee",
          6804 => x"a8",
          6805 => x"15",
          6806 => x"2e",
          6807 => x"10",
          6808 => x"2a",
          6809 => x"05",
          6810 => x"ff",
          6811 => x"53",
          6812 => x"9c",
          6813 => x"81",
          6814 => x"0b",
          6815 => x"ff",
          6816 => x"0c",
          6817 => x"84",
          6818 => x"83",
          6819 => x"06",
          6820 => x"80",
          6821 => x"d8",
          6822 => x"b5",
          6823 => x"ff",
          6824 => x"72",
          6825 => x"81",
          6826 => x"38",
          6827 => x"73",
          6828 => x"3f",
          6829 => x"08",
          6830 => x"82",
          6831 => x"84",
          6832 => x"b2",
          6833 => x"87",
          6834 => x"c8",
          6835 => x"ff",
          6836 => x"82",
          6837 => x"09",
          6838 => x"c8",
          6839 => x"51",
          6840 => x"82",
          6841 => x"84",
          6842 => x"d2",
          6843 => x"06",
          6844 => x"98",
          6845 => x"ee",
          6846 => x"c8",
          6847 => x"85",
          6848 => x"09",
          6849 => x"38",
          6850 => x"51",
          6851 => x"82",
          6852 => x"90",
          6853 => x"a0",
          6854 => x"ca",
          6855 => x"c8",
          6856 => x"0c",
          6857 => x"82",
          6858 => x"81",
          6859 => x"82",
          6860 => x"72",
          6861 => x"80",
          6862 => x"0c",
          6863 => x"82",
          6864 => x"90",
          6865 => x"fb",
          6866 => x"54",
          6867 => x"80",
          6868 => x"73",
          6869 => x"80",
          6870 => x"72",
          6871 => x"80",
          6872 => x"86",
          6873 => x"15",
          6874 => x"71",
          6875 => x"81",
          6876 => x"81",
          6877 => x"d0",
          6878 => x"b5",
          6879 => x"06",
          6880 => x"38",
          6881 => x"54",
          6882 => x"80",
          6883 => x"71",
          6884 => x"82",
          6885 => x"87",
          6886 => x"fa",
          6887 => x"ab",
          6888 => x"58",
          6889 => x"05",
          6890 => x"e6",
          6891 => x"80",
          6892 => x"c8",
          6893 => x"38",
          6894 => x"08",
          6895 => x"cd",
          6896 => x"08",
          6897 => x"80",
          6898 => x"80",
          6899 => x"54",
          6900 => x"84",
          6901 => x"34",
          6902 => x"75",
          6903 => x"2e",
          6904 => x"53",
          6905 => x"53",
          6906 => x"f7",
          6907 => x"b5",
          6908 => x"73",
          6909 => x"0c",
          6910 => x"04",
          6911 => x"67",
          6912 => x"80",
          6913 => x"59",
          6914 => x"78",
          6915 => x"c8",
          6916 => x"06",
          6917 => x"3d",
          6918 => x"99",
          6919 => x"52",
          6920 => x"3f",
          6921 => x"08",
          6922 => x"c8",
          6923 => x"38",
          6924 => x"52",
          6925 => x"52",
          6926 => x"3f",
          6927 => x"08",
          6928 => x"c8",
          6929 => x"02",
          6930 => x"33",
          6931 => x"55",
          6932 => x"25",
          6933 => x"55",
          6934 => x"54",
          6935 => x"81",
          6936 => x"80",
          6937 => x"74",
          6938 => x"81",
          6939 => x"75",
          6940 => x"3f",
          6941 => x"08",
          6942 => x"02",
          6943 => x"91",
          6944 => x"81",
          6945 => x"82",
          6946 => x"06",
          6947 => x"80",
          6948 => x"88",
          6949 => x"39",
          6950 => x"58",
          6951 => x"38",
          6952 => x"70",
          6953 => x"54",
          6954 => x"81",
          6955 => x"52",
          6956 => x"a5",
          6957 => x"c8",
          6958 => x"88",
          6959 => x"62",
          6960 => x"d4",
          6961 => x"54",
          6962 => x"15",
          6963 => x"62",
          6964 => x"e8",
          6965 => x"52",
          6966 => x"51",
          6967 => x"7a",
          6968 => x"83",
          6969 => x"80",
          6970 => x"38",
          6971 => x"08",
          6972 => x"53",
          6973 => x"3d",
          6974 => x"dd",
          6975 => x"b5",
          6976 => x"82",
          6977 => x"82",
          6978 => x"39",
          6979 => x"38",
          6980 => x"33",
          6981 => x"70",
          6982 => x"55",
          6983 => x"2e",
          6984 => x"55",
          6985 => x"77",
          6986 => x"81",
          6987 => x"73",
          6988 => x"38",
          6989 => x"54",
          6990 => x"a0",
          6991 => x"82",
          6992 => x"52",
          6993 => x"a3",
          6994 => x"c8",
          6995 => x"18",
          6996 => x"55",
          6997 => x"c8",
          6998 => x"38",
          6999 => x"70",
          7000 => x"54",
          7001 => x"86",
          7002 => x"c0",
          7003 => x"b0",
          7004 => x"1b",
          7005 => x"1b",
          7006 => x"70",
          7007 => x"d9",
          7008 => x"c8",
          7009 => x"c8",
          7010 => x"0c",
          7011 => x"52",
          7012 => x"3f",
          7013 => x"08",
          7014 => x"08",
          7015 => x"77",
          7016 => x"86",
          7017 => x"1a",
          7018 => x"1a",
          7019 => x"91",
          7020 => x"0b",
          7021 => x"80",
          7022 => x"0c",
          7023 => x"70",
          7024 => x"54",
          7025 => x"81",
          7026 => x"b5",
          7027 => x"2e",
          7028 => x"82",
          7029 => x"94",
          7030 => x"17",
          7031 => x"2b",
          7032 => x"57",
          7033 => x"52",
          7034 => x"9f",
          7035 => x"c8",
          7036 => x"b5",
          7037 => x"26",
          7038 => x"55",
          7039 => x"08",
          7040 => x"81",
          7041 => x"79",
          7042 => x"31",
          7043 => x"70",
          7044 => x"25",
          7045 => x"76",
          7046 => x"81",
          7047 => x"55",
          7048 => x"38",
          7049 => x"0c",
          7050 => x"75",
          7051 => x"54",
          7052 => x"a2",
          7053 => x"7a",
          7054 => x"3f",
          7055 => x"08",
          7056 => x"55",
          7057 => x"89",
          7058 => x"c8",
          7059 => x"1a",
          7060 => x"80",
          7061 => x"54",
          7062 => x"c8",
          7063 => x"0d",
          7064 => x"0d",
          7065 => x"64",
          7066 => x"59",
          7067 => x"90",
          7068 => x"52",
          7069 => x"cf",
          7070 => x"c8",
          7071 => x"b5",
          7072 => x"38",
          7073 => x"55",
          7074 => x"86",
          7075 => x"82",
          7076 => x"19",
          7077 => x"55",
          7078 => x"80",
          7079 => x"38",
          7080 => x"0b",
          7081 => x"82",
          7082 => x"39",
          7083 => x"1a",
          7084 => x"82",
          7085 => x"19",
          7086 => x"08",
          7087 => x"7c",
          7088 => x"74",
          7089 => x"2e",
          7090 => x"94",
          7091 => x"83",
          7092 => x"56",
          7093 => x"38",
          7094 => x"22",
          7095 => x"89",
          7096 => x"55",
          7097 => x"75",
          7098 => x"19",
          7099 => x"39",
          7100 => x"52",
          7101 => x"93",
          7102 => x"c8",
          7103 => x"75",
          7104 => x"38",
          7105 => x"ff",
          7106 => x"98",
          7107 => x"19",
          7108 => x"51",
          7109 => x"82",
          7110 => x"80",
          7111 => x"38",
          7112 => x"08",
          7113 => x"2a",
          7114 => x"80",
          7115 => x"38",
          7116 => x"8a",
          7117 => x"5c",
          7118 => x"27",
          7119 => x"7a",
          7120 => x"54",
          7121 => x"52",
          7122 => x"51",
          7123 => x"82",
          7124 => x"fe",
          7125 => x"83",
          7126 => x"56",
          7127 => x"9f",
          7128 => x"08",
          7129 => x"74",
          7130 => x"38",
          7131 => x"b4",
          7132 => x"16",
          7133 => x"89",
          7134 => x"51",
          7135 => x"77",
          7136 => x"b9",
          7137 => x"1a",
          7138 => x"08",
          7139 => x"84",
          7140 => x"57",
          7141 => x"27",
          7142 => x"56",
          7143 => x"52",
          7144 => x"c7",
          7145 => x"c8",
          7146 => x"38",
          7147 => x"19",
          7148 => x"06",
          7149 => x"52",
          7150 => x"a2",
          7151 => x"31",
          7152 => x"7f",
          7153 => x"94",
          7154 => x"94",
          7155 => x"5c",
          7156 => x"80",
          7157 => x"b5",
          7158 => x"3d",
          7159 => x"3d",
          7160 => x"65",
          7161 => x"5d",
          7162 => x"0c",
          7163 => x"05",
          7164 => x"f6",
          7165 => x"b5",
          7166 => x"82",
          7167 => x"8a",
          7168 => x"33",
          7169 => x"2e",
          7170 => x"56",
          7171 => x"90",
          7172 => x"81",
          7173 => x"06",
          7174 => x"87",
          7175 => x"2e",
          7176 => x"95",
          7177 => x"91",
          7178 => x"56",
          7179 => x"81",
          7180 => x"34",
          7181 => x"8e",
          7182 => x"08",
          7183 => x"56",
          7184 => x"84",
          7185 => x"5c",
          7186 => x"82",
          7187 => x"18",
          7188 => x"ff",
          7189 => x"74",
          7190 => x"7e",
          7191 => x"ff",
          7192 => x"2a",
          7193 => x"7a",
          7194 => x"8c",
          7195 => x"08",
          7196 => x"38",
          7197 => x"39",
          7198 => x"52",
          7199 => x"e7",
          7200 => x"c8",
          7201 => x"b5",
          7202 => x"2e",
          7203 => x"74",
          7204 => x"91",
          7205 => x"2e",
          7206 => x"74",
          7207 => x"88",
          7208 => x"38",
          7209 => x"0c",
          7210 => x"15",
          7211 => x"08",
          7212 => x"06",
          7213 => x"51",
          7214 => x"82",
          7215 => x"fe",
          7216 => x"18",
          7217 => x"51",
          7218 => x"82",
          7219 => x"80",
          7220 => x"38",
          7221 => x"08",
          7222 => x"2a",
          7223 => x"80",
          7224 => x"38",
          7225 => x"8a",
          7226 => x"5b",
          7227 => x"27",
          7228 => x"7b",
          7229 => x"54",
          7230 => x"52",
          7231 => x"51",
          7232 => x"82",
          7233 => x"fe",
          7234 => x"b0",
          7235 => x"31",
          7236 => x"79",
          7237 => x"84",
          7238 => x"16",
          7239 => x"89",
          7240 => x"52",
          7241 => x"cc",
          7242 => x"55",
          7243 => x"16",
          7244 => x"2b",
          7245 => x"39",
          7246 => x"94",
          7247 => x"93",
          7248 => x"cd",
          7249 => x"b5",
          7250 => x"e3",
          7251 => x"b0",
          7252 => x"76",
          7253 => x"94",
          7254 => x"ff",
          7255 => x"71",
          7256 => x"7b",
          7257 => x"38",
          7258 => x"18",
          7259 => x"51",
          7260 => x"82",
          7261 => x"fd",
          7262 => x"53",
          7263 => x"18",
          7264 => x"06",
          7265 => x"51",
          7266 => x"7e",
          7267 => x"83",
          7268 => x"76",
          7269 => x"17",
          7270 => x"1e",
          7271 => x"18",
          7272 => x"0c",
          7273 => x"58",
          7274 => x"74",
          7275 => x"38",
          7276 => x"8c",
          7277 => x"90",
          7278 => x"33",
          7279 => x"55",
          7280 => x"34",
          7281 => x"82",
          7282 => x"90",
          7283 => x"f8",
          7284 => x"8b",
          7285 => x"53",
          7286 => x"f2",
          7287 => x"b5",
          7288 => x"82",
          7289 => x"80",
          7290 => x"16",
          7291 => x"2a",
          7292 => x"51",
          7293 => x"80",
          7294 => x"38",
          7295 => x"52",
          7296 => x"e7",
          7297 => x"c8",
          7298 => x"b5",
          7299 => x"d4",
          7300 => x"08",
          7301 => x"a0",
          7302 => x"73",
          7303 => x"88",
          7304 => x"74",
          7305 => x"51",
          7306 => x"8c",
          7307 => x"9c",
          7308 => x"fb",
          7309 => x"b2",
          7310 => x"15",
          7311 => x"3f",
          7312 => x"15",
          7313 => x"3f",
          7314 => x"0b",
          7315 => x"78",
          7316 => x"3f",
          7317 => x"08",
          7318 => x"81",
          7319 => x"57",
          7320 => x"34",
          7321 => x"c8",
          7322 => x"0d",
          7323 => x"0d",
          7324 => x"54",
          7325 => x"82",
          7326 => x"53",
          7327 => x"08",
          7328 => x"3d",
          7329 => x"73",
          7330 => x"3f",
          7331 => x"08",
          7332 => x"c8",
          7333 => x"82",
          7334 => x"74",
          7335 => x"b5",
          7336 => x"3d",
          7337 => x"3d",
          7338 => x"51",
          7339 => x"8b",
          7340 => x"82",
          7341 => x"24",
          7342 => x"b5",
          7343 => x"cd",
          7344 => x"52",
          7345 => x"c8",
          7346 => x"0d",
          7347 => x"0d",
          7348 => x"3d",
          7349 => x"94",
          7350 => x"c1",
          7351 => x"c8",
          7352 => x"b5",
          7353 => x"e0",
          7354 => x"63",
          7355 => x"d4",
          7356 => x"8d",
          7357 => x"c8",
          7358 => x"b5",
          7359 => x"38",
          7360 => x"05",
          7361 => x"2b",
          7362 => x"80",
          7363 => x"76",
          7364 => x"0c",
          7365 => x"02",
          7366 => x"70",
          7367 => x"81",
          7368 => x"56",
          7369 => x"9e",
          7370 => x"53",
          7371 => x"db",
          7372 => x"b5",
          7373 => x"15",
          7374 => x"82",
          7375 => x"84",
          7376 => x"06",
          7377 => x"55",
          7378 => x"c8",
          7379 => x"0d",
          7380 => x"0d",
          7381 => x"5b",
          7382 => x"80",
          7383 => x"ff",
          7384 => x"9f",
          7385 => x"b5",
          7386 => x"c8",
          7387 => x"b5",
          7388 => x"fc",
          7389 => x"7a",
          7390 => x"08",
          7391 => x"64",
          7392 => x"2e",
          7393 => x"a0",
          7394 => x"70",
          7395 => x"ea",
          7396 => x"c8",
          7397 => x"b5",
          7398 => x"d4",
          7399 => x"7b",
          7400 => x"3f",
          7401 => x"08",
          7402 => x"c8",
          7403 => x"38",
          7404 => x"51",
          7405 => x"82",
          7406 => x"45",
          7407 => x"51",
          7408 => x"82",
          7409 => x"57",
          7410 => x"08",
          7411 => x"80",
          7412 => x"da",
          7413 => x"b5",
          7414 => x"82",
          7415 => x"a4",
          7416 => x"7b",
          7417 => x"3f",
          7418 => x"c8",
          7419 => x"38",
          7420 => x"51",
          7421 => x"82",
          7422 => x"57",
          7423 => x"08",
          7424 => x"38",
          7425 => x"09",
          7426 => x"38",
          7427 => x"e0",
          7428 => x"dc",
          7429 => x"ff",
          7430 => x"74",
          7431 => x"3f",
          7432 => x"78",
          7433 => x"33",
          7434 => x"56",
          7435 => x"91",
          7436 => x"05",
          7437 => x"81",
          7438 => x"56",
          7439 => x"f5",
          7440 => x"54",
          7441 => x"81",
          7442 => x"80",
          7443 => x"78",
          7444 => x"55",
          7445 => x"11",
          7446 => x"18",
          7447 => x"58",
          7448 => x"34",
          7449 => x"ff",
          7450 => x"55",
          7451 => x"34",
          7452 => x"77",
          7453 => x"81",
          7454 => x"ff",
          7455 => x"55",
          7456 => x"34",
          7457 => x"cd",
          7458 => x"84",
          7459 => x"80",
          7460 => x"70",
          7461 => x"56",
          7462 => x"76",
          7463 => x"81",
          7464 => x"70",
          7465 => x"56",
          7466 => x"82",
          7467 => x"78",
          7468 => x"80",
          7469 => x"27",
          7470 => x"19",
          7471 => x"7a",
          7472 => x"5c",
          7473 => x"55",
          7474 => x"7a",
          7475 => x"5c",
          7476 => x"2e",
          7477 => x"85",
          7478 => x"94",
          7479 => x"81",
          7480 => x"73",
          7481 => x"81",
          7482 => x"7a",
          7483 => x"38",
          7484 => x"76",
          7485 => x"0c",
          7486 => x"04",
          7487 => x"7b",
          7488 => x"fc",
          7489 => x"53",
          7490 => x"bb",
          7491 => x"c8",
          7492 => x"b5",
          7493 => x"fa",
          7494 => x"33",
          7495 => x"f2",
          7496 => x"08",
          7497 => x"27",
          7498 => x"15",
          7499 => x"2a",
          7500 => x"51",
          7501 => x"83",
          7502 => x"94",
          7503 => x"80",
          7504 => x"0c",
          7505 => x"2e",
          7506 => x"79",
          7507 => x"70",
          7508 => x"51",
          7509 => x"2e",
          7510 => x"52",
          7511 => x"fe",
          7512 => x"82",
          7513 => x"ff",
          7514 => x"70",
          7515 => x"fe",
          7516 => x"82",
          7517 => x"73",
          7518 => x"76",
          7519 => x"06",
          7520 => x"0c",
          7521 => x"98",
          7522 => x"58",
          7523 => x"39",
          7524 => x"54",
          7525 => x"73",
          7526 => x"cd",
          7527 => x"b5",
          7528 => x"82",
          7529 => x"81",
          7530 => x"38",
          7531 => x"08",
          7532 => x"9b",
          7533 => x"c8",
          7534 => x"0c",
          7535 => x"0c",
          7536 => x"81",
          7537 => x"76",
          7538 => x"38",
          7539 => x"94",
          7540 => x"94",
          7541 => x"16",
          7542 => x"2a",
          7543 => x"51",
          7544 => x"72",
          7545 => x"38",
          7546 => x"51",
          7547 => x"82",
          7548 => x"54",
          7549 => x"08",
          7550 => x"b5",
          7551 => x"a7",
          7552 => x"74",
          7553 => x"3f",
          7554 => x"08",
          7555 => x"2e",
          7556 => x"74",
          7557 => x"79",
          7558 => x"14",
          7559 => x"38",
          7560 => x"0c",
          7561 => x"94",
          7562 => x"94",
          7563 => x"83",
          7564 => x"72",
          7565 => x"38",
          7566 => x"51",
          7567 => x"82",
          7568 => x"94",
          7569 => x"91",
          7570 => x"53",
          7571 => x"81",
          7572 => x"34",
          7573 => x"39",
          7574 => x"82",
          7575 => x"05",
          7576 => x"08",
          7577 => x"08",
          7578 => x"38",
          7579 => x"0c",
          7580 => x"80",
          7581 => x"72",
          7582 => x"73",
          7583 => x"53",
          7584 => x"8c",
          7585 => x"16",
          7586 => x"38",
          7587 => x"0c",
          7588 => x"82",
          7589 => x"8b",
          7590 => x"f9",
          7591 => x"56",
          7592 => x"80",
          7593 => x"38",
          7594 => x"3d",
          7595 => x"8a",
          7596 => x"51",
          7597 => x"82",
          7598 => x"55",
          7599 => x"08",
          7600 => x"77",
          7601 => x"52",
          7602 => x"b5",
          7603 => x"c8",
          7604 => x"b5",
          7605 => x"c3",
          7606 => x"33",
          7607 => x"55",
          7608 => x"24",
          7609 => x"16",
          7610 => x"2a",
          7611 => x"51",
          7612 => x"80",
          7613 => x"9c",
          7614 => x"77",
          7615 => x"3f",
          7616 => x"08",
          7617 => x"77",
          7618 => x"22",
          7619 => x"74",
          7620 => x"ce",
          7621 => x"b5",
          7622 => x"74",
          7623 => x"81",
          7624 => x"85",
          7625 => x"74",
          7626 => x"38",
          7627 => x"74",
          7628 => x"b5",
          7629 => x"3d",
          7630 => x"3d",
          7631 => x"3d",
          7632 => x"70",
          7633 => x"ff",
          7634 => x"c8",
          7635 => x"82",
          7636 => x"73",
          7637 => x"0d",
          7638 => x"0d",
          7639 => x"3d",
          7640 => x"71",
          7641 => x"e7",
          7642 => x"b5",
          7643 => x"82",
          7644 => x"80",
          7645 => x"93",
          7646 => x"c8",
          7647 => x"51",
          7648 => x"82",
          7649 => x"53",
          7650 => x"82",
          7651 => x"52",
          7652 => x"ac",
          7653 => x"c8",
          7654 => x"b5",
          7655 => x"2e",
          7656 => x"85",
          7657 => x"87",
          7658 => x"c8",
          7659 => x"74",
          7660 => x"d5",
          7661 => x"52",
          7662 => x"89",
          7663 => x"c8",
          7664 => x"70",
          7665 => x"07",
          7666 => x"82",
          7667 => x"06",
          7668 => x"54",
          7669 => x"c8",
          7670 => x"0d",
          7671 => x"0d",
          7672 => x"53",
          7673 => x"53",
          7674 => x"56",
          7675 => x"82",
          7676 => x"55",
          7677 => x"08",
          7678 => x"52",
          7679 => x"81",
          7680 => x"c8",
          7681 => x"b5",
          7682 => x"38",
          7683 => x"05",
          7684 => x"2b",
          7685 => x"80",
          7686 => x"86",
          7687 => x"76",
          7688 => x"38",
          7689 => x"51",
          7690 => x"74",
          7691 => x"0c",
          7692 => x"04",
          7693 => x"63",
          7694 => x"80",
          7695 => x"ec",
          7696 => x"3d",
          7697 => x"3f",
          7698 => x"08",
          7699 => x"c8",
          7700 => x"38",
          7701 => x"73",
          7702 => x"08",
          7703 => x"13",
          7704 => x"58",
          7705 => x"26",
          7706 => x"7c",
          7707 => x"39",
          7708 => x"cc",
          7709 => x"81",
          7710 => x"b5",
          7711 => x"33",
          7712 => x"81",
          7713 => x"06",
          7714 => x"75",
          7715 => x"52",
          7716 => x"05",
          7717 => x"3f",
          7718 => x"08",
          7719 => x"38",
          7720 => x"08",
          7721 => x"38",
          7722 => x"08",
          7723 => x"b5",
          7724 => x"80",
          7725 => x"81",
          7726 => x"59",
          7727 => x"14",
          7728 => x"ca",
          7729 => x"39",
          7730 => x"82",
          7731 => x"57",
          7732 => x"38",
          7733 => x"18",
          7734 => x"ff",
          7735 => x"82",
          7736 => x"5b",
          7737 => x"08",
          7738 => x"7c",
          7739 => x"12",
          7740 => x"52",
          7741 => x"82",
          7742 => x"06",
          7743 => x"14",
          7744 => x"cb",
          7745 => x"c8",
          7746 => x"ff",
          7747 => x"70",
          7748 => x"82",
          7749 => x"51",
          7750 => x"b4",
          7751 => x"bb",
          7752 => x"b5",
          7753 => x"0a",
          7754 => x"70",
          7755 => x"84",
          7756 => x"51",
          7757 => x"ff",
          7758 => x"56",
          7759 => x"38",
          7760 => x"7c",
          7761 => x"0c",
          7762 => x"81",
          7763 => x"74",
          7764 => x"7a",
          7765 => x"0c",
          7766 => x"04",
          7767 => x"79",
          7768 => x"05",
          7769 => x"57",
          7770 => x"82",
          7771 => x"56",
          7772 => x"08",
          7773 => x"91",
          7774 => x"75",
          7775 => x"90",
          7776 => x"81",
          7777 => x"06",
          7778 => x"87",
          7779 => x"2e",
          7780 => x"94",
          7781 => x"73",
          7782 => x"27",
          7783 => x"73",
          7784 => x"b5",
          7785 => x"88",
          7786 => x"76",
          7787 => x"3f",
          7788 => x"08",
          7789 => x"0c",
          7790 => x"39",
          7791 => x"52",
          7792 => x"bf",
          7793 => x"b5",
          7794 => x"2e",
          7795 => x"83",
          7796 => x"82",
          7797 => x"81",
          7798 => x"06",
          7799 => x"56",
          7800 => x"a0",
          7801 => x"82",
          7802 => x"98",
          7803 => x"94",
          7804 => x"08",
          7805 => x"c8",
          7806 => x"51",
          7807 => x"82",
          7808 => x"56",
          7809 => x"8c",
          7810 => x"17",
          7811 => x"07",
          7812 => x"18",
          7813 => x"2e",
          7814 => x"91",
          7815 => x"55",
          7816 => x"c8",
          7817 => x"0d",
          7818 => x"0d",
          7819 => x"3d",
          7820 => x"52",
          7821 => x"da",
          7822 => x"b5",
          7823 => x"82",
          7824 => x"81",
          7825 => x"45",
          7826 => x"52",
          7827 => x"52",
          7828 => x"3f",
          7829 => x"08",
          7830 => x"c8",
          7831 => x"38",
          7832 => x"05",
          7833 => x"2a",
          7834 => x"51",
          7835 => x"55",
          7836 => x"38",
          7837 => x"54",
          7838 => x"81",
          7839 => x"80",
          7840 => x"70",
          7841 => x"54",
          7842 => x"81",
          7843 => x"52",
          7844 => x"c5",
          7845 => x"c8",
          7846 => x"2a",
          7847 => x"51",
          7848 => x"80",
          7849 => x"38",
          7850 => x"b5",
          7851 => x"15",
          7852 => x"86",
          7853 => x"82",
          7854 => x"5c",
          7855 => x"3d",
          7856 => x"c7",
          7857 => x"b5",
          7858 => x"82",
          7859 => x"80",
          7860 => x"b5",
          7861 => x"73",
          7862 => x"3f",
          7863 => x"08",
          7864 => x"c8",
          7865 => x"87",
          7866 => x"39",
          7867 => x"08",
          7868 => x"38",
          7869 => x"08",
          7870 => x"77",
          7871 => x"3f",
          7872 => x"08",
          7873 => x"08",
          7874 => x"b5",
          7875 => x"80",
          7876 => x"55",
          7877 => x"94",
          7878 => x"2e",
          7879 => x"53",
          7880 => x"51",
          7881 => x"82",
          7882 => x"55",
          7883 => x"78",
          7884 => x"fe",
          7885 => x"c8",
          7886 => x"82",
          7887 => x"a0",
          7888 => x"e9",
          7889 => x"53",
          7890 => x"05",
          7891 => x"51",
          7892 => x"82",
          7893 => x"54",
          7894 => x"08",
          7895 => x"78",
          7896 => x"8e",
          7897 => x"58",
          7898 => x"82",
          7899 => x"54",
          7900 => x"08",
          7901 => x"54",
          7902 => x"82",
          7903 => x"84",
          7904 => x"06",
          7905 => x"02",
          7906 => x"33",
          7907 => x"81",
          7908 => x"86",
          7909 => x"f6",
          7910 => x"74",
          7911 => x"70",
          7912 => x"c3",
          7913 => x"c8",
          7914 => x"56",
          7915 => x"08",
          7916 => x"54",
          7917 => x"08",
          7918 => x"81",
          7919 => x"82",
          7920 => x"c8",
          7921 => x"09",
          7922 => x"38",
          7923 => x"b4",
          7924 => x"b0",
          7925 => x"c8",
          7926 => x"51",
          7927 => x"82",
          7928 => x"54",
          7929 => x"08",
          7930 => x"8b",
          7931 => x"b4",
          7932 => x"b7",
          7933 => x"54",
          7934 => x"15",
          7935 => x"90",
          7936 => x"34",
          7937 => x"0a",
          7938 => x"19",
          7939 => x"9f",
          7940 => x"78",
          7941 => x"51",
          7942 => x"a0",
          7943 => x"11",
          7944 => x"05",
          7945 => x"b6",
          7946 => x"ae",
          7947 => x"15",
          7948 => x"78",
          7949 => x"53",
          7950 => x"3f",
          7951 => x"0b",
          7952 => x"77",
          7953 => x"3f",
          7954 => x"08",
          7955 => x"c8",
          7956 => x"82",
          7957 => x"52",
          7958 => x"51",
          7959 => x"3f",
          7960 => x"52",
          7961 => x"aa",
          7962 => x"90",
          7963 => x"34",
          7964 => x"0b",
          7965 => x"78",
          7966 => x"b6",
          7967 => x"c8",
          7968 => x"39",
          7969 => x"52",
          7970 => x"be",
          7971 => x"82",
          7972 => x"99",
          7973 => x"da",
          7974 => x"3d",
          7975 => x"d2",
          7976 => x"53",
          7977 => x"84",
          7978 => x"3d",
          7979 => x"3f",
          7980 => x"08",
          7981 => x"c8",
          7982 => x"38",
          7983 => x"3d",
          7984 => x"3d",
          7985 => x"cc",
          7986 => x"b5",
          7987 => x"82",
          7988 => x"82",
          7989 => x"81",
          7990 => x"81",
          7991 => x"86",
          7992 => x"aa",
          7993 => x"a4",
          7994 => x"a8",
          7995 => x"05",
          7996 => x"ea",
          7997 => x"77",
          7998 => x"70",
          7999 => x"b4",
          8000 => x"3d",
          8001 => x"51",
          8002 => x"82",
          8003 => x"55",
          8004 => x"08",
          8005 => x"6f",
          8006 => x"06",
          8007 => x"a2",
          8008 => x"92",
          8009 => x"81",
          8010 => x"b5",
          8011 => x"2e",
          8012 => x"81",
          8013 => x"51",
          8014 => x"82",
          8015 => x"55",
          8016 => x"08",
          8017 => x"68",
          8018 => x"a8",
          8019 => x"05",
          8020 => x"51",
          8021 => x"3f",
          8022 => x"33",
          8023 => x"8b",
          8024 => x"84",
          8025 => x"06",
          8026 => x"73",
          8027 => x"a0",
          8028 => x"8b",
          8029 => x"54",
          8030 => x"15",
          8031 => x"33",
          8032 => x"70",
          8033 => x"55",
          8034 => x"2e",
          8035 => x"6e",
          8036 => x"df",
          8037 => x"78",
          8038 => x"3f",
          8039 => x"08",
          8040 => x"ff",
          8041 => x"82",
          8042 => x"c8",
          8043 => x"80",
          8044 => x"b5",
          8045 => x"78",
          8046 => x"af",
          8047 => x"c8",
          8048 => x"d4",
          8049 => x"55",
          8050 => x"08",
          8051 => x"81",
          8052 => x"73",
          8053 => x"81",
          8054 => x"63",
          8055 => x"76",
          8056 => x"3f",
          8057 => x"0b",
          8058 => x"87",
          8059 => x"c8",
          8060 => x"77",
          8061 => x"3f",
          8062 => x"08",
          8063 => x"c8",
          8064 => x"78",
          8065 => x"aa",
          8066 => x"c8",
          8067 => x"82",
          8068 => x"a8",
          8069 => x"ed",
          8070 => x"80",
          8071 => x"02",
          8072 => x"df",
          8073 => x"57",
          8074 => x"3d",
          8075 => x"96",
          8076 => x"e9",
          8077 => x"c8",
          8078 => x"b5",
          8079 => x"cf",
          8080 => x"65",
          8081 => x"d4",
          8082 => x"b5",
          8083 => x"c8",
          8084 => x"b5",
          8085 => x"38",
          8086 => x"05",
          8087 => x"06",
          8088 => x"73",
          8089 => x"a7",
          8090 => x"09",
          8091 => x"71",
          8092 => x"06",
          8093 => x"55",
          8094 => x"15",
          8095 => x"81",
          8096 => x"34",
          8097 => x"b4",
          8098 => x"b5",
          8099 => x"74",
          8100 => x"0c",
          8101 => x"04",
          8102 => x"64",
          8103 => x"93",
          8104 => x"52",
          8105 => x"d1",
          8106 => x"b5",
          8107 => x"82",
          8108 => x"80",
          8109 => x"58",
          8110 => x"3d",
          8111 => x"c8",
          8112 => x"b5",
          8113 => x"82",
          8114 => x"b4",
          8115 => x"c7",
          8116 => x"a0",
          8117 => x"55",
          8118 => x"84",
          8119 => x"17",
          8120 => x"2b",
          8121 => x"96",
          8122 => x"b0",
          8123 => x"54",
          8124 => x"15",
          8125 => x"ff",
          8126 => x"82",
          8127 => x"55",
          8128 => x"c8",
          8129 => x"0d",
          8130 => x"0d",
          8131 => x"5a",
          8132 => x"3d",
          8133 => x"99",
          8134 => x"81",
          8135 => x"c8",
          8136 => x"c8",
          8137 => x"82",
          8138 => x"07",
          8139 => x"55",
          8140 => x"2e",
          8141 => x"81",
          8142 => x"55",
          8143 => x"2e",
          8144 => x"7b",
          8145 => x"80",
          8146 => x"70",
          8147 => x"be",
          8148 => x"b5",
          8149 => x"82",
          8150 => x"80",
          8151 => x"52",
          8152 => x"dc",
          8153 => x"c8",
          8154 => x"b5",
          8155 => x"38",
          8156 => x"08",
          8157 => x"08",
          8158 => x"56",
          8159 => x"19",
          8160 => x"59",
          8161 => x"74",
          8162 => x"56",
          8163 => x"ec",
          8164 => x"75",
          8165 => x"74",
          8166 => x"2e",
          8167 => x"16",
          8168 => x"33",
          8169 => x"73",
          8170 => x"38",
          8171 => x"84",
          8172 => x"06",
          8173 => x"7a",
          8174 => x"76",
          8175 => x"07",
          8176 => x"54",
          8177 => x"80",
          8178 => x"80",
          8179 => x"7b",
          8180 => x"53",
          8181 => x"93",
          8182 => x"c8",
          8183 => x"b5",
          8184 => x"38",
          8185 => x"55",
          8186 => x"56",
          8187 => x"8b",
          8188 => x"56",
          8189 => x"83",
          8190 => x"75",
          8191 => x"51",
          8192 => x"3f",
          8193 => x"08",
          8194 => x"82",
          8195 => x"98",
          8196 => x"e6",
          8197 => x"53",
          8198 => x"b8",
          8199 => x"3d",
          8200 => x"3f",
          8201 => x"08",
          8202 => x"08",
          8203 => x"b5",
          8204 => x"98",
          8205 => x"a0",
          8206 => x"70",
          8207 => x"ae",
          8208 => x"6d",
          8209 => x"81",
          8210 => x"57",
          8211 => x"74",
          8212 => x"38",
          8213 => x"81",
          8214 => x"81",
          8215 => x"52",
          8216 => x"89",
          8217 => x"c8",
          8218 => x"a5",
          8219 => x"33",
          8220 => x"54",
          8221 => x"3f",
          8222 => x"08",
          8223 => x"38",
          8224 => x"76",
          8225 => x"05",
          8226 => x"39",
          8227 => x"08",
          8228 => x"15",
          8229 => x"ff",
          8230 => x"73",
          8231 => x"38",
          8232 => x"83",
          8233 => x"56",
          8234 => x"75",
          8235 => x"82",
          8236 => x"33",
          8237 => x"2e",
          8238 => x"52",
          8239 => x"51",
          8240 => x"3f",
          8241 => x"08",
          8242 => x"ff",
          8243 => x"38",
          8244 => x"88",
          8245 => x"8a",
          8246 => x"38",
          8247 => x"ec",
          8248 => x"75",
          8249 => x"74",
          8250 => x"73",
          8251 => x"05",
          8252 => x"17",
          8253 => x"70",
          8254 => x"34",
          8255 => x"70",
          8256 => x"ff",
          8257 => x"55",
          8258 => x"26",
          8259 => x"8b",
          8260 => x"86",
          8261 => x"e5",
          8262 => x"38",
          8263 => x"99",
          8264 => x"05",
          8265 => x"70",
          8266 => x"73",
          8267 => x"81",
          8268 => x"ff",
          8269 => x"ed",
          8270 => x"80",
          8271 => x"91",
          8272 => x"55",
          8273 => x"3f",
          8274 => x"08",
          8275 => x"c8",
          8276 => x"38",
          8277 => x"51",
          8278 => x"3f",
          8279 => x"08",
          8280 => x"c8",
          8281 => x"76",
          8282 => x"67",
          8283 => x"34",
          8284 => x"82",
          8285 => x"84",
          8286 => x"06",
          8287 => x"80",
          8288 => x"2e",
          8289 => x"81",
          8290 => x"ff",
          8291 => x"82",
          8292 => x"54",
          8293 => x"08",
          8294 => x"53",
          8295 => x"08",
          8296 => x"ff",
          8297 => x"67",
          8298 => x"8b",
          8299 => x"53",
          8300 => x"51",
          8301 => x"3f",
          8302 => x"0b",
          8303 => x"79",
          8304 => x"ee",
          8305 => x"c8",
          8306 => x"55",
          8307 => x"c8",
          8308 => x"0d",
          8309 => x"0d",
          8310 => x"88",
          8311 => x"05",
          8312 => x"fc",
          8313 => x"54",
          8314 => x"d2",
          8315 => x"b5",
          8316 => x"82",
          8317 => x"82",
          8318 => x"1a",
          8319 => x"82",
          8320 => x"80",
          8321 => x"8c",
          8322 => x"78",
          8323 => x"1a",
          8324 => x"2a",
          8325 => x"51",
          8326 => x"90",
          8327 => x"82",
          8328 => x"58",
          8329 => x"81",
          8330 => x"39",
          8331 => x"22",
          8332 => x"70",
          8333 => x"56",
          8334 => x"c2",
          8335 => x"14",
          8336 => x"30",
          8337 => x"9f",
          8338 => x"c8",
          8339 => x"19",
          8340 => x"5a",
          8341 => x"81",
          8342 => x"38",
          8343 => x"77",
          8344 => x"82",
          8345 => x"56",
          8346 => x"74",
          8347 => x"ff",
          8348 => x"81",
          8349 => x"55",
          8350 => x"75",
          8351 => x"82",
          8352 => x"c8",
          8353 => x"ff",
          8354 => x"b5",
          8355 => x"2e",
          8356 => x"82",
          8357 => x"8e",
          8358 => x"56",
          8359 => x"09",
          8360 => x"38",
          8361 => x"59",
          8362 => x"77",
          8363 => x"06",
          8364 => x"87",
          8365 => x"39",
          8366 => x"ba",
          8367 => x"55",
          8368 => x"2e",
          8369 => x"15",
          8370 => x"2e",
          8371 => x"83",
          8372 => x"75",
          8373 => x"7e",
          8374 => x"a8",
          8375 => x"c8",
          8376 => x"b5",
          8377 => x"ce",
          8378 => x"16",
          8379 => x"56",
          8380 => x"38",
          8381 => x"19",
          8382 => x"8c",
          8383 => x"7d",
          8384 => x"38",
          8385 => x"0c",
          8386 => x"0c",
          8387 => x"80",
          8388 => x"73",
          8389 => x"98",
          8390 => x"05",
          8391 => x"57",
          8392 => x"26",
          8393 => x"7b",
          8394 => x"0c",
          8395 => x"81",
          8396 => x"84",
          8397 => x"54",
          8398 => x"c8",
          8399 => x"0d",
          8400 => x"0d",
          8401 => x"88",
          8402 => x"05",
          8403 => x"54",
          8404 => x"c5",
          8405 => x"56",
          8406 => x"b5",
          8407 => x"8b",
          8408 => x"b5",
          8409 => x"29",
          8410 => x"05",
          8411 => x"55",
          8412 => x"84",
          8413 => x"34",
          8414 => x"08",
          8415 => x"5f",
          8416 => x"51",
          8417 => x"3f",
          8418 => x"08",
          8419 => x"70",
          8420 => x"57",
          8421 => x"8b",
          8422 => x"82",
          8423 => x"06",
          8424 => x"56",
          8425 => x"38",
          8426 => x"05",
          8427 => x"7e",
          8428 => x"f0",
          8429 => x"c8",
          8430 => x"67",
          8431 => x"2e",
          8432 => x"82",
          8433 => x"8b",
          8434 => x"75",
          8435 => x"80",
          8436 => x"81",
          8437 => x"2e",
          8438 => x"80",
          8439 => x"38",
          8440 => x"0a",
          8441 => x"ff",
          8442 => x"55",
          8443 => x"86",
          8444 => x"8a",
          8445 => x"89",
          8446 => x"2a",
          8447 => x"77",
          8448 => x"59",
          8449 => x"81",
          8450 => x"70",
          8451 => x"07",
          8452 => x"56",
          8453 => x"38",
          8454 => x"05",
          8455 => x"7e",
          8456 => x"80",
          8457 => x"82",
          8458 => x"8a",
          8459 => x"83",
          8460 => x"06",
          8461 => x"08",
          8462 => x"74",
          8463 => x"41",
          8464 => x"56",
          8465 => x"8a",
          8466 => x"61",
          8467 => x"55",
          8468 => x"27",
          8469 => x"93",
          8470 => x"80",
          8471 => x"38",
          8472 => x"70",
          8473 => x"43",
          8474 => x"95",
          8475 => x"06",
          8476 => x"2e",
          8477 => x"77",
          8478 => x"74",
          8479 => x"83",
          8480 => x"06",
          8481 => x"82",
          8482 => x"2e",
          8483 => x"78",
          8484 => x"2e",
          8485 => x"80",
          8486 => x"ae",
          8487 => x"2a",
          8488 => x"82",
          8489 => x"56",
          8490 => x"2e",
          8491 => x"77",
          8492 => x"82",
          8493 => x"79",
          8494 => x"70",
          8495 => x"5a",
          8496 => x"86",
          8497 => x"27",
          8498 => x"52",
          8499 => x"bd",
          8500 => x"b5",
          8501 => x"29",
          8502 => x"70",
          8503 => x"55",
          8504 => x"0b",
          8505 => x"08",
          8506 => x"05",
          8507 => x"ff",
          8508 => x"27",
          8509 => x"88",
          8510 => x"ae",
          8511 => x"2a",
          8512 => x"82",
          8513 => x"56",
          8514 => x"2e",
          8515 => x"77",
          8516 => x"82",
          8517 => x"79",
          8518 => x"70",
          8519 => x"5a",
          8520 => x"86",
          8521 => x"27",
          8522 => x"52",
          8523 => x"bc",
          8524 => x"b5",
          8525 => x"84",
          8526 => x"b5",
          8527 => x"f5",
          8528 => x"81",
          8529 => x"c8",
          8530 => x"b5",
          8531 => x"71",
          8532 => x"83",
          8533 => x"5e",
          8534 => x"89",
          8535 => x"5c",
          8536 => x"1c",
          8537 => x"05",
          8538 => x"ff",
          8539 => x"70",
          8540 => x"31",
          8541 => x"57",
          8542 => x"83",
          8543 => x"06",
          8544 => x"1c",
          8545 => x"5c",
          8546 => x"1d",
          8547 => x"29",
          8548 => x"31",
          8549 => x"55",
          8550 => x"87",
          8551 => x"7c",
          8552 => x"7a",
          8553 => x"31",
          8554 => x"bb",
          8555 => x"b5",
          8556 => x"7d",
          8557 => x"81",
          8558 => x"82",
          8559 => x"83",
          8560 => x"80",
          8561 => x"87",
          8562 => x"81",
          8563 => x"fd",
          8564 => x"f8",
          8565 => x"2e",
          8566 => x"80",
          8567 => x"ff",
          8568 => x"b5",
          8569 => x"a0",
          8570 => x"38",
          8571 => x"74",
          8572 => x"86",
          8573 => x"fd",
          8574 => x"81",
          8575 => x"80",
          8576 => x"83",
          8577 => x"39",
          8578 => x"08",
          8579 => x"92",
          8580 => x"b8",
          8581 => x"59",
          8582 => x"27",
          8583 => x"86",
          8584 => x"55",
          8585 => x"09",
          8586 => x"38",
          8587 => x"f5",
          8588 => x"38",
          8589 => x"55",
          8590 => x"86",
          8591 => x"80",
          8592 => x"7a",
          8593 => x"b9",
          8594 => x"82",
          8595 => x"7a",
          8596 => x"8a",
          8597 => x"52",
          8598 => x"ff",
          8599 => x"79",
          8600 => x"7b",
          8601 => x"06",
          8602 => x"51",
          8603 => x"3f",
          8604 => x"1c",
          8605 => x"32",
          8606 => x"96",
          8607 => x"06",
          8608 => x"91",
          8609 => x"a1",
          8610 => x"55",
          8611 => x"ff",
          8612 => x"74",
          8613 => x"06",
          8614 => x"51",
          8615 => x"3f",
          8616 => x"52",
          8617 => x"ff",
          8618 => x"f8",
          8619 => x"34",
          8620 => x"1b",
          8621 => x"d9",
          8622 => x"52",
          8623 => x"ff",
          8624 => x"60",
          8625 => x"51",
          8626 => x"3f",
          8627 => x"09",
          8628 => x"cb",
          8629 => x"b2",
          8630 => x"c3",
          8631 => x"a0",
          8632 => x"52",
          8633 => x"ff",
          8634 => x"82",
          8635 => x"51",
          8636 => x"3f",
          8637 => x"1b",
          8638 => x"95",
          8639 => x"b2",
          8640 => x"a0",
          8641 => x"80",
          8642 => x"1c",
          8643 => x"80",
          8644 => x"93",
          8645 => x"d8",
          8646 => x"1b",
          8647 => x"82",
          8648 => x"52",
          8649 => x"ff",
          8650 => x"7c",
          8651 => x"06",
          8652 => x"51",
          8653 => x"3f",
          8654 => x"a4",
          8655 => x"0b",
          8656 => x"93",
          8657 => x"ec",
          8658 => x"51",
          8659 => x"3f",
          8660 => x"52",
          8661 => x"70",
          8662 => x"9f",
          8663 => x"54",
          8664 => x"52",
          8665 => x"9b",
          8666 => x"56",
          8667 => x"08",
          8668 => x"7d",
          8669 => x"81",
          8670 => x"38",
          8671 => x"86",
          8672 => x"52",
          8673 => x"9b",
          8674 => x"80",
          8675 => x"7a",
          8676 => x"ed",
          8677 => x"85",
          8678 => x"7a",
          8679 => x"8f",
          8680 => x"85",
          8681 => x"83",
          8682 => x"ff",
          8683 => x"ff",
          8684 => x"e8",
          8685 => x"9e",
          8686 => x"52",
          8687 => x"51",
          8688 => x"3f",
          8689 => x"52",
          8690 => x"9e",
          8691 => x"54",
          8692 => x"53",
          8693 => x"51",
          8694 => x"3f",
          8695 => x"16",
          8696 => x"7e",
          8697 => x"d8",
          8698 => x"80",
          8699 => x"ff",
          8700 => x"7f",
          8701 => x"7d",
          8702 => x"81",
          8703 => x"f8",
          8704 => x"ff",
          8705 => x"ff",
          8706 => x"51",
          8707 => x"3f",
          8708 => x"88",
          8709 => x"39",
          8710 => x"f8",
          8711 => x"2e",
          8712 => x"55",
          8713 => x"51",
          8714 => x"3f",
          8715 => x"57",
          8716 => x"83",
          8717 => x"76",
          8718 => x"7a",
          8719 => x"ff",
          8720 => x"82",
          8721 => x"82",
          8722 => x"80",
          8723 => x"c8",
          8724 => x"51",
          8725 => x"3f",
          8726 => x"78",
          8727 => x"74",
          8728 => x"18",
          8729 => x"2e",
          8730 => x"79",
          8731 => x"2e",
          8732 => x"55",
          8733 => x"62",
          8734 => x"74",
          8735 => x"75",
          8736 => x"7e",
          8737 => x"b8",
          8738 => x"c8",
          8739 => x"38",
          8740 => x"78",
          8741 => x"74",
          8742 => x"56",
          8743 => x"93",
          8744 => x"66",
          8745 => x"26",
          8746 => x"56",
          8747 => x"83",
          8748 => x"64",
          8749 => x"77",
          8750 => x"84",
          8751 => x"52",
          8752 => x"9d",
          8753 => x"d4",
          8754 => x"51",
          8755 => x"3f",
          8756 => x"55",
          8757 => x"81",
          8758 => x"34",
          8759 => x"16",
          8760 => x"16",
          8761 => x"16",
          8762 => x"05",
          8763 => x"c1",
          8764 => x"fe",
          8765 => x"fe",
          8766 => x"34",
          8767 => x"08",
          8768 => x"07",
          8769 => x"16",
          8770 => x"c8",
          8771 => x"34",
          8772 => x"c6",
          8773 => x"9c",
          8774 => x"52",
          8775 => x"51",
          8776 => x"3f",
          8777 => x"53",
          8778 => x"51",
          8779 => x"3f",
          8780 => x"b5",
          8781 => x"38",
          8782 => x"52",
          8783 => x"99",
          8784 => x"56",
          8785 => x"08",
          8786 => x"39",
          8787 => x"39",
          8788 => x"39",
          8789 => x"08",
          8790 => x"b5",
          8791 => x"3d",
          8792 => x"3d",
          8793 => x"5b",
          8794 => x"60",
          8795 => x"57",
          8796 => x"25",
          8797 => x"3d",
          8798 => x"55",
          8799 => x"15",
          8800 => x"c9",
          8801 => x"81",
          8802 => x"06",
          8803 => x"3d",
          8804 => x"8d",
          8805 => x"74",
          8806 => x"05",
          8807 => x"17",
          8808 => x"2e",
          8809 => x"c9",
          8810 => x"34",
          8811 => x"83",
          8812 => x"74",
          8813 => x"0c",
          8814 => x"04",
          8815 => x"7b",
          8816 => x"b3",
          8817 => x"57",
          8818 => x"09",
          8819 => x"38",
          8820 => x"51",
          8821 => x"17",
          8822 => x"76",
          8823 => x"88",
          8824 => x"17",
          8825 => x"59",
          8826 => x"81",
          8827 => x"76",
          8828 => x"8b",
          8829 => x"54",
          8830 => x"17",
          8831 => x"51",
          8832 => x"79",
          8833 => x"30",
          8834 => x"9f",
          8835 => x"53",
          8836 => x"75",
          8837 => x"81",
          8838 => x"0c",
          8839 => x"04",
          8840 => x"79",
          8841 => x"56",
          8842 => x"24",
          8843 => x"3d",
          8844 => x"74",
          8845 => x"52",
          8846 => x"cb",
          8847 => x"b5",
          8848 => x"38",
          8849 => x"78",
          8850 => x"06",
          8851 => x"16",
          8852 => x"39",
          8853 => x"82",
          8854 => x"89",
          8855 => x"fd",
          8856 => x"54",
          8857 => x"80",
          8858 => x"ff",
          8859 => x"76",
          8860 => x"3d",
          8861 => x"3d",
          8862 => x"e3",
          8863 => x"53",
          8864 => x"53",
          8865 => x"3f",
          8866 => x"51",
          8867 => x"72",
          8868 => x"3f",
          8869 => x"04",
          8870 => x"ff",
          8871 => x"ff",
          8872 => x"ff",
          8873 => x"00",
          8874 => x"aa",
          8875 => x"2e",
          8876 => x"35",
          8877 => x"3c",
          8878 => x"43",
          8879 => x"4a",
          8880 => x"51",
          8881 => x"58",
          8882 => x"5f",
          8883 => x"66",
          8884 => x"6d",
          8885 => x"74",
          8886 => x"7a",
          8887 => x"80",
          8888 => x"86",
          8889 => x"8c",
          8890 => x"92",
          8891 => x"98",
          8892 => x"9e",
          8893 => x"a4",
          8894 => x"4f",
          8895 => x"55",
          8896 => x"5b",
          8897 => x"61",
          8898 => x"67",
          8899 => x"45",
          8900 => x"45",
          8901 => x"56",
          8902 => x"ae",
          8903 => x"2d",
          8904 => x"1a",
          8905 => x"1e",
          8906 => x"7f",
          8907 => x"61",
          8908 => x"f7",
          8909 => x"7d",
          8910 => x"00",
          8911 => x"1a",
          8912 => x"56",
          8913 => x"7f",
          8914 => x"1e",
          8915 => x"1a",
          8916 => x"1a",
          8917 => x"7d",
          8918 => x"f7",
          8919 => x"7f",
          8920 => x"ae",
          8921 => x"31",
          8922 => x"1a",
          8923 => x"1a",
          8924 => x"60",
          8925 => x"1a",
          8926 => x"1a",
          8927 => x"1a",
          8928 => x"1a",
          8929 => x"1a",
          8930 => x"1a",
          8931 => x"1a",
          8932 => x"1d",
          8933 => x"1a",
          8934 => x"48",
          8935 => x"78",
          8936 => x"1a",
          8937 => x"1a",
          8938 => x"1a",
          8939 => x"1a",
          8940 => x"1a",
          8941 => x"1a",
          8942 => x"1a",
          8943 => x"1a",
          8944 => x"1a",
          8945 => x"1a",
          8946 => x"1a",
          8947 => x"1a",
          8948 => x"1a",
          8949 => x"1a",
          8950 => x"1a",
          8951 => x"1a",
          8952 => x"1a",
          8953 => x"1a",
          8954 => x"1a",
          8955 => x"1a",
          8956 => x"1a",
          8957 => x"1a",
          8958 => x"1a",
          8959 => x"1a",
          8960 => x"1a",
          8961 => x"1a",
          8962 => x"1a",
          8963 => x"1a",
          8964 => x"1a",
          8965 => x"1a",
          8966 => x"1a",
          8967 => x"1a",
          8968 => x"1a",
          8969 => x"1a",
          8970 => x"1a",
          8971 => x"1a",
          8972 => x"a8",
          8973 => x"1a",
          8974 => x"1a",
          8975 => x"1a",
          8976 => x"1a",
          8977 => x"16",
          8978 => x"1a",
          8979 => x"1a",
          8980 => x"1a",
          8981 => x"1a",
          8982 => x"1a",
          8983 => x"1a",
          8984 => x"1a",
          8985 => x"1a",
          8986 => x"1a",
          8987 => x"1a",
          8988 => x"d8",
          8989 => x"3f",
          8990 => x"af",
          8991 => x"af",
          8992 => x"af",
          8993 => x"1a",
          8994 => x"3f",
          8995 => x"1a",
          8996 => x"1a",
          8997 => x"98",
          8998 => x"1a",
          8999 => x"1a",
          9000 => x"ec",
          9001 => x"f7",
          9002 => x"1a",
          9003 => x"1a",
          9004 => x"11",
          9005 => x"1a",
          9006 => x"1f",
          9007 => x"1a",
          9008 => x"1a",
          9009 => x"16",
          9010 => x"69",
          9011 => x"00",
          9012 => x"63",
          9013 => x"00",
          9014 => x"69",
          9015 => x"00",
          9016 => x"61",
          9017 => x"00",
          9018 => x"65",
          9019 => x"00",
          9020 => x"65",
          9021 => x"00",
          9022 => x"70",
          9023 => x"00",
          9024 => x"66",
          9025 => x"00",
          9026 => x"6d",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"6c",
          9036 => x"00",
          9037 => x"00",
          9038 => x"74",
          9039 => x"00",
          9040 => x"65",
          9041 => x"00",
          9042 => x"6f",
          9043 => x"00",
          9044 => x"74",
          9045 => x"00",
          9046 => x"73",
          9047 => x"00",
          9048 => x"73",
          9049 => x"00",
          9050 => x"6f",
          9051 => x"00",
          9052 => x"00",
          9053 => x"6b",
          9054 => x"72",
          9055 => x"00",
          9056 => x"65",
          9057 => x"6c",
          9058 => x"72",
          9059 => x"00",
          9060 => x"6b",
          9061 => x"74",
          9062 => x"61",
          9063 => x"00",
          9064 => x"66",
          9065 => x"20",
          9066 => x"6e",
          9067 => x"00",
          9068 => x"70",
          9069 => x"20",
          9070 => x"6e",
          9071 => x"00",
          9072 => x"61",
          9073 => x"20",
          9074 => x"65",
          9075 => x"65",
          9076 => x"00",
          9077 => x"65",
          9078 => x"64",
          9079 => x"65",
          9080 => x"00",
          9081 => x"65",
          9082 => x"72",
          9083 => x"79",
          9084 => x"69",
          9085 => x"2e",
          9086 => x"00",
          9087 => x"65",
          9088 => x"6e",
          9089 => x"20",
          9090 => x"61",
          9091 => x"2e",
          9092 => x"00",
          9093 => x"69",
          9094 => x"72",
          9095 => x"20",
          9096 => x"74",
          9097 => x"65",
          9098 => x"00",
          9099 => x"76",
          9100 => x"75",
          9101 => x"72",
          9102 => x"20",
          9103 => x"61",
          9104 => x"2e",
          9105 => x"00",
          9106 => x"6b",
          9107 => x"74",
          9108 => x"61",
          9109 => x"64",
          9110 => x"00",
          9111 => x"63",
          9112 => x"61",
          9113 => x"6c",
          9114 => x"69",
          9115 => x"79",
          9116 => x"6d",
          9117 => x"75",
          9118 => x"6f",
          9119 => x"69",
          9120 => x"00",
          9121 => x"6d",
          9122 => x"61",
          9123 => x"74",
          9124 => x"00",
          9125 => x"65",
          9126 => x"2c",
          9127 => x"65",
          9128 => x"69",
          9129 => x"63",
          9130 => x"65",
          9131 => x"64",
          9132 => x"00",
          9133 => x"65",
          9134 => x"20",
          9135 => x"6b",
          9136 => x"00",
          9137 => x"75",
          9138 => x"63",
          9139 => x"74",
          9140 => x"6d",
          9141 => x"2e",
          9142 => x"00",
          9143 => x"20",
          9144 => x"79",
          9145 => x"65",
          9146 => x"69",
          9147 => x"2e",
          9148 => x"00",
          9149 => x"61",
          9150 => x"65",
          9151 => x"69",
          9152 => x"72",
          9153 => x"74",
          9154 => x"00",
          9155 => x"63",
          9156 => x"2e",
          9157 => x"00",
          9158 => x"6e",
          9159 => x"20",
          9160 => x"6f",
          9161 => x"00",
          9162 => x"75",
          9163 => x"74",
          9164 => x"25",
          9165 => x"74",
          9166 => x"75",
          9167 => x"74",
          9168 => x"73",
          9169 => x"0a",
          9170 => x"00",
          9171 => x"64",
          9172 => x"00",
          9173 => x"6c",
          9174 => x"00",
          9175 => x"00",
          9176 => x"58",
          9177 => x"00",
          9178 => x"20",
          9179 => x"20",
          9180 => x"00",
          9181 => x"58",
          9182 => x"00",
          9183 => x"00",
          9184 => x"00",
          9185 => x"00",
          9186 => x"00",
          9187 => x"20",
          9188 => x"28",
          9189 => x"00",
          9190 => x"30",
          9191 => x"30",
          9192 => x"00",
          9193 => x"30",
          9194 => x"00",
          9195 => x"55",
          9196 => x"65",
          9197 => x"30",
          9198 => x"20",
          9199 => x"25",
          9200 => x"2a",
          9201 => x"00",
          9202 => x"20",
          9203 => x"65",
          9204 => x"70",
          9205 => x"61",
          9206 => x"65",
          9207 => x"00",
          9208 => x"65",
          9209 => x"6e",
          9210 => x"72",
          9211 => x"00",
          9212 => x"20",
          9213 => x"65",
          9214 => x"70",
          9215 => x"00",
          9216 => x"54",
          9217 => x"44",
          9218 => x"74",
          9219 => x"75",
          9220 => x"00",
          9221 => x"54",
          9222 => x"52",
          9223 => x"74",
          9224 => x"75",
          9225 => x"00",
          9226 => x"54",
          9227 => x"58",
          9228 => x"74",
          9229 => x"75",
          9230 => x"00",
          9231 => x"54",
          9232 => x"58",
          9233 => x"74",
          9234 => x"75",
          9235 => x"00",
          9236 => x"54",
          9237 => x"58",
          9238 => x"74",
          9239 => x"75",
          9240 => x"00",
          9241 => x"54",
          9242 => x"58",
          9243 => x"74",
          9244 => x"75",
          9245 => x"00",
          9246 => x"74",
          9247 => x"20",
          9248 => x"74",
          9249 => x"72",
          9250 => x"00",
          9251 => x"62",
          9252 => x"67",
          9253 => x"6d",
          9254 => x"2e",
          9255 => x"00",
          9256 => x"6f",
          9257 => x"63",
          9258 => x"74",
          9259 => x"00",
          9260 => x"2e",
          9261 => x"00",
          9262 => x"00",
          9263 => x"6c",
          9264 => x"74",
          9265 => x"6e",
          9266 => x"61",
          9267 => x"65",
          9268 => x"20",
          9269 => x"64",
          9270 => x"20",
          9271 => x"61",
          9272 => x"69",
          9273 => x"20",
          9274 => x"75",
          9275 => x"79",
          9276 => x"00",
          9277 => x"00",
          9278 => x"61",
          9279 => x"67",
          9280 => x"2e",
          9281 => x"00",
          9282 => x"79",
          9283 => x"2e",
          9284 => x"00",
          9285 => x"70",
          9286 => x"6e",
          9287 => x"2e",
          9288 => x"00",
          9289 => x"6c",
          9290 => x"30",
          9291 => x"2d",
          9292 => x"38",
          9293 => x"25",
          9294 => x"29",
          9295 => x"00",
          9296 => x"70",
          9297 => x"6d",
          9298 => x"00",
          9299 => x"6d",
          9300 => x"74",
          9301 => x"00",
          9302 => x"6c",
          9303 => x"30",
          9304 => x"00",
          9305 => x"00",
          9306 => x"6c",
          9307 => x"30",
          9308 => x"00",
          9309 => x"6c",
          9310 => x"30",
          9311 => x"2d",
          9312 => x"00",
          9313 => x"63",
          9314 => x"6e",
          9315 => x"6f",
          9316 => x"40",
          9317 => x"38",
          9318 => x"2e",
          9319 => x"00",
          9320 => x"6c",
          9321 => x"20",
          9322 => x"65",
          9323 => x"25",
          9324 => x"78",
          9325 => x"2e",
          9326 => x"00",
          9327 => x"6c",
          9328 => x"74",
          9329 => x"65",
          9330 => x"6f",
          9331 => x"28",
          9332 => x"2e",
          9333 => x"00",
          9334 => x"74",
          9335 => x"69",
          9336 => x"61",
          9337 => x"69",
          9338 => x"69",
          9339 => x"2e",
          9340 => x"00",
          9341 => x"64",
          9342 => x"62",
          9343 => x"69",
          9344 => x"2e",
          9345 => x"00",
          9346 => x"00",
          9347 => x"00",
          9348 => x"5c",
          9349 => x"25",
          9350 => x"73",
          9351 => x"00",
          9352 => x"5c",
          9353 => x"25",
          9354 => x"00",
          9355 => x"5c",
          9356 => x"00",
          9357 => x"20",
          9358 => x"6d",
          9359 => x"2e",
          9360 => x"00",
          9361 => x"6e",
          9362 => x"2e",
          9363 => x"00",
          9364 => x"62",
          9365 => x"67",
          9366 => x"74",
          9367 => x"75",
          9368 => x"2e",
          9369 => x"00",
          9370 => x"25",
          9371 => x"64",
          9372 => x"3a",
          9373 => x"25",
          9374 => x"64",
          9375 => x"00",
          9376 => x"20",
          9377 => x"66",
          9378 => x"72",
          9379 => x"6f",
          9380 => x"00",
          9381 => x"72",
          9382 => x"53",
          9383 => x"63",
          9384 => x"69",
          9385 => x"00",
          9386 => x"65",
          9387 => x"65",
          9388 => x"6d",
          9389 => x"6d",
          9390 => x"65",
          9391 => x"00",
          9392 => x"20",
          9393 => x"53",
          9394 => x"4d",
          9395 => x"25",
          9396 => x"3a",
          9397 => x"58",
          9398 => x"00",
          9399 => x"20",
          9400 => x"41",
          9401 => x"20",
          9402 => x"25",
          9403 => x"3a",
          9404 => x"58",
          9405 => x"00",
          9406 => x"20",
          9407 => x"4e",
          9408 => x"41",
          9409 => x"25",
          9410 => x"3a",
          9411 => x"58",
          9412 => x"00",
          9413 => x"20",
          9414 => x"4d",
          9415 => x"20",
          9416 => x"25",
          9417 => x"3a",
          9418 => x"58",
          9419 => x"00",
          9420 => x"20",
          9421 => x"20",
          9422 => x"20",
          9423 => x"25",
          9424 => x"3a",
          9425 => x"58",
          9426 => x"00",
          9427 => x"20",
          9428 => x"43",
          9429 => x"20",
          9430 => x"44",
          9431 => x"63",
          9432 => x"3d",
          9433 => x"64",
          9434 => x"00",
          9435 => x"20",
          9436 => x"45",
          9437 => x"20",
          9438 => x"54",
          9439 => x"72",
          9440 => x"3d",
          9441 => x"64",
          9442 => x"00",
          9443 => x"20",
          9444 => x"52",
          9445 => x"52",
          9446 => x"43",
          9447 => x"6e",
          9448 => x"3d",
          9449 => x"64",
          9450 => x"00",
          9451 => x"20",
          9452 => x"48",
          9453 => x"45",
          9454 => x"53",
          9455 => x"00",
          9456 => x"20",
          9457 => x"49",
          9458 => x"00",
          9459 => x"20",
          9460 => x"54",
          9461 => x"00",
          9462 => x"20",
          9463 => x"0a",
          9464 => x"00",
          9465 => x"20",
          9466 => x"0a",
          9467 => x"00",
          9468 => x"72",
          9469 => x"65",
          9470 => x"00",
          9471 => x"20",
          9472 => x"20",
          9473 => x"65",
          9474 => x"65",
          9475 => x"72",
          9476 => x"64",
          9477 => x"73",
          9478 => x"25",
          9479 => x"0a",
          9480 => x"00",
          9481 => x"20",
          9482 => x"20",
          9483 => x"6f",
          9484 => x"53",
          9485 => x"74",
          9486 => x"64",
          9487 => x"73",
          9488 => x"25",
          9489 => x"0a",
          9490 => x"00",
          9491 => x"20",
          9492 => x"63",
          9493 => x"74",
          9494 => x"20",
          9495 => x"72",
          9496 => x"20",
          9497 => x"20",
          9498 => x"25",
          9499 => x"0a",
          9500 => x"00",
          9501 => x"63",
          9502 => x"00",
          9503 => x"20",
          9504 => x"20",
          9505 => x"20",
          9506 => x"20",
          9507 => x"20",
          9508 => x"20",
          9509 => x"20",
          9510 => x"25",
          9511 => x"0a",
          9512 => x"00",
          9513 => x"20",
          9514 => x"74",
          9515 => x"43",
          9516 => x"6b",
          9517 => x"65",
          9518 => x"20",
          9519 => x"20",
          9520 => x"25",
          9521 => x"30",
          9522 => x"48",
          9523 => x"00",
          9524 => x"20",
          9525 => x"41",
          9526 => x"6c",
          9527 => x"20",
          9528 => x"71",
          9529 => x"20",
          9530 => x"20",
          9531 => x"25",
          9532 => x"30",
          9533 => x"48",
          9534 => x"00",
          9535 => x"20",
          9536 => x"68",
          9537 => x"65",
          9538 => x"52",
          9539 => x"43",
          9540 => x"6b",
          9541 => x"65",
          9542 => x"25",
          9543 => x"30",
          9544 => x"48",
          9545 => x"00",
          9546 => x"6c",
          9547 => x"00",
          9548 => x"69",
          9549 => x"00",
          9550 => x"78",
          9551 => x"00",
          9552 => x"00",
          9553 => x"6d",
          9554 => x"00",
          9555 => x"6e",
          9556 => x"00",
          9557 => x"b0",
          9558 => x"00",
          9559 => x"02",
          9560 => x"ac",
          9561 => x"00",
          9562 => x"03",
          9563 => x"a8",
          9564 => x"00",
          9565 => x"04",
          9566 => x"a4",
          9567 => x"00",
          9568 => x"05",
          9569 => x"a0",
          9570 => x"00",
          9571 => x"06",
          9572 => x"9c",
          9573 => x"00",
          9574 => x"07",
          9575 => x"98",
          9576 => x"00",
          9577 => x"01",
          9578 => x"94",
          9579 => x"00",
          9580 => x"08",
          9581 => x"90",
          9582 => x"00",
          9583 => x"0b",
          9584 => x"8c",
          9585 => x"00",
          9586 => x"09",
          9587 => x"88",
          9588 => x"00",
          9589 => x"0a",
          9590 => x"84",
          9591 => x"00",
          9592 => x"0d",
          9593 => x"80",
          9594 => x"00",
          9595 => x"0c",
          9596 => x"7c",
          9597 => x"00",
          9598 => x"0e",
          9599 => x"78",
          9600 => x"00",
          9601 => x"0f",
          9602 => x"74",
          9603 => x"00",
          9604 => x"0f",
          9605 => x"70",
          9606 => x"00",
          9607 => x"10",
          9608 => x"6c",
          9609 => x"00",
          9610 => x"11",
          9611 => x"68",
          9612 => x"00",
          9613 => x"12",
          9614 => x"64",
          9615 => x"00",
          9616 => x"13",
          9617 => x"60",
          9618 => x"00",
          9619 => x"14",
          9620 => x"5c",
          9621 => x"00",
          9622 => x"15",
          9623 => x"00",
          9624 => x"00",
          9625 => x"00",
          9626 => x"00",
          9627 => x"7e",
          9628 => x"7e",
          9629 => x"7e",
          9630 => x"00",
          9631 => x"7e",
          9632 => x"7e",
          9633 => x"7e",
          9634 => x"00",
          9635 => x"00",
          9636 => x"00",
          9637 => x"00",
          9638 => x"00",
          9639 => x"00",
          9640 => x"00",
          9641 => x"00",
          9642 => x"00",
          9643 => x"00",
          9644 => x"00",
          9645 => x"74",
          9646 => x"00",
          9647 => x"74",
          9648 => x"00",
          9649 => x"00",
          9650 => x"6c",
          9651 => x"25",
          9652 => x"00",
          9653 => x"6c",
          9654 => x"74",
          9655 => x"65",
          9656 => x"20",
          9657 => x"20",
          9658 => x"74",
          9659 => x"20",
          9660 => x"65",
          9661 => x"20",
          9662 => x"2e",
          9663 => x"00",
          9664 => x"6e",
          9665 => x"6f",
          9666 => x"2f",
          9667 => x"61",
          9668 => x"68",
          9669 => x"6f",
          9670 => x"66",
          9671 => x"2c",
          9672 => x"73",
          9673 => x"69",
          9674 => x"00",
          9675 => x"00",
          9676 => x"2c",
          9677 => x"3d",
          9678 => x"5d",
          9679 => x"00",
          9680 => x"00",
          9681 => x"33",
          9682 => x"00",
          9683 => x"4d",
          9684 => x"53",
          9685 => x"00",
          9686 => x"4e",
          9687 => x"20",
          9688 => x"46",
          9689 => x"32",
          9690 => x"00",
          9691 => x"4e",
          9692 => x"20",
          9693 => x"46",
          9694 => x"20",
          9695 => x"00",
          9696 => x"2c",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"41",
          9701 => x"80",
          9702 => x"49",
          9703 => x"8f",
          9704 => x"4f",
          9705 => x"55",
          9706 => x"9b",
          9707 => x"9f",
          9708 => x"55",
          9709 => x"a7",
          9710 => x"ab",
          9711 => x"af",
          9712 => x"b3",
          9713 => x"b7",
          9714 => x"bb",
          9715 => x"bf",
          9716 => x"c3",
          9717 => x"c7",
          9718 => x"cb",
          9719 => x"cf",
          9720 => x"d3",
          9721 => x"d7",
          9722 => x"db",
          9723 => x"df",
          9724 => x"e3",
          9725 => x"e7",
          9726 => x"eb",
          9727 => x"ef",
          9728 => x"f3",
          9729 => x"f7",
          9730 => x"fb",
          9731 => x"ff",
          9732 => x"3b",
          9733 => x"2f",
          9734 => x"3a",
          9735 => x"7c",
          9736 => x"00",
          9737 => x"04",
          9738 => x"40",
          9739 => x"00",
          9740 => x"00",
          9741 => x"02",
          9742 => x"08",
          9743 => x"20",
          9744 => x"00",
          9745 => x"00",
          9746 => x"c8",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"d0",
          9751 => x"00",
          9752 => x"00",
          9753 => x"00",
          9754 => x"d8",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"e0",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"e8",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"f0",
          9767 => x"00",
          9768 => x"00",
          9769 => x"00",
          9770 => x"f8",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"00",
          9776 => x"00",
          9777 => x"00",
          9778 => x"08",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"10",
          9783 => x"00",
          9784 => x"00",
          9785 => x"00",
          9786 => x"14",
          9787 => x"00",
          9788 => x"00",
          9789 => x"00",
          9790 => x"18",
          9791 => x"00",
          9792 => x"00",
          9793 => x"00",
          9794 => x"1c",
          9795 => x"00",
          9796 => x"00",
          9797 => x"00",
          9798 => x"20",
          9799 => x"00",
          9800 => x"00",
          9801 => x"00",
          9802 => x"24",
          9803 => x"00",
          9804 => x"00",
          9805 => x"00",
          9806 => x"28",
          9807 => x"00",
          9808 => x"00",
          9809 => x"00",
          9810 => x"2c",
          9811 => x"00",
          9812 => x"00",
          9813 => x"00",
          9814 => x"34",
          9815 => x"00",
          9816 => x"00",
          9817 => x"00",
          9818 => x"38",
          9819 => x"00",
          9820 => x"00",
          9821 => x"00",
          9822 => x"40",
          9823 => x"00",
          9824 => x"00",
          9825 => x"00",
          9826 => x"48",
          9827 => x"00",
          9828 => x"00",
          9829 => x"00",
          9830 => x"50",
          9831 => x"00",
          9832 => x"00",
          9833 => x"00",
          9834 => x"58",
          9835 => x"00",
          9836 => x"00",
          9837 => x"00",
          9838 => x"60",
          9839 => x"00",
          9840 => x"00",
          9841 => x"00",
          9842 => x"68",
          9843 => x"00",
          9844 => x"00",
          9845 => x"00",
          9846 => x"70",
          9847 => x"00",
          9848 => x"00",
          9849 => x"00",
          9850 => x"00",
          9851 => x"00",
          9852 => x"ff",
          9853 => x"00",
          9854 => x"ff",
          9855 => x"00",
          9856 => x"ff",
          9857 => x"00",
          9858 => x"00",
          9859 => x"00",
          9860 => x"ff",
          9861 => x"00",
          9862 => x"00",
          9863 => x"00",
          9864 => x"00",
          9865 => x"00",
          9866 => x"00",
          9867 => x"00",
          9868 => x"00",
          9869 => x"01",
          9870 => x"01",
          9871 => x"01",
          9872 => x"00",
          9873 => x"00",
          9874 => x"00",
          9875 => x"00",
          9876 => x"00",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"00",
          9881 => x"00",
          9882 => x"00",
          9883 => x"00",
          9884 => x"00",
          9885 => x"00",
          9886 => x"00",
          9887 => x"00",
          9888 => x"00",
          9889 => x"00",
          9890 => x"00",
          9891 => x"00",
          9892 => x"00",
          9893 => x"00",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"b4",
          9898 => x"00",
          9899 => x"bc",
          9900 => x"00",
          9901 => x"c4",
          9902 => x"00",
          9903 => x"00",
          9904 => x"00",
          9905 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"83",
             1 => x"0b",
             2 => x"b9",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"82",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"80",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"80",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a4",
           270 => x"0b",
           271 => x"0b",
           272 => x"c2",
           273 => x"0b",
           274 => x"0b",
           275 => x"e0",
           276 => x"0b",
           277 => x"0b",
           278 => x"80",
           279 => x"0b",
           280 => x"0b",
           281 => x"9e",
           282 => x"0b",
           283 => x"0b",
           284 => x"bd",
           285 => x"0b",
           286 => x"0b",
           287 => x"dd",
           288 => x"0b",
           289 => x"0b",
           290 => x"fd",
           291 => x"0b",
           292 => x"0b",
           293 => x"9d",
           294 => x"0b",
           295 => x"0b",
           296 => x"bd",
           297 => x"0b",
           298 => x"0b",
           299 => x"dd",
           300 => x"0b",
           301 => x"0b",
           302 => x"fd",
           303 => x"0b",
           304 => x"0b",
           305 => x"9d",
           306 => x"0b",
           307 => x"0b",
           308 => x"bd",
           309 => x"0b",
           310 => x"0b",
           311 => x"dd",
           312 => x"0b",
           313 => x"0b",
           314 => x"fd",
           315 => x"0b",
           316 => x"0b",
           317 => x"9d",
           318 => x"0b",
           319 => x"0b",
           320 => x"bd",
           321 => x"0b",
           322 => x"0b",
           323 => x"dd",
           324 => x"0b",
           325 => x"0b",
           326 => x"fd",
           327 => x"0b",
           328 => x"0b",
           329 => x"9d",
           330 => x"0b",
           331 => x"0b",
           332 => x"bd",
           333 => x"0b",
           334 => x"0b",
           335 => x"dd",
           336 => x"0b",
           337 => x"0b",
           338 => x"fd",
           339 => x"0b",
           340 => x"0b",
           341 => x"9d",
           342 => x"0b",
           343 => x"0b",
           344 => x"bd",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"b5",
           386 => x"f4",
           387 => x"b5",
           388 => x"d0",
           389 => x"b5",
           390 => x"b2",
           391 => x"d4",
           392 => x"90",
           393 => x"d4",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"82",
           399 => x"82",
           400 => x"82",
           401 => x"94",
           402 => x"b5",
           403 => x"d0",
           404 => x"b5",
           405 => x"c2",
           406 => x"d4",
           407 => x"90",
           408 => x"d4",
           409 => x"cc",
           410 => x"d4",
           411 => x"90",
           412 => x"d4",
           413 => x"fb",
           414 => x"d4",
           415 => x"90",
           416 => x"d4",
           417 => x"2d",
           418 => x"08",
           419 => x"04",
           420 => x"0c",
           421 => x"82",
           422 => x"82",
           423 => x"82",
           424 => x"97",
           425 => x"b5",
           426 => x"d0",
           427 => x"b5",
           428 => x"f8",
           429 => x"b5",
           430 => x"d0",
           431 => x"b5",
           432 => x"f8",
           433 => x"b5",
           434 => x"d0",
           435 => x"b5",
           436 => x"f0",
           437 => x"b5",
           438 => x"d0",
           439 => x"b5",
           440 => x"f2",
           441 => x"b5",
           442 => x"d0",
           443 => x"b5",
           444 => x"f3",
           445 => x"b5",
           446 => x"d0",
           447 => x"b5",
           448 => x"d7",
           449 => x"b5",
           450 => x"d0",
           451 => x"b5",
           452 => x"e4",
           453 => x"b5",
           454 => x"d0",
           455 => x"b5",
           456 => x"dc",
           457 => x"b5",
           458 => x"d0",
           459 => x"b5",
           460 => x"df",
           461 => x"b5",
           462 => x"d0",
           463 => x"b5",
           464 => x"e9",
           465 => x"b5",
           466 => x"d0",
           467 => x"b5",
           468 => x"f2",
           469 => x"b5",
           470 => x"d0",
           471 => x"b5",
           472 => x"e3",
           473 => x"b5",
           474 => x"d0",
           475 => x"b5",
           476 => x"ed",
           477 => x"b5",
           478 => x"d0",
           479 => x"b5",
           480 => x"ee",
           481 => x"b5",
           482 => x"d0",
           483 => x"b5",
           484 => x"ee",
           485 => x"b5",
           486 => x"d0",
           487 => x"b5",
           488 => x"f6",
           489 => x"b5",
           490 => x"d0",
           491 => x"b5",
           492 => x"f4",
           493 => x"b5",
           494 => x"d0",
           495 => x"b5",
           496 => x"f9",
           497 => x"b5",
           498 => x"d0",
           499 => x"b5",
           500 => x"ef",
           501 => x"b5",
           502 => x"d0",
           503 => x"b5",
           504 => x"fc",
           505 => x"b5",
           506 => x"d0",
           507 => x"b5",
           508 => x"fd",
           509 => x"b5",
           510 => x"d0",
           511 => x"b5",
           512 => x"e5",
           513 => x"b5",
           514 => x"d0",
           515 => x"b5",
           516 => x"e5",
           517 => x"b5",
           518 => x"d0",
           519 => x"b5",
           520 => x"e6",
           521 => x"b5",
           522 => x"d0",
           523 => x"b5",
           524 => x"f0",
           525 => x"b5",
           526 => x"d0",
           527 => x"b5",
           528 => x"fe",
           529 => x"b5",
           530 => x"d0",
           531 => x"b5",
           532 => x"80",
           533 => x"b5",
           534 => x"d0",
           535 => x"b5",
           536 => x"83",
           537 => x"b5",
           538 => x"d0",
           539 => x"b5",
           540 => x"d7",
           541 => x"b5",
           542 => x"d0",
           543 => x"b5",
           544 => x"86",
           545 => x"b5",
           546 => x"d0",
           547 => x"b5",
           548 => x"94",
           549 => x"b5",
           550 => x"d0",
           551 => x"b5",
           552 => x"92",
           553 => x"b5",
           554 => x"d0",
           555 => x"b5",
           556 => x"a8",
           557 => x"b5",
           558 => x"d0",
           559 => x"b5",
           560 => x"aa",
           561 => x"b5",
           562 => x"d0",
           563 => x"b5",
           564 => x"ac",
           565 => x"b5",
           566 => x"d0",
           567 => x"b5",
           568 => x"f0",
           569 => x"b5",
           570 => x"d0",
           571 => x"b5",
           572 => x"f1",
           573 => x"b5",
           574 => x"d0",
           575 => x"b5",
           576 => x"f5",
           577 => x"b5",
           578 => x"d0",
           579 => x"b5",
           580 => x"d6",
           581 => x"b5",
           582 => x"d0",
           583 => x"b5",
           584 => x"a2",
           585 => x"b5",
           586 => x"d0",
           587 => x"b5",
           588 => x"a3",
           589 => x"b5",
           590 => x"d0",
           591 => x"b5",
           592 => x"a7",
           593 => x"b5",
           594 => x"d0",
           595 => x"b5",
           596 => x"9f",
           597 => x"b5",
           598 => x"d0",
           599 => x"04",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"04",
           609 => x"81",
           610 => x"83",
           611 => x"05",
           612 => x"10",
           613 => x"72",
           614 => x"51",
           615 => x"72",
           616 => x"06",
           617 => x"72",
           618 => x"10",
           619 => x"10",
           620 => x"ed",
           621 => x"53",
           622 => x"b5",
           623 => x"cd",
           624 => x"38",
           625 => x"84",
           626 => x"0b",
           627 => x"bc",
           628 => x"51",
           629 => x"04",
           630 => x"d4",
           631 => x"b5",
           632 => x"3d",
           633 => x"d4",
           634 => x"70",
           635 => x"08",
           636 => x"82",
           637 => x"fc",
           638 => x"82",
           639 => x"88",
           640 => x"82",
           641 => x"52",
           642 => x"3f",
           643 => x"08",
           644 => x"d4",
           645 => x"0c",
           646 => x"08",
           647 => x"70",
           648 => x"0c",
           649 => x"3d",
           650 => x"d4",
           651 => x"b5",
           652 => x"82",
           653 => x"fb",
           654 => x"b5",
           655 => x"05",
           656 => x"33",
           657 => x"70",
           658 => x"51",
           659 => x"8f",
           660 => x"82",
           661 => x"8c",
           662 => x"83",
           663 => x"80",
           664 => x"d4",
           665 => x"0c",
           666 => x"82",
           667 => x"8c",
           668 => x"05",
           669 => x"08",
           670 => x"80",
           671 => x"d4",
           672 => x"0c",
           673 => x"08",
           674 => x"82",
           675 => x"fc",
           676 => x"b5",
           677 => x"05",
           678 => x"80",
           679 => x"0b",
           680 => x"08",
           681 => x"25",
           682 => x"82",
           683 => x"90",
           684 => x"a0",
           685 => x"b5",
           686 => x"82",
           687 => x"f8",
           688 => x"82",
           689 => x"f8",
           690 => x"2e",
           691 => x"8d",
           692 => x"82",
           693 => x"f4",
           694 => x"d2",
           695 => x"d4",
           696 => x"08",
           697 => x"08",
           698 => x"53",
           699 => x"34",
           700 => x"08",
           701 => x"ff",
           702 => x"d4",
           703 => x"0c",
           704 => x"08",
           705 => x"81",
           706 => x"d4",
           707 => x"0c",
           708 => x"82",
           709 => x"fc",
           710 => x"80",
           711 => x"b5",
           712 => x"05",
           713 => x"b5",
           714 => x"05",
           715 => x"b5",
           716 => x"05",
           717 => x"c8",
           718 => x"0d",
           719 => x"0c",
           720 => x"d4",
           721 => x"b5",
           722 => x"3d",
           723 => x"82",
           724 => x"e5",
           725 => x"b5",
           726 => x"05",
           727 => x"d4",
           728 => x"0c",
           729 => x"82",
           730 => x"e8",
           731 => x"b5",
           732 => x"05",
           733 => x"d4",
           734 => x"0c",
           735 => x"08",
           736 => x"54",
           737 => x"08",
           738 => x"53",
           739 => x"08",
           740 => x"53",
           741 => x"8d",
           742 => x"c8",
           743 => x"b5",
           744 => x"05",
           745 => x"d4",
           746 => x"08",
           747 => x"08",
           748 => x"05",
           749 => x"74",
           750 => x"d4",
           751 => x"08",
           752 => x"c8",
           753 => x"3d",
           754 => x"d4",
           755 => x"b5",
           756 => x"82",
           757 => x"fb",
           758 => x"b5",
           759 => x"05",
           760 => x"d4",
           761 => x"0c",
           762 => x"08",
           763 => x"54",
           764 => x"08",
           765 => x"53",
           766 => x"08",
           767 => x"52",
           768 => x"82",
           769 => x"70",
           770 => x"08",
           771 => x"82",
           772 => x"f8",
           773 => x"82",
           774 => x"51",
           775 => x"0d",
           776 => x"0c",
           777 => x"d4",
           778 => x"b5",
           779 => x"3d",
           780 => x"82",
           781 => x"e4",
           782 => x"b5",
           783 => x"05",
           784 => x"0b",
           785 => x"82",
           786 => x"88",
           787 => x"11",
           788 => x"2a",
           789 => x"70",
           790 => x"51",
           791 => x"72",
           792 => x"38",
           793 => x"b5",
           794 => x"05",
           795 => x"39",
           796 => x"08",
           797 => x"53",
           798 => x"72",
           799 => x"08",
           800 => x"72",
           801 => x"53",
           802 => x"95",
           803 => x"b5",
           804 => x"05",
           805 => x"82",
           806 => x"8c",
           807 => x"b5",
           808 => x"05",
           809 => x"06",
           810 => x"80",
           811 => x"38",
           812 => x"08",
           813 => x"53",
           814 => x"81",
           815 => x"b5",
           816 => x"05",
           817 => x"b9",
           818 => x"38",
           819 => x"08",
           820 => x"53",
           821 => x"09",
           822 => x"c5",
           823 => x"d4",
           824 => x"33",
           825 => x"70",
           826 => x"51",
           827 => x"38",
           828 => x"08",
           829 => x"70",
           830 => x"81",
           831 => x"06",
           832 => x"53",
           833 => x"99",
           834 => x"d4",
           835 => x"22",
           836 => x"07",
           837 => x"82",
           838 => x"e4",
           839 => x"d0",
           840 => x"d4",
           841 => x"33",
           842 => x"70",
           843 => x"70",
           844 => x"11",
           845 => x"51",
           846 => x"55",
           847 => x"b5",
           848 => x"05",
           849 => x"d4",
           850 => x"33",
           851 => x"d4",
           852 => x"33",
           853 => x"11",
           854 => x"72",
           855 => x"08",
           856 => x"82",
           857 => x"e8",
           858 => x"98",
           859 => x"2c",
           860 => x"72",
           861 => x"38",
           862 => x"82",
           863 => x"e8",
           864 => x"b5",
           865 => x"05",
           866 => x"2a",
           867 => x"51",
           868 => x"fd",
           869 => x"b5",
           870 => x"05",
           871 => x"2b",
           872 => x"70",
           873 => x"88",
           874 => x"51",
           875 => x"82",
           876 => x"ec",
           877 => x"b8",
           878 => x"d4",
           879 => x"22",
           880 => x"70",
           881 => x"51",
           882 => x"2e",
           883 => x"b5",
           884 => x"05",
           885 => x"2b",
           886 => x"51",
           887 => x"8a",
           888 => x"82",
           889 => x"e8",
           890 => x"b5",
           891 => x"05",
           892 => x"82",
           893 => x"c4",
           894 => x"82",
           895 => x"c4",
           896 => x"d8",
           897 => x"38",
           898 => x"08",
           899 => x"70",
           900 => x"96",
           901 => x"08",
           902 => x"53",
           903 => x"b5",
           904 => x"05",
           905 => x"07",
           906 => x"82",
           907 => x"e4",
           908 => x"b5",
           909 => x"05",
           910 => x"07",
           911 => x"82",
           912 => x"e4",
           913 => x"a8",
           914 => x"d4",
           915 => x"22",
           916 => x"07",
           917 => x"82",
           918 => x"e4",
           919 => x"90",
           920 => x"d4",
           921 => x"22",
           922 => x"07",
           923 => x"82",
           924 => x"e4",
           925 => x"f8",
           926 => x"d4",
           927 => x"22",
           928 => x"51",
           929 => x"b5",
           930 => x"05",
           931 => x"82",
           932 => x"e8",
           933 => x"d8",
           934 => x"d4",
           935 => x"22",
           936 => x"51",
           937 => x"b5",
           938 => x"05",
           939 => x"39",
           940 => x"b5",
           941 => x"05",
           942 => x"d4",
           943 => x"22",
           944 => x"53",
           945 => x"d4",
           946 => x"23",
           947 => x"82",
           948 => x"f8",
           949 => x"a8",
           950 => x"d4",
           951 => x"08",
           952 => x"08",
           953 => x"84",
           954 => x"d4",
           955 => x"0c",
           956 => x"53",
           957 => x"d4",
           958 => x"34",
           959 => x"08",
           960 => x"ff",
           961 => x"72",
           962 => x"08",
           963 => x"8c",
           964 => x"b5",
           965 => x"05",
           966 => x"d4",
           967 => x"08",
           968 => x"b5",
           969 => x"05",
           970 => x"82",
           971 => x"fc",
           972 => x"b5",
           973 => x"05",
           974 => x"2a",
           975 => x"51",
           976 => x"72",
           977 => x"38",
           978 => x"08",
           979 => x"70",
           980 => x"72",
           981 => x"82",
           982 => x"fc",
           983 => x"53",
           984 => x"82",
           985 => x"53",
           986 => x"d4",
           987 => x"23",
           988 => x"b5",
           989 => x"05",
           990 => x"8a",
           991 => x"c8",
           992 => x"82",
           993 => x"f4",
           994 => x"b5",
           995 => x"05",
           996 => x"b5",
           997 => x"05",
           998 => x"31",
           999 => x"82",
          1000 => x"ec",
          1001 => x"d8",
          1002 => x"d4",
          1003 => x"08",
          1004 => x"08",
          1005 => x"84",
          1006 => x"d4",
          1007 => x"0c",
          1008 => x"b5",
          1009 => x"05",
          1010 => x"d4",
          1011 => x"22",
          1012 => x"70",
          1013 => x"51",
          1014 => x"80",
          1015 => x"82",
          1016 => x"e8",
          1017 => x"98",
          1018 => x"98",
          1019 => x"b5",
          1020 => x"05",
          1021 => x"a1",
          1022 => x"b5",
          1023 => x"72",
          1024 => x"08",
          1025 => x"99",
          1026 => x"d4",
          1027 => x"08",
          1028 => x"3f",
          1029 => x"08",
          1030 => x"b5",
          1031 => x"05",
          1032 => x"d4",
          1033 => x"22",
          1034 => x"d4",
          1035 => x"22",
          1036 => x"54",
          1037 => x"b5",
          1038 => x"05",
          1039 => x"39",
          1040 => x"08",
          1041 => x"70",
          1042 => x"81",
          1043 => x"53",
          1044 => x"a4",
          1045 => x"d4",
          1046 => x"08",
          1047 => x"08",
          1048 => x"84",
          1049 => x"d4",
          1050 => x"0c",
          1051 => x"b5",
          1052 => x"05",
          1053 => x"39",
          1054 => x"08",
          1055 => x"82",
          1056 => x"90",
          1057 => x"05",
          1058 => x"08",
          1059 => x"70",
          1060 => x"d4",
          1061 => x"0c",
          1062 => x"d4",
          1063 => x"08",
          1064 => x"08",
          1065 => x"82",
          1066 => x"fc",
          1067 => x"25",
          1068 => x"b5",
          1069 => x"05",
          1070 => x"07",
          1071 => x"82",
          1072 => x"e4",
          1073 => x"b5",
          1074 => x"05",
          1075 => x"b5",
          1076 => x"05",
          1077 => x"d4",
          1078 => x"22",
          1079 => x"06",
          1080 => x"82",
          1081 => x"e4",
          1082 => x"af",
          1083 => x"82",
          1084 => x"f4",
          1085 => x"39",
          1086 => x"08",
          1087 => x"70",
          1088 => x"51",
          1089 => x"b5",
          1090 => x"05",
          1091 => x"0b",
          1092 => x"08",
          1093 => x"90",
          1094 => x"d4",
          1095 => x"23",
          1096 => x"08",
          1097 => x"70",
          1098 => x"81",
          1099 => x"53",
          1100 => x"a4",
          1101 => x"d4",
          1102 => x"08",
          1103 => x"08",
          1104 => x"84",
          1105 => x"d4",
          1106 => x"0c",
          1107 => x"b5",
          1108 => x"05",
          1109 => x"39",
          1110 => x"08",
          1111 => x"82",
          1112 => x"90",
          1113 => x"05",
          1114 => x"08",
          1115 => x"70",
          1116 => x"d4",
          1117 => x"0c",
          1118 => x"d4",
          1119 => x"08",
          1120 => x"08",
          1121 => x"82",
          1122 => x"e4",
          1123 => x"cf",
          1124 => x"72",
          1125 => x"08",
          1126 => x"82",
          1127 => x"82",
          1128 => x"f0",
          1129 => x"b5",
          1130 => x"05",
          1131 => x"d4",
          1132 => x"22",
          1133 => x"08",
          1134 => x"71",
          1135 => x"56",
          1136 => x"f3",
          1137 => x"c8",
          1138 => x"75",
          1139 => x"d4",
          1140 => x"08",
          1141 => x"08",
          1142 => x"82",
          1143 => x"f0",
          1144 => x"33",
          1145 => x"73",
          1146 => x"82",
          1147 => x"f0",
          1148 => x"72",
          1149 => x"b5",
          1150 => x"05",
          1151 => x"df",
          1152 => x"53",
          1153 => x"d4",
          1154 => x"34",
          1155 => x"b5",
          1156 => x"05",
          1157 => x"33",
          1158 => x"53",
          1159 => x"d4",
          1160 => x"34",
          1161 => x"08",
          1162 => x"53",
          1163 => x"08",
          1164 => x"73",
          1165 => x"d4",
          1166 => x"08",
          1167 => x"b5",
          1168 => x"05",
          1169 => x"d4",
          1170 => x"22",
          1171 => x"b5",
          1172 => x"05",
          1173 => x"a2",
          1174 => x"b5",
          1175 => x"82",
          1176 => x"fc",
          1177 => x"82",
          1178 => x"fc",
          1179 => x"2e",
          1180 => x"b2",
          1181 => x"d4",
          1182 => x"08",
          1183 => x"54",
          1184 => x"74",
          1185 => x"51",
          1186 => x"b5",
          1187 => x"05",
          1188 => x"d4",
          1189 => x"22",
          1190 => x"51",
          1191 => x"2e",
          1192 => x"b5",
          1193 => x"05",
          1194 => x"51",
          1195 => x"b5",
          1196 => x"05",
          1197 => x"d4",
          1198 => x"22",
          1199 => x"70",
          1200 => x"51",
          1201 => x"2e",
          1202 => x"82",
          1203 => x"ec",
          1204 => x"90",
          1205 => x"d4",
          1206 => x"0c",
          1207 => x"08",
          1208 => x"90",
          1209 => x"d4",
          1210 => x"0c",
          1211 => x"08",
          1212 => x"51",
          1213 => x"2e",
          1214 => x"95",
          1215 => x"d4",
          1216 => x"08",
          1217 => x"72",
          1218 => x"08",
          1219 => x"93",
          1220 => x"d4",
          1221 => x"08",
          1222 => x"72",
          1223 => x"08",
          1224 => x"82",
          1225 => x"c8",
          1226 => x"b5",
          1227 => x"05",
          1228 => x"d4",
          1229 => x"22",
          1230 => x"70",
          1231 => x"51",
          1232 => x"2e",
          1233 => x"82",
          1234 => x"e8",
          1235 => x"98",
          1236 => x"2c",
          1237 => x"08",
          1238 => x"57",
          1239 => x"72",
          1240 => x"38",
          1241 => x"08",
          1242 => x"70",
          1243 => x"53",
          1244 => x"d4",
          1245 => x"23",
          1246 => x"b5",
          1247 => x"05",
          1248 => x"b5",
          1249 => x"05",
          1250 => x"31",
          1251 => x"82",
          1252 => x"e8",
          1253 => x"b5",
          1254 => x"05",
          1255 => x"2a",
          1256 => x"51",
          1257 => x"80",
          1258 => x"82",
          1259 => x"e8",
          1260 => x"88",
          1261 => x"2b",
          1262 => x"70",
          1263 => x"51",
          1264 => x"72",
          1265 => x"d4",
          1266 => x"22",
          1267 => x"51",
          1268 => x"b5",
          1269 => x"05",
          1270 => x"82",
          1271 => x"fc",
          1272 => x"88",
          1273 => x"2b",
          1274 => x"70",
          1275 => x"51",
          1276 => x"72",
          1277 => x"d4",
          1278 => x"22",
          1279 => x"51",
          1280 => x"b5",
          1281 => x"05",
          1282 => x"d4",
          1283 => x"22",
          1284 => x"06",
          1285 => x"b0",
          1286 => x"d4",
          1287 => x"22",
          1288 => x"54",
          1289 => x"d4",
          1290 => x"23",
          1291 => x"70",
          1292 => x"53",
          1293 => x"90",
          1294 => x"d4",
          1295 => x"08",
          1296 => x"8a",
          1297 => x"39",
          1298 => x"08",
          1299 => x"70",
          1300 => x"81",
          1301 => x"53",
          1302 => x"91",
          1303 => x"d4",
          1304 => x"08",
          1305 => x"8a",
          1306 => x"c7",
          1307 => x"d4",
          1308 => x"22",
          1309 => x"70",
          1310 => x"51",
          1311 => x"2e",
          1312 => x"b5",
          1313 => x"05",
          1314 => x"51",
          1315 => x"a3",
          1316 => x"d4",
          1317 => x"22",
          1318 => x"70",
          1319 => x"51",
          1320 => x"2e",
          1321 => x"b5",
          1322 => x"05",
          1323 => x"51",
          1324 => x"82",
          1325 => x"e4",
          1326 => x"86",
          1327 => x"06",
          1328 => x"72",
          1329 => x"38",
          1330 => x"08",
          1331 => x"52",
          1332 => x"df",
          1333 => x"d4",
          1334 => x"22",
          1335 => x"2e",
          1336 => x"94",
          1337 => x"d4",
          1338 => x"08",
          1339 => x"d4",
          1340 => x"33",
          1341 => x"3f",
          1342 => x"08",
          1343 => x"70",
          1344 => x"81",
          1345 => x"53",
          1346 => x"b0",
          1347 => x"d4",
          1348 => x"22",
          1349 => x"54",
          1350 => x"d4",
          1351 => x"23",
          1352 => x"70",
          1353 => x"53",
          1354 => x"90",
          1355 => x"d4",
          1356 => x"08",
          1357 => x"88",
          1358 => x"39",
          1359 => x"08",
          1360 => x"70",
          1361 => x"81",
          1362 => x"53",
          1363 => x"b0",
          1364 => x"d4",
          1365 => x"33",
          1366 => x"54",
          1367 => x"d4",
          1368 => x"34",
          1369 => x"70",
          1370 => x"53",
          1371 => x"90",
          1372 => x"d4",
          1373 => x"08",
          1374 => x"88",
          1375 => x"39",
          1376 => x"08",
          1377 => x"70",
          1378 => x"81",
          1379 => x"53",
          1380 => x"82",
          1381 => x"ec",
          1382 => x"11",
          1383 => x"82",
          1384 => x"ec",
          1385 => x"90",
          1386 => x"2c",
          1387 => x"73",
          1388 => x"82",
          1389 => x"88",
          1390 => x"a0",
          1391 => x"3f",
          1392 => x"b5",
          1393 => x"05",
          1394 => x"80",
          1395 => x"81",
          1396 => x"82",
          1397 => x"88",
          1398 => x"82",
          1399 => x"fc",
          1400 => x"87",
          1401 => x"ee",
          1402 => x"d4",
          1403 => x"33",
          1404 => x"f3",
          1405 => x"06",
          1406 => x"82",
          1407 => x"f4",
          1408 => x"11",
          1409 => x"82",
          1410 => x"f4",
          1411 => x"83",
          1412 => x"53",
          1413 => x"ff",
          1414 => x"38",
          1415 => x"08",
          1416 => x"52",
          1417 => x"08",
          1418 => x"70",
          1419 => x"b5",
          1420 => x"05",
          1421 => x"82",
          1422 => x"fc",
          1423 => x"86",
          1424 => x"b7",
          1425 => x"d4",
          1426 => x"33",
          1427 => x"d3",
          1428 => x"06",
          1429 => x"82",
          1430 => x"f4",
          1431 => x"11",
          1432 => x"82",
          1433 => x"f4",
          1434 => x"83",
          1435 => x"53",
          1436 => x"ff",
          1437 => x"38",
          1438 => x"08",
          1439 => x"52",
          1440 => x"08",
          1441 => x"70",
          1442 => x"86",
          1443 => x"b5",
          1444 => x"05",
          1445 => x"82",
          1446 => x"fc",
          1447 => x"b7",
          1448 => x"d4",
          1449 => x"08",
          1450 => x"2e",
          1451 => x"b5",
          1452 => x"05",
          1453 => x"b5",
          1454 => x"05",
          1455 => x"82",
          1456 => x"f0",
          1457 => x"b5",
          1458 => x"05",
          1459 => x"52",
          1460 => x"3f",
          1461 => x"b5",
          1462 => x"05",
          1463 => x"2a",
          1464 => x"51",
          1465 => x"80",
          1466 => x"38",
          1467 => x"08",
          1468 => x"ff",
          1469 => x"72",
          1470 => x"08",
          1471 => x"73",
          1472 => x"90",
          1473 => x"80",
          1474 => x"38",
          1475 => x"08",
          1476 => x"52",
          1477 => x"9b",
          1478 => x"82",
          1479 => x"88",
          1480 => x"82",
          1481 => x"f8",
          1482 => x"85",
          1483 => x"0b",
          1484 => x"08",
          1485 => x"ea",
          1486 => x"b5",
          1487 => x"05",
          1488 => x"a5",
          1489 => x"06",
          1490 => x"0b",
          1491 => x"08",
          1492 => x"80",
          1493 => x"d4",
          1494 => x"23",
          1495 => x"b5",
          1496 => x"05",
          1497 => x"82",
          1498 => x"f4",
          1499 => x"80",
          1500 => x"d4",
          1501 => x"08",
          1502 => x"d4",
          1503 => x"33",
          1504 => x"3f",
          1505 => x"82",
          1506 => x"88",
          1507 => x"11",
          1508 => x"b5",
          1509 => x"05",
          1510 => x"82",
          1511 => x"e0",
          1512 => x"b5",
          1513 => x"3d",
          1514 => x"d4",
          1515 => x"b5",
          1516 => x"82",
          1517 => x"fd",
          1518 => x"cd",
          1519 => x"82",
          1520 => x"8c",
          1521 => x"82",
          1522 => x"88",
          1523 => x"e4",
          1524 => x"b5",
          1525 => x"82",
          1526 => x"54",
          1527 => x"82",
          1528 => x"04",
          1529 => x"08",
          1530 => x"d4",
          1531 => x"0d",
          1532 => x"b5",
          1533 => x"05",
          1534 => x"9c",
          1535 => x"33",
          1536 => x"70",
          1537 => x"81",
          1538 => x"51",
          1539 => x"80",
          1540 => x"ff",
          1541 => x"d4",
          1542 => x"0c",
          1543 => x"82",
          1544 => x"88",
          1545 => x"72",
          1546 => x"d4",
          1547 => x"08",
          1548 => x"b5",
          1549 => x"05",
          1550 => x"82",
          1551 => x"fc",
          1552 => x"81",
          1553 => x"72",
          1554 => x"38",
          1555 => x"08",
          1556 => x"08",
          1557 => x"d4",
          1558 => x"33",
          1559 => x"08",
          1560 => x"2d",
          1561 => x"08",
          1562 => x"2e",
          1563 => x"ff",
          1564 => x"d4",
          1565 => x"0c",
          1566 => x"82",
          1567 => x"82",
          1568 => x"53",
          1569 => x"90",
          1570 => x"72",
          1571 => x"c8",
          1572 => x"80",
          1573 => x"ff",
          1574 => x"d4",
          1575 => x"0c",
          1576 => x"08",
          1577 => x"70",
          1578 => x"08",
          1579 => x"53",
          1580 => x"08",
          1581 => x"82",
          1582 => x"87",
          1583 => x"b5",
          1584 => x"82",
          1585 => x"02",
          1586 => x"0c",
          1587 => x"80",
          1588 => x"d4",
          1589 => x"0c",
          1590 => x"08",
          1591 => x"85",
          1592 => x"81",
          1593 => x"32",
          1594 => x"51",
          1595 => x"53",
          1596 => x"8d",
          1597 => x"82",
          1598 => x"f4",
          1599 => x"f3",
          1600 => x"d4",
          1601 => x"08",
          1602 => x"82",
          1603 => x"88",
          1604 => x"05",
          1605 => x"08",
          1606 => x"53",
          1607 => x"d4",
          1608 => x"34",
          1609 => x"06",
          1610 => x"2e",
          1611 => x"b5",
          1612 => x"05",
          1613 => x"d4",
          1614 => x"08",
          1615 => x"d4",
          1616 => x"33",
          1617 => x"08",
          1618 => x"2d",
          1619 => x"08",
          1620 => x"2e",
          1621 => x"ff",
          1622 => x"d4",
          1623 => x"0c",
          1624 => x"82",
          1625 => x"f8",
          1626 => x"82",
          1627 => x"f4",
          1628 => x"82",
          1629 => x"f4",
          1630 => x"b5",
          1631 => x"3d",
          1632 => x"d4",
          1633 => x"b5",
          1634 => x"82",
          1635 => x"fe",
          1636 => x"cd",
          1637 => x"82",
          1638 => x"88",
          1639 => x"93",
          1640 => x"c8",
          1641 => x"b5",
          1642 => x"84",
          1643 => x"b5",
          1644 => x"82",
          1645 => x"02",
          1646 => x"0c",
          1647 => x"82",
          1648 => x"8c",
          1649 => x"11",
          1650 => x"2a",
          1651 => x"70",
          1652 => x"51",
          1653 => x"72",
          1654 => x"38",
          1655 => x"b5",
          1656 => x"05",
          1657 => x"39",
          1658 => x"08",
          1659 => x"85",
          1660 => x"82",
          1661 => x"06",
          1662 => x"53",
          1663 => x"80",
          1664 => x"b5",
          1665 => x"05",
          1666 => x"d4",
          1667 => x"08",
          1668 => x"14",
          1669 => x"08",
          1670 => x"82",
          1671 => x"8c",
          1672 => x"08",
          1673 => x"d4",
          1674 => x"08",
          1675 => x"54",
          1676 => x"73",
          1677 => x"74",
          1678 => x"d4",
          1679 => x"08",
          1680 => x"81",
          1681 => x"0c",
          1682 => x"08",
          1683 => x"70",
          1684 => x"08",
          1685 => x"51",
          1686 => x"39",
          1687 => x"08",
          1688 => x"82",
          1689 => x"8c",
          1690 => x"82",
          1691 => x"88",
          1692 => x"81",
          1693 => x"90",
          1694 => x"54",
          1695 => x"82",
          1696 => x"53",
          1697 => x"82",
          1698 => x"8c",
          1699 => x"11",
          1700 => x"8c",
          1701 => x"b5",
          1702 => x"05",
          1703 => x"b5",
          1704 => x"05",
          1705 => x"8a",
          1706 => x"82",
          1707 => x"fc",
          1708 => x"b5",
          1709 => x"05",
          1710 => x"c8",
          1711 => x"0d",
          1712 => x"0c",
          1713 => x"d4",
          1714 => x"b5",
          1715 => x"3d",
          1716 => x"d4",
          1717 => x"08",
          1718 => x"70",
          1719 => x"81",
          1720 => x"51",
          1721 => x"2e",
          1722 => x"0b",
          1723 => x"08",
          1724 => x"83",
          1725 => x"b5",
          1726 => x"05",
          1727 => x"33",
          1728 => x"70",
          1729 => x"51",
          1730 => x"80",
          1731 => x"38",
          1732 => x"08",
          1733 => x"82",
          1734 => x"88",
          1735 => x"53",
          1736 => x"70",
          1737 => x"51",
          1738 => x"14",
          1739 => x"d4",
          1740 => x"08",
          1741 => x"81",
          1742 => x"0c",
          1743 => x"08",
          1744 => x"84",
          1745 => x"82",
          1746 => x"f8",
          1747 => x"51",
          1748 => x"39",
          1749 => x"08",
          1750 => x"85",
          1751 => x"82",
          1752 => x"06",
          1753 => x"52",
          1754 => x"80",
          1755 => x"b5",
          1756 => x"05",
          1757 => x"70",
          1758 => x"d4",
          1759 => x"0c",
          1760 => x"b5",
          1761 => x"05",
          1762 => x"82",
          1763 => x"88",
          1764 => x"b5",
          1765 => x"05",
          1766 => x"85",
          1767 => x"a0",
          1768 => x"71",
          1769 => x"ff",
          1770 => x"d4",
          1771 => x"0c",
          1772 => x"82",
          1773 => x"88",
          1774 => x"08",
          1775 => x"0c",
          1776 => x"39",
          1777 => x"08",
          1778 => x"82",
          1779 => x"88",
          1780 => x"94",
          1781 => x"52",
          1782 => x"b5",
          1783 => x"82",
          1784 => x"fc",
          1785 => x"82",
          1786 => x"fc",
          1787 => x"25",
          1788 => x"82",
          1789 => x"88",
          1790 => x"b5",
          1791 => x"05",
          1792 => x"d4",
          1793 => x"08",
          1794 => x"82",
          1795 => x"f0",
          1796 => x"82",
          1797 => x"fc",
          1798 => x"2e",
          1799 => x"95",
          1800 => x"d4",
          1801 => x"08",
          1802 => x"71",
          1803 => x"08",
          1804 => x"93",
          1805 => x"d4",
          1806 => x"08",
          1807 => x"71",
          1808 => x"08",
          1809 => x"82",
          1810 => x"f4",
          1811 => x"82",
          1812 => x"ec",
          1813 => x"13",
          1814 => x"82",
          1815 => x"f8",
          1816 => x"39",
          1817 => x"08",
          1818 => x"8c",
          1819 => x"05",
          1820 => x"82",
          1821 => x"fc",
          1822 => x"81",
          1823 => x"82",
          1824 => x"f8",
          1825 => x"51",
          1826 => x"d4",
          1827 => x"08",
          1828 => x"0c",
          1829 => x"82",
          1830 => x"04",
          1831 => x"08",
          1832 => x"d4",
          1833 => x"0d",
          1834 => x"08",
          1835 => x"82",
          1836 => x"fc",
          1837 => x"b5",
          1838 => x"05",
          1839 => x"d4",
          1840 => x"0c",
          1841 => x"08",
          1842 => x"80",
          1843 => x"38",
          1844 => x"08",
          1845 => x"82",
          1846 => x"fc",
          1847 => x"81",
          1848 => x"b5",
          1849 => x"05",
          1850 => x"d4",
          1851 => x"08",
          1852 => x"b5",
          1853 => x"05",
          1854 => x"81",
          1855 => x"b5",
          1856 => x"05",
          1857 => x"d4",
          1858 => x"08",
          1859 => x"d4",
          1860 => x"0c",
          1861 => x"08",
          1862 => x"82",
          1863 => x"90",
          1864 => x"82",
          1865 => x"f8",
          1866 => x"b5",
          1867 => x"05",
          1868 => x"82",
          1869 => x"90",
          1870 => x"b5",
          1871 => x"05",
          1872 => x"82",
          1873 => x"90",
          1874 => x"b5",
          1875 => x"05",
          1876 => x"81",
          1877 => x"b5",
          1878 => x"05",
          1879 => x"82",
          1880 => x"fc",
          1881 => x"b5",
          1882 => x"05",
          1883 => x"82",
          1884 => x"f8",
          1885 => x"b5",
          1886 => x"05",
          1887 => x"d4",
          1888 => x"08",
          1889 => x"33",
          1890 => x"ae",
          1891 => x"d4",
          1892 => x"08",
          1893 => x"b5",
          1894 => x"05",
          1895 => x"d4",
          1896 => x"08",
          1897 => x"b5",
          1898 => x"05",
          1899 => x"d4",
          1900 => x"08",
          1901 => x"38",
          1902 => x"08",
          1903 => x"51",
          1904 => x"b5",
          1905 => x"05",
          1906 => x"82",
          1907 => x"f8",
          1908 => x"b5",
          1909 => x"05",
          1910 => x"71",
          1911 => x"b5",
          1912 => x"05",
          1913 => x"82",
          1914 => x"fc",
          1915 => x"ad",
          1916 => x"d4",
          1917 => x"08",
          1918 => x"c8",
          1919 => x"3d",
          1920 => x"d4",
          1921 => x"b5",
          1922 => x"82",
          1923 => x"fe",
          1924 => x"b5",
          1925 => x"05",
          1926 => x"d4",
          1927 => x"0c",
          1928 => x"08",
          1929 => x"52",
          1930 => x"b5",
          1931 => x"05",
          1932 => x"82",
          1933 => x"fc",
          1934 => x"81",
          1935 => x"51",
          1936 => x"83",
          1937 => x"82",
          1938 => x"fc",
          1939 => x"05",
          1940 => x"08",
          1941 => x"82",
          1942 => x"fc",
          1943 => x"b5",
          1944 => x"05",
          1945 => x"82",
          1946 => x"51",
          1947 => x"82",
          1948 => x"04",
          1949 => x"08",
          1950 => x"d4",
          1951 => x"0d",
          1952 => x"08",
          1953 => x"82",
          1954 => x"fc",
          1955 => x"b5",
          1956 => x"05",
          1957 => x"33",
          1958 => x"08",
          1959 => x"81",
          1960 => x"d4",
          1961 => x"0c",
          1962 => x"08",
          1963 => x"53",
          1964 => x"34",
          1965 => x"08",
          1966 => x"81",
          1967 => x"d4",
          1968 => x"0c",
          1969 => x"06",
          1970 => x"2e",
          1971 => x"be",
          1972 => x"d4",
          1973 => x"08",
          1974 => x"c8",
          1975 => x"3d",
          1976 => x"d4",
          1977 => x"b5",
          1978 => x"82",
          1979 => x"fd",
          1980 => x"b5",
          1981 => x"05",
          1982 => x"d4",
          1983 => x"0c",
          1984 => x"08",
          1985 => x"82",
          1986 => x"f8",
          1987 => x"b5",
          1988 => x"05",
          1989 => x"80",
          1990 => x"b5",
          1991 => x"05",
          1992 => x"82",
          1993 => x"90",
          1994 => x"b5",
          1995 => x"05",
          1996 => x"82",
          1997 => x"90",
          1998 => x"b5",
          1999 => x"05",
          2000 => x"ba",
          2001 => x"d4",
          2002 => x"08",
          2003 => x"82",
          2004 => x"f8",
          2005 => x"05",
          2006 => x"08",
          2007 => x"82",
          2008 => x"fc",
          2009 => x"52",
          2010 => x"82",
          2011 => x"fc",
          2012 => x"05",
          2013 => x"08",
          2014 => x"ff",
          2015 => x"b5",
          2016 => x"05",
          2017 => x"b5",
          2018 => x"85",
          2019 => x"b5",
          2020 => x"82",
          2021 => x"02",
          2022 => x"0c",
          2023 => x"82",
          2024 => x"90",
          2025 => x"2e",
          2026 => x"82",
          2027 => x"8c",
          2028 => x"71",
          2029 => x"d4",
          2030 => x"08",
          2031 => x"b5",
          2032 => x"05",
          2033 => x"d4",
          2034 => x"08",
          2035 => x"81",
          2036 => x"54",
          2037 => x"71",
          2038 => x"80",
          2039 => x"b5",
          2040 => x"05",
          2041 => x"33",
          2042 => x"08",
          2043 => x"81",
          2044 => x"d4",
          2045 => x"0c",
          2046 => x"06",
          2047 => x"8d",
          2048 => x"82",
          2049 => x"fc",
          2050 => x"9b",
          2051 => x"d4",
          2052 => x"08",
          2053 => x"b5",
          2054 => x"05",
          2055 => x"d4",
          2056 => x"08",
          2057 => x"38",
          2058 => x"82",
          2059 => x"90",
          2060 => x"2e",
          2061 => x"82",
          2062 => x"88",
          2063 => x"33",
          2064 => x"8d",
          2065 => x"82",
          2066 => x"fc",
          2067 => x"d7",
          2068 => x"d4",
          2069 => x"08",
          2070 => x"b5",
          2071 => x"05",
          2072 => x"d4",
          2073 => x"08",
          2074 => x"52",
          2075 => x"81",
          2076 => x"d4",
          2077 => x"0c",
          2078 => x"b5",
          2079 => x"05",
          2080 => x"82",
          2081 => x"8c",
          2082 => x"33",
          2083 => x"70",
          2084 => x"08",
          2085 => x"53",
          2086 => x"53",
          2087 => x"0b",
          2088 => x"08",
          2089 => x"82",
          2090 => x"fc",
          2091 => x"b5",
          2092 => x"3d",
          2093 => x"d4",
          2094 => x"b5",
          2095 => x"82",
          2096 => x"fd",
          2097 => x"b5",
          2098 => x"05",
          2099 => x"d4",
          2100 => x"0c",
          2101 => x"08",
          2102 => x"8d",
          2103 => x"82",
          2104 => x"fc",
          2105 => x"ec",
          2106 => x"d4",
          2107 => x"08",
          2108 => x"82",
          2109 => x"f8",
          2110 => x"05",
          2111 => x"08",
          2112 => x"70",
          2113 => x"51",
          2114 => x"2e",
          2115 => x"b5",
          2116 => x"05",
          2117 => x"82",
          2118 => x"8c",
          2119 => x"b5",
          2120 => x"05",
          2121 => x"84",
          2122 => x"39",
          2123 => x"08",
          2124 => x"ff",
          2125 => x"d4",
          2126 => x"0c",
          2127 => x"08",
          2128 => x"82",
          2129 => x"88",
          2130 => x"70",
          2131 => x"08",
          2132 => x"51",
          2133 => x"08",
          2134 => x"82",
          2135 => x"85",
          2136 => x"b5",
          2137 => x"82",
          2138 => x"02",
          2139 => x"0c",
          2140 => x"82",
          2141 => x"88",
          2142 => x"b5",
          2143 => x"05",
          2144 => x"d4",
          2145 => x"08",
          2146 => x"d4",
          2147 => x"d4",
          2148 => x"08",
          2149 => x"b5",
          2150 => x"05",
          2151 => x"d4",
          2152 => x"08",
          2153 => x"b5",
          2154 => x"05",
          2155 => x"d4",
          2156 => x"08",
          2157 => x"38",
          2158 => x"08",
          2159 => x"51",
          2160 => x"d4",
          2161 => x"08",
          2162 => x"71",
          2163 => x"d4",
          2164 => x"08",
          2165 => x"b5",
          2166 => x"05",
          2167 => x"39",
          2168 => x"08",
          2169 => x"70",
          2170 => x"0c",
          2171 => x"0d",
          2172 => x"0c",
          2173 => x"d4",
          2174 => x"b5",
          2175 => x"3d",
          2176 => x"82",
          2177 => x"fc",
          2178 => x"b5",
          2179 => x"05",
          2180 => x"b9",
          2181 => x"d4",
          2182 => x"08",
          2183 => x"d4",
          2184 => x"0c",
          2185 => x"b5",
          2186 => x"05",
          2187 => x"d4",
          2188 => x"08",
          2189 => x"0b",
          2190 => x"08",
          2191 => x"82",
          2192 => x"f4",
          2193 => x"b5",
          2194 => x"05",
          2195 => x"d4",
          2196 => x"08",
          2197 => x"38",
          2198 => x"08",
          2199 => x"30",
          2200 => x"08",
          2201 => x"80",
          2202 => x"d4",
          2203 => x"0c",
          2204 => x"08",
          2205 => x"8a",
          2206 => x"82",
          2207 => x"f0",
          2208 => x"b5",
          2209 => x"05",
          2210 => x"d4",
          2211 => x"0c",
          2212 => x"b5",
          2213 => x"05",
          2214 => x"b5",
          2215 => x"05",
          2216 => x"c5",
          2217 => x"c8",
          2218 => x"b5",
          2219 => x"05",
          2220 => x"b5",
          2221 => x"05",
          2222 => x"90",
          2223 => x"d4",
          2224 => x"08",
          2225 => x"d4",
          2226 => x"0c",
          2227 => x"08",
          2228 => x"70",
          2229 => x"0c",
          2230 => x"0d",
          2231 => x"0c",
          2232 => x"d4",
          2233 => x"b5",
          2234 => x"3d",
          2235 => x"82",
          2236 => x"fc",
          2237 => x"b5",
          2238 => x"05",
          2239 => x"99",
          2240 => x"d4",
          2241 => x"08",
          2242 => x"d4",
          2243 => x"0c",
          2244 => x"b5",
          2245 => x"05",
          2246 => x"d4",
          2247 => x"08",
          2248 => x"38",
          2249 => x"08",
          2250 => x"30",
          2251 => x"08",
          2252 => x"81",
          2253 => x"d4",
          2254 => x"08",
          2255 => x"d4",
          2256 => x"08",
          2257 => x"3f",
          2258 => x"08",
          2259 => x"d4",
          2260 => x"0c",
          2261 => x"d4",
          2262 => x"08",
          2263 => x"38",
          2264 => x"08",
          2265 => x"30",
          2266 => x"08",
          2267 => x"82",
          2268 => x"f8",
          2269 => x"82",
          2270 => x"54",
          2271 => x"82",
          2272 => x"04",
          2273 => x"08",
          2274 => x"d4",
          2275 => x"0d",
          2276 => x"b5",
          2277 => x"05",
          2278 => x"b5",
          2279 => x"05",
          2280 => x"c5",
          2281 => x"c8",
          2282 => x"b5",
          2283 => x"85",
          2284 => x"b5",
          2285 => x"82",
          2286 => x"02",
          2287 => x"0c",
          2288 => x"81",
          2289 => x"d4",
          2290 => x"08",
          2291 => x"d4",
          2292 => x"08",
          2293 => x"82",
          2294 => x"70",
          2295 => x"0c",
          2296 => x"0d",
          2297 => x"0c",
          2298 => x"d4",
          2299 => x"b5",
          2300 => x"3d",
          2301 => x"82",
          2302 => x"fc",
          2303 => x"0b",
          2304 => x"08",
          2305 => x"82",
          2306 => x"8c",
          2307 => x"b5",
          2308 => x"05",
          2309 => x"38",
          2310 => x"08",
          2311 => x"80",
          2312 => x"80",
          2313 => x"d4",
          2314 => x"08",
          2315 => x"82",
          2316 => x"8c",
          2317 => x"82",
          2318 => x"8c",
          2319 => x"b5",
          2320 => x"05",
          2321 => x"b5",
          2322 => x"05",
          2323 => x"39",
          2324 => x"08",
          2325 => x"80",
          2326 => x"38",
          2327 => x"08",
          2328 => x"82",
          2329 => x"88",
          2330 => x"ad",
          2331 => x"d4",
          2332 => x"08",
          2333 => x"08",
          2334 => x"31",
          2335 => x"08",
          2336 => x"82",
          2337 => x"f8",
          2338 => x"b5",
          2339 => x"05",
          2340 => x"b5",
          2341 => x"05",
          2342 => x"d4",
          2343 => x"08",
          2344 => x"b5",
          2345 => x"05",
          2346 => x"d4",
          2347 => x"08",
          2348 => x"b5",
          2349 => x"05",
          2350 => x"39",
          2351 => x"08",
          2352 => x"80",
          2353 => x"82",
          2354 => x"88",
          2355 => x"82",
          2356 => x"f4",
          2357 => x"91",
          2358 => x"d4",
          2359 => x"08",
          2360 => x"d4",
          2361 => x"0c",
          2362 => x"d4",
          2363 => x"08",
          2364 => x"0c",
          2365 => x"82",
          2366 => x"04",
          2367 => x"08",
          2368 => x"d4",
          2369 => x"0d",
          2370 => x"b5",
          2371 => x"05",
          2372 => x"d4",
          2373 => x"08",
          2374 => x"0c",
          2375 => x"08",
          2376 => x"70",
          2377 => x"72",
          2378 => x"82",
          2379 => x"f8",
          2380 => x"81",
          2381 => x"72",
          2382 => x"81",
          2383 => x"82",
          2384 => x"88",
          2385 => x"08",
          2386 => x"0c",
          2387 => x"82",
          2388 => x"f8",
          2389 => x"72",
          2390 => x"81",
          2391 => x"81",
          2392 => x"d4",
          2393 => x"34",
          2394 => x"08",
          2395 => x"70",
          2396 => x"71",
          2397 => x"51",
          2398 => x"82",
          2399 => x"f8",
          2400 => x"b5",
          2401 => x"05",
          2402 => x"b0",
          2403 => x"06",
          2404 => x"82",
          2405 => x"88",
          2406 => x"08",
          2407 => x"0c",
          2408 => x"53",
          2409 => x"b5",
          2410 => x"05",
          2411 => x"d4",
          2412 => x"33",
          2413 => x"08",
          2414 => x"82",
          2415 => x"e8",
          2416 => x"e2",
          2417 => x"82",
          2418 => x"e8",
          2419 => x"f8",
          2420 => x"80",
          2421 => x"0b",
          2422 => x"08",
          2423 => x"82",
          2424 => x"88",
          2425 => x"08",
          2426 => x"0c",
          2427 => x"53",
          2428 => x"b5",
          2429 => x"05",
          2430 => x"39",
          2431 => x"b5",
          2432 => x"05",
          2433 => x"d4",
          2434 => x"08",
          2435 => x"05",
          2436 => x"08",
          2437 => x"33",
          2438 => x"08",
          2439 => x"80",
          2440 => x"b5",
          2441 => x"05",
          2442 => x"a0",
          2443 => x"81",
          2444 => x"d4",
          2445 => x"0c",
          2446 => x"82",
          2447 => x"f8",
          2448 => x"af",
          2449 => x"38",
          2450 => x"08",
          2451 => x"53",
          2452 => x"83",
          2453 => x"80",
          2454 => x"d4",
          2455 => x"0c",
          2456 => x"88",
          2457 => x"d4",
          2458 => x"34",
          2459 => x"b5",
          2460 => x"05",
          2461 => x"73",
          2462 => x"82",
          2463 => x"f8",
          2464 => x"72",
          2465 => x"38",
          2466 => x"0b",
          2467 => x"08",
          2468 => x"82",
          2469 => x"0b",
          2470 => x"08",
          2471 => x"80",
          2472 => x"d4",
          2473 => x"0c",
          2474 => x"08",
          2475 => x"53",
          2476 => x"81",
          2477 => x"b5",
          2478 => x"05",
          2479 => x"e0",
          2480 => x"38",
          2481 => x"08",
          2482 => x"e0",
          2483 => x"72",
          2484 => x"08",
          2485 => x"82",
          2486 => x"f8",
          2487 => x"11",
          2488 => x"82",
          2489 => x"f8",
          2490 => x"b5",
          2491 => x"05",
          2492 => x"73",
          2493 => x"82",
          2494 => x"f8",
          2495 => x"11",
          2496 => x"82",
          2497 => x"f8",
          2498 => x"b5",
          2499 => x"05",
          2500 => x"89",
          2501 => x"80",
          2502 => x"d4",
          2503 => x"0c",
          2504 => x"82",
          2505 => x"f8",
          2506 => x"b5",
          2507 => x"05",
          2508 => x"72",
          2509 => x"38",
          2510 => x"b5",
          2511 => x"05",
          2512 => x"39",
          2513 => x"08",
          2514 => x"70",
          2515 => x"08",
          2516 => x"29",
          2517 => x"08",
          2518 => x"70",
          2519 => x"d4",
          2520 => x"0c",
          2521 => x"08",
          2522 => x"70",
          2523 => x"71",
          2524 => x"51",
          2525 => x"53",
          2526 => x"b5",
          2527 => x"05",
          2528 => x"39",
          2529 => x"08",
          2530 => x"53",
          2531 => x"90",
          2532 => x"d4",
          2533 => x"08",
          2534 => x"d4",
          2535 => x"0c",
          2536 => x"08",
          2537 => x"82",
          2538 => x"fc",
          2539 => x"0c",
          2540 => x"82",
          2541 => x"ec",
          2542 => x"b5",
          2543 => x"05",
          2544 => x"c8",
          2545 => x"0d",
          2546 => x"0c",
          2547 => x"d4",
          2548 => x"b5",
          2549 => x"3d",
          2550 => x"82",
          2551 => x"f0",
          2552 => x"b5",
          2553 => x"05",
          2554 => x"73",
          2555 => x"d4",
          2556 => x"08",
          2557 => x"53",
          2558 => x"72",
          2559 => x"08",
          2560 => x"72",
          2561 => x"53",
          2562 => x"09",
          2563 => x"38",
          2564 => x"08",
          2565 => x"70",
          2566 => x"71",
          2567 => x"39",
          2568 => x"08",
          2569 => x"53",
          2570 => x"09",
          2571 => x"38",
          2572 => x"b5",
          2573 => x"05",
          2574 => x"d4",
          2575 => x"08",
          2576 => x"05",
          2577 => x"08",
          2578 => x"33",
          2579 => x"08",
          2580 => x"82",
          2581 => x"f8",
          2582 => x"72",
          2583 => x"81",
          2584 => x"38",
          2585 => x"08",
          2586 => x"70",
          2587 => x"71",
          2588 => x"51",
          2589 => x"82",
          2590 => x"f8",
          2591 => x"b5",
          2592 => x"05",
          2593 => x"d4",
          2594 => x"0c",
          2595 => x"08",
          2596 => x"80",
          2597 => x"38",
          2598 => x"08",
          2599 => x"80",
          2600 => x"38",
          2601 => x"90",
          2602 => x"d4",
          2603 => x"34",
          2604 => x"08",
          2605 => x"70",
          2606 => x"71",
          2607 => x"51",
          2608 => x"82",
          2609 => x"f8",
          2610 => x"a4",
          2611 => x"82",
          2612 => x"f4",
          2613 => x"b5",
          2614 => x"05",
          2615 => x"81",
          2616 => x"70",
          2617 => x"72",
          2618 => x"d4",
          2619 => x"34",
          2620 => x"82",
          2621 => x"f8",
          2622 => x"72",
          2623 => x"38",
          2624 => x"b5",
          2625 => x"05",
          2626 => x"39",
          2627 => x"08",
          2628 => x"53",
          2629 => x"90",
          2630 => x"d4",
          2631 => x"33",
          2632 => x"26",
          2633 => x"39",
          2634 => x"b5",
          2635 => x"05",
          2636 => x"39",
          2637 => x"b5",
          2638 => x"05",
          2639 => x"82",
          2640 => x"f8",
          2641 => x"af",
          2642 => x"38",
          2643 => x"08",
          2644 => x"53",
          2645 => x"83",
          2646 => x"80",
          2647 => x"d4",
          2648 => x"0c",
          2649 => x"8a",
          2650 => x"d4",
          2651 => x"34",
          2652 => x"b5",
          2653 => x"05",
          2654 => x"d4",
          2655 => x"33",
          2656 => x"27",
          2657 => x"82",
          2658 => x"f8",
          2659 => x"80",
          2660 => x"94",
          2661 => x"d4",
          2662 => x"33",
          2663 => x"53",
          2664 => x"d4",
          2665 => x"34",
          2666 => x"08",
          2667 => x"d0",
          2668 => x"72",
          2669 => x"08",
          2670 => x"82",
          2671 => x"f8",
          2672 => x"90",
          2673 => x"38",
          2674 => x"08",
          2675 => x"f9",
          2676 => x"72",
          2677 => x"08",
          2678 => x"82",
          2679 => x"f8",
          2680 => x"72",
          2681 => x"38",
          2682 => x"b5",
          2683 => x"05",
          2684 => x"39",
          2685 => x"08",
          2686 => x"82",
          2687 => x"f4",
          2688 => x"54",
          2689 => x"8d",
          2690 => x"82",
          2691 => x"ec",
          2692 => x"f7",
          2693 => x"d4",
          2694 => x"33",
          2695 => x"d4",
          2696 => x"08",
          2697 => x"d4",
          2698 => x"33",
          2699 => x"b5",
          2700 => x"05",
          2701 => x"d4",
          2702 => x"08",
          2703 => x"05",
          2704 => x"08",
          2705 => x"55",
          2706 => x"82",
          2707 => x"f8",
          2708 => x"a5",
          2709 => x"d4",
          2710 => x"33",
          2711 => x"2e",
          2712 => x"b5",
          2713 => x"05",
          2714 => x"b5",
          2715 => x"05",
          2716 => x"d4",
          2717 => x"08",
          2718 => x"08",
          2719 => x"71",
          2720 => x"0b",
          2721 => x"08",
          2722 => x"82",
          2723 => x"ec",
          2724 => x"b5",
          2725 => x"3d",
          2726 => x"d4",
          2727 => x"3d",
          2728 => x"08",
          2729 => x"58",
          2730 => x"80",
          2731 => x"39",
          2732 => x"e6",
          2733 => x"b5",
          2734 => x"78",
          2735 => x"33",
          2736 => x"39",
          2737 => x"73",
          2738 => x"81",
          2739 => x"81",
          2740 => x"39",
          2741 => x"90",
          2742 => x"c8",
          2743 => x"52",
          2744 => x"3f",
          2745 => x"08",
          2746 => x"75",
          2747 => x"a3",
          2748 => x"c8",
          2749 => x"84",
          2750 => x"73",
          2751 => x"b0",
          2752 => x"70",
          2753 => x"58",
          2754 => x"27",
          2755 => x"54",
          2756 => x"c8",
          2757 => x"0d",
          2758 => x"0d",
          2759 => x"93",
          2760 => x"38",
          2761 => x"82",
          2762 => x"52",
          2763 => x"82",
          2764 => x"81",
          2765 => x"9b",
          2766 => x"f9",
          2767 => x"90",
          2768 => x"39",
          2769 => x"51",
          2770 => x"82",
          2771 => x"80",
          2772 => x"9b",
          2773 => x"dd",
          2774 => x"d4",
          2775 => x"39",
          2776 => x"51",
          2777 => x"82",
          2778 => x"80",
          2779 => x"9c",
          2780 => x"c1",
          2781 => x"ac",
          2782 => x"82",
          2783 => x"b5",
          2784 => x"dc",
          2785 => x"82",
          2786 => x"a9",
          2787 => x"94",
          2788 => x"82",
          2789 => x"9d",
          2790 => x"c4",
          2791 => x"82",
          2792 => x"91",
          2793 => x"f4",
          2794 => x"82",
          2795 => x"85",
          2796 => x"98",
          2797 => x"3f",
          2798 => x"04",
          2799 => x"77",
          2800 => x"74",
          2801 => x"8a",
          2802 => x"75",
          2803 => x"51",
          2804 => x"e8",
          2805 => x"ef",
          2806 => x"b5",
          2807 => x"75",
          2808 => x"3f",
          2809 => x"08",
          2810 => x"75",
          2811 => x"a8",
          2812 => x"e5",
          2813 => x"0d",
          2814 => x"0d",
          2815 => x"05",
          2816 => x"33",
          2817 => x"68",
          2818 => x"7a",
          2819 => x"51",
          2820 => x"78",
          2821 => x"ff",
          2822 => x"81",
          2823 => x"07",
          2824 => x"06",
          2825 => x"56",
          2826 => x"38",
          2827 => x"52",
          2828 => x"52",
          2829 => x"c5",
          2830 => x"c8",
          2831 => x"b5",
          2832 => x"38",
          2833 => x"08",
          2834 => x"88",
          2835 => x"c8",
          2836 => x"3d",
          2837 => x"84",
          2838 => x"52",
          2839 => x"84",
          2840 => x"b5",
          2841 => x"82",
          2842 => x"90",
          2843 => x"74",
          2844 => x"38",
          2845 => x"19",
          2846 => x"39",
          2847 => x"05",
          2848 => x"ea",
          2849 => x"70",
          2850 => x"25",
          2851 => x"9f",
          2852 => x"51",
          2853 => x"74",
          2854 => x"38",
          2855 => x"53",
          2856 => x"88",
          2857 => x"51",
          2858 => x"76",
          2859 => x"b5",
          2860 => x"3d",
          2861 => x"3d",
          2862 => x"84",
          2863 => x"33",
          2864 => x"58",
          2865 => x"52",
          2866 => x"ad",
          2867 => x"c8",
          2868 => x"76",
          2869 => x"38",
          2870 => x"9c",
          2871 => x"82",
          2872 => x"61",
          2873 => x"82",
          2874 => x"7f",
          2875 => x"78",
          2876 => x"c8",
          2877 => x"39",
          2878 => x"82",
          2879 => x"8a",
          2880 => x"f3",
          2881 => x"61",
          2882 => x"05",
          2883 => x"33",
          2884 => x"68",
          2885 => x"5c",
          2886 => x"7a",
          2887 => x"d4",
          2888 => x"b5",
          2889 => x"dc",
          2890 => x"ad",
          2891 => x"74",
          2892 => x"80",
          2893 => x"2e",
          2894 => x"a0",
          2895 => x"80",
          2896 => x"18",
          2897 => x"27",
          2898 => x"22",
          2899 => x"e0",
          2900 => x"85",
          2901 => x"82",
          2902 => x"ff",
          2903 => x"82",
          2904 => x"c3",
          2905 => x"53",
          2906 => x"8e",
          2907 => x"52",
          2908 => x"51",
          2909 => x"3f",
          2910 => x"9e",
          2911 => x"b8",
          2912 => x"15",
          2913 => x"74",
          2914 => x"7a",
          2915 => x"72",
          2916 => x"9e",
          2917 => x"b8",
          2918 => x"39",
          2919 => x"51",
          2920 => x"3f",
          2921 => x"82",
          2922 => x"52",
          2923 => x"83",
          2924 => x"39",
          2925 => x"51",
          2926 => x"3f",
          2927 => x"79",
          2928 => x"38",
          2929 => x"33",
          2930 => x"56",
          2931 => x"83",
          2932 => x"80",
          2933 => x"27",
          2934 => x"53",
          2935 => x"70",
          2936 => x"51",
          2937 => x"2e",
          2938 => x"80",
          2939 => x"38",
          2940 => x"08",
          2941 => x"88",
          2942 => x"9c",
          2943 => x"51",
          2944 => x"81",
          2945 => x"b6",
          2946 => x"84",
          2947 => x"3f",
          2948 => x"1c",
          2949 => x"cb",
          2950 => x"c8",
          2951 => x"70",
          2952 => x"57",
          2953 => x"09",
          2954 => x"38",
          2955 => x"82",
          2956 => x"98",
          2957 => x"2c",
          2958 => x"70",
          2959 => x"32",
          2960 => x"72",
          2961 => x"07",
          2962 => x"58",
          2963 => x"57",
          2964 => x"d8",
          2965 => x"2e",
          2966 => x"85",
          2967 => x"8c",
          2968 => x"53",
          2969 => x"fd",
          2970 => x"53",
          2971 => x"c8",
          2972 => x"0d",
          2973 => x"0d",
          2974 => x"33",
          2975 => x"53",
          2976 => x"52",
          2977 => x"d1",
          2978 => x"a0",
          2979 => x"a6",
          2980 => x"98",
          2981 => x"a4",
          2982 => x"a1",
          2983 => x"9f",
          2984 => x"b6",
          2985 => x"80",
          2986 => x"a0",
          2987 => x"3d",
          2988 => x"3d",
          2989 => x"96",
          2990 => x"a5",
          2991 => x"51",
          2992 => x"82",
          2993 => x"99",
          2994 => x"51",
          2995 => x"72",
          2996 => x"81",
          2997 => x"71",
          2998 => x"38",
          2999 => x"f0",
          3000 => x"e0",
          3001 => x"3f",
          3002 => x"e4",
          3003 => x"2a",
          3004 => x"51",
          3005 => x"2e",
          3006 => x"51",
          3007 => x"82",
          3008 => x"98",
          3009 => x"51",
          3010 => x"72",
          3011 => x"81",
          3012 => x"71",
          3013 => x"38",
          3014 => x"b4",
          3015 => x"80",
          3016 => x"3f",
          3017 => x"a8",
          3018 => x"2a",
          3019 => x"51",
          3020 => x"2e",
          3021 => x"51",
          3022 => x"82",
          3023 => x"98",
          3024 => x"51",
          3025 => x"72",
          3026 => x"81",
          3027 => x"71",
          3028 => x"38",
          3029 => x"f8",
          3030 => x"a8",
          3031 => x"3f",
          3032 => x"ec",
          3033 => x"2a",
          3034 => x"51",
          3035 => x"2e",
          3036 => x"51",
          3037 => x"82",
          3038 => x"97",
          3039 => x"51",
          3040 => x"72",
          3041 => x"81",
          3042 => x"71",
          3043 => x"38",
          3044 => x"bc",
          3045 => x"d0",
          3046 => x"3f",
          3047 => x"b0",
          3048 => x"2a",
          3049 => x"51",
          3050 => x"2e",
          3051 => x"51",
          3052 => x"82",
          3053 => x"97",
          3054 => x"51",
          3055 => x"a3",
          3056 => x"3d",
          3057 => x"3d",
          3058 => x"84",
          3059 => x"33",
          3060 => x"56",
          3061 => x"51",
          3062 => x"0b",
          3063 => x"c4",
          3064 => x"a9",
          3065 => x"82",
          3066 => x"82",
          3067 => x"80",
          3068 => x"82",
          3069 => x"30",
          3070 => x"c8",
          3071 => x"25",
          3072 => x"51",
          3073 => x"0b",
          3074 => x"c4",
          3075 => x"82",
          3076 => x"54",
          3077 => x"09",
          3078 => x"38",
          3079 => x"53",
          3080 => x"51",
          3081 => x"3f",
          3082 => x"08",
          3083 => x"38",
          3084 => x"08",
          3085 => x"3f",
          3086 => x"cc",
          3087 => x"84",
          3088 => x"0b",
          3089 => x"b0",
          3090 => x"0b",
          3091 => x"33",
          3092 => x"2e",
          3093 => x"8c",
          3094 => x"b0",
          3095 => x"75",
          3096 => x"3f",
          3097 => x"b5",
          3098 => x"3d",
          3099 => x"3d",
          3100 => x"71",
          3101 => x"0c",
          3102 => x"52",
          3103 => x"c6",
          3104 => x"b5",
          3105 => x"ff",
          3106 => x"7d",
          3107 => x"06",
          3108 => x"3d",
          3109 => x"82",
          3110 => x"78",
          3111 => x"3f",
          3112 => x"52",
          3113 => x"51",
          3114 => x"3f",
          3115 => x"08",
          3116 => x"38",
          3117 => x"51",
          3118 => x"81",
          3119 => x"82",
          3120 => x"ff",
          3121 => x"96",
          3122 => x"5a",
          3123 => x"79",
          3124 => x"3f",
          3125 => x"84",
          3126 => x"c2",
          3127 => x"c8",
          3128 => x"70",
          3129 => x"59",
          3130 => x"2e",
          3131 => x"78",
          3132 => x"b2",
          3133 => x"2e",
          3134 => x"78",
          3135 => x"38",
          3136 => x"ff",
          3137 => x"bc",
          3138 => x"38",
          3139 => x"78",
          3140 => x"83",
          3141 => x"80",
          3142 => x"cd",
          3143 => x"2e",
          3144 => x"8a",
          3145 => x"80",
          3146 => x"d9",
          3147 => x"f9",
          3148 => x"78",
          3149 => x"88",
          3150 => x"80",
          3151 => x"a1",
          3152 => x"39",
          3153 => x"2e",
          3154 => x"78",
          3155 => x"8b",
          3156 => x"82",
          3157 => x"38",
          3158 => x"78",
          3159 => x"89",
          3160 => x"fe",
          3161 => x"ff",
          3162 => x"ff",
          3163 => x"ec",
          3164 => x"b5",
          3165 => x"2e",
          3166 => x"b4",
          3167 => x"11",
          3168 => x"05",
          3169 => x"3f",
          3170 => x"08",
          3171 => x"af",
          3172 => x"fe",
          3173 => x"ff",
          3174 => x"ec",
          3175 => x"b5",
          3176 => x"38",
          3177 => x"08",
          3178 => x"f8",
          3179 => x"a9",
          3180 => x"5c",
          3181 => x"27",
          3182 => x"61",
          3183 => x"70",
          3184 => x"0c",
          3185 => x"f5",
          3186 => x"39",
          3187 => x"80",
          3188 => x"84",
          3189 => x"f5",
          3190 => x"c8",
          3191 => x"fd",
          3192 => x"3d",
          3193 => x"53",
          3194 => x"51",
          3195 => x"82",
          3196 => x"80",
          3197 => x"38",
          3198 => x"f8",
          3199 => x"84",
          3200 => x"c9",
          3201 => x"c8",
          3202 => x"fd",
          3203 => x"a2",
          3204 => x"af",
          3205 => x"5a",
          3206 => x"81",
          3207 => x"59",
          3208 => x"05",
          3209 => x"34",
          3210 => x"42",
          3211 => x"3d",
          3212 => x"53",
          3213 => x"51",
          3214 => x"82",
          3215 => x"80",
          3216 => x"38",
          3217 => x"fc",
          3218 => x"84",
          3219 => x"fd",
          3220 => x"c8",
          3221 => x"fc",
          3222 => x"3d",
          3223 => x"53",
          3224 => x"51",
          3225 => x"82",
          3226 => x"80",
          3227 => x"38",
          3228 => x"51",
          3229 => x"3f",
          3230 => x"63",
          3231 => x"61",
          3232 => x"33",
          3233 => x"78",
          3234 => x"38",
          3235 => x"54",
          3236 => x"79",
          3237 => x"a4",
          3238 => x"bd",
          3239 => x"62",
          3240 => x"5a",
          3241 => x"51",
          3242 => x"fc",
          3243 => x"3d",
          3244 => x"53",
          3245 => x"51",
          3246 => x"82",
          3247 => x"80",
          3248 => x"b4",
          3249 => x"78",
          3250 => x"38",
          3251 => x"08",
          3252 => x"39",
          3253 => x"33",
          3254 => x"2e",
          3255 => x"b3",
          3256 => x"bc",
          3257 => x"b6",
          3258 => x"80",
          3259 => x"82",
          3260 => x"44",
          3261 => x"b4",
          3262 => x"78",
          3263 => x"38",
          3264 => x"08",
          3265 => x"82",
          3266 => x"59",
          3267 => x"88",
          3268 => x"8c",
          3269 => x"39",
          3270 => x"08",
          3271 => x"44",
          3272 => x"fc",
          3273 => x"84",
          3274 => x"a1",
          3275 => x"c8",
          3276 => x"38",
          3277 => x"33",
          3278 => x"2e",
          3279 => x"b3",
          3280 => x"80",
          3281 => x"b4",
          3282 => x"78",
          3283 => x"38",
          3284 => x"08",
          3285 => x"82",
          3286 => x"59",
          3287 => x"88",
          3288 => x"80",
          3289 => x"39",
          3290 => x"33",
          3291 => x"2e",
          3292 => x"b4",
          3293 => x"99",
          3294 => x"b2",
          3295 => x"80",
          3296 => x"82",
          3297 => x"43",
          3298 => x"b4",
          3299 => x"05",
          3300 => x"fe",
          3301 => x"ff",
          3302 => x"e8",
          3303 => x"b5",
          3304 => x"2e",
          3305 => x"62",
          3306 => x"88",
          3307 => x"81",
          3308 => x"32",
          3309 => x"72",
          3310 => x"70",
          3311 => x"51",
          3312 => x"80",
          3313 => x"7a",
          3314 => x"38",
          3315 => x"a2",
          3316 => x"90",
          3317 => x"63",
          3318 => x"62",
          3319 => x"f2",
          3320 => x"a2",
          3321 => x"f5",
          3322 => x"ff",
          3323 => x"ff",
          3324 => x"e7",
          3325 => x"b5",
          3326 => x"2e",
          3327 => x"b4",
          3328 => x"11",
          3329 => x"05",
          3330 => x"3f",
          3331 => x"08",
          3332 => x"38",
          3333 => x"80",
          3334 => x"79",
          3335 => x"05",
          3336 => x"fe",
          3337 => x"ff",
          3338 => x"e7",
          3339 => x"b5",
          3340 => x"38",
          3341 => x"63",
          3342 => x"52",
          3343 => x"51",
          3344 => x"3f",
          3345 => x"08",
          3346 => x"52",
          3347 => x"ab",
          3348 => x"45",
          3349 => x"78",
          3350 => x"e3",
          3351 => x"27",
          3352 => x"3d",
          3353 => x"53",
          3354 => x"51",
          3355 => x"82",
          3356 => x"80",
          3357 => x"63",
          3358 => x"cb",
          3359 => x"34",
          3360 => x"44",
          3361 => x"82",
          3362 => x"c6",
          3363 => x"a7",
          3364 => x"fe",
          3365 => x"ff",
          3366 => x"e0",
          3367 => x"b5",
          3368 => x"2e",
          3369 => x"b4",
          3370 => x"11",
          3371 => x"05",
          3372 => x"3f",
          3373 => x"08",
          3374 => x"38",
          3375 => x"be",
          3376 => x"70",
          3377 => x"23",
          3378 => x"3d",
          3379 => x"53",
          3380 => x"51",
          3381 => x"82",
          3382 => x"e0",
          3383 => x"39",
          3384 => x"54",
          3385 => x"e8",
          3386 => x"ed",
          3387 => x"98",
          3388 => x"f8",
          3389 => x"ff",
          3390 => x"79",
          3391 => x"59",
          3392 => x"f7",
          3393 => x"9f",
          3394 => x"60",
          3395 => x"d0",
          3396 => x"fe",
          3397 => x"ff",
          3398 => x"df",
          3399 => x"b5",
          3400 => x"2e",
          3401 => x"59",
          3402 => x"22",
          3403 => x"05",
          3404 => x"41",
          3405 => x"82",
          3406 => x"c5",
          3407 => x"a0",
          3408 => x"fe",
          3409 => x"ff",
          3410 => x"df",
          3411 => x"b5",
          3412 => x"2e",
          3413 => x"b4",
          3414 => x"11",
          3415 => x"05",
          3416 => x"3f",
          3417 => x"08",
          3418 => x"38",
          3419 => x"0c",
          3420 => x"05",
          3421 => x"fe",
          3422 => x"ff",
          3423 => x"de",
          3424 => x"b5",
          3425 => x"38",
          3426 => x"60",
          3427 => x"52",
          3428 => x"51",
          3429 => x"3f",
          3430 => x"08",
          3431 => x"52",
          3432 => x"a9",
          3433 => x"45",
          3434 => x"78",
          3435 => x"8f",
          3436 => x"27",
          3437 => x"3d",
          3438 => x"53",
          3439 => x"51",
          3440 => x"82",
          3441 => x"80",
          3442 => x"60",
          3443 => x"59",
          3444 => x"41",
          3445 => x"82",
          3446 => x"c4",
          3447 => x"ab",
          3448 => x"ff",
          3449 => x"ff",
          3450 => x"e3",
          3451 => x"b5",
          3452 => x"2e",
          3453 => x"63",
          3454 => x"84",
          3455 => x"d9",
          3456 => x"78",
          3457 => x"ff",
          3458 => x"ff",
          3459 => x"e3",
          3460 => x"b5",
          3461 => x"2e",
          3462 => x"63",
          3463 => x"a0",
          3464 => x"b5",
          3465 => x"78",
          3466 => x"c8",
          3467 => x"f5",
          3468 => x"b5",
          3469 => x"82",
          3470 => x"ff",
          3471 => x"f4",
          3472 => x"a3",
          3473 => x"9c",
          3474 => x"ee",
          3475 => x"39",
          3476 => x"51",
          3477 => x"80",
          3478 => x"39",
          3479 => x"f4",
          3480 => x"45",
          3481 => x"78",
          3482 => x"d3",
          3483 => x"06",
          3484 => x"2e",
          3485 => x"b4",
          3486 => x"05",
          3487 => x"3f",
          3488 => x"08",
          3489 => x"7a",
          3490 => x"38",
          3491 => x"89",
          3492 => x"2e",
          3493 => x"ca",
          3494 => x"2e",
          3495 => x"c2",
          3496 => x"88",
          3497 => x"82",
          3498 => x"80",
          3499 => x"90",
          3500 => x"ff",
          3501 => x"ff",
          3502 => x"b8",
          3503 => x"b4",
          3504 => x"05",
          3505 => x"3f",
          3506 => x"55",
          3507 => x"54",
          3508 => x"a4",
          3509 => x"3d",
          3510 => x"51",
          3511 => x"3f",
          3512 => x"54",
          3513 => x"a4",
          3514 => x"3d",
          3515 => x"51",
          3516 => x"3f",
          3517 => x"58",
          3518 => x"57",
          3519 => x"55",
          3520 => x"d0",
          3521 => x"d0",
          3522 => x"3d",
          3523 => x"51",
          3524 => x"82",
          3525 => x"82",
          3526 => x"09",
          3527 => x"72",
          3528 => x"51",
          3529 => x"80",
          3530 => x"26",
          3531 => x"5a",
          3532 => x"59",
          3533 => x"8d",
          3534 => x"70",
          3535 => x"5c",
          3536 => x"c3",
          3537 => x"32",
          3538 => x"07",
          3539 => x"38",
          3540 => x"09",
          3541 => x"e7",
          3542 => x"b4",
          3543 => x"3f",
          3544 => x"f5",
          3545 => x"0b",
          3546 => x"34",
          3547 => x"8c",
          3548 => x"55",
          3549 => x"52",
          3550 => x"88",
          3551 => x"c8",
          3552 => x"75",
          3553 => x"87",
          3554 => x"73",
          3555 => x"3f",
          3556 => x"c8",
          3557 => x"0c",
          3558 => x"9c",
          3559 => x"55",
          3560 => x"52",
          3561 => x"dc",
          3562 => x"c8",
          3563 => x"75",
          3564 => x"87",
          3565 => x"73",
          3566 => x"3f",
          3567 => x"c8",
          3568 => x"0c",
          3569 => x"0b",
          3570 => x"84",
          3571 => x"83",
          3572 => x"94",
          3573 => x"f5",
          3574 => x"f8",
          3575 => x"02",
          3576 => x"05",
          3577 => x"82",
          3578 => x"87",
          3579 => x"13",
          3580 => x"0c",
          3581 => x"0c",
          3582 => x"3f",
          3583 => x"82",
          3584 => x"ff",
          3585 => x"82",
          3586 => x"ff",
          3587 => x"80",
          3588 => x"92",
          3589 => x"51",
          3590 => x"f0",
          3591 => x"04",
          3592 => x"80",
          3593 => x"71",
          3594 => x"87",
          3595 => x"b5",
          3596 => x"ff",
          3597 => x"ff",
          3598 => x"72",
          3599 => x"38",
          3600 => x"c8",
          3601 => x"0d",
          3602 => x"0d",
          3603 => x"54",
          3604 => x"52",
          3605 => x"2e",
          3606 => x"72",
          3607 => x"a0",
          3608 => x"06",
          3609 => x"13",
          3610 => x"72",
          3611 => x"a2",
          3612 => x"06",
          3613 => x"13",
          3614 => x"72",
          3615 => x"2e",
          3616 => x"9f",
          3617 => x"81",
          3618 => x"72",
          3619 => x"70",
          3620 => x"38",
          3621 => x"80",
          3622 => x"73",
          3623 => x"39",
          3624 => x"80",
          3625 => x"54",
          3626 => x"83",
          3627 => x"70",
          3628 => x"38",
          3629 => x"80",
          3630 => x"54",
          3631 => x"09",
          3632 => x"38",
          3633 => x"a2",
          3634 => x"70",
          3635 => x"07",
          3636 => x"70",
          3637 => x"38",
          3638 => x"81",
          3639 => x"71",
          3640 => x"51",
          3641 => x"c8",
          3642 => x"0d",
          3643 => x"0d",
          3644 => x"08",
          3645 => x"38",
          3646 => x"05",
          3647 => x"d7",
          3648 => x"b5",
          3649 => x"38",
          3650 => x"39",
          3651 => x"82",
          3652 => x"86",
          3653 => x"fc",
          3654 => x"82",
          3655 => x"05",
          3656 => x"52",
          3657 => x"81",
          3658 => x"13",
          3659 => x"51",
          3660 => x"9e",
          3661 => x"38",
          3662 => x"51",
          3663 => x"97",
          3664 => x"38",
          3665 => x"51",
          3666 => x"bb",
          3667 => x"38",
          3668 => x"51",
          3669 => x"bb",
          3670 => x"38",
          3671 => x"55",
          3672 => x"87",
          3673 => x"d9",
          3674 => x"22",
          3675 => x"73",
          3676 => x"80",
          3677 => x"0b",
          3678 => x"9c",
          3679 => x"87",
          3680 => x"0c",
          3681 => x"87",
          3682 => x"0c",
          3683 => x"87",
          3684 => x"0c",
          3685 => x"87",
          3686 => x"0c",
          3687 => x"87",
          3688 => x"0c",
          3689 => x"87",
          3690 => x"0c",
          3691 => x"98",
          3692 => x"87",
          3693 => x"0c",
          3694 => x"c0",
          3695 => x"80",
          3696 => x"b5",
          3697 => x"3d",
          3698 => x"3d",
          3699 => x"87",
          3700 => x"5d",
          3701 => x"87",
          3702 => x"08",
          3703 => x"23",
          3704 => x"b8",
          3705 => x"82",
          3706 => x"c0",
          3707 => x"5a",
          3708 => x"34",
          3709 => x"b0",
          3710 => x"84",
          3711 => x"c0",
          3712 => x"5a",
          3713 => x"34",
          3714 => x"a8",
          3715 => x"86",
          3716 => x"c0",
          3717 => x"5c",
          3718 => x"23",
          3719 => x"a0",
          3720 => x"8a",
          3721 => x"7d",
          3722 => x"ff",
          3723 => x"7b",
          3724 => x"06",
          3725 => x"33",
          3726 => x"33",
          3727 => x"33",
          3728 => x"33",
          3729 => x"33",
          3730 => x"ff",
          3731 => x"82",
          3732 => x"ff",
          3733 => x"8f",
          3734 => x"fb",
          3735 => x"9f",
          3736 => x"b3",
          3737 => x"81",
          3738 => x"55",
          3739 => x"94",
          3740 => x"80",
          3741 => x"87",
          3742 => x"51",
          3743 => x"96",
          3744 => x"06",
          3745 => x"70",
          3746 => x"38",
          3747 => x"70",
          3748 => x"51",
          3749 => x"72",
          3750 => x"81",
          3751 => x"70",
          3752 => x"38",
          3753 => x"70",
          3754 => x"51",
          3755 => x"38",
          3756 => x"06",
          3757 => x"94",
          3758 => x"80",
          3759 => x"87",
          3760 => x"52",
          3761 => x"74",
          3762 => x"0c",
          3763 => x"04",
          3764 => x"02",
          3765 => x"70",
          3766 => x"2a",
          3767 => x"70",
          3768 => x"34",
          3769 => x"04",
          3770 => x"02",
          3771 => x"58",
          3772 => x"09",
          3773 => x"38",
          3774 => x"51",
          3775 => x"b3",
          3776 => x"81",
          3777 => x"56",
          3778 => x"84",
          3779 => x"2e",
          3780 => x"c0",
          3781 => x"72",
          3782 => x"2a",
          3783 => x"55",
          3784 => x"80",
          3785 => x"73",
          3786 => x"81",
          3787 => x"72",
          3788 => x"81",
          3789 => x"06",
          3790 => x"80",
          3791 => x"73",
          3792 => x"81",
          3793 => x"72",
          3794 => x"75",
          3795 => x"53",
          3796 => x"80",
          3797 => x"2e",
          3798 => x"c0",
          3799 => x"77",
          3800 => x"0b",
          3801 => x"0c",
          3802 => x"04",
          3803 => x"79",
          3804 => x"33",
          3805 => x"06",
          3806 => x"70",
          3807 => x"fc",
          3808 => x"ff",
          3809 => x"82",
          3810 => x"70",
          3811 => x"59",
          3812 => x"87",
          3813 => x"51",
          3814 => x"86",
          3815 => x"94",
          3816 => x"08",
          3817 => x"70",
          3818 => x"54",
          3819 => x"2e",
          3820 => x"91",
          3821 => x"06",
          3822 => x"d7",
          3823 => x"32",
          3824 => x"51",
          3825 => x"2e",
          3826 => x"93",
          3827 => x"06",
          3828 => x"ff",
          3829 => x"81",
          3830 => x"87",
          3831 => x"52",
          3832 => x"86",
          3833 => x"94",
          3834 => x"72",
          3835 => x"74",
          3836 => x"ff",
          3837 => x"57",
          3838 => x"38",
          3839 => x"c8",
          3840 => x"0d",
          3841 => x"0d",
          3842 => x"33",
          3843 => x"06",
          3844 => x"c0",
          3845 => x"72",
          3846 => x"38",
          3847 => x"94",
          3848 => x"70",
          3849 => x"81",
          3850 => x"51",
          3851 => x"e2",
          3852 => x"ff",
          3853 => x"c0",
          3854 => x"70",
          3855 => x"38",
          3856 => x"90",
          3857 => x"70",
          3858 => x"82",
          3859 => x"51",
          3860 => x"04",
          3861 => x"82",
          3862 => x"81",
          3863 => x"b5",
          3864 => x"fe",
          3865 => x"b3",
          3866 => x"81",
          3867 => x"53",
          3868 => x"84",
          3869 => x"2e",
          3870 => x"c0",
          3871 => x"71",
          3872 => x"2a",
          3873 => x"51",
          3874 => x"52",
          3875 => x"a0",
          3876 => x"ff",
          3877 => x"c0",
          3878 => x"70",
          3879 => x"38",
          3880 => x"90",
          3881 => x"70",
          3882 => x"98",
          3883 => x"51",
          3884 => x"c8",
          3885 => x"0d",
          3886 => x"0d",
          3887 => x"80",
          3888 => x"2a",
          3889 => x"51",
          3890 => x"84",
          3891 => x"c0",
          3892 => x"82",
          3893 => x"87",
          3894 => x"08",
          3895 => x"0c",
          3896 => x"94",
          3897 => x"f4",
          3898 => x"9e",
          3899 => x"b3",
          3900 => x"c0",
          3901 => x"82",
          3902 => x"87",
          3903 => x"08",
          3904 => x"0c",
          3905 => x"ac",
          3906 => x"84",
          3907 => x"9e",
          3908 => x"b4",
          3909 => x"c0",
          3910 => x"82",
          3911 => x"87",
          3912 => x"08",
          3913 => x"0c",
          3914 => x"bc",
          3915 => x"94",
          3916 => x"9e",
          3917 => x"b4",
          3918 => x"c0",
          3919 => x"82",
          3920 => x"87",
          3921 => x"08",
          3922 => x"b4",
          3923 => x"c0",
          3924 => x"82",
          3925 => x"87",
          3926 => x"08",
          3927 => x"0c",
          3928 => x"8c",
          3929 => x"ac",
          3930 => x"82",
          3931 => x"80",
          3932 => x"9e",
          3933 => x"84",
          3934 => x"51",
          3935 => x"80",
          3936 => x"81",
          3937 => x"b4",
          3938 => x"0b",
          3939 => x"90",
          3940 => x"80",
          3941 => x"52",
          3942 => x"2e",
          3943 => x"52",
          3944 => x"b2",
          3945 => x"87",
          3946 => x"08",
          3947 => x"0a",
          3948 => x"52",
          3949 => x"83",
          3950 => x"71",
          3951 => x"34",
          3952 => x"c0",
          3953 => x"70",
          3954 => x"06",
          3955 => x"70",
          3956 => x"38",
          3957 => x"82",
          3958 => x"80",
          3959 => x"9e",
          3960 => x"a0",
          3961 => x"51",
          3962 => x"80",
          3963 => x"81",
          3964 => x"b4",
          3965 => x"0b",
          3966 => x"90",
          3967 => x"80",
          3968 => x"52",
          3969 => x"2e",
          3970 => x"52",
          3971 => x"b6",
          3972 => x"87",
          3973 => x"08",
          3974 => x"80",
          3975 => x"52",
          3976 => x"83",
          3977 => x"71",
          3978 => x"34",
          3979 => x"c0",
          3980 => x"70",
          3981 => x"06",
          3982 => x"70",
          3983 => x"38",
          3984 => x"82",
          3985 => x"80",
          3986 => x"9e",
          3987 => x"81",
          3988 => x"51",
          3989 => x"80",
          3990 => x"81",
          3991 => x"b4",
          3992 => x"0b",
          3993 => x"90",
          3994 => x"c0",
          3995 => x"52",
          3996 => x"2e",
          3997 => x"52",
          3998 => x"ba",
          3999 => x"87",
          4000 => x"08",
          4001 => x"06",
          4002 => x"70",
          4003 => x"38",
          4004 => x"82",
          4005 => x"87",
          4006 => x"08",
          4007 => x"06",
          4008 => x"51",
          4009 => x"82",
          4010 => x"80",
          4011 => x"9e",
          4012 => x"84",
          4013 => x"52",
          4014 => x"2e",
          4015 => x"52",
          4016 => x"bd",
          4017 => x"9e",
          4018 => x"83",
          4019 => x"84",
          4020 => x"51",
          4021 => x"be",
          4022 => x"87",
          4023 => x"08",
          4024 => x"51",
          4025 => x"80",
          4026 => x"81",
          4027 => x"b4",
          4028 => x"c0",
          4029 => x"70",
          4030 => x"51",
          4031 => x"c0",
          4032 => x"0d",
          4033 => x"0d",
          4034 => x"51",
          4035 => x"3f",
          4036 => x"33",
          4037 => x"2e",
          4038 => x"a5",
          4039 => x"b1",
          4040 => x"a5",
          4041 => x"b1",
          4042 => x"b4",
          4043 => x"73",
          4044 => x"38",
          4045 => x"08",
          4046 => x"08",
          4047 => x"82",
          4048 => x"ff",
          4049 => x"82",
          4050 => x"54",
          4051 => x"94",
          4052 => x"84",
          4053 => x"88",
          4054 => x"52",
          4055 => x"51",
          4056 => x"3f",
          4057 => x"33",
          4058 => x"2e",
          4059 => x"b3",
          4060 => x"b3",
          4061 => x"54",
          4062 => x"f8",
          4063 => x"d9",
          4064 => x"b5",
          4065 => x"80",
          4066 => x"82",
          4067 => x"82",
          4068 => x"11",
          4069 => x"a6",
          4070 => x"94",
          4071 => x"b4",
          4072 => x"73",
          4073 => x"38",
          4074 => x"08",
          4075 => x"08",
          4076 => x"82",
          4077 => x"ff",
          4078 => x"82",
          4079 => x"54",
          4080 => x"8e",
          4081 => x"bc",
          4082 => x"a6",
          4083 => x"94",
          4084 => x"b4",
          4085 => x"73",
          4086 => x"38",
          4087 => x"33",
          4088 => x"ec",
          4089 => x"f1",
          4090 => x"bd",
          4091 => x"80",
          4092 => x"82",
          4093 => x"52",
          4094 => x"51",
          4095 => x"3f",
          4096 => x"33",
          4097 => x"2e",
          4098 => x"a7",
          4099 => x"af",
          4100 => x"b4",
          4101 => x"73",
          4102 => x"38",
          4103 => x"51",
          4104 => x"3f",
          4105 => x"33",
          4106 => x"2e",
          4107 => x"a7",
          4108 => x"af",
          4109 => x"b4",
          4110 => x"73",
          4111 => x"38",
          4112 => x"51",
          4113 => x"3f",
          4114 => x"33",
          4115 => x"2e",
          4116 => x"a7",
          4117 => x"af",
          4118 => x"a7",
          4119 => x"af",
          4120 => x"b4",
          4121 => x"82",
          4122 => x"ff",
          4123 => x"82",
          4124 => x"52",
          4125 => x"51",
          4126 => x"3f",
          4127 => x"08",
          4128 => x"cc",
          4129 => x"d1",
          4130 => x"f4",
          4131 => x"d4",
          4132 => x"a0",
          4133 => x"a8",
          4134 => x"92",
          4135 => x"b4",
          4136 => x"bd",
          4137 => x"75",
          4138 => x"3f",
          4139 => x"08",
          4140 => x"29",
          4141 => x"54",
          4142 => x"c8",
          4143 => x"a9",
          4144 => x"92",
          4145 => x"b4",
          4146 => x"73",
          4147 => x"38",
          4148 => x"08",
          4149 => x"c0",
          4150 => x"c5",
          4151 => x"b5",
          4152 => x"84",
          4153 => x"71",
          4154 => x"82",
          4155 => x"52",
          4156 => x"51",
          4157 => x"3f",
          4158 => x"33",
          4159 => x"2e",
          4160 => x"b4",
          4161 => x"bd",
          4162 => x"75",
          4163 => x"3f",
          4164 => x"08",
          4165 => x"29",
          4166 => x"54",
          4167 => x"c8",
          4168 => x"a9",
          4169 => x"91",
          4170 => x"a2",
          4171 => x"ad",
          4172 => x"3d",
          4173 => x"3d",
          4174 => x"05",
          4175 => x"52",
          4176 => x"aa",
          4177 => x"29",
          4178 => x"05",
          4179 => x"04",
          4180 => x"51",
          4181 => x"aa",
          4182 => x"39",
          4183 => x"51",
          4184 => x"aa",
          4185 => x"39",
          4186 => x"51",
          4187 => x"aa",
          4188 => x"ac",
          4189 => x"3d",
          4190 => x"88",
          4191 => x"80",
          4192 => x"96",
          4193 => x"82",
          4194 => x"87",
          4195 => x"0c",
          4196 => x"0d",
          4197 => x"70",
          4198 => x"98",
          4199 => x"2c",
          4200 => x"70",
          4201 => x"53",
          4202 => x"51",
          4203 => x"aa",
          4204 => x"55",
          4205 => x"25",
          4206 => x"aa",
          4207 => x"12",
          4208 => x"97",
          4209 => x"33",
          4210 => x"70",
          4211 => x"81",
          4212 => x"81",
          4213 => x"b5",
          4214 => x"3d",
          4215 => x"3d",
          4216 => x"84",
          4217 => x"33",
          4218 => x"56",
          4219 => x"2e",
          4220 => x"cd",
          4221 => x"88",
          4222 => x"b7",
          4223 => x"9c",
          4224 => x"51",
          4225 => x"3f",
          4226 => x"08",
          4227 => x"ff",
          4228 => x"73",
          4229 => x"53",
          4230 => x"72",
          4231 => x"53",
          4232 => x"51",
          4233 => x"3f",
          4234 => x"87",
          4235 => x"f6",
          4236 => x"02",
          4237 => x"05",
          4238 => x"05",
          4239 => x"82",
          4240 => x"70",
          4241 => x"b4",
          4242 => x"08",
          4243 => x"5a",
          4244 => x"80",
          4245 => x"74",
          4246 => x"3f",
          4247 => x"33",
          4248 => x"82",
          4249 => x"81",
          4250 => x"58",
          4251 => x"fb",
          4252 => x"c8",
          4253 => x"82",
          4254 => x"70",
          4255 => x"b4",
          4256 => x"08",
          4257 => x"74",
          4258 => x"38",
          4259 => x"52",
          4260 => x"b8",
          4261 => x"b5",
          4262 => x"05",
          4263 => x"b5",
          4264 => x"81",
          4265 => x"93",
          4266 => x"38",
          4267 => x"b5",
          4268 => x"80",
          4269 => x"82",
          4270 => x"56",
          4271 => x"ac",
          4272 => x"98",
          4273 => x"a4",
          4274 => x"fc",
          4275 => x"53",
          4276 => x"51",
          4277 => x"3f",
          4278 => x"08",
          4279 => x"81",
          4280 => x"82",
          4281 => x"51",
          4282 => x"3f",
          4283 => x"04",
          4284 => x"82",
          4285 => x"93",
          4286 => x"52",
          4287 => x"89",
          4288 => x"99",
          4289 => x"73",
          4290 => x"84",
          4291 => x"73",
          4292 => x"38",
          4293 => x"b5",
          4294 => x"b5",
          4295 => x"71",
          4296 => x"38",
          4297 => x"de",
          4298 => x"b5",
          4299 => x"99",
          4300 => x"0b",
          4301 => x"0c",
          4302 => x"04",
          4303 => x"81",
          4304 => x"82",
          4305 => x"51",
          4306 => x"3f",
          4307 => x"08",
          4308 => x"82",
          4309 => x"53",
          4310 => x"88",
          4311 => x"56",
          4312 => x"3f",
          4313 => x"08",
          4314 => x"38",
          4315 => x"b5",
          4316 => x"b5",
          4317 => x"80",
          4318 => x"c8",
          4319 => x"38",
          4320 => x"08",
          4321 => x"17",
          4322 => x"74",
          4323 => x"76",
          4324 => x"82",
          4325 => x"57",
          4326 => x"3f",
          4327 => x"09",
          4328 => x"af",
          4329 => x"0d",
          4330 => x"0d",
          4331 => x"ad",
          4332 => x"5a",
          4333 => x"58",
          4334 => x"b5",
          4335 => x"80",
          4336 => x"82",
          4337 => x"81",
          4338 => x"0b",
          4339 => x"08",
          4340 => x"f8",
          4341 => x"70",
          4342 => x"8b",
          4343 => x"b5",
          4344 => x"2e",
          4345 => x"51",
          4346 => x"3f",
          4347 => x"08",
          4348 => x"55",
          4349 => x"b5",
          4350 => x"8e",
          4351 => x"c8",
          4352 => x"70",
          4353 => x"80",
          4354 => x"09",
          4355 => x"72",
          4356 => x"51",
          4357 => x"77",
          4358 => x"73",
          4359 => x"82",
          4360 => x"8c",
          4361 => x"51",
          4362 => x"3f",
          4363 => x"08",
          4364 => x"38",
          4365 => x"51",
          4366 => x"3f",
          4367 => x"09",
          4368 => x"38",
          4369 => x"51",
          4370 => x"3f",
          4371 => x"b3",
          4372 => x"3d",
          4373 => x"b5",
          4374 => x"34",
          4375 => x"82",
          4376 => x"a9",
          4377 => x"f6",
          4378 => x"7e",
          4379 => x"72",
          4380 => x"5a",
          4381 => x"2e",
          4382 => x"a2",
          4383 => x"78",
          4384 => x"76",
          4385 => x"81",
          4386 => x"70",
          4387 => x"58",
          4388 => x"2e",
          4389 => x"86",
          4390 => x"26",
          4391 => x"54",
          4392 => x"82",
          4393 => x"70",
          4394 => x"ff",
          4395 => x"82",
          4396 => x"53",
          4397 => x"08",
          4398 => x"d7",
          4399 => x"c8",
          4400 => x"38",
          4401 => x"55",
          4402 => x"88",
          4403 => x"2e",
          4404 => x"39",
          4405 => x"ac",
          4406 => x"5a",
          4407 => x"11",
          4408 => x"51",
          4409 => x"82",
          4410 => x"80",
          4411 => x"ff",
          4412 => x"52",
          4413 => x"b1",
          4414 => x"c8",
          4415 => x"06",
          4416 => x"38",
          4417 => x"39",
          4418 => x"81",
          4419 => x"54",
          4420 => x"ff",
          4421 => x"54",
          4422 => x"c8",
          4423 => x"0d",
          4424 => x"0d",
          4425 => x"b2",
          4426 => x"3d",
          4427 => x"5a",
          4428 => x"3d",
          4429 => x"a0",
          4430 => x"9c",
          4431 => x"73",
          4432 => x"73",
          4433 => x"33",
          4434 => x"83",
          4435 => x"76",
          4436 => x"bc",
          4437 => x"76",
          4438 => x"73",
          4439 => x"ad",
          4440 => x"98",
          4441 => x"b5",
          4442 => x"b5",
          4443 => x"b5",
          4444 => x"2e",
          4445 => x"93",
          4446 => x"82",
          4447 => x"51",
          4448 => x"3f",
          4449 => x"08",
          4450 => x"38",
          4451 => x"51",
          4452 => x"3f",
          4453 => x"82",
          4454 => x"5b",
          4455 => x"08",
          4456 => x"52",
          4457 => x"52",
          4458 => x"b7",
          4459 => x"c8",
          4460 => x"b5",
          4461 => x"2e",
          4462 => x"80",
          4463 => x"b5",
          4464 => x"ff",
          4465 => x"82",
          4466 => x"55",
          4467 => x"b5",
          4468 => x"a9",
          4469 => x"c8",
          4470 => x"70",
          4471 => x"80",
          4472 => x"53",
          4473 => x"06",
          4474 => x"f8",
          4475 => x"1b",
          4476 => x"06",
          4477 => x"7b",
          4478 => x"80",
          4479 => x"2e",
          4480 => x"ff",
          4481 => x"39",
          4482 => x"98",
          4483 => x"38",
          4484 => x"08",
          4485 => x"38",
          4486 => x"8f",
          4487 => x"c3",
          4488 => x"c8",
          4489 => x"70",
          4490 => x"59",
          4491 => x"ee",
          4492 => x"ff",
          4493 => x"f4",
          4494 => x"2b",
          4495 => x"82",
          4496 => x"70",
          4497 => x"97",
          4498 => x"2c",
          4499 => x"29",
          4500 => x"05",
          4501 => x"70",
          4502 => x"51",
          4503 => x"51",
          4504 => x"81",
          4505 => x"2e",
          4506 => x"77",
          4507 => x"38",
          4508 => x"0a",
          4509 => x"0a",
          4510 => x"2c",
          4511 => x"75",
          4512 => x"38",
          4513 => x"52",
          4514 => x"85",
          4515 => x"c8",
          4516 => x"06",
          4517 => x"2e",
          4518 => x"82",
          4519 => x"81",
          4520 => x"74",
          4521 => x"29",
          4522 => x"05",
          4523 => x"70",
          4524 => x"56",
          4525 => x"95",
          4526 => x"76",
          4527 => x"77",
          4528 => x"3f",
          4529 => x"08",
          4530 => x"54",
          4531 => x"d3",
          4532 => x"75",
          4533 => x"ca",
          4534 => x"55",
          4535 => x"f4",
          4536 => x"2b",
          4537 => x"82",
          4538 => x"70",
          4539 => x"98",
          4540 => x"11",
          4541 => x"82",
          4542 => x"33",
          4543 => x"51",
          4544 => x"55",
          4545 => x"09",
          4546 => x"92",
          4547 => x"dc",
          4548 => x"0c",
          4549 => x"cc",
          4550 => x"0b",
          4551 => x"34",
          4552 => x"82",
          4553 => x"75",
          4554 => x"34",
          4555 => x"34",
          4556 => x"7e",
          4557 => x"26",
          4558 => x"73",
          4559 => x"96",
          4560 => x"73",
          4561 => x"cc",
          4562 => x"73",
          4563 => x"cb",
          4564 => x"f8",
          4565 => x"75",
          4566 => x"74",
          4567 => x"98",
          4568 => x"73",
          4569 => x"38",
          4570 => x"73",
          4571 => x"34",
          4572 => x"0a",
          4573 => x"0a",
          4574 => x"2c",
          4575 => x"33",
          4576 => x"df",
          4577 => x"fc",
          4578 => x"56",
          4579 => x"cc",
          4580 => x"1a",
          4581 => x"33",
          4582 => x"cc",
          4583 => x"73",
          4584 => x"38",
          4585 => x"73",
          4586 => x"34",
          4587 => x"33",
          4588 => x"0a",
          4589 => x"0a",
          4590 => x"2c",
          4591 => x"33",
          4592 => x"56",
          4593 => x"a8",
          4594 => x"9c",
          4595 => x"1a",
          4596 => x"54",
          4597 => x"3f",
          4598 => x"0a",
          4599 => x"0a",
          4600 => x"2c",
          4601 => x"33",
          4602 => x"73",
          4603 => x"38",
          4604 => x"33",
          4605 => x"70",
          4606 => x"cc",
          4607 => x"51",
          4608 => x"77",
          4609 => x"38",
          4610 => x"08",
          4611 => x"ff",
          4612 => x"74",
          4613 => x"29",
          4614 => x"05",
          4615 => x"82",
          4616 => x"56",
          4617 => x"75",
          4618 => x"fb",
          4619 => x"7a",
          4620 => x"81",
          4621 => x"cc",
          4622 => x"52",
          4623 => x"51",
          4624 => x"81",
          4625 => x"cc",
          4626 => x"81",
          4627 => x"55",
          4628 => x"fb",
          4629 => x"cc",
          4630 => x"05",
          4631 => x"cc",
          4632 => x"15",
          4633 => x"cc",
          4634 => x"cd",
          4635 => x"88",
          4636 => x"bf",
          4637 => x"fc",
          4638 => x"2b",
          4639 => x"82",
          4640 => x"57",
          4641 => x"74",
          4642 => x"38",
          4643 => x"81",
          4644 => x"34",
          4645 => x"08",
          4646 => x"51",
          4647 => x"3f",
          4648 => x"0a",
          4649 => x"0a",
          4650 => x"2c",
          4651 => x"33",
          4652 => x"75",
          4653 => x"38",
          4654 => x"08",
          4655 => x"ff",
          4656 => x"82",
          4657 => x"70",
          4658 => x"98",
          4659 => x"f8",
          4660 => x"56",
          4661 => x"24",
          4662 => x"82",
          4663 => x"52",
          4664 => x"a1",
          4665 => x"81",
          4666 => x"81",
          4667 => x"70",
          4668 => x"cc",
          4669 => x"51",
          4670 => x"25",
          4671 => x"9b",
          4672 => x"f8",
          4673 => x"54",
          4674 => x"82",
          4675 => x"52",
          4676 => x"a1",
          4677 => x"cc",
          4678 => x"51",
          4679 => x"82",
          4680 => x"81",
          4681 => x"73",
          4682 => x"cc",
          4683 => x"73",
          4684 => x"38",
          4685 => x"52",
          4686 => x"f3",
          4687 => x"80",
          4688 => x"0b",
          4689 => x"34",
          4690 => x"cc",
          4691 => x"82",
          4692 => x"af",
          4693 => x"82",
          4694 => x"54",
          4695 => x"f9",
          4696 => x"cd",
          4697 => x"88",
          4698 => x"c7",
          4699 => x"fc",
          4700 => x"54",
          4701 => x"fc",
          4702 => x"ff",
          4703 => x"39",
          4704 => x"33",
          4705 => x"33",
          4706 => x"75",
          4707 => x"38",
          4708 => x"73",
          4709 => x"34",
          4710 => x"70",
          4711 => x"81",
          4712 => x"51",
          4713 => x"25",
          4714 => x"1a",
          4715 => x"33",
          4716 => x"cd",
          4717 => x"73",
          4718 => x"9f",
          4719 => x"81",
          4720 => x"81",
          4721 => x"70",
          4722 => x"cc",
          4723 => x"51",
          4724 => x"24",
          4725 => x"cd",
          4726 => x"a0",
          4727 => x"d3",
          4728 => x"fc",
          4729 => x"2b",
          4730 => x"82",
          4731 => x"57",
          4732 => x"74",
          4733 => x"a3",
          4734 => x"9c",
          4735 => x"51",
          4736 => x"3f",
          4737 => x"0a",
          4738 => x"0a",
          4739 => x"2c",
          4740 => x"33",
          4741 => x"75",
          4742 => x"38",
          4743 => x"82",
          4744 => x"70",
          4745 => x"82",
          4746 => x"59",
          4747 => x"77",
          4748 => x"38",
          4749 => x"08",
          4750 => x"54",
          4751 => x"fc",
          4752 => x"70",
          4753 => x"ff",
          4754 => x"82",
          4755 => x"70",
          4756 => x"82",
          4757 => x"58",
          4758 => x"75",
          4759 => x"f7",
          4760 => x"cc",
          4761 => x"52",
          4762 => x"51",
          4763 => x"80",
          4764 => x"fc",
          4765 => x"82",
          4766 => x"f7",
          4767 => x"b0",
          4768 => x"94",
          4769 => x"80",
          4770 => x"74",
          4771 => x"f6",
          4772 => x"c8",
          4773 => x"f8",
          4774 => x"c8",
          4775 => x"06",
          4776 => x"74",
          4777 => x"ff",
          4778 => x"93",
          4779 => x"39",
          4780 => x"82",
          4781 => x"fc",
          4782 => x"54",
          4783 => x"a7",
          4784 => x"ff",
          4785 => x"82",
          4786 => x"82",
          4787 => x"82",
          4788 => x"81",
          4789 => x"05",
          4790 => x"79",
          4791 => x"86",
          4792 => x"54",
          4793 => x"73",
          4794 => x"80",
          4795 => x"38",
          4796 => x"a6",
          4797 => x"39",
          4798 => x"09",
          4799 => x"38",
          4800 => x"08",
          4801 => x"2e",
          4802 => x"51",
          4803 => x"3f",
          4804 => x"08",
          4805 => x"34",
          4806 => x"08",
          4807 => x"81",
          4808 => x"52",
          4809 => x"a7",
          4810 => x"c3",
          4811 => x"29",
          4812 => x"05",
          4813 => x"54",
          4814 => x"ab",
          4815 => x"ff",
          4816 => x"82",
          4817 => x"82",
          4818 => x"82",
          4819 => x"81",
          4820 => x"05",
          4821 => x"79",
          4822 => x"8a",
          4823 => x"54",
          4824 => x"06",
          4825 => x"74",
          4826 => x"34",
          4827 => x"82",
          4828 => x"82",
          4829 => x"52",
          4830 => x"e2",
          4831 => x"39",
          4832 => x"33",
          4833 => x"06",
          4834 => x"33",
          4835 => x"74",
          4836 => x"87",
          4837 => x"9c",
          4838 => x"14",
          4839 => x"cc",
          4840 => x"1a",
          4841 => x"54",
          4842 => x"3f",
          4843 => x"82",
          4844 => x"54",
          4845 => x"f4",
          4846 => x"cd",
          4847 => x"88",
          4848 => x"ef",
          4849 => x"fc",
          4850 => x"54",
          4851 => x"fc",
          4852 => x"39",
          4853 => x"83",
          4854 => x"82",
          4855 => x"84",
          4856 => x"b5",
          4857 => x"80",
          4858 => x"83",
          4859 => x"ff",
          4860 => x"82",
          4861 => x"54",
          4862 => x"74",
          4863 => x"76",
          4864 => x"82",
          4865 => x"54",
          4866 => x"34",
          4867 => x"34",
          4868 => x"08",
          4869 => x"15",
          4870 => x"15",
          4871 => x"c0",
          4872 => x"bc",
          4873 => x"fe",
          4874 => x"70",
          4875 => x"06",
          4876 => x"58",
          4877 => x"74",
          4878 => x"73",
          4879 => x"82",
          4880 => x"70",
          4881 => x"b5",
          4882 => x"f8",
          4883 => x"55",
          4884 => x"34",
          4885 => x"34",
          4886 => x"04",
          4887 => x"73",
          4888 => x"84",
          4889 => x"38",
          4890 => x"2a",
          4891 => x"83",
          4892 => x"51",
          4893 => x"82",
          4894 => x"83",
          4895 => x"f9",
          4896 => x"a6",
          4897 => x"84",
          4898 => x"22",
          4899 => x"b5",
          4900 => x"83",
          4901 => x"74",
          4902 => x"11",
          4903 => x"12",
          4904 => x"2b",
          4905 => x"05",
          4906 => x"71",
          4907 => x"06",
          4908 => x"2a",
          4909 => x"59",
          4910 => x"57",
          4911 => x"71",
          4912 => x"81",
          4913 => x"b5",
          4914 => x"75",
          4915 => x"54",
          4916 => x"34",
          4917 => x"34",
          4918 => x"08",
          4919 => x"33",
          4920 => x"71",
          4921 => x"70",
          4922 => x"ff",
          4923 => x"52",
          4924 => x"05",
          4925 => x"ff",
          4926 => x"2a",
          4927 => x"71",
          4928 => x"72",
          4929 => x"53",
          4930 => x"34",
          4931 => x"08",
          4932 => x"76",
          4933 => x"17",
          4934 => x"0d",
          4935 => x"0d",
          4936 => x"08",
          4937 => x"9e",
          4938 => x"83",
          4939 => x"86",
          4940 => x"12",
          4941 => x"2b",
          4942 => x"07",
          4943 => x"52",
          4944 => x"05",
          4945 => x"85",
          4946 => x"88",
          4947 => x"88",
          4948 => x"56",
          4949 => x"13",
          4950 => x"13",
          4951 => x"c0",
          4952 => x"84",
          4953 => x"12",
          4954 => x"2b",
          4955 => x"07",
          4956 => x"52",
          4957 => x"12",
          4958 => x"33",
          4959 => x"07",
          4960 => x"54",
          4961 => x"70",
          4962 => x"73",
          4963 => x"82",
          4964 => x"13",
          4965 => x"12",
          4966 => x"2b",
          4967 => x"ff",
          4968 => x"88",
          4969 => x"53",
          4970 => x"73",
          4971 => x"14",
          4972 => x"0d",
          4973 => x"0d",
          4974 => x"22",
          4975 => x"08",
          4976 => x"71",
          4977 => x"81",
          4978 => x"88",
          4979 => x"88",
          4980 => x"33",
          4981 => x"71",
          4982 => x"90",
          4983 => x"5f",
          4984 => x"5a",
          4985 => x"54",
          4986 => x"80",
          4987 => x"51",
          4988 => x"82",
          4989 => x"70",
          4990 => x"81",
          4991 => x"8b",
          4992 => x"2b",
          4993 => x"70",
          4994 => x"33",
          4995 => x"07",
          4996 => x"8f",
          4997 => x"51",
          4998 => x"53",
          4999 => x"72",
          5000 => x"2a",
          5001 => x"82",
          5002 => x"83",
          5003 => x"b5",
          5004 => x"16",
          5005 => x"12",
          5006 => x"2b",
          5007 => x"07",
          5008 => x"55",
          5009 => x"33",
          5010 => x"71",
          5011 => x"70",
          5012 => x"06",
          5013 => x"57",
          5014 => x"52",
          5015 => x"71",
          5016 => x"88",
          5017 => x"fb",
          5018 => x"b5",
          5019 => x"84",
          5020 => x"22",
          5021 => x"72",
          5022 => x"33",
          5023 => x"71",
          5024 => x"83",
          5025 => x"5b",
          5026 => x"52",
          5027 => x"33",
          5028 => x"71",
          5029 => x"02",
          5030 => x"05",
          5031 => x"70",
          5032 => x"51",
          5033 => x"71",
          5034 => x"81",
          5035 => x"b5",
          5036 => x"15",
          5037 => x"12",
          5038 => x"2b",
          5039 => x"07",
          5040 => x"52",
          5041 => x"12",
          5042 => x"33",
          5043 => x"07",
          5044 => x"54",
          5045 => x"70",
          5046 => x"72",
          5047 => x"82",
          5048 => x"14",
          5049 => x"83",
          5050 => x"88",
          5051 => x"b5",
          5052 => x"54",
          5053 => x"04",
          5054 => x"7b",
          5055 => x"08",
          5056 => x"70",
          5057 => x"06",
          5058 => x"53",
          5059 => x"82",
          5060 => x"76",
          5061 => x"11",
          5062 => x"83",
          5063 => x"8b",
          5064 => x"2b",
          5065 => x"70",
          5066 => x"33",
          5067 => x"71",
          5068 => x"53",
          5069 => x"53",
          5070 => x"59",
          5071 => x"25",
          5072 => x"80",
          5073 => x"51",
          5074 => x"81",
          5075 => x"14",
          5076 => x"33",
          5077 => x"71",
          5078 => x"76",
          5079 => x"2a",
          5080 => x"58",
          5081 => x"14",
          5082 => x"ff",
          5083 => x"87",
          5084 => x"b5",
          5085 => x"19",
          5086 => x"85",
          5087 => x"88",
          5088 => x"88",
          5089 => x"5b",
          5090 => x"84",
          5091 => x"85",
          5092 => x"b5",
          5093 => x"53",
          5094 => x"14",
          5095 => x"87",
          5096 => x"b5",
          5097 => x"76",
          5098 => x"75",
          5099 => x"82",
          5100 => x"18",
          5101 => x"12",
          5102 => x"2b",
          5103 => x"80",
          5104 => x"88",
          5105 => x"55",
          5106 => x"74",
          5107 => x"15",
          5108 => x"0d",
          5109 => x"0d",
          5110 => x"b5",
          5111 => x"38",
          5112 => x"71",
          5113 => x"38",
          5114 => x"8c",
          5115 => x"0d",
          5116 => x"0d",
          5117 => x"58",
          5118 => x"82",
          5119 => x"83",
          5120 => x"82",
          5121 => x"84",
          5122 => x"12",
          5123 => x"2b",
          5124 => x"59",
          5125 => x"81",
          5126 => x"75",
          5127 => x"cb",
          5128 => x"29",
          5129 => x"81",
          5130 => x"88",
          5131 => x"81",
          5132 => x"79",
          5133 => x"ff",
          5134 => x"7f",
          5135 => x"51",
          5136 => x"77",
          5137 => x"38",
          5138 => x"85",
          5139 => x"5a",
          5140 => x"33",
          5141 => x"71",
          5142 => x"57",
          5143 => x"38",
          5144 => x"ff",
          5145 => x"7a",
          5146 => x"80",
          5147 => x"82",
          5148 => x"11",
          5149 => x"12",
          5150 => x"2b",
          5151 => x"ff",
          5152 => x"52",
          5153 => x"55",
          5154 => x"83",
          5155 => x"80",
          5156 => x"26",
          5157 => x"74",
          5158 => x"2e",
          5159 => x"77",
          5160 => x"81",
          5161 => x"75",
          5162 => x"3f",
          5163 => x"82",
          5164 => x"79",
          5165 => x"f7",
          5166 => x"b5",
          5167 => x"1c",
          5168 => x"87",
          5169 => x"8b",
          5170 => x"2b",
          5171 => x"5e",
          5172 => x"7a",
          5173 => x"ff",
          5174 => x"88",
          5175 => x"56",
          5176 => x"15",
          5177 => x"ff",
          5178 => x"85",
          5179 => x"b5",
          5180 => x"83",
          5181 => x"72",
          5182 => x"33",
          5183 => x"71",
          5184 => x"70",
          5185 => x"5b",
          5186 => x"56",
          5187 => x"19",
          5188 => x"19",
          5189 => x"c0",
          5190 => x"84",
          5191 => x"12",
          5192 => x"2b",
          5193 => x"07",
          5194 => x"55",
          5195 => x"78",
          5196 => x"76",
          5197 => x"82",
          5198 => x"70",
          5199 => x"84",
          5200 => x"12",
          5201 => x"2b",
          5202 => x"2a",
          5203 => x"52",
          5204 => x"84",
          5205 => x"85",
          5206 => x"b5",
          5207 => x"84",
          5208 => x"82",
          5209 => x"8d",
          5210 => x"fe",
          5211 => x"52",
          5212 => x"08",
          5213 => x"dc",
          5214 => x"71",
          5215 => x"38",
          5216 => x"ed",
          5217 => x"c8",
          5218 => x"82",
          5219 => x"84",
          5220 => x"ee",
          5221 => x"66",
          5222 => x"70",
          5223 => x"b5",
          5224 => x"2e",
          5225 => x"84",
          5226 => x"3f",
          5227 => x"7e",
          5228 => x"3f",
          5229 => x"08",
          5230 => x"39",
          5231 => x"7b",
          5232 => x"3f",
          5233 => x"ba",
          5234 => x"f5",
          5235 => x"b5",
          5236 => x"ff",
          5237 => x"b5",
          5238 => x"71",
          5239 => x"70",
          5240 => x"06",
          5241 => x"73",
          5242 => x"81",
          5243 => x"88",
          5244 => x"75",
          5245 => x"ff",
          5246 => x"88",
          5247 => x"73",
          5248 => x"70",
          5249 => x"33",
          5250 => x"07",
          5251 => x"53",
          5252 => x"48",
          5253 => x"54",
          5254 => x"56",
          5255 => x"80",
          5256 => x"76",
          5257 => x"06",
          5258 => x"83",
          5259 => x"42",
          5260 => x"33",
          5261 => x"71",
          5262 => x"70",
          5263 => x"70",
          5264 => x"33",
          5265 => x"71",
          5266 => x"53",
          5267 => x"56",
          5268 => x"25",
          5269 => x"75",
          5270 => x"ff",
          5271 => x"54",
          5272 => x"81",
          5273 => x"18",
          5274 => x"2e",
          5275 => x"8f",
          5276 => x"f6",
          5277 => x"83",
          5278 => x"58",
          5279 => x"7f",
          5280 => x"74",
          5281 => x"78",
          5282 => x"3f",
          5283 => x"7f",
          5284 => x"75",
          5285 => x"38",
          5286 => x"11",
          5287 => x"33",
          5288 => x"07",
          5289 => x"f4",
          5290 => x"52",
          5291 => x"b7",
          5292 => x"c8",
          5293 => x"ff",
          5294 => x"7c",
          5295 => x"2b",
          5296 => x"08",
          5297 => x"53",
          5298 => x"93",
          5299 => x"b5",
          5300 => x"84",
          5301 => x"ff",
          5302 => x"5c",
          5303 => x"60",
          5304 => x"74",
          5305 => x"38",
          5306 => x"c9",
          5307 => x"c0",
          5308 => x"11",
          5309 => x"33",
          5310 => x"07",
          5311 => x"f4",
          5312 => x"52",
          5313 => x"df",
          5314 => x"c8",
          5315 => x"ff",
          5316 => x"7c",
          5317 => x"2b",
          5318 => x"08",
          5319 => x"53",
          5320 => x"92",
          5321 => x"b5",
          5322 => x"84",
          5323 => x"05",
          5324 => x"73",
          5325 => x"06",
          5326 => x"7b",
          5327 => x"f9",
          5328 => x"b5",
          5329 => x"82",
          5330 => x"80",
          5331 => x"7d",
          5332 => x"82",
          5333 => x"51",
          5334 => x"3f",
          5335 => x"98",
          5336 => x"7a",
          5337 => x"38",
          5338 => x"52",
          5339 => x"8f",
          5340 => x"83",
          5341 => x"c0",
          5342 => x"05",
          5343 => x"3f",
          5344 => x"82",
          5345 => x"94",
          5346 => x"fc",
          5347 => x"77",
          5348 => x"54",
          5349 => x"82",
          5350 => x"55",
          5351 => x"08",
          5352 => x"38",
          5353 => x"52",
          5354 => x"08",
          5355 => x"b7",
          5356 => x"b5",
          5357 => x"3d",
          5358 => x"3d",
          5359 => x"05",
          5360 => x"52",
          5361 => x"87",
          5362 => x"c4",
          5363 => x"71",
          5364 => x"0c",
          5365 => x"04",
          5366 => x"02",
          5367 => x"02",
          5368 => x"05",
          5369 => x"83",
          5370 => x"26",
          5371 => x"72",
          5372 => x"c0",
          5373 => x"53",
          5374 => x"74",
          5375 => x"38",
          5376 => x"73",
          5377 => x"c0",
          5378 => x"51",
          5379 => x"85",
          5380 => x"98",
          5381 => x"52",
          5382 => x"82",
          5383 => x"70",
          5384 => x"38",
          5385 => x"8c",
          5386 => x"ec",
          5387 => x"fc",
          5388 => x"52",
          5389 => x"87",
          5390 => x"08",
          5391 => x"2e",
          5392 => x"82",
          5393 => x"34",
          5394 => x"13",
          5395 => x"82",
          5396 => x"86",
          5397 => x"f3",
          5398 => x"62",
          5399 => x"05",
          5400 => x"57",
          5401 => x"83",
          5402 => x"fe",
          5403 => x"b5",
          5404 => x"06",
          5405 => x"71",
          5406 => x"71",
          5407 => x"2b",
          5408 => x"80",
          5409 => x"92",
          5410 => x"c0",
          5411 => x"41",
          5412 => x"5a",
          5413 => x"87",
          5414 => x"0c",
          5415 => x"84",
          5416 => x"08",
          5417 => x"70",
          5418 => x"53",
          5419 => x"2e",
          5420 => x"08",
          5421 => x"70",
          5422 => x"34",
          5423 => x"80",
          5424 => x"53",
          5425 => x"2e",
          5426 => x"53",
          5427 => x"26",
          5428 => x"80",
          5429 => x"87",
          5430 => x"08",
          5431 => x"38",
          5432 => x"8c",
          5433 => x"80",
          5434 => x"78",
          5435 => x"99",
          5436 => x"0c",
          5437 => x"8c",
          5438 => x"08",
          5439 => x"51",
          5440 => x"38",
          5441 => x"8d",
          5442 => x"17",
          5443 => x"81",
          5444 => x"53",
          5445 => x"2e",
          5446 => x"fc",
          5447 => x"52",
          5448 => x"7d",
          5449 => x"ed",
          5450 => x"80",
          5451 => x"71",
          5452 => x"38",
          5453 => x"53",
          5454 => x"c8",
          5455 => x"0d",
          5456 => x"0d",
          5457 => x"02",
          5458 => x"05",
          5459 => x"58",
          5460 => x"80",
          5461 => x"fc",
          5462 => x"b5",
          5463 => x"06",
          5464 => x"71",
          5465 => x"81",
          5466 => x"38",
          5467 => x"2b",
          5468 => x"80",
          5469 => x"92",
          5470 => x"c0",
          5471 => x"40",
          5472 => x"5a",
          5473 => x"c0",
          5474 => x"76",
          5475 => x"76",
          5476 => x"75",
          5477 => x"2a",
          5478 => x"51",
          5479 => x"80",
          5480 => x"7a",
          5481 => x"5c",
          5482 => x"81",
          5483 => x"81",
          5484 => x"06",
          5485 => x"80",
          5486 => x"87",
          5487 => x"08",
          5488 => x"38",
          5489 => x"8c",
          5490 => x"80",
          5491 => x"77",
          5492 => x"99",
          5493 => x"0c",
          5494 => x"8c",
          5495 => x"08",
          5496 => x"51",
          5497 => x"38",
          5498 => x"8d",
          5499 => x"70",
          5500 => x"84",
          5501 => x"5b",
          5502 => x"2e",
          5503 => x"fc",
          5504 => x"52",
          5505 => x"7d",
          5506 => x"f8",
          5507 => x"80",
          5508 => x"71",
          5509 => x"38",
          5510 => x"53",
          5511 => x"c8",
          5512 => x"0d",
          5513 => x"0d",
          5514 => x"05",
          5515 => x"02",
          5516 => x"05",
          5517 => x"54",
          5518 => x"fe",
          5519 => x"c8",
          5520 => x"53",
          5521 => x"80",
          5522 => x"0b",
          5523 => x"8c",
          5524 => x"71",
          5525 => x"dc",
          5526 => x"24",
          5527 => x"84",
          5528 => x"92",
          5529 => x"54",
          5530 => x"8d",
          5531 => x"39",
          5532 => x"80",
          5533 => x"cb",
          5534 => x"70",
          5535 => x"81",
          5536 => x"52",
          5537 => x"8a",
          5538 => x"98",
          5539 => x"71",
          5540 => x"c0",
          5541 => x"52",
          5542 => x"81",
          5543 => x"c0",
          5544 => x"53",
          5545 => x"82",
          5546 => x"71",
          5547 => x"39",
          5548 => x"39",
          5549 => x"77",
          5550 => x"81",
          5551 => x"72",
          5552 => x"84",
          5553 => x"73",
          5554 => x"0c",
          5555 => x"04",
          5556 => x"74",
          5557 => x"71",
          5558 => x"2b",
          5559 => x"c8",
          5560 => x"84",
          5561 => x"fd",
          5562 => x"83",
          5563 => x"12",
          5564 => x"2b",
          5565 => x"07",
          5566 => x"70",
          5567 => x"2b",
          5568 => x"07",
          5569 => x"0c",
          5570 => x"56",
          5571 => x"3d",
          5572 => x"3d",
          5573 => x"84",
          5574 => x"22",
          5575 => x"72",
          5576 => x"54",
          5577 => x"2a",
          5578 => x"34",
          5579 => x"04",
          5580 => x"73",
          5581 => x"70",
          5582 => x"05",
          5583 => x"88",
          5584 => x"72",
          5585 => x"54",
          5586 => x"2a",
          5587 => x"70",
          5588 => x"34",
          5589 => x"51",
          5590 => x"83",
          5591 => x"fe",
          5592 => x"75",
          5593 => x"51",
          5594 => x"92",
          5595 => x"81",
          5596 => x"73",
          5597 => x"55",
          5598 => x"51",
          5599 => x"3d",
          5600 => x"3d",
          5601 => x"76",
          5602 => x"72",
          5603 => x"05",
          5604 => x"11",
          5605 => x"38",
          5606 => x"04",
          5607 => x"78",
          5608 => x"56",
          5609 => x"81",
          5610 => x"74",
          5611 => x"56",
          5612 => x"31",
          5613 => x"52",
          5614 => x"80",
          5615 => x"71",
          5616 => x"38",
          5617 => x"c8",
          5618 => x"0d",
          5619 => x"0d",
          5620 => x"51",
          5621 => x"73",
          5622 => x"81",
          5623 => x"33",
          5624 => x"38",
          5625 => x"b5",
          5626 => x"3d",
          5627 => x"0b",
          5628 => x"0c",
          5629 => x"82",
          5630 => x"04",
          5631 => x"7b",
          5632 => x"83",
          5633 => x"5a",
          5634 => x"80",
          5635 => x"54",
          5636 => x"53",
          5637 => x"53",
          5638 => x"52",
          5639 => x"3f",
          5640 => x"08",
          5641 => x"81",
          5642 => x"82",
          5643 => x"83",
          5644 => x"16",
          5645 => x"18",
          5646 => x"18",
          5647 => x"58",
          5648 => x"9f",
          5649 => x"33",
          5650 => x"2e",
          5651 => x"93",
          5652 => x"76",
          5653 => x"52",
          5654 => x"51",
          5655 => x"83",
          5656 => x"79",
          5657 => x"0c",
          5658 => x"04",
          5659 => x"78",
          5660 => x"80",
          5661 => x"17",
          5662 => x"38",
          5663 => x"fc",
          5664 => x"c8",
          5665 => x"b5",
          5666 => x"38",
          5667 => x"53",
          5668 => x"81",
          5669 => x"f7",
          5670 => x"b5",
          5671 => x"2e",
          5672 => x"55",
          5673 => x"b0",
          5674 => x"82",
          5675 => x"88",
          5676 => x"f8",
          5677 => x"70",
          5678 => x"c0",
          5679 => x"c8",
          5680 => x"b5",
          5681 => x"91",
          5682 => x"55",
          5683 => x"09",
          5684 => x"f0",
          5685 => x"33",
          5686 => x"2e",
          5687 => x"80",
          5688 => x"80",
          5689 => x"c8",
          5690 => x"17",
          5691 => x"fd",
          5692 => x"d4",
          5693 => x"b2",
          5694 => x"96",
          5695 => x"85",
          5696 => x"75",
          5697 => x"3f",
          5698 => x"e4",
          5699 => x"98",
          5700 => x"9c",
          5701 => x"08",
          5702 => x"17",
          5703 => x"3f",
          5704 => x"52",
          5705 => x"51",
          5706 => x"a0",
          5707 => x"05",
          5708 => x"0c",
          5709 => x"75",
          5710 => x"33",
          5711 => x"3f",
          5712 => x"34",
          5713 => x"52",
          5714 => x"51",
          5715 => x"82",
          5716 => x"80",
          5717 => x"81",
          5718 => x"b5",
          5719 => x"3d",
          5720 => x"3d",
          5721 => x"1a",
          5722 => x"fe",
          5723 => x"54",
          5724 => x"73",
          5725 => x"8a",
          5726 => x"71",
          5727 => x"08",
          5728 => x"75",
          5729 => x"0c",
          5730 => x"04",
          5731 => x"7a",
          5732 => x"56",
          5733 => x"77",
          5734 => x"38",
          5735 => x"08",
          5736 => x"38",
          5737 => x"54",
          5738 => x"2e",
          5739 => x"72",
          5740 => x"38",
          5741 => x"8d",
          5742 => x"39",
          5743 => x"81",
          5744 => x"b6",
          5745 => x"2a",
          5746 => x"2a",
          5747 => x"05",
          5748 => x"55",
          5749 => x"82",
          5750 => x"81",
          5751 => x"83",
          5752 => x"b4",
          5753 => x"17",
          5754 => x"a4",
          5755 => x"55",
          5756 => x"57",
          5757 => x"3f",
          5758 => x"08",
          5759 => x"74",
          5760 => x"14",
          5761 => x"70",
          5762 => x"07",
          5763 => x"71",
          5764 => x"52",
          5765 => x"72",
          5766 => x"75",
          5767 => x"58",
          5768 => x"76",
          5769 => x"15",
          5770 => x"73",
          5771 => x"3f",
          5772 => x"08",
          5773 => x"76",
          5774 => x"06",
          5775 => x"05",
          5776 => x"3f",
          5777 => x"08",
          5778 => x"06",
          5779 => x"76",
          5780 => x"15",
          5781 => x"73",
          5782 => x"3f",
          5783 => x"08",
          5784 => x"82",
          5785 => x"06",
          5786 => x"05",
          5787 => x"3f",
          5788 => x"08",
          5789 => x"58",
          5790 => x"58",
          5791 => x"c8",
          5792 => x"0d",
          5793 => x"0d",
          5794 => x"5a",
          5795 => x"59",
          5796 => x"82",
          5797 => x"98",
          5798 => x"82",
          5799 => x"33",
          5800 => x"2e",
          5801 => x"72",
          5802 => x"38",
          5803 => x"8d",
          5804 => x"39",
          5805 => x"81",
          5806 => x"f7",
          5807 => x"2a",
          5808 => x"2a",
          5809 => x"05",
          5810 => x"55",
          5811 => x"82",
          5812 => x"59",
          5813 => x"08",
          5814 => x"74",
          5815 => x"16",
          5816 => x"16",
          5817 => x"59",
          5818 => x"53",
          5819 => x"8f",
          5820 => x"2b",
          5821 => x"74",
          5822 => x"71",
          5823 => x"72",
          5824 => x"0b",
          5825 => x"74",
          5826 => x"17",
          5827 => x"75",
          5828 => x"3f",
          5829 => x"08",
          5830 => x"c8",
          5831 => x"38",
          5832 => x"06",
          5833 => x"78",
          5834 => x"54",
          5835 => x"77",
          5836 => x"33",
          5837 => x"71",
          5838 => x"51",
          5839 => x"34",
          5840 => x"76",
          5841 => x"17",
          5842 => x"75",
          5843 => x"3f",
          5844 => x"08",
          5845 => x"c8",
          5846 => x"38",
          5847 => x"ff",
          5848 => x"10",
          5849 => x"76",
          5850 => x"51",
          5851 => x"be",
          5852 => x"2a",
          5853 => x"05",
          5854 => x"f9",
          5855 => x"b5",
          5856 => x"82",
          5857 => x"ab",
          5858 => x"0a",
          5859 => x"2b",
          5860 => x"70",
          5861 => x"70",
          5862 => x"54",
          5863 => x"82",
          5864 => x"8f",
          5865 => x"07",
          5866 => x"f7",
          5867 => x"0b",
          5868 => x"78",
          5869 => x"0c",
          5870 => x"04",
          5871 => x"7a",
          5872 => x"08",
          5873 => x"59",
          5874 => x"a4",
          5875 => x"17",
          5876 => x"38",
          5877 => x"aa",
          5878 => x"73",
          5879 => x"fd",
          5880 => x"b5",
          5881 => x"82",
          5882 => x"80",
          5883 => x"39",
          5884 => x"eb",
          5885 => x"80",
          5886 => x"b5",
          5887 => x"80",
          5888 => x"52",
          5889 => x"84",
          5890 => x"c8",
          5891 => x"b5",
          5892 => x"2e",
          5893 => x"82",
          5894 => x"81",
          5895 => x"82",
          5896 => x"ff",
          5897 => x"80",
          5898 => x"75",
          5899 => x"3f",
          5900 => x"08",
          5901 => x"16",
          5902 => x"90",
          5903 => x"55",
          5904 => x"27",
          5905 => x"15",
          5906 => x"84",
          5907 => x"07",
          5908 => x"17",
          5909 => x"76",
          5910 => x"a6",
          5911 => x"73",
          5912 => x"0c",
          5913 => x"04",
          5914 => x"7c",
          5915 => x"59",
          5916 => x"95",
          5917 => x"08",
          5918 => x"2e",
          5919 => x"17",
          5920 => x"b2",
          5921 => x"ae",
          5922 => x"7a",
          5923 => x"3f",
          5924 => x"82",
          5925 => x"27",
          5926 => x"82",
          5927 => x"55",
          5928 => x"08",
          5929 => x"d2",
          5930 => x"08",
          5931 => x"08",
          5932 => x"38",
          5933 => x"17",
          5934 => x"54",
          5935 => x"82",
          5936 => x"7a",
          5937 => x"06",
          5938 => x"81",
          5939 => x"17",
          5940 => x"83",
          5941 => x"75",
          5942 => x"f9",
          5943 => x"59",
          5944 => x"08",
          5945 => x"81",
          5946 => x"82",
          5947 => x"59",
          5948 => x"08",
          5949 => x"70",
          5950 => x"25",
          5951 => x"82",
          5952 => x"54",
          5953 => x"55",
          5954 => x"38",
          5955 => x"08",
          5956 => x"38",
          5957 => x"54",
          5958 => x"90",
          5959 => x"18",
          5960 => x"38",
          5961 => x"39",
          5962 => x"38",
          5963 => x"16",
          5964 => x"08",
          5965 => x"38",
          5966 => x"78",
          5967 => x"38",
          5968 => x"51",
          5969 => x"82",
          5970 => x"80",
          5971 => x"80",
          5972 => x"c8",
          5973 => x"09",
          5974 => x"38",
          5975 => x"08",
          5976 => x"c8",
          5977 => x"30",
          5978 => x"80",
          5979 => x"07",
          5980 => x"55",
          5981 => x"38",
          5982 => x"09",
          5983 => x"ae",
          5984 => x"80",
          5985 => x"53",
          5986 => x"51",
          5987 => x"82",
          5988 => x"82",
          5989 => x"30",
          5990 => x"c8",
          5991 => x"25",
          5992 => x"79",
          5993 => x"38",
          5994 => x"8f",
          5995 => x"79",
          5996 => x"f9",
          5997 => x"b5",
          5998 => x"74",
          5999 => x"8c",
          6000 => x"17",
          6001 => x"90",
          6002 => x"54",
          6003 => x"86",
          6004 => x"90",
          6005 => x"17",
          6006 => x"54",
          6007 => x"34",
          6008 => x"56",
          6009 => x"90",
          6010 => x"80",
          6011 => x"82",
          6012 => x"55",
          6013 => x"56",
          6014 => x"82",
          6015 => x"8c",
          6016 => x"f8",
          6017 => x"70",
          6018 => x"f0",
          6019 => x"c8",
          6020 => x"56",
          6021 => x"08",
          6022 => x"7b",
          6023 => x"f6",
          6024 => x"b5",
          6025 => x"b5",
          6026 => x"17",
          6027 => x"80",
          6028 => x"b4",
          6029 => x"57",
          6030 => x"77",
          6031 => x"81",
          6032 => x"15",
          6033 => x"78",
          6034 => x"81",
          6035 => x"53",
          6036 => x"15",
          6037 => x"e9",
          6038 => x"c8",
          6039 => x"df",
          6040 => x"22",
          6041 => x"30",
          6042 => x"70",
          6043 => x"51",
          6044 => x"82",
          6045 => x"8a",
          6046 => x"f8",
          6047 => x"7c",
          6048 => x"56",
          6049 => x"80",
          6050 => x"f1",
          6051 => x"06",
          6052 => x"e9",
          6053 => x"18",
          6054 => x"08",
          6055 => x"38",
          6056 => x"82",
          6057 => x"38",
          6058 => x"54",
          6059 => x"74",
          6060 => x"82",
          6061 => x"22",
          6062 => x"79",
          6063 => x"38",
          6064 => x"98",
          6065 => x"cd",
          6066 => x"22",
          6067 => x"54",
          6068 => x"26",
          6069 => x"52",
          6070 => x"b0",
          6071 => x"c8",
          6072 => x"b5",
          6073 => x"2e",
          6074 => x"0b",
          6075 => x"08",
          6076 => x"98",
          6077 => x"b5",
          6078 => x"85",
          6079 => x"bd",
          6080 => x"31",
          6081 => x"73",
          6082 => x"f4",
          6083 => x"b5",
          6084 => x"18",
          6085 => x"18",
          6086 => x"08",
          6087 => x"72",
          6088 => x"38",
          6089 => x"58",
          6090 => x"89",
          6091 => x"18",
          6092 => x"ff",
          6093 => x"05",
          6094 => x"80",
          6095 => x"b5",
          6096 => x"3d",
          6097 => x"3d",
          6098 => x"08",
          6099 => x"a0",
          6100 => x"54",
          6101 => x"77",
          6102 => x"80",
          6103 => x"0c",
          6104 => x"53",
          6105 => x"80",
          6106 => x"38",
          6107 => x"06",
          6108 => x"b5",
          6109 => x"98",
          6110 => x"14",
          6111 => x"92",
          6112 => x"2a",
          6113 => x"56",
          6114 => x"26",
          6115 => x"80",
          6116 => x"16",
          6117 => x"77",
          6118 => x"53",
          6119 => x"38",
          6120 => x"51",
          6121 => x"82",
          6122 => x"53",
          6123 => x"0b",
          6124 => x"08",
          6125 => x"38",
          6126 => x"b5",
          6127 => x"2e",
          6128 => x"98",
          6129 => x"b5",
          6130 => x"80",
          6131 => x"8a",
          6132 => x"15",
          6133 => x"80",
          6134 => x"14",
          6135 => x"51",
          6136 => x"82",
          6137 => x"53",
          6138 => x"b5",
          6139 => x"2e",
          6140 => x"82",
          6141 => x"c8",
          6142 => x"ba",
          6143 => x"82",
          6144 => x"ff",
          6145 => x"82",
          6146 => x"52",
          6147 => x"f3",
          6148 => x"c8",
          6149 => x"72",
          6150 => x"72",
          6151 => x"f2",
          6152 => x"b5",
          6153 => x"15",
          6154 => x"15",
          6155 => x"b4",
          6156 => x"0c",
          6157 => x"82",
          6158 => x"8a",
          6159 => x"f7",
          6160 => x"7d",
          6161 => x"5b",
          6162 => x"76",
          6163 => x"3f",
          6164 => x"08",
          6165 => x"c8",
          6166 => x"38",
          6167 => x"08",
          6168 => x"08",
          6169 => x"f0",
          6170 => x"b5",
          6171 => x"82",
          6172 => x"80",
          6173 => x"b5",
          6174 => x"18",
          6175 => x"51",
          6176 => x"81",
          6177 => x"81",
          6178 => x"81",
          6179 => x"c8",
          6180 => x"83",
          6181 => x"77",
          6182 => x"72",
          6183 => x"38",
          6184 => x"75",
          6185 => x"81",
          6186 => x"a5",
          6187 => x"c8",
          6188 => x"52",
          6189 => x"8e",
          6190 => x"c8",
          6191 => x"b5",
          6192 => x"2e",
          6193 => x"73",
          6194 => x"81",
          6195 => x"87",
          6196 => x"b5",
          6197 => x"3d",
          6198 => x"3d",
          6199 => x"11",
          6200 => x"ec",
          6201 => x"c8",
          6202 => x"ff",
          6203 => x"33",
          6204 => x"71",
          6205 => x"81",
          6206 => x"94",
          6207 => x"d0",
          6208 => x"c8",
          6209 => x"73",
          6210 => x"82",
          6211 => x"85",
          6212 => x"fc",
          6213 => x"79",
          6214 => x"ff",
          6215 => x"12",
          6216 => x"eb",
          6217 => x"70",
          6218 => x"72",
          6219 => x"81",
          6220 => x"73",
          6221 => x"94",
          6222 => x"d6",
          6223 => x"0d",
          6224 => x"0d",
          6225 => x"55",
          6226 => x"5a",
          6227 => x"08",
          6228 => x"8a",
          6229 => x"08",
          6230 => x"ee",
          6231 => x"b5",
          6232 => x"82",
          6233 => x"80",
          6234 => x"15",
          6235 => x"55",
          6236 => x"38",
          6237 => x"e6",
          6238 => x"33",
          6239 => x"70",
          6240 => x"58",
          6241 => x"86",
          6242 => x"b5",
          6243 => x"73",
          6244 => x"83",
          6245 => x"73",
          6246 => x"38",
          6247 => x"06",
          6248 => x"80",
          6249 => x"75",
          6250 => x"38",
          6251 => x"08",
          6252 => x"54",
          6253 => x"2e",
          6254 => x"83",
          6255 => x"73",
          6256 => x"38",
          6257 => x"51",
          6258 => x"82",
          6259 => x"58",
          6260 => x"08",
          6261 => x"15",
          6262 => x"38",
          6263 => x"0b",
          6264 => x"77",
          6265 => x"0c",
          6266 => x"04",
          6267 => x"77",
          6268 => x"54",
          6269 => x"51",
          6270 => x"82",
          6271 => x"55",
          6272 => x"08",
          6273 => x"14",
          6274 => x"51",
          6275 => x"82",
          6276 => x"55",
          6277 => x"08",
          6278 => x"53",
          6279 => x"08",
          6280 => x"08",
          6281 => x"3f",
          6282 => x"14",
          6283 => x"08",
          6284 => x"3f",
          6285 => x"17",
          6286 => x"b5",
          6287 => x"3d",
          6288 => x"3d",
          6289 => x"08",
          6290 => x"54",
          6291 => x"53",
          6292 => x"82",
          6293 => x"8d",
          6294 => x"08",
          6295 => x"34",
          6296 => x"15",
          6297 => x"0d",
          6298 => x"0d",
          6299 => x"57",
          6300 => x"17",
          6301 => x"08",
          6302 => x"82",
          6303 => x"89",
          6304 => x"55",
          6305 => x"14",
          6306 => x"16",
          6307 => x"71",
          6308 => x"38",
          6309 => x"09",
          6310 => x"38",
          6311 => x"73",
          6312 => x"81",
          6313 => x"ae",
          6314 => x"05",
          6315 => x"15",
          6316 => x"70",
          6317 => x"34",
          6318 => x"8a",
          6319 => x"38",
          6320 => x"05",
          6321 => x"81",
          6322 => x"17",
          6323 => x"12",
          6324 => x"34",
          6325 => x"9c",
          6326 => x"e8",
          6327 => x"b5",
          6328 => x"0c",
          6329 => x"e7",
          6330 => x"b5",
          6331 => x"17",
          6332 => x"51",
          6333 => x"82",
          6334 => x"84",
          6335 => x"3d",
          6336 => x"3d",
          6337 => x"08",
          6338 => x"61",
          6339 => x"55",
          6340 => x"2e",
          6341 => x"55",
          6342 => x"2e",
          6343 => x"80",
          6344 => x"94",
          6345 => x"1c",
          6346 => x"81",
          6347 => x"61",
          6348 => x"56",
          6349 => x"2e",
          6350 => x"83",
          6351 => x"73",
          6352 => x"70",
          6353 => x"25",
          6354 => x"51",
          6355 => x"38",
          6356 => x"0c",
          6357 => x"51",
          6358 => x"26",
          6359 => x"80",
          6360 => x"34",
          6361 => x"51",
          6362 => x"82",
          6363 => x"55",
          6364 => x"91",
          6365 => x"1d",
          6366 => x"8b",
          6367 => x"79",
          6368 => x"3f",
          6369 => x"57",
          6370 => x"55",
          6371 => x"2e",
          6372 => x"80",
          6373 => x"18",
          6374 => x"1a",
          6375 => x"70",
          6376 => x"2a",
          6377 => x"07",
          6378 => x"5a",
          6379 => x"8c",
          6380 => x"54",
          6381 => x"81",
          6382 => x"39",
          6383 => x"70",
          6384 => x"2a",
          6385 => x"75",
          6386 => x"8c",
          6387 => x"2e",
          6388 => x"a0",
          6389 => x"38",
          6390 => x"0c",
          6391 => x"76",
          6392 => x"38",
          6393 => x"b8",
          6394 => x"70",
          6395 => x"5a",
          6396 => x"76",
          6397 => x"38",
          6398 => x"70",
          6399 => x"dc",
          6400 => x"72",
          6401 => x"80",
          6402 => x"51",
          6403 => x"73",
          6404 => x"38",
          6405 => x"18",
          6406 => x"1a",
          6407 => x"55",
          6408 => x"2e",
          6409 => x"83",
          6410 => x"73",
          6411 => x"70",
          6412 => x"25",
          6413 => x"51",
          6414 => x"38",
          6415 => x"75",
          6416 => x"81",
          6417 => x"81",
          6418 => x"27",
          6419 => x"73",
          6420 => x"38",
          6421 => x"70",
          6422 => x"32",
          6423 => x"80",
          6424 => x"2a",
          6425 => x"56",
          6426 => x"81",
          6427 => x"57",
          6428 => x"f5",
          6429 => x"2b",
          6430 => x"25",
          6431 => x"80",
          6432 => x"af",
          6433 => x"57",
          6434 => x"e6",
          6435 => x"b5",
          6436 => x"2e",
          6437 => x"18",
          6438 => x"1a",
          6439 => x"56",
          6440 => x"3f",
          6441 => x"08",
          6442 => x"e8",
          6443 => x"54",
          6444 => x"80",
          6445 => x"17",
          6446 => x"34",
          6447 => x"11",
          6448 => x"74",
          6449 => x"75",
          6450 => x"b0",
          6451 => x"3f",
          6452 => x"08",
          6453 => x"9f",
          6454 => x"99",
          6455 => x"e0",
          6456 => x"ff",
          6457 => x"79",
          6458 => x"74",
          6459 => x"57",
          6460 => x"77",
          6461 => x"76",
          6462 => x"38",
          6463 => x"73",
          6464 => x"09",
          6465 => x"38",
          6466 => x"84",
          6467 => x"27",
          6468 => x"39",
          6469 => x"f2",
          6470 => x"80",
          6471 => x"54",
          6472 => x"34",
          6473 => x"58",
          6474 => x"f2",
          6475 => x"b5",
          6476 => x"82",
          6477 => x"80",
          6478 => x"1b",
          6479 => x"51",
          6480 => x"82",
          6481 => x"56",
          6482 => x"08",
          6483 => x"9c",
          6484 => x"33",
          6485 => x"80",
          6486 => x"38",
          6487 => x"bf",
          6488 => x"86",
          6489 => x"15",
          6490 => x"2a",
          6491 => x"51",
          6492 => x"92",
          6493 => x"79",
          6494 => x"e4",
          6495 => x"b5",
          6496 => x"2e",
          6497 => x"52",
          6498 => x"ba",
          6499 => x"39",
          6500 => x"33",
          6501 => x"80",
          6502 => x"74",
          6503 => x"81",
          6504 => x"38",
          6505 => x"70",
          6506 => x"82",
          6507 => x"54",
          6508 => x"96",
          6509 => x"06",
          6510 => x"2e",
          6511 => x"ff",
          6512 => x"1c",
          6513 => x"80",
          6514 => x"81",
          6515 => x"ba",
          6516 => x"b6",
          6517 => x"2a",
          6518 => x"51",
          6519 => x"38",
          6520 => x"70",
          6521 => x"81",
          6522 => x"55",
          6523 => x"e1",
          6524 => x"08",
          6525 => x"1d",
          6526 => x"7c",
          6527 => x"3f",
          6528 => x"08",
          6529 => x"fa",
          6530 => x"82",
          6531 => x"8f",
          6532 => x"f6",
          6533 => x"5b",
          6534 => x"70",
          6535 => x"59",
          6536 => x"73",
          6537 => x"c6",
          6538 => x"81",
          6539 => x"70",
          6540 => x"52",
          6541 => x"8d",
          6542 => x"38",
          6543 => x"09",
          6544 => x"a5",
          6545 => x"d0",
          6546 => x"ff",
          6547 => x"53",
          6548 => x"91",
          6549 => x"73",
          6550 => x"d0",
          6551 => x"71",
          6552 => x"f7",
          6553 => x"82",
          6554 => x"55",
          6555 => x"55",
          6556 => x"81",
          6557 => x"74",
          6558 => x"56",
          6559 => x"12",
          6560 => x"70",
          6561 => x"38",
          6562 => x"81",
          6563 => x"51",
          6564 => x"51",
          6565 => x"89",
          6566 => x"70",
          6567 => x"53",
          6568 => x"70",
          6569 => x"51",
          6570 => x"09",
          6571 => x"38",
          6572 => x"38",
          6573 => x"77",
          6574 => x"70",
          6575 => x"2a",
          6576 => x"07",
          6577 => x"51",
          6578 => x"8f",
          6579 => x"84",
          6580 => x"83",
          6581 => x"94",
          6582 => x"74",
          6583 => x"38",
          6584 => x"0c",
          6585 => x"86",
          6586 => x"94",
          6587 => x"82",
          6588 => x"8c",
          6589 => x"fa",
          6590 => x"56",
          6591 => x"17",
          6592 => x"b0",
          6593 => x"52",
          6594 => x"e0",
          6595 => x"82",
          6596 => x"81",
          6597 => x"b2",
          6598 => x"b4",
          6599 => x"c8",
          6600 => x"ff",
          6601 => x"55",
          6602 => x"d5",
          6603 => x"06",
          6604 => x"80",
          6605 => x"33",
          6606 => x"81",
          6607 => x"81",
          6608 => x"81",
          6609 => x"eb",
          6610 => x"70",
          6611 => x"07",
          6612 => x"73",
          6613 => x"81",
          6614 => x"81",
          6615 => x"83",
          6616 => x"c0",
          6617 => x"16",
          6618 => x"3f",
          6619 => x"08",
          6620 => x"c8",
          6621 => x"9d",
          6622 => x"82",
          6623 => x"81",
          6624 => x"e0",
          6625 => x"b5",
          6626 => x"82",
          6627 => x"80",
          6628 => x"82",
          6629 => x"b5",
          6630 => x"3d",
          6631 => x"3d",
          6632 => x"84",
          6633 => x"05",
          6634 => x"80",
          6635 => x"51",
          6636 => x"82",
          6637 => x"58",
          6638 => x"0b",
          6639 => x"08",
          6640 => x"38",
          6641 => x"08",
          6642 => x"cd",
          6643 => x"08",
          6644 => x"56",
          6645 => x"86",
          6646 => x"75",
          6647 => x"fe",
          6648 => x"54",
          6649 => x"2e",
          6650 => x"14",
          6651 => x"ca",
          6652 => x"c8",
          6653 => x"06",
          6654 => x"54",
          6655 => x"38",
          6656 => x"86",
          6657 => x"82",
          6658 => x"06",
          6659 => x"56",
          6660 => x"38",
          6661 => x"80",
          6662 => x"81",
          6663 => x"52",
          6664 => x"51",
          6665 => x"82",
          6666 => x"81",
          6667 => x"81",
          6668 => x"83",
          6669 => x"87",
          6670 => x"2e",
          6671 => x"82",
          6672 => x"06",
          6673 => x"56",
          6674 => x"38",
          6675 => x"74",
          6676 => x"a3",
          6677 => x"c8",
          6678 => x"06",
          6679 => x"2e",
          6680 => x"80",
          6681 => x"3d",
          6682 => x"83",
          6683 => x"15",
          6684 => x"53",
          6685 => x"8d",
          6686 => x"15",
          6687 => x"3f",
          6688 => x"08",
          6689 => x"70",
          6690 => x"0c",
          6691 => x"16",
          6692 => x"80",
          6693 => x"80",
          6694 => x"54",
          6695 => x"84",
          6696 => x"5b",
          6697 => x"80",
          6698 => x"7a",
          6699 => x"fc",
          6700 => x"b5",
          6701 => x"ff",
          6702 => x"77",
          6703 => x"81",
          6704 => x"76",
          6705 => x"81",
          6706 => x"2e",
          6707 => x"8d",
          6708 => x"26",
          6709 => x"bf",
          6710 => x"f4",
          6711 => x"c8",
          6712 => x"ff",
          6713 => x"84",
          6714 => x"81",
          6715 => x"38",
          6716 => x"51",
          6717 => x"82",
          6718 => x"83",
          6719 => x"58",
          6720 => x"80",
          6721 => x"db",
          6722 => x"b5",
          6723 => x"77",
          6724 => x"80",
          6725 => x"82",
          6726 => x"c4",
          6727 => x"11",
          6728 => x"06",
          6729 => x"8d",
          6730 => x"26",
          6731 => x"74",
          6732 => x"78",
          6733 => x"c1",
          6734 => x"59",
          6735 => x"15",
          6736 => x"2e",
          6737 => x"13",
          6738 => x"72",
          6739 => x"38",
          6740 => x"eb",
          6741 => x"14",
          6742 => x"3f",
          6743 => x"08",
          6744 => x"c8",
          6745 => x"23",
          6746 => x"57",
          6747 => x"83",
          6748 => x"c7",
          6749 => x"d8",
          6750 => x"c8",
          6751 => x"ff",
          6752 => x"8d",
          6753 => x"14",
          6754 => x"3f",
          6755 => x"08",
          6756 => x"14",
          6757 => x"3f",
          6758 => x"08",
          6759 => x"06",
          6760 => x"72",
          6761 => x"97",
          6762 => x"22",
          6763 => x"84",
          6764 => x"5a",
          6765 => x"83",
          6766 => x"14",
          6767 => x"79",
          6768 => x"f3",
          6769 => x"b5",
          6770 => x"82",
          6771 => x"80",
          6772 => x"38",
          6773 => x"08",
          6774 => x"ff",
          6775 => x"38",
          6776 => x"83",
          6777 => x"83",
          6778 => x"74",
          6779 => x"85",
          6780 => x"89",
          6781 => x"76",
          6782 => x"c3",
          6783 => x"70",
          6784 => x"7b",
          6785 => x"73",
          6786 => x"17",
          6787 => x"ac",
          6788 => x"55",
          6789 => x"09",
          6790 => x"38",
          6791 => x"51",
          6792 => x"82",
          6793 => x"83",
          6794 => x"53",
          6795 => x"82",
          6796 => x"82",
          6797 => x"e0",
          6798 => x"ab",
          6799 => x"c8",
          6800 => x"0c",
          6801 => x"53",
          6802 => x"56",
          6803 => x"81",
          6804 => x"13",
          6805 => x"74",
          6806 => x"82",
          6807 => x"74",
          6808 => x"81",
          6809 => x"06",
          6810 => x"83",
          6811 => x"2a",
          6812 => x"72",
          6813 => x"26",
          6814 => x"ff",
          6815 => x"0c",
          6816 => x"15",
          6817 => x"0b",
          6818 => x"76",
          6819 => x"81",
          6820 => x"38",
          6821 => x"51",
          6822 => x"82",
          6823 => x"83",
          6824 => x"53",
          6825 => x"09",
          6826 => x"f9",
          6827 => x"52",
          6828 => x"b8",
          6829 => x"c8",
          6830 => x"38",
          6831 => x"08",
          6832 => x"84",
          6833 => x"d8",
          6834 => x"b5",
          6835 => x"ff",
          6836 => x"72",
          6837 => x"2e",
          6838 => x"80",
          6839 => x"14",
          6840 => x"3f",
          6841 => x"08",
          6842 => x"a4",
          6843 => x"81",
          6844 => x"84",
          6845 => x"d7",
          6846 => x"b5",
          6847 => x"8a",
          6848 => x"2e",
          6849 => x"9d",
          6850 => x"14",
          6851 => x"3f",
          6852 => x"08",
          6853 => x"84",
          6854 => x"d7",
          6855 => x"b5",
          6856 => x"15",
          6857 => x"34",
          6858 => x"22",
          6859 => x"72",
          6860 => x"23",
          6861 => x"23",
          6862 => x"15",
          6863 => x"75",
          6864 => x"0c",
          6865 => x"04",
          6866 => x"77",
          6867 => x"73",
          6868 => x"38",
          6869 => x"72",
          6870 => x"38",
          6871 => x"71",
          6872 => x"38",
          6873 => x"84",
          6874 => x"52",
          6875 => x"09",
          6876 => x"38",
          6877 => x"51",
          6878 => x"82",
          6879 => x"81",
          6880 => x"88",
          6881 => x"08",
          6882 => x"39",
          6883 => x"73",
          6884 => x"74",
          6885 => x"0c",
          6886 => x"04",
          6887 => x"02",
          6888 => x"7a",
          6889 => x"fc",
          6890 => x"f4",
          6891 => x"54",
          6892 => x"b5",
          6893 => x"bc",
          6894 => x"c8",
          6895 => x"82",
          6896 => x"70",
          6897 => x"73",
          6898 => x"38",
          6899 => x"78",
          6900 => x"2e",
          6901 => x"74",
          6902 => x"0c",
          6903 => x"80",
          6904 => x"80",
          6905 => x"70",
          6906 => x"51",
          6907 => x"82",
          6908 => x"54",
          6909 => x"c8",
          6910 => x"0d",
          6911 => x"0d",
          6912 => x"05",
          6913 => x"33",
          6914 => x"54",
          6915 => x"84",
          6916 => x"bf",
          6917 => x"98",
          6918 => x"53",
          6919 => x"05",
          6920 => x"fa",
          6921 => x"c8",
          6922 => x"b5",
          6923 => x"a4",
          6924 => x"68",
          6925 => x"70",
          6926 => x"c6",
          6927 => x"c8",
          6928 => x"b5",
          6929 => x"38",
          6930 => x"05",
          6931 => x"2b",
          6932 => x"80",
          6933 => x"86",
          6934 => x"06",
          6935 => x"2e",
          6936 => x"74",
          6937 => x"38",
          6938 => x"09",
          6939 => x"38",
          6940 => x"f8",
          6941 => x"c8",
          6942 => x"39",
          6943 => x"33",
          6944 => x"73",
          6945 => x"77",
          6946 => x"81",
          6947 => x"73",
          6948 => x"38",
          6949 => x"bc",
          6950 => x"07",
          6951 => x"b4",
          6952 => x"2a",
          6953 => x"51",
          6954 => x"2e",
          6955 => x"62",
          6956 => x"e8",
          6957 => x"b5",
          6958 => x"82",
          6959 => x"52",
          6960 => x"51",
          6961 => x"62",
          6962 => x"8b",
          6963 => x"53",
          6964 => x"51",
          6965 => x"80",
          6966 => x"05",
          6967 => x"3f",
          6968 => x"0b",
          6969 => x"75",
          6970 => x"f1",
          6971 => x"11",
          6972 => x"80",
          6973 => x"97",
          6974 => x"51",
          6975 => x"82",
          6976 => x"55",
          6977 => x"08",
          6978 => x"b7",
          6979 => x"c4",
          6980 => x"05",
          6981 => x"2a",
          6982 => x"51",
          6983 => x"80",
          6984 => x"84",
          6985 => x"39",
          6986 => x"70",
          6987 => x"54",
          6988 => x"a9",
          6989 => x"06",
          6990 => x"2e",
          6991 => x"55",
          6992 => x"73",
          6993 => x"d6",
          6994 => x"b5",
          6995 => x"ff",
          6996 => x"0c",
          6997 => x"b5",
          6998 => x"f8",
          6999 => x"2a",
          7000 => x"51",
          7001 => x"2e",
          7002 => x"80",
          7003 => x"7a",
          7004 => x"a0",
          7005 => x"a4",
          7006 => x"53",
          7007 => x"e6",
          7008 => x"b5",
          7009 => x"b5",
          7010 => x"1b",
          7011 => x"05",
          7012 => x"d3",
          7013 => x"c8",
          7014 => x"c8",
          7015 => x"0c",
          7016 => x"56",
          7017 => x"84",
          7018 => x"90",
          7019 => x"0b",
          7020 => x"80",
          7021 => x"0c",
          7022 => x"1a",
          7023 => x"2a",
          7024 => x"51",
          7025 => x"2e",
          7026 => x"82",
          7027 => x"80",
          7028 => x"38",
          7029 => x"08",
          7030 => x"8a",
          7031 => x"89",
          7032 => x"59",
          7033 => x"76",
          7034 => x"d7",
          7035 => x"b5",
          7036 => x"82",
          7037 => x"81",
          7038 => x"82",
          7039 => x"c8",
          7040 => x"09",
          7041 => x"38",
          7042 => x"78",
          7043 => x"30",
          7044 => x"80",
          7045 => x"77",
          7046 => x"38",
          7047 => x"06",
          7048 => x"c3",
          7049 => x"1a",
          7050 => x"38",
          7051 => x"06",
          7052 => x"2e",
          7053 => x"52",
          7054 => x"a6",
          7055 => x"c8",
          7056 => x"82",
          7057 => x"75",
          7058 => x"b5",
          7059 => x"9c",
          7060 => x"39",
          7061 => x"74",
          7062 => x"b5",
          7063 => x"3d",
          7064 => x"3d",
          7065 => x"65",
          7066 => x"5d",
          7067 => x"0c",
          7068 => x"05",
          7069 => x"f9",
          7070 => x"b5",
          7071 => x"82",
          7072 => x"8a",
          7073 => x"33",
          7074 => x"2e",
          7075 => x"56",
          7076 => x"90",
          7077 => x"06",
          7078 => x"74",
          7079 => x"b6",
          7080 => x"82",
          7081 => x"34",
          7082 => x"aa",
          7083 => x"91",
          7084 => x"56",
          7085 => x"8c",
          7086 => x"1a",
          7087 => x"74",
          7088 => x"38",
          7089 => x"80",
          7090 => x"38",
          7091 => x"70",
          7092 => x"56",
          7093 => x"b2",
          7094 => x"11",
          7095 => x"77",
          7096 => x"5b",
          7097 => x"38",
          7098 => x"88",
          7099 => x"8f",
          7100 => x"08",
          7101 => x"d5",
          7102 => x"b5",
          7103 => x"81",
          7104 => x"9f",
          7105 => x"2e",
          7106 => x"74",
          7107 => x"98",
          7108 => x"7e",
          7109 => x"3f",
          7110 => x"08",
          7111 => x"83",
          7112 => x"c8",
          7113 => x"89",
          7114 => x"77",
          7115 => x"d6",
          7116 => x"7f",
          7117 => x"58",
          7118 => x"75",
          7119 => x"75",
          7120 => x"77",
          7121 => x"7c",
          7122 => x"33",
          7123 => x"3f",
          7124 => x"08",
          7125 => x"7e",
          7126 => x"56",
          7127 => x"2e",
          7128 => x"16",
          7129 => x"55",
          7130 => x"94",
          7131 => x"53",
          7132 => x"b0",
          7133 => x"31",
          7134 => x"05",
          7135 => x"3f",
          7136 => x"56",
          7137 => x"9c",
          7138 => x"19",
          7139 => x"06",
          7140 => x"31",
          7141 => x"76",
          7142 => x"7b",
          7143 => x"08",
          7144 => x"d1",
          7145 => x"b5",
          7146 => x"81",
          7147 => x"94",
          7148 => x"ff",
          7149 => x"05",
          7150 => x"cf",
          7151 => x"76",
          7152 => x"17",
          7153 => x"1e",
          7154 => x"18",
          7155 => x"5e",
          7156 => x"39",
          7157 => x"82",
          7158 => x"90",
          7159 => x"f2",
          7160 => x"63",
          7161 => x"40",
          7162 => x"7e",
          7163 => x"fc",
          7164 => x"51",
          7165 => x"82",
          7166 => x"55",
          7167 => x"08",
          7168 => x"18",
          7169 => x"80",
          7170 => x"74",
          7171 => x"39",
          7172 => x"70",
          7173 => x"81",
          7174 => x"56",
          7175 => x"80",
          7176 => x"38",
          7177 => x"0b",
          7178 => x"82",
          7179 => x"39",
          7180 => x"19",
          7181 => x"83",
          7182 => x"18",
          7183 => x"56",
          7184 => x"27",
          7185 => x"09",
          7186 => x"2e",
          7187 => x"94",
          7188 => x"83",
          7189 => x"56",
          7190 => x"38",
          7191 => x"22",
          7192 => x"89",
          7193 => x"55",
          7194 => x"75",
          7195 => x"18",
          7196 => x"9c",
          7197 => x"85",
          7198 => x"08",
          7199 => x"d7",
          7200 => x"b5",
          7201 => x"82",
          7202 => x"80",
          7203 => x"38",
          7204 => x"ff",
          7205 => x"ff",
          7206 => x"38",
          7207 => x"0c",
          7208 => x"85",
          7209 => x"19",
          7210 => x"b0",
          7211 => x"19",
          7212 => x"81",
          7213 => x"74",
          7214 => x"3f",
          7215 => x"08",
          7216 => x"98",
          7217 => x"7e",
          7218 => x"3f",
          7219 => x"08",
          7220 => x"d2",
          7221 => x"c8",
          7222 => x"89",
          7223 => x"78",
          7224 => x"d5",
          7225 => x"7f",
          7226 => x"58",
          7227 => x"75",
          7228 => x"75",
          7229 => x"78",
          7230 => x"7c",
          7231 => x"33",
          7232 => x"3f",
          7233 => x"08",
          7234 => x"7e",
          7235 => x"78",
          7236 => x"74",
          7237 => x"38",
          7238 => x"b0",
          7239 => x"31",
          7240 => x"05",
          7241 => x"51",
          7242 => x"7e",
          7243 => x"83",
          7244 => x"89",
          7245 => x"db",
          7246 => x"08",
          7247 => x"26",
          7248 => x"51",
          7249 => x"82",
          7250 => x"fd",
          7251 => x"77",
          7252 => x"55",
          7253 => x"0c",
          7254 => x"83",
          7255 => x"80",
          7256 => x"55",
          7257 => x"83",
          7258 => x"9c",
          7259 => x"7e",
          7260 => x"3f",
          7261 => x"08",
          7262 => x"75",
          7263 => x"94",
          7264 => x"ff",
          7265 => x"05",
          7266 => x"3f",
          7267 => x"0b",
          7268 => x"7b",
          7269 => x"08",
          7270 => x"76",
          7271 => x"08",
          7272 => x"1c",
          7273 => x"08",
          7274 => x"5c",
          7275 => x"83",
          7276 => x"74",
          7277 => x"fd",
          7278 => x"18",
          7279 => x"07",
          7280 => x"19",
          7281 => x"75",
          7282 => x"0c",
          7283 => x"04",
          7284 => x"7a",
          7285 => x"05",
          7286 => x"56",
          7287 => x"82",
          7288 => x"57",
          7289 => x"08",
          7290 => x"90",
          7291 => x"86",
          7292 => x"06",
          7293 => x"73",
          7294 => x"e9",
          7295 => x"08",
          7296 => x"cc",
          7297 => x"b5",
          7298 => x"82",
          7299 => x"80",
          7300 => x"16",
          7301 => x"33",
          7302 => x"55",
          7303 => x"34",
          7304 => x"53",
          7305 => x"08",
          7306 => x"3f",
          7307 => x"52",
          7308 => x"c9",
          7309 => x"88",
          7310 => x"96",
          7311 => x"f0",
          7312 => x"92",
          7313 => x"ca",
          7314 => x"81",
          7315 => x"34",
          7316 => x"df",
          7317 => x"c8",
          7318 => x"33",
          7319 => x"55",
          7320 => x"17",
          7321 => x"b5",
          7322 => x"3d",
          7323 => x"3d",
          7324 => x"52",
          7325 => x"3f",
          7326 => x"08",
          7327 => x"c8",
          7328 => x"86",
          7329 => x"52",
          7330 => x"bc",
          7331 => x"c8",
          7332 => x"b5",
          7333 => x"38",
          7334 => x"08",
          7335 => x"82",
          7336 => x"86",
          7337 => x"ff",
          7338 => x"3d",
          7339 => x"3f",
          7340 => x"0b",
          7341 => x"08",
          7342 => x"82",
          7343 => x"82",
          7344 => x"80",
          7345 => x"b5",
          7346 => x"3d",
          7347 => x"3d",
          7348 => x"93",
          7349 => x"52",
          7350 => x"e9",
          7351 => x"b5",
          7352 => x"82",
          7353 => x"80",
          7354 => x"58",
          7355 => x"3d",
          7356 => x"e0",
          7357 => x"b5",
          7358 => x"82",
          7359 => x"bc",
          7360 => x"c7",
          7361 => x"98",
          7362 => x"73",
          7363 => x"38",
          7364 => x"12",
          7365 => x"39",
          7366 => x"33",
          7367 => x"70",
          7368 => x"55",
          7369 => x"2e",
          7370 => x"7f",
          7371 => x"54",
          7372 => x"82",
          7373 => x"94",
          7374 => x"39",
          7375 => x"08",
          7376 => x"81",
          7377 => x"85",
          7378 => x"b5",
          7379 => x"3d",
          7380 => x"3d",
          7381 => x"5b",
          7382 => x"34",
          7383 => x"3d",
          7384 => x"52",
          7385 => x"e8",
          7386 => x"b5",
          7387 => x"82",
          7388 => x"82",
          7389 => x"43",
          7390 => x"11",
          7391 => x"58",
          7392 => x"80",
          7393 => x"38",
          7394 => x"3d",
          7395 => x"d5",
          7396 => x"b5",
          7397 => x"82",
          7398 => x"82",
          7399 => x"52",
          7400 => x"c8",
          7401 => x"c8",
          7402 => x"b5",
          7403 => x"c1",
          7404 => x"7b",
          7405 => x"3f",
          7406 => x"08",
          7407 => x"74",
          7408 => x"3f",
          7409 => x"08",
          7410 => x"c8",
          7411 => x"38",
          7412 => x"51",
          7413 => x"82",
          7414 => x"57",
          7415 => x"08",
          7416 => x"52",
          7417 => x"f2",
          7418 => x"b5",
          7419 => x"a6",
          7420 => x"74",
          7421 => x"3f",
          7422 => x"08",
          7423 => x"c8",
          7424 => x"cc",
          7425 => x"2e",
          7426 => x"86",
          7427 => x"81",
          7428 => x"81",
          7429 => x"3d",
          7430 => x"52",
          7431 => x"c9",
          7432 => x"3d",
          7433 => x"11",
          7434 => x"5a",
          7435 => x"2e",
          7436 => x"b9",
          7437 => x"16",
          7438 => x"33",
          7439 => x"73",
          7440 => x"16",
          7441 => x"26",
          7442 => x"75",
          7443 => x"38",
          7444 => x"05",
          7445 => x"6f",
          7446 => x"ff",
          7447 => x"55",
          7448 => x"74",
          7449 => x"38",
          7450 => x"11",
          7451 => x"74",
          7452 => x"39",
          7453 => x"09",
          7454 => x"38",
          7455 => x"11",
          7456 => x"74",
          7457 => x"82",
          7458 => x"70",
          7459 => x"af",
          7460 => x"08",
          7461 => x"5c",
          7462 => x"73",
          7463 => x"38",
          7464 => x"1a",
          7465 => x"55",
          7466 => x"38",
          7467 => x"73",
          7468 => x"38",
          7469 => x"76",
          7470 => x"74",
          7471 => x"33",
          7472 => x"05",
          7473 => x"15",
          7474 => x"ba",
          7475 => x"05",
          7476 => x"ff",
          7477 => x"06",
          7478 => x"57",
          7479 => x"18",
          7480 => x"54",
          7481 => x"70",
          7482 => x"34",
          7483 => x"ee",
          7484 => x"34",
          7485 => x"c8",
          7486 => x"0d",
          7487 => x"0d",
          7488 => x"3d",
          7489 => x"71",
          7490 => x"ec",
          7491 => x"b5",
          7492 => x"82",
          7493 => x"82",
          7494 => x"15",
          7495 => x"82",
          7496 => x"15",
          7497 => x"76",
          7498 => x"90",
          7499 => x"81",
          7500 => x"06",
          7501 => x"72",
          7502 => x"56",
          7503 => x"54",
          7504 => x"17",
          7505 => x"78",
          7506 => x"38",
          7507 => x"22",
          7508 => x"59",
          7509 => x"78",
          7510 => x"76",
          7511 => x"51",
          7512 => x"3f",
          7513 => x"08",
          7514 => x"54",
          7515 => x"53",
          7516 => x"3f",
          7517 => x"08",
          7518 => x"38",
          7519 => x"75",
          7520 => x"18",
          7521 => x"31",
          7522 => x"57",
          7523 => x"b1",
          7524 => x"08",
          7525 => x"38",
          7526 => x"51",
          7527 => x"82",
          7528 => x"54",
          7529 => x"08",
          7530 => x"9a",
          7531 => x"c8",
          7532 => x"81",
          7533 => x"b5",
          7534 => x"16",
          7535 => x"16",
          7536 => x"2e",
          7537 => x"76",
          7538 => x"dc",
          7539 => x"31",
          7540 => x"18",
          7541 => x"90",
          7542 => x"81",
          7543 => x"06",
          7544 => x"56",
          7545 => x"9a",
          7546 => x"74",
          7547 => x"3f",
          7548 => x"08",
          7549 => x"c8",
          7550 => x"82",
          7551 => x"56",
          7552 => x"52",
          7553 => x"84",
          7554 => x"c8",
          7555 => x"ff",
          7556 => x"81",
          7557 => x"38",
          7558 => x"98",
          7559 => x"a6",
          7560 => x"16",
          7561 => x"39",
          7562 => x"16",
          7563 => x"75",
          7564 => x"53",
          7565 => x"aa",
          7566 => x"79",
          7567 => x"3f",
          7568 => x"08",
          7569 => x"0b",
          7570 => x"82",
          7571 => x"39",
          7572 => x"16",
          7573 => x"bb",
          7574 => x"2a",
          7575 => x"08",
          7576 => x"15",
          7577 => x"15",
          7578 => x"90",
          7579 => x"16",
          7580 => x"33",
          7581 => x"53",
          7582 => x"34",
          7583 => x"06",
          7584 => x"2e",
          7585 => x"9c",
          7586 => x"85",
          7587 => x"16",
          7588 => x"72",
          7589 => x"0c",
          7590 => x"04",
          7591 => x"79",
          7592 => x"75",
          7593 => x"8a",
          7594 => x"89",
          7595 => x"52",
          7596 => x"05",
          7597 => x"3f",
          7598 => x"08",
          7599 => x"c8",
          7600 => x"38",
          7601 => x"7a",
          7602 => x"d8",
          7603 => x"b5",
          7604 => x"82",
          7605 => x"80",
          7606 => x"16",
          7607 => x"2b",
          7608 => x"74",
          7609 => x"86",
          7610 => x"84",
          7611 => x"06",
          7612 => x"73",
          7613 => x"38",
          7614 => x"52",
          7615 => x"da",
          7616 => x"c8",
          7617 => x"0c",
          7618 => x"14",
          7619 => x"23",
          7620 => x"51",
          7621 => x"82",
          7622 => x"55",
          7623 => x"09",
          7624 => x"38",
          7625 => x"39",
          7626 => x"84",
          7627 => x"0c",
          7628 => x"82",
          7629 => x"89",
          7630 => x"fc",
          7631 => x"87",
          7632 => x"53",
          7633 => x"e7",
          7634 => x"b5",
          7635 => x"38",
          7636 => x"08",
          7637 => x"3d",
          7638 => x"3d",
          7639 => x"89",
          7640 => x"54",
          7641 => x"54",
          7642 => x"82",
          7643 => x"53",
          7644 => x"08",
          7645 => x"74",
          7646 => x"b5",
          7647 => x"73",
          7648 => x"3f",
          7649 => x"08",
          7650 => x"39",
          7651 => x"08",
          7652 => x"d3",
          7653 => x"b5",
          7654 => x"82",
          7655 => x"84",
          7656 => x"06",
          7657 => x"53",
          7658 => x"b5",
          7659 => x"38",
          7660 => x"51",
          7661 => x"72",
          7662 => x"cf",
          7663 => x"b5",
          7664 => x"32",
          7665 => x"72",
          7666 => x"70",
          7667 => x"08",
          7668 => x"54",
          7669 => x"b5",
          7670 => x"3d",
          7671 => x"3d",
          7672 => x"80",
          7673 => x"70",
          7674 => x"52",
          7675 => x"3f",
          7676 => x"08",
          7677 => x"c8",
          7678 => x"64",
          7679 => x"d6",
          7680 => x"b5",
          7681 => x"82",
          7682 => x"a0",
          7683 => x"cb",
          7684 => x"98",
          7685 => x"73",
          7686 => x"38",
          7687 => x"39",
          7688 => x"88",
          7689 => x"75",
          7690 => x"3f",
          7691 => x"c8",
          7692 => x"0d",
          7693 => x"0d",
          7694 => x"5c",
          7695 => x"3d",
          7696 => x"93",
          7697 => x"d6",
          7698 => x"c8",
          7699 => x"b5",
          7700 => x"80",
          7701 => x"0c",
          7702 => x"11",
          7703 => x"90",
          7704 => x"56",
          7705 => x"74",
          7706 => x"75",
          7707 => x"e4",
          7708 => x"81",
          7709 => x"5b",
          7710 => x"82",
          7711 => x"75",
          7712 => x"73",
          7713 => x"81",
          7714 => x"82",
          7715 => x"76",
          7716 => x"f0",
          7717 => x"f4",
          7718 => x"c8",
          7719 => x"d1",
          7720 => x"c8",
          7721 => x"ce",
          7722 => x"c8",
          7723 => x"82",
          7724 => x"07",
          7725 => x"05",
          7726 => x"53",
          7727 => x"98",
          7728 => x"26",
          7729 => x"f9",
          7730 => x"08",
          7731 => x"08",
          7732 => x"98",
          7733 => x"81",
          7734 => x"58",
          7735 => x"3f",
          7736 => x"08",
          7737 => x"c8",
          7738 => x"38",
          7739 => x"77",
          7740 => x"5d",
          7741 => x"74",
          7742 => x"81",
          7743 => x"b4",
          7744 => x"bb",
          7745 => x"b5",
          7746 => x"ff",
          7747 => x"30",
          7748 => x"1b",
          7749 => x"5b",
          7750 => x"39",
          7751 => x"ff",
          7752 => x"82",
          7753 => x"f0",
          7754 => x"30",
          7755 => x"1b",
          7756 => x"5b",
          7757 => x"83",
          7758 => x"58",
          7759 => x"92",
          7760 => x"0c",
          7761 => x"12",
          7762 => x"33",
          7763 => x"54",
          7764 => x"34",
          7765 => x"c8",
          7766 => x"0d",
          7767 => x"0d",
          7768 => x"fc",
          7769 => x"52",
          7770 => x"3f",
          7771 => x"08",
          7772 => x"c8",
          7773 => x"38",
          7774 => x"56",
          7775 => x"38",
          7776 => x"70",
          7777 => x"81",
          7778 => x"55",
          7779 => x"80",
          7780 => x"38",
          7781 => x"54",
          7782 => x"08",
          7783 => x"38",
          7784 => x"82",
          7785 => x"53",
          7786 => x"52",
          7787 => x"8c",
          7788 => x"c8",
          7789 => x"19",
          7790 => x"c9",
          7791 => x"08",
          7792 => x"ff",
          7793 => x"82",
          7794 => x"ff",
          7795 => x"06",
          7796 => x"56",
          7797 => x"08",
          7798 => x"81",
          7799 => x"82",
          7800 => x"75",
          7801 => x"54",
          7802 => x"08",
          7803 => x"27",
          7804 => x"17",
          7805 => x"b5",
          7806 => x"76",
          7807 => x"3f",
          7808 => x"08",
          7809 => x"08",
          7810 => x"90",
          7811 => x"c0",
          7812 => x"90",
          7813 => x"80",
          7814 => x"75",
          7815 => x"75",
          7816 => x"b5",
          7817 => x"3d",
          7818 => x"3d",
          7819 => x"a0",
          7820 => x"05",
          7821 => x"51",
          7822 => x"82",
          7823 => x"55",
          7824 => x"08",
          7825 => x"78",
          7826 => x"08",
          7827 => x"70",
          7828 => x"ae",
          7829 => x"c8",
          7830 => x"b5",
          7831 => x"db",
          7832 => x"fb",
          7833 => x"85",
          7834 => x"06",
          7835 => x"86",
          7836 => x"c7",
          7837 => x"2b",
          7838 => x"24",
          7839 => x"02",
          7840 => x"33",
          7841 => x"58",
          7842 => x"76",
          7843 => x"6b",
          7844 => x"cc",
          7845 => x"b5",
          7846 => x"84",
          7847 => x"06",
          7848 => x"73",
          7849 => x"d4",
          7850 => x"82",
          7851 => x"94",
          7852 => x"81",
          7853 => x"5a",
          7854 => x"08",
          7855 => x"8a",
          7856 => x"54",
          7857 => x"82",
          7858 => x"55",
          7859 => x"08",
          7860 => x"82",
          7861 => x"52",
          7862 => x"e5",
          7863 => x"c8",
          7864 => x"b5",
          7865 => x"38",
          7866 => x"cf",
          7867 => x"c8",
          7868 => x"88",
          7869 => x"c8",
          7870 => x"38",
          7871 => x"c2",
          7872 => x"c8",
          7873 => x"c8",
          7874 => x"82",
          7875 => x"07",
          7876 => x"55",
          7877 => x"2e",
          7878 => x"80",
          7879 => x"80",
          7880 => x"77",
          7881 => x"3f",
          7882 => x"08",
          7883 => x"38",
          7884 => x"ba",
          7885 => x"b5",
          7886 => x"74",
          7887 => x"0c",
          7888 => x"04",
          7889 => x"82",
          7890 => x"c0",
          7891 => x"3d",
          7892 => x"3f",
          7893 => x"08",
          7894 => x"c8",
          7895 => x"38",
          7896 => x"52",
          7897 => x"52",
          7898 => x"3f",
          7899 => x"08",
          7900 => x"c8",
          7901 => x"88",
          7902 => x"39",
          7903 => x"08",
          7904 => x"81",
          7905 => x"38",
          7906 => x"05",
          7907 => x"2a",
          7908 => x"55",
          7909 => x"81",
          7910 => x"5a",
          7911 => x"3d",
          7912 => x"c1",
          7913 => x"b5",
          7914 => x"55",
          7915 => x"c8",
          7916 => x"87",
          7917 => x"c8",
          7918 => x"09",
          7919 => x"38",
          7920 => x"b5",
          7921 => x"2e",
          7922 => x"86",
          7923 => x"81",
          7924 => x"81",
          7925 => x"b5",
          7926 => x"78",
          7927 => x"3f",
          7928 => x"08",
          7929 => x"c8",
          7930 => x"38",
          7931 => x"52",
          7932 => x"ff",
          7933 => x"78",
          7934 => x"b4",
          7935 => x"54",
          7936 => x"15",
          7937 => x"b2",
          7938 => x"ca",
          7939 => x"b6",
          7940 => x"53",
          7941 => x"53",
          7942 => x"3f",
          7943 => x"b4",
          7944 => x"d4",
          7945 => x"b6",
          7946 => x"54",
          7947 => x"d5",
          7948 => x"53",
          7949 => x"11",
          7950 => x"d7",
          7951 => x"81",
          7952 => x"34",
          7953 => x"a4",
          7954 => x"c8",
          7955 => x"b5",
          7956 => x"38",
          7957 => x"0a",
          7958 => x"05",
          7959 => x"d0",
          7960 => x"64",
          7961 => x"c9",
          7962 => x"54",
          7963 => x"15",
          7964 => x"81",
          7965 => x"34",
          7966 => x"b8",
          7967 => x"b5",
          7968 => x"8b",
          7969 => x"75",
          7970 => x"ff",
          7971 => x"73",
          7972 => x"0c",
          7973 => x"04",
          7974 => x"a9",
          7975 => x"51",
          7976 => x"82",
          7977 => x"ff",
          7978 => x"a9",
          7979 => x"ee",
          7980 => x"c8",
          7981 => x"b5",
          7982 => x"d3",
          7983 => x"a9",
          7984 => x"9d",
          7985 => x"58",
          7986 => x"82",
          7987 => x"55",
          7988 => x"08",
          7989 => x"02",
          7990 => x"33",
          7991 => x"54",
          7992 => x"82",
          7993 => x"53",
          7994 => x"52",
          7995 => x"88",
          7996 => x"b4",
          7997 => x"53",
          7998 => x"3d",
          7999 => x"ff",
          8000 => x"aa",
          8001 => x"73",
          8002 => x"3f",
          8003 => x"08",
          8004 => x"c8",
          8005 => x"63",
          8006 => x"81",
          8007 => x"65",
          8008 => x"2e",
          8009 => x"55",
          8010 => x"82",
          8011 => x"84",
          8012 => x"06",
          8013 => x"73",
          8014 => x"3f",
          8015 => x"08",
          8016 => x"c8",
          8017 => x"38",
          8018 => x"53",
          8019 => x"95",
          8020 => x"16",
          8021 => x"87",
          8022 => x"05",
          8023 => x"34",
          8024 => x"70",
          8025 => x"81",
          8026 => x"55",
          8027 => x"74",
          8028 => x"73",
          8029 => x"78",
          8030 => x"83",
          8031 => x"16",
          8032 => x"2a",
          8033 => x"51",
          8034 => x"80",
          8035 => x"38",
          8036 => x"80",
          8037 => x"52",
          8038 => x"be",
          8039 => x"c8",
          8040 => x"51",
          8041 => x"3f",
          8042 => x"b5",
          8043 => x"2e",
          8044 => x"82",
          8045 => x"52",
          8046 => x"b5",
          8047 => x"b5",
          8048 => x"80",
          8049 => x"58",
          8050 => x"c8",
          8051 => x"38",
          8052 => x"54",
          8053 => x"09",
          8054 => x"38",
          8055 => x"52",
          8056 => x"af",
          8057 => x"81",
          8058 => x"34",
          8059 => x"b5",
          8060 => x"38",
          8061 => x"ca",
          8062 => x"c8",
          8063 => x"b5",
          8064 => x"38",
          8065 => x"b5",
          8066 => x"b5",
          8067 => x"74",
          8068 => x"0c",
          8069 => x"04",
          8070 => x"02",
          8071 => x"33",
          8072 => x"80",
          8073 => x"57",
          8074 => x"95",
          8075 => x"52",
          8076 => x"d2",
          8077 => x"b5",
          8078 => x"82",
          8079 => x"80",
          8080 => x"5a",
          8081 => x"3d",
          8082 => x"c9",
          8083 => x"b5",
          8084 => x"82",
          8085 => x"b8",
          8086 => x"cf",
          8087 => x"a0",
          8088 => x"55",
          8089 => x"75",
          8090 => x"71",
          8091 => x"33",
          8092 => x"74",
          8093 => x"57",
          8094 => x"8b",
          8095 => x"54",
          8096 => x"15",
          8097 => x"ff",
          8098 => x"82",
          8099 => x"55",
          8100 => x"c8",
          8101 => x"0d",
          8102 => x"0d",
          8103 => x"53",
          8104 => x"05",
          8105 => x"51",
          8106 => x"82",
          8107 => x"55",
          8108 => x"08",
          8109 => x"76",
          8110 => x"93",
          8111 => x"51",
          8112 => x"82",
          8113 => x"55",
          8114 => x"08",
          8115 => x"80",
          8116 => x"81",
          8117 => x"86",
          8118 => x"38",
          8119 => x"86",
          8120 => x"90",
          8121 => x"54",
          8122 => x"ff",
          8123 => x"76",
          8124 => x"83",
          8125 => x"51",
          8126 => x"3f",
          8127 => x"08",
          8128 => x"b5",
          8129 => x"3d",
          8130 => x"3d",
          8131 => x"5c",
          8132 => x"98",
          8133 => x"52",
          8134 => x"d1",
          8135 => x"b5",
          8136 => x"b5",
          8137 => x"70",
          8138 => x"08",
          8139 => x"51",
          8140 => x"80",
          8141 => x"38",
          8142 => x"06",
          8143 => x"80",
          8144 => x"38",
          8145 => x"5f",
          8146 => x"3d",
          8147 => x"ff",
          8148 => x"82",
          8149 => x"57",
          8150 => x"08",
          8151 => x"74",
          8152 => x"c3",
          8153 => x"b5",
          8154 => x"82",
          8155 => x"bf",
          8156 => x"c8",
          8157 => x"c8",
          8158 => x"59",
          8159 => x"81",
          8160 => x"56",
          8161 => x"33",
          8162 => x"16",
          8163 => x"27",
          8164 => x"56",
          8165 => x"80",
          8166 => x"80",
          8167 => x"ff",
          8168 => x"70",
          8169 => x"56",
          8170 => x"e8",
          8171 => x"76",
          8172 => x"81",
          8173 => x"80",
          8174 => x"57",
          8175 => x"78",
          8176 => x"51",
          8177 => x"2e",
          8178 => x"73",
          8179 => x"38",
          8180 => x"08",
          8181 => x"b1",
          8182 => x"b5",
          8183 => x"82",
          8184 => x"a7",
          8185 => x"33",
          8186 => x"c3",
          8187 => x"2e",
          8188 => x"e4",
          8189 => x"2e",
          8190 => x"56",
          8191 => x"05",
          8192 => x"e3",
          8193 => x"c8",
          8194 => x"76",
          8195 => x"0c",
          8196 => x"04",
          8197 => x"82",
          8198 => x"ff",
          8199 => x"9d",
          8200 => x"fa",
          8201 => x"c8",
          8202 => x"c8",
          8203 => x"82",
          8204 => x"83",
          8205 => x"53",
          8206 => x"3d",
          8207 => x"ff",
          8208 => x"73",
          8209 => x"70",
          8210 => x"52",
          8211 => x"9f",
          8212 => x"bc",
          8213 => x"74",
          8214 => x"6d",
          8215 => x"70",
          8216 => x"af",
          8217 => x"b5",
          8218 => x"2e",
          8219 => x"70",
          8220 => x"57",
          8221 => x"fd",
          8222 => x"c8",
          8223 => x"8d",
          8224 => x"2b",
          8225 => x"81",
          8226 => x"86",
          8227 => x"c8",
          8228 => x"9f",
          8229 => x"ff",
          8230 => x"54",
          8231 => x"8a",
          8232 => x"70",
          8233 => x"06",
          8234 => x"ff",
          8235 => x"38",
          8236 => x"15",
          8237 => x"80",
          8238 => x"74",
          8239 => x"90",
          8240 => x"89",
          8241 => x"c8",
          8242 => x"81",
          8243 => x"88",
          8244 => x"26",
          8245 => x"39",
          8246 => x"86",
          8247 => x"81",
          8248 => x"ff",
          8249 => x"38",
          8250 => x"54",
          8251 => x"81",
          8252 => x"81",
          8253 => x"78",
          8254 => x"5a",
          8255 => x"6d",
          8256 => x"81",
          8257 => x"57",
          8258 => x"9f",
          8259 => x"38",
          8260 => x"54",
          8261 => x"81",
          8262 => x"b1",
          8263 => x"2e",
          8264 => x"a7",
          8265 => x"15",
          8266 => x"54",
          8267 => x"09",
          8268 => x"38",
          8269 => x"76",
          8270 => x"41",
          8271 => x"52",
          8272 => x"52",
          8273 => x"b3",
          8274 => x"c8",
          8275 => x"b5",
          8276 => x"f7",
          8277 => x"74",
          8278 => x"e5",
          8279 => x"c8",
          8280 => x"b5",
          8281 => x"38",
          8282 => x"38",
          8283 => x"74",
          8284 => x"39",
          8285 => x"08",
          8286 => x"81",
          8287 => x"38",
          8288 => x"74",
          8289 => x"38",
          8290 => x"51",
          8291 => x"3f",
          8292 => x"08",
          8293 => x"c8",
          8294 => x"a0",
          8295 => x"c8",
          8296 => x"51",
          8297 => x"3f",
          8298 => x"0b",
          8299 => x"8b",
          8300 => x"67",
          8301 => x"a7",
          8302 => x"81",
          8303 => x"34",
          8304 => x"ad",
          8305 => x"b5",
          8306 => x"73",
          8307 => x"b5",
          8308 => x"3d",
          8309 => x"3d",
          8310 => x"02",
          8311 => x"cb",
          8312 => x"3d",
          8313 => x"72",
          8314 => x"5a",
          8315 => x"82",
          8316 => x"58",
          8317 => x"08",
          8318 => x"91",
          8319 => x"77",
          8320 => x"7c",
          8321 => x"38",
          8322 => x"59",
          8323 => x"90",
          8324 => x"81",
          8325 => x"06",
          8326 => x"73",
          8327 => x"54",
          8328 => x"82",
          8329 => x"39",
          8330 => x"8b",
          8331 => x"11",
          8332 => x"2b",
          8333 => x"54",
          8334 => x"fe",
          8335 => x"ff",
          8336 => x"70",
          8337 => x"07",
          8338 => x"b5",
          8339 => x"8c",
          8340 => x"40",
          8341 => x"55",
          8342 => x"88",
          8343 => x"08",
          8344 => x"38",
          8345 => x"77",
          8346 => x"56",
          8347 => x"51",
          8348 => x"3f",
          8349 => x"55",
          8350 => x"08",
          8351 => x"38",
          8352 => x"b5",
          8353 => x"2e",
          8354 => x"82",
          8355 => x"ff",
          8356 => x"38",
          8357 => x"08",
          8358 => x"16",
          8359 => x"2e",
          8360 => x"87",
          8361 => x"74",
          8362 => x"74",
          8363 => x"81",
          8364 => x"38",
          8365 => x"ff",
          8366 => x"2e",
          8367 => x"7b",
          8368 => x"80",
          8369 => x"81",
          8370 => x"81",
          8371 => x"06",
          8372 => x"56",
          8373 => x"52",
          8374 => x"af",
          8375 => x"b5",
          8376 => x"82",
          8377 => x"80",
          8378 => x"81",
          8379 => x"56",
          8380 => x"d3",
          8381 => x"ff",
          8382 => x"7c",
          8383 => x"55",
          8384 => x"b3",
          8385 => x"1b",
          8386 => x"1b",
          8387 => x"33",
          8388 => x"54",
          8389 => x"34",
          8390 => x"fe",
          8391 => x"08",
          8392 => x"74",
          8393 => x"75",
          8394 => x"16",
          8395 => x"33",
          8396 => x"73",
          8397 => x"77",
          8398 => x"b5",
          8399 => x"3d",
          8400 => x"3d",
          8401 => x"02",
          8402 => x"eb",
          8403 => x"3d",
          8404 => x"59",
          8405 => x"8b",
          8406 => x"82",
          8407 => x"24",
          8408 => x"82",
          8409 => x"84",
          8410 => x"80",
          8411 => x"51",
          8412 => x"2e",
          8413 => x"75",
          8414 => x"c8",
          8415 => x"06",
          8416 => x"7e",
          8417 => x"d0",
          8418 => x"c8",
          8419 => x"06",
          8420 => x"56",
          8421 => x"74",
          8422 => x"76",
          8423 => x"81",
          8424 => x"8a",
          8425 => x"b2",
          8426 => x"fc",
          8427 => x"52",
          8428 => x"a4",
          8429 => x"b5",
          8430 => x"38",
          8431 => x"80",
          8432 => x"74",
          8433 => x"26",
          8434 => x"15",
          8435 => x"74",
          8436 => x"38",
          8437 => x"80",
          8438 => x"84",
          8439 => x"92",
          8440 => x"80",
          8441 => x"38",
          8442 => x"06",
          8443 => x"2e",
          8444 => x"56",
          8445 => x"78",
          8446 => x"89",
          8447 => x"2b",
          8448 => x"43",
          8449 => x"38",
          8450 => x"30",
          8451 => x"77",
          8452 => x"91",
          8453 => x"c2",
          8454 => x"f8",
          8455 => x"52",
          8456 => x"a4",
          8457 => x"56",
          8458 => x"08",
          8459 => x"77",
          8460 => x"77",
          8461 => x"c8",
          8462 => x"45",
          8463 => x"bf",
          8464 => x"8e",
          8465 => x"26",
          8466 => x"74",
          8467 => x"48",
          8468 => x"75",
          8469 => x"38",
          8470 => x"81",
          8471 => x"fa",
          8472 => x"2a",
          8473 => x"56",
          8474 => x"2e",
          8475 => x"87",
          8476 => x"82",
          8477 => x"38",
          8478 => x"55",
          8479 => x"83",
          8480 => x"81",
          8481 => x"56",
          8482 => x"80",
          8483 => x"38",
          8484 => x"83",
          8485 => x"06",
          8486 => x"78",
          8487 => x"91",
          8488 => x"0b",
          8489 => x"22",
          8490 => x"80",
          8491 => x"74",
          8492 => x"38",
          8493 => x"56",
          8494 => x"17",
          8495 => x"57",
          8496 => x"2e",
          8497 => x"75",
          8498 => x"79",
          8499 => x"fe",
          8500 => x"82",
          8501 => x"84",
          8502 => x"05",
          8503 => x"5e",
          8504 => x"80",
          8505 => x"c8",
          8506 => x"8a",
          8507 => x"fd",
          8508 => x"75",
          8509 => x"38",
          8510 => x"78",
          8511 => x"8c",
          8512 => x"0b",
          8513 => x"22",
          8514 => x"80",
          8515 => x"74",
          8516 => x"38",
          8517 => x"56",
          8518 => x"17",
          8519 => x"57",
          8520 => x"2e",
          8521 => x"75",
          8522 => x"79",
          8523 => x"fe",
          8524 => x"82",
          8525 => x"10",
          8526 => x"82",
          8527 => x"9f",
          8528 => x"38",
          8529 => x"b5",
          8530 => x"82",
          8531 => x"05",
          8532 => x"2a",
          8533 => x"56",
          8534 => x"17",
          8535 => x"81",
          8536 => x"60",
          8537 => x"65",
          8538 => x"12",
          8539 => x"30",
          8540 => x"74",
          8541 => x"59",
          8542 => x"7d",
          8543 => x"81",
          8544 => x"76",
          8545 => x"41",
          8546 => x"76",
          8547 => x"90",
          8548 => x"62",
          8549 => x"51",
          8550 => x"26",
          8551 => x"75",
          8552 => x"31",
          8553 => x"65",
          8554 => x"fe",
          8555 => x"82",
          8556 => x"58",
          8557 => x"09",
          8558 => x"38",
          8559 => x"08",
          8560 => x"26",
          8561 => x"78",
          8562 => x"79",
          8563 => x"78",
          8564 => x"86",
          8565 => x"82",
          8566 => x"06",
          8567 => x"83",
          8568 => x"82",
          8569 => x"27",
          8570 => x"8f",
          8571 => x"55",
          8572 => x"26",
          8573 => x"59",
          8574 => x"62",
          8575 => x"74",
          8576 => x"38",
          8577 => x"88",
          8578 => x"c8",
          8579 => x"26",
          8580 => x"86",
          8581 => x"1a",
          8582 => x"79",
          8583 => x"38",
          8584 => x"80",
          8585 => x"2e",
          8586 => x"83",
          8587 => x"9f",
          8588 => x"8b",
          8589 => x"06",
          8590 => x"74",
          8591 => x"84",
          8592 => x"52",
          8593 => x"a2",
          8594 => x"53",
          8595 => x"52",
          8596 => x"a2",
          8597 => x"80",
          8598 => x"51",
          8599 => x"3f",
          8600 => x"34",
          8601 => x"ff",
          8602 => x"1b",
          8603 => x"a2",
          8604 => x"90",
          8605 => x"83",
          8606 => x"70",
          8607 => x"80",
          8608 => x"55",
          8609 => x"ff",
          8610 => x"66",
          8611 => x"ff",
          8612 => x"38",
          8613 => x"ff",
          8614 => x"1b",
          8615 => x"f2",
          8616 => x"74",
          8617 => x"51",
          8618 => x"3f",
          8619 => x"1c",
          8620 => x"98",
          8621 => x"a0",
          8622 => x"ff",
          8623 => x"51",
          8624 => x"3f",
          8625 => x"1b",
          8626 => x"e4",
          8627 => x"2e",
          8628 => x"80",
          8629 => x"88",
          8630 => x"80",
          8631 => x"ff",
          8632 => x"7c",
          8633 => x"51",
          8634 => x"3f",
          8635 => x"1b",
          8636 => x"bc",
          8637 => x"b0",
          8638 => x"a0",
          8639 => x"52",
          8640 => x"ff",
          8641 => x"ff",
          8642 => x"c0",
          8643 => x"0b",
          8644 => x"34",
          8645 => x"ae",
          8646 => x"c7",
          8647 => x"39",
          8648 => x"0a",
          8649 => x"51",
          8650 => x"3f",
          8651 => x"ff",
          8652 => x"1b",
          8653 => x"da",
          8654 => x"0b",
          8655 => x"a9",
          8656 => x"34",
          8657 => x"ae",
          8658 => x"1b",
          8659 => x"8f",
          8660 => x"d5",
          8661 => x"1b",
          8662 => x"ff",
          8663 => x"81",
          8664 => x"7a",
          8665 => x"ff",
          8666 => x"81",
          8667 => x"c8",
          8668 => x"38",
          8669 => x"09",
          8670 => x"ee",
          8671 => x"60",
          8672 => x"7a",
          8673 => x"ff",
          8674 => x"84",
          8675 => x"52",
          8676 => x"9f",
          8677 => x"8b",
          8678 => x"52",
          8679 => x"9f",
          8680 => x"8a",
          8681 => x"52",
          8682 => x"51",
          8683 => x"3f",
          8684 => x"83",
          8685 => x"ff",
          8686 => x"82",
          8687 => x"1b",
          8688 => x"ec",
          8689 => x"d5",
          8690 => x"ff",
          8691 => x"75",
          8692 => x"05",
          8693 => x"7e",
          8694 => x"e5",
          8695 => x"60",
          8696 => x"52",
          8697 => x"9a",
          8698 => x"53",
          8699 => x"51",
          8700 => x"3f",
          8701 => x"58",
          8702 => x"09",
          8703 => x"38",
          8704 => x"51",
          8705 => x"3f",
          8706 => x"1b",
          8707 => x"a0",
          8708 => x"52",
          8709 => x"91",
          8710 => x"ff",
          8711 => x"81",
          8712 => x"f8",
          8713 => x"7a",
          8714 => x"84",
          8715 => x"61",
          8716 => x"26",
          8717 => x"57",
          8718 => x"53",
          8719 => x"51",
          8720 => x"3f",
          8721 => x"08",
          8722 => x"84",
          8723 => x"b5",
          8724 => x"7a",
          8725 => x"aa",
          8726 => x"75",
          8727 => x"56",
          8728 => x"81",
          8729 => x"80",
          8730 => x"38",
          8731 => x"83",
          8732 => x"63",
          8733 => x"74",
          8734 => x"38",
          8735 => x"54",
          8736 => x"52",
          8737 => x"99",
          8738 => x"b5",
          8739 => x"c1",
          8740 => x"75",
          8741 => x"56",
          8742 => x"8c",
          8743 => x"2e",
          8744 => x"56",
          8745 => x"ff",
          8746 => x"84",
          8747 => x"2e",
          8748 => x"56",
          8749 => x"58",
          8750 => x"38",
          8751 => x"77",
          8752 => x"ff",
          8753 => x"82",
          8754 => x"78",
          8755 => x"c2",
          8756 => x"1b",
          8757 => x"34",
          8758 => x"16",
          8759 => x"82",
          8760 => x"83",
          8761 => x"84",
          8762 => x"67",
          8763 => x"fd",
          8764 => x"51",
          8765 => x"3f",
          8766 => x"16",
          8767 => x"c8",
          8768 => x"bf",
          8769 => x"86",
          8770 => x"b5",
          8771 => x"16",
          8772 => x"83",
          8773 => x"ff",
          8774 => x"66",
          8775 => x"1b",
          8776 => x"8c",
          8777 => x"77",
          8778 => x"7e",
          8779 => x"91",
          8780 => x"82",
          8781 => x"a2",
          8782 => x"80",
          8783 => x"ff",
          8784 => x"81",
          8785 => x"c8",
          8786 => x"89",
          8787 => x"8a",
          8788 => x"86",
          8789 => x"c8",
          8790 => x"82",
          8791 => x"99",
          8792 => x"f5",
          8793 => x"60",
          8794 => x"79",
          8795 => x"5a",
          8796 => x"78",
          8797 => x"8d",
          8798 => x"55",
          8799 => x"fc",
          8800 => x"51",
          8801 => x"7a",
          8802 => x"81",
          8803 => x"8c",
          8804 => x"74",
          8805 => x"38",
          8806 => x"81",
          8807 => x"81",
          8808 => x"8a",
          8809 => x"06",
          8810 => x"76",
          8811 => x"76",
          8812 => x"55",
          8813 => x"c8",
          8814 => x"0d",
          8815 => x"0d",
          8816 => x"05",
          8817 => x"59",
          8818 => x"2e",
          8819 => x"87",
          8820 => x"76",
          8821 => x"84",
          8822 => x"80",
          8823 => x"38",
          8824 => x"77",
          8825 => x"56",
          8826 => x"34",
          8827 => x"bb",
          8828 => x"38",
          8829 => x"05",
          8830 => x"8c",
          8831 => x"08",
          8832 => x"3f",
          8833 => x"70",
          8834 => x"07",
          8835 => x"30",
          8836 => x"56",
          8837 => x"0c",
          8838 => x"18",
          8839 => x"0d",
          8840 => x"0d",
          8841 => x"08",
          8842 => x"75",
          8843 => x"89",
          8844 => x"54",
          8845 => x"16",
          8846 => x"51",
          8847 => x"82",
          8848 => x"91",
          8849 => x"08",
          8850 => x"81",
          8851 => x"88",
          8852 => x"83",
          8853 => x"74",
          8854 => x"0c",
          8855 => x"04",
          8856 => x"75",
          8857 => x"53",
          8858 => x"51",
          8859 => x"3f",
          8860 => x"85",
          8861 => x"ea",
          8862 => x"80",
          8863 => x"6a",
          8864 => x"70",
          8865 => x"d8",
          8866 => x"72",
          8867 => x"3f",
          8868 => x"8d",
          8869 => x"0d",
          8870 => x"ff",
          8871 => x"ff",
          8872 => x"00",
          8873 => x"ff",
          8874 => x"2b",
          8875 => x"2b",
          8876 => x"2b",
          8877 => x"2b",
          8878 => x"2b",
          8879 => x"2b",
          8880 => x"2b",
          8881 => x"2b",
          8882 => x"2b",
          8883 => x"2b",
          8884 => x"2b",
          8885 => x"2b",
          8886 => x"2b",
          8887 => x"2b",
          8888 => x"2b",
          8889 => x"2b",
          8890 => x"2b",
          8891 => x"2b",
          8892 => x"2b",
          8893 => x"2b",
          8894 => x"41",
          8895 => x"41",
          8896 => x"41",
          8897 => x"41",
          8898 => x"41",
          8899 => x"47",
          8900 => x"48",
          8901 => x"49",
          8902 => x"4b",
          8903 => x"48",
          8904 => x"46",
          8905 => x"4a",
          8906 => x"4b",
          8907 => x"4a",
          8908 => x"4a",
          8909 => x"4a",
          8910 => x"49",
          8911 => x"46",
          8912 => x"49",
          8913 => x"49",
          8914 => x"4a",
          8915 => x"46",
          8916 => x"46",
          8917 => x"4a",
          8918 => x"4a",
          8919 => x"4b",
          8920 => x"4b",
          8921 => x"0e",
          8922 => x"17",
          8923 => x"17",
          8924 => x"0e",
          8925 => x"17",
          8926 => x"17",
          8927 => x"17",
          8928 => x"17",
          8929 => x"17",
          8930 => x"17",
          8931 => x"17",
          8932 => x"0e",
          8933 => x"17",
          8934 => x"0e",
          8935 => x"0e",
          8936 => x"17",
          8937 => x"17",
          8938 => x"17",
          8939 => x"17",
          8940 => x"17",
          8941 => x"17",
          8942 => x"17",
          8943 => x"17",
          8944 => x"17",
          8945 => x"17",
          8946 => x"17",
          8947 => x"17",
          8948 => x"17",
          8949 => x"17",
          8950 => x"17",
          8951 => x"17",
          8952 => x"17",
          8953 => x"17",
          8954 => x"17",
          8955 => x"17",
          8956 => x"17",
          8957 => x"17",
          8958 => x"17",
          8959 => x"17",
          8960 => x"17",
          8961 => x"17",
          8962 => x"17",
          8963 => x"17",
          8964 => x"17",
          8965 => x"17",
          8966 => x"17",
          8967 => x"17",
          8968 => x"17",
          8969 => x"17",
          8970 => x"17",
          8971 => x"17",
          8972 => x"0f",
          8973 => x"17",
          8974 => x"17",
          8975 => x"17",
          8976 => x"17",
          8977 => x"11",
          8978 => x"17",
          8979 => x"17",
          8980 => x"17",
          8981 => x"17",
          8982 => x"17",
          8983 => x"17",
          8984 => x"17",
          8985 => x"17",
          8986 => x"17",
          8987 => x"17",
          8988 => x"0e",
          8989 => x"10",
          8990 => x"0e",
          8991 => x"0e",
          8992 => x"0e",
          8993 => x"17",
          8994 => x"10",
          8995 => x"17",
          8996 => x"17",
          8997 => x"0e",
          8998 => x"17",
          8999 => x"17",
          9000 => x"10",
          9001 => x"10",
          9002 => x"17",
          9003 => x"17",
          9004 => x"0f",
          9005 => x"17",
          9006 => x"11",
          9007 => x"17",
          9008 => x"17",
          9009 => x"11",
          9010 => x"6e",
          9011 => x"00",
          9012 => x"6f",
          9013 => x"00",
          9014 => x"6e",
          9015 => x"00",
          9016 => x"6f",
          9017 => x"00",
          9018 => x"78",
          9019 => x"00",
          9020 => x"6c",
          9021 => x"00",
          9022 => x"6f",
          9023 => x"00",
          9024 => x"69",
          9025 => x"00",
          9026 => x"75",
          9027 => x"00",
          9028 => x"62",
          9029 => x"68",
          9030 => x"77",
          9031 => x"64",
          9032 => x"65",
          9033 => x"64",
          9034 => x"65",
          9035 => x"6c",
          9036 => x"00",
          9037 => x"70",
          9038 => x"73",
          9039 => x"74",
          9040 => x"73",
          9041 => x"00",
          9042 => x"66",
          9043 => x"00",
          9044 => x"73",
          9045 => x"00",
          9046 => x"61",
          9047 => x"00",
          9048 => x"61",
          9049 => x"00",
          9050 => x"6c",
          9051 => x"00",
          9052 => x"00",
          9053 => x"73",
          9054 => x"72",
          9055 => x"00",
          9056 => x"74",
          9057 => x"61",
          9058 => x"72",
          9059 => x"2e",
          9060 => x"73",
          9061 => x"6f",
          9062 => x"65",
          9063 => x"2e",
          9064 => x"20",
          9065 => x"65",
          9066 => x"75",
          9067 => x"00",
          9068 => x"20",
          9069 => x"68",
          9070 => x"75",
          9071 => x"00",
          9072 => x"76",
          9073 => x"64",
          9074 => x"6c",
          9075 => x"6d",
          9076 => x"00",
          9077 => x"63",
          9078 => x"20",
          9079 => x"69",
          9080 => x"00",
          9081 => x"6c",
          9082 => x"6c",
          9083 => x"64",
          9084 => x"78",
          9085 => x"73",
          9086 => x"00",
          9087 => x"6c",
          9088 => x"61",
          9089 => x"65",
          9090 => x"76",
          9091 => x"64",
          9092 => x"00",
          9093 => x"20",
          9094 => x"77",
          9095 => x"65",
          9096 => x"6f",
          9097 => x"74",
          9098 => x"00",
          9099 => x"69",
          9100 => x"6e",
          9101 => x"65",
          9102 => x"73",
          9103 => x"76",
          9104 => x"64",
          9105 => x"00",
          9106 => x"73",
          9107 => x"6f",
          9108 => x"6e",
          9109 => x"65",
          9110 => x"00",
          9111 => x"20",
          9112 => x"70",
          9113 => x"62",
          9114 => x"66",
          9115 => x"73",
          9116 => x"65",
          9117 => x"6f",
          9118 => x"20",
          9119 => x"64",
          9120 => x"2e",
          9121 => x"72",
          9122 => x"20",
          9123 => x"72",
          9124 => x"2e",
          9125 => x"6d",
          9126 => x"74",
          9127 => x"70",
          9128 => x"74",
          9129 => x"20",
          9130 => x"63",
          9131 => x"65",
          9132 => x"00",
          9133 => x"6c",
          9134 => x"73",
          9135 => x"63",
          9136 => x"2e",
          9137 => x"73",
          9138 => x"69",
          9139 => x"6e",
          9140 => x"65",
          9141 => x"79",
          9142 => x"00",
          9143 => x"6f",
          9144 => x"6e",
          9145 => x"70",
          9146 => x"66",
          9147 => x"73",
          9148 => x"00",
          9149 => x"72",
          9150 => x"74",
          9151 => x"20",
          9152 => x"6f",
          9153 => x"63",
          9154 => x"00",
          9155 => x"63",
          9156 => x"73",
          9157 => x"00",
          9158 => x"6b",
          9159 => x"6e",
          9160 => x"72",
          9161 => x"00",
          9162 => x"6c",
          9163 => x"79",
          9164 => x"20",
          9165 => x"61",
          9166 => x"6c",
          9167 => x"79",
          9168 => x"2f",
          9169 => x"2e",
          9170 => x"00",
          9171 => x"61",
          9172 => x"00",
          9173 => x"38",
          9174 => x"00",
          9175 => x"20",
          9176 => x"34",
          9177 => x"00",
          9178 => x"20",
          9179 => x"20",
          9180 => x"00",
          9181 => x"32",
          9182 => x"00",
          9183 => x"00",
          9184 => x"00",
          9185 => x"00",
          9186 => x"53",
          9187 => x"2a",
          9188 => x"20",
          9189 => x"00",
          9190 => x"2f",
          9191 => x"32",
          9192 => x"00",
          9193 => x"2e",
          9194 => x"00",
          9195 => x"50",
          9196 => x"72",
          9197 => x"25",
          9198 => x"29",
          9199 => x"20",
          9200 => x"2a",
          9201 => x"00",
          9202 => x"55",
          9203 => x"74",
          9204 => x"75",
          9205 => x"48",
          9206 => x"6c",
          9207 => x"00",
          9208 => x"6d",
          9209 => x"69",
          9210 => x"72",
          9211 => x"74",
          9212 => x"32",
          9213 => x"74",
          9214 => x"75",
          9215 => x"00",
          9216 => x"43",
          9217 => x"52",
          9218 => x"6e",
          9219 => x"72",
          9220 => x"00",
          9221 => x"43",
          9222 => x"57",
          9223 => x"6e",
          9224 => x"72",
          9225 => x"00",
          9226 => x"52",
          9227 => x"52",
          9228 => x"6e",
          9229 => x"72",
          9230 => x"00",
          9231 => x"52",
          9232 => x"54",
          9233 => x"6e",
          9234 => x"72",
          9235 => x"00",
          9236 => x"52",
          9237 => x"52",
          9238 => x"6e",
          9239 => x"72",
          9240 => x"00",
          9241 => x"52",
          9242 => x"54",
          9243 => x"6e",
          9244 => x"72",
          9245 => x"00",
          9246 => x"74",
          9247 => x"67",
          9248 => x"20",
          9249 => x"65",
          9250 => x"2e",
          9251 => x"61",
          9252 => x"6e",
          9253 => x"69",
          9254 => x"2e",
          9255 => x"00",
          9256 => x"74",
          9257 => x"65",
          9258 => x"61",
          9259 => x"00",
          9260 => x"53",
          9261 => x"74",
          9262 => x"00",
          9263 => x"69",
          9264 => x"20",
          9265 => x"69",
          9266 => x"69",
          9267 => x"73",
          9268 => x"64",
          9269 => x"72",
          9270 => x"2c",
          9271 => x"65",
          9272 => x"20",
          9273 => x"74",
          9274 => x"6e",
          9275 => x"6c",
          9276 => x"00",
          9277 => x"00",
          9278 => x"65",
          9279 => x"6e",
          9280 => x"2e",
          9281 => x"00",
          9282 => x"70",
          9283 => x"67",
          9284 => x"00",
          9285 => x"6d",
          9286 => x"69",
          9287 => x"2e",
          9288 => x"00",
          9289 => x"38",
          9290 => x"25",
          9291 => x"29",
          9292 => x"30",
          9293 => x"28",
          9294 => x"78",
          9295 => x"00",
          9296 => x"6d",
          9297 => x"65",
          9298 => x"79",
          9299 => x"6f",
          9300 => x"65",
          9301 => x"00",
          9302 => x"38",
          9303 => x"25",
          9304 => x"2d",
          9305 => x"3f",
          9306 => x"38",
          9307 => x"25",
          9308 => x"2d",
          9309 => x"38",
          9310 => x"25",
          9311 => x"58",
          9312 => x"00",
          9313 => x"65",
          9314 => x"69",
          9315 => x"63",
          9316 => x"20",
          9317 => x"30",
          9318 => x"20",
          9319 => x"0a",
          9320 => x"6c",
          9321 => x"67",
          9322 => x"64",
          9323 => x"20",
          9324 => x"6c",
          9325 => x"2e",
          9326 => x"00",
          9327 => x"6c",
          9328 => x"65",
          9329 => x"6e",
          9330 => x"63",
          9331 => x"20",
          9332 => x"29",
          9333 => x"00",
          9334 => x"73",
          9335 => x"74",
          9336 => x"20",
          9337 => x"6c",
          9338 => x"74",
          9339 => x"2e",
          9340 => x"00",
          9341 => x"6c",
          9342 => x"65",
          9343 => x"74",
          9344 => x"2e",
          9345 => x"00",
          9346 => x"55",
          9347 => x"6e",
          9348 => x"3a",
          9349 => x"5c",
          9350 => x"25",
          9351 => x"00",
          9352 => x"3a",
          9353 => x"5c",
          9354 => x"00",
          9355 => x"3a",
          9356 => x"00",
          9357 => x"64",
          9358 => x"6d",
          9359 => x"64",
          9360 => x"00",
          9361 => x"6e",
          9362 => x"67",
          9363 => x"00",
          9364 => x"61",
          9365 => x"6e",
          9366 => x"6e",
          9367 => x"72",
          9368 => x"73",
          9369 => x"00",
          9370 => x"2f",
          9371 => x"25",
          9372 => x"64",
          9373 => x"3a",
          9374 => x"25",
          9375 => x"0a",
          9376 => x"43",
          9377 => x"6e",
          9378 => x"75",
          9379 => x"69",
          9380 => x"00",
          9381 => x"66",
          9382 => x"20",
          9383 => x"20",
          9384 => x"66",
          9385 => x"00",
          9386 => x"44",
          9387 => x"63",
          9388 => x"69",
          9389 => x"65",
          9390 => x"74",
          9391 => x"0a",
          9392 => x"20",
          9393 => x"20",
          9394 => x"41",
          9395 => x"28",
          9396 => x"58",
          9397 => x"38",
          9398 => x"0a",
          9399 => x"20",
          9400 => x"52",
          9401 => x"20",
          9402 => x"28",
          9403 => x"58",
          9404 => x"38",
          9405 => x"0a",
          9406 => x"20",
          9407 => x"53",
          9408 => x"52",
          9409 => x"28",
          9410 => x"58",
          9411 => x"38",
          9412 => x"0a",
          9413 => x"20",
          9414 => x"41",
          9415 => x"20",
          9416 => x"28",
          9417 => x"58",
          9418 => x"38",
          9419 => x"0a",
          9420 => x"20",
          9421 => x"4d",
          9422 => x"20",
          9423 => x"28",
          9424 => x"58",
          9425 => x"38",
          9426 => x"0a",
          9427 => x"20",
          9428 => x"20",
          9429 => x"44",
          9430 => x"28",
          9431 => x"69",
          9432 => x"20",
          9433 => x"32",
          9434 => x"0a",
          9435 => x"20",
          9436 => x"4d",
          9437 => x"20",
          9438 => x"28",
          9439 => x"65",
          9440 => x"20",
          9441 => x"32",
          9442 => x"0a",
          9443 => x"20",
          9444 => x"54",
          9445 => x"54",
          9446 => x"28",
          9447 => x"6e",
          9448 => x"73",
          9449 => x"32",
          9450 => x"0a",
          9451 => x"20",
          9452 => x"53",
          9453 => x"4e",
          9454 => x"55",
          9455 => x"00",
          9456 => x"20",
          9457 => x"20",
          9458 => x"0a",
          9459 => x"20",
          9460 => x"43",
          9461 => x"00",
          9462 => x"20",
          9463 => x"32",
          9464 => x"00",
          9465 => x"20",
          9466 => x"49",
          9467 => x"00",
          9468 => x"64",
          9469 => x"73",
          9470 => x"0a",
          9471 => x"20",
          9472 => x"55",
          9473 => x"73",
          9474 => x"56",
          9475 => x"6f",
          9476 => x"64",
          9477 => x"73",
          9478 => x"20",
          9479 => x"58",
          9480 => x"00",
          9481 => x"20",
          9482 => x"55",
          9483 => x"6d",
          9484 => x"20",
          9485 => x"72",
          9486 => x"64",
          9487 => x"73",
          9488 => x"20",
          9489 => x"58",
          9490 => x"00",
          9491 => x"20",
          9492 => x"61",
          9493 => x"53",
          9494 => x"74",
          9495 => x"64",
          9496 => x"73",
          9497 => x"20",
          9498 => x"20",
          9499 => x"58",
          9500 => x"00",
          9501 => x"73",
          9502 => x"00",
          9503 => x"20",
          9504 => x"55",
          9505 => x"20",
          9506 => x"20",
          9507 => x"20",
          9508 => x"20",
          9509 => x"20",
          9510 => x"20",
          9511 => x"58",
          9512 => x"00",
          9513 => x"20",
          9514 => x"73",
          9515 => x"20",
          9516 => x"63",
          9517 => x"72",
          9518 => x"20",
          9519 => x"20",
          9520 => x"20",
          9521 => x"25",
          9522 => x"4d",
          9523 => x"00",
          9524 => x"20",
          9525 => x"52",
          9526 => x"43",
          9527 => x"6b",
          9528 => x"65",
          9529 => x"20",
          9530 => x"20",
          9531 => x"20",
          9532 => x"25",
          9533 => x"4d",
          9534 => x"00",
          9535 => x"20",
          9536 => x"73",
          9537 => x"6e",
          9538 => x"44",
          9539 => x"20",
          9540 => x"63",
          9541 => x"72",
          9542 => x"20",
          9543 => x"25",
          9544 => x"4d",
          9545 => x"00",
          9546 => x"61",
          9547 => x"00",
          9548 => x"64",
          9549 => x"00",
          9550 => x"65",
          9551 => x"00",
          9552 => x"4f",
          9553 => x"4f",
          9554 => x"00",
          9555 => x"6b",
          9556 => x"6e",
          9557 => x"96",
          9558 => x"00",
          9559 => x"00",
          9560 => x"96",
          9561 => x"00",
          9562 => x"00",
          9563 => x"96",
          9564 => x"00",
          9565 => x"00",
          9566 => x"96",
          9567 => x"00",
          9568 => x"00",
          9569 => x"96",
          9570 => x"00",
          9571 => x"00",
          9572 => x"96",
          9573 => x"00",
          9574 => x"00",
          9575 => x"96",
          9576 => x"00",
          9577 => x"00",
          9578 => x"96",
          9579 => x"00",
          9580 => x"00",
          9581 => x"96",
          9582 => x"00",
          9583 => x"00",
          9584 => x"96",
          9585 => x"00",
          9586 => x"00",
          9587 => x"96",
          9588 => x"00",
          9589 => x"00",
          9590 => x"96",
          9591 => x"00",
          9592 => x"00",
          9593 => x"96",
          9594 => x"00",
          9595 => x"00",
          9596 => x"96",
          9597 => x"00",
          9598 => x"00",
          9599 => x"96",
          9600 => x"00",
          9601 => x"00",
          9602 => x"96",
          9603 => x"00",
          9604 => x"00",
          9605 => x"96",
          9606 => x"00",
          9607 => x"00",
          9608 => x"96",
          9609 => x"00",
          9610 => x"00",
          9611 => x"96",
          9612 => x"00",
          9613 => x"00",
          9614 => x"96",
          9615 => x"00",
          9616 => x"00",
          9617 => x"96",
          9618 => x"00",
          9619 => x"00",
          9620 => x"96",
          9621 => x"00",
          9622 => x"00",
          9623 => x"44",
          9624 => x"43",
          9625 => x"42",
          9626 => x"41",
          9627 => x"36",
          9628 => x"35",
          9629 => x"34",
          9630 => x"46",
          9631 => x"33",
          9632 => x"32",
          9633 => x"31",
          9634 => x"00",
          9635 => x"00",
          9636 => x"00",
          9637 => x"00",
          9638 => x"00",
          9639 => x"00",
          9640 => x"00",
          9641 => x"00",
          9642 => x"00",
          9643 => x"00",
          9644 => x"00",
          9645 => x"73",
          9646 => x"79",
          9647 => x"73",
          9648 => x"00",
          9649 => x"00",
          9650 => x"34",
          9651 => x"20",
          9652 => x"00",
          9653 => x"69",
          9654 => x"20",
          9655 => x"72",
          9656 => x"74",
          9657 => x"65",
          9658 => x"73",
          9659 => x"79",
          9660 => x"6c",
          9661 => x"6f",
          9662 => x"46",
          9663 => x"00",
          9664 => x"6e",
          9665 => x"20",
          9666 => x"6e",
          9667 => x"65",
          9668 => x"20",
          9669 => x"74",
          9670 => x"20",
          9671 => x"65",
          9672 => x"69",
          9673 => x"6c",
          9674 => x"2e",
          9675 => x"00",
          9676 => x"2b",
          9677 => x"3c",
          9678 => x"5b",
          9679 => x"00",
          9680 => x"54",
          9681 => x"54",
          9682 => x"00",
          9683 => x"90",
          9684 => x"4f",
          9685 => x"30",
          9686 => x"20",
          9687 => x"45",
          9688 => x"20",
          9689 => x"33",
          9690 => x"20",
          9691 => x"20",
          9692 => x"45",
          9693 => x"20",
          9694 => x"20",
          9695 => x"20",
          9696 => x"97",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"45",
          9701 => x"8f",
          9702 => x"45",
          9703 => x"8e",
          9704 => x"92",
          9705 => x"55",
          9706 => x"9a",
          9707 => x"9e",
          9708 => x"4f",
          9709 => x"a6",
          9710 => x"aa",
          9711 => x"ae",
          9712 => x"b2",
          9713 => x"b6",
          9714 => x"ba",
          9715 => x"be",
          9716 => x"c2",
          9717 => x"c6",
          9718 => x"ca",
          9719 => x"ce",
          9720 => x"d2",
          9721 => x"d6",
          9722 => x"da",
          9723 => x"de",
          9724 => x"e2",
          9725 => x"e6",
          9726 => x"ea",
          9727 => x"ee",
          9728 => x"f2",
          9729 => x"f6",
          9730 => x"fa",
          9731 => x"fe",
          9732 => x"2c",
          9733 => x"5d",
          9734 => x"2a",
          9735 => x"3f",
          9736 => x"00",
          9737 => x"00",
          9738 => x"00",
          9739 => x"02",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"8c",
          9747 => x"01",
          9748 => x"00",
          9749 => x"00",
          9750 => x"8c",
          9751 => x"01",
          9752 => x"00",
          9753 => x"00",
          9754 => x"8c",
          9755 => x"03",
          9756 => x"00",
          9757 => x"00",
          9758 => x"8c",
          9759 => x"03",
          9760 => x"00",
          9761 => x"00",
          9762 => x"8c",
          9763 => x"03",
          9764 => x"00",
          9765 => x"00",
          9766 => x"8c",
          9767 => x"04",
          9768 => x"00",
          9769 => x"00",
          9770 => x"8c",
          9771 => x"04",
          9772 => x"00",
          9773 => x"00",
          9774 => x"8d",
          9775 => x"04",
          9776 => x"00",
          9777 => x"00",
          9778 => x"8d",
          9779 => x"04",
          9780 => x"00",
          9781 => x"00",
          9782 => x"8d",
          9783 => x"04",
          9784 => x"00",
          9785 => x"00",
          9786 => x"8d",
          9787 => x"04",
          9788 => x"00",
          9789 => x"00",
          9790 => x"8d",
          9791 => x"04",
          9792 => x"00",
          9793 => x"00",
          9794 => x"8d",
          9795 => x"05",
          9796 => x"00",
          9797 => x"00",
          9798 => x"8d",
          9799 => x"05",
          9800 => x"00",
          9801 => x"00",
          9802 => x"8d",
          9803 => x"05",
          9804 => x"00",
          9805 => x"00",
          9806 => x"8d",
          9807 => x"05",
          9808 => x"00",
          9809 => x"00",
          9810 => x"8d",
          9811 => x"07",
          9812 => x"00",
          9813 => x"00",
          9814 => x"8d",
          9815 => x"07",
          9816 => x"00",
          9817 => x"00",
          9818 => x"8d",
          9819 => x"08",
          9820 => x"00",
          9821 => x"00",
          9822 => x"8d",
          9823 => x"08",
          9824 => x"00",
          9825 => x"00",
          9826 => x"8d",
          9827 => x"08",
          9828 => x"00",
          9829 => x"00",
          9830 => x"8d",
          9831 => x"08",
          9832 => x"00",
          9833 => x"00",
          9834 => x"8d",
          9835 => x"09",
          9836 => x"00",
          9837 => x"00",
          9838 => x"8d",
          9839 => x"09",
          9840 => x"00",
          9841 => x"00",
          9842 => x"8d",
          9843 => x"09",
          9844 => x"00",
          9845 => x"00",
          9846 => x"8d",
          9847 => x"09",
          9848 => x"00",
          9849 => x"00",
          9850 => x"00",
          9851 => x"00",
          9852 => x"7f",
          9853 => x"00",
          9854 => x"7f",
          9855 => x"00",
          9856 => x"7f",
          9857 => x"00",
          9858 => x"00",
          9859 => x"00",
          9860 => x"ff",
          9861 => x"00",
          9862 => x"00",
          9863 => x"78",
          9864 => x"00",
          9865 => x"e1",
          9866 => x"e1",
          9867 => x"e1",
          9868 => x"00",
          9869 => x"01",
          9870 => x"01",
          9871 => x"10",
          9872 => x"00",
          9873 => x"00",
          9874 => x"00",
          9875 => x"00",
          9876 => x"00",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"00",
          9881 => x"00",
          9882 => x"00",
          9883 => x"00",
          9884 => x"00",
          9885 => x"00",
          9886 => x"00",
          9887 => x"00",
          9888 => x"00",
          9889 => x"00",
          9890 => x"00",
          9891 => x"00",
          9892 => x"00",
          9893 => x"00",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"96",
          9898 => x"00",
          9899 => x"96",
          9900 => x"00",
          9901 => x"96",
          9902 => x"00",
          9903 => x"00",
          9904 => x"00",
          9905 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"85",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"80",
           387 => x"82",
           388 => x"82",
           389 => x"82",
           390 => x"b3",
           391 => x"b5",
           392 => x"d0",
           393 => x"b5",
           394 => x"e3",
           395 => x"d4",
           396 => x"90",
           397 => x"d4",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"82",
           403 => x"82",
           404 => x"82",
           405 => x"b1",
           406 => x"b5",
           407 => x"d0",
           408 => x"b5",
           409 => x"cf",
           410 => x"b5",
           411 => x"d0",
           412 => x"b5",
           413 => x"c9",
           414 => x"b5",
           415 => x"d0",
           416 => x"b5",
           417 => x"d8",
           418 => x"d4",
           419 => x"90",
           420 => x"d4",
           421 => x"2d",
           422 => x"08",
           423 => x"04",
           424 => x"0c",
           425 => x"82",
           426 => x"82",
           427 => x"82",
           428 => x"80",
           429 => x"82",
           430 => x"82",
           431 => x"82",
           432 => x"80",
           433 => x"82",
           434 => x"82",
           435 => x"82",
           436 => x"80",
           437 => x"82",
           438 => x"82",
           439 => x"82",
           440 => x"80",
           441 => x"82",
           442 => x"82",
           443 => x"82",
           444 => x"80",
           445 => x"82",
           446 => x"82",
           447 => x"82",
           448 => x"81",
           449 => x"82",
           450 => x"82",
           451 => x"82",
           452 => x"81",
           453 => x"82",
           454 => x"82",
           455 => x"82",
           456 => x"81",
           457 => x"82",
           458 => x"82",
           459 => x"82",
           460 => x"81",
           461 => x"82",
           462 => x"82",
           463 => x"82",
           464 => x"81",
           465 => x"82",
           466 => x"82",
           467 => x"82",
           468 => x"81",
           469 => x"82",
           470 => x"82",
           471 => x"82",
           472 => x"81",
           473 => x"82",
           474 => x"82",
           475 => x"82",
           476 => x"81",
           477 => x"82",
           478 => x"82",
           479 => x"82",
           480 => x"81",
           481 => x"82",
           482 => x"82",
           483 => x"82",
           484 => x"81",
           485 => x"82",
           486 => x"82",
           487 => x"82",
           488 => x"81",
           489 => x"82",
           490 => x"82",
           491 => x"82",
           492 => x"81",
           493 => x"82",
           494 => x"82",
           495 => x"82",
           496 => x"81",
           497 => x"82",
           498 => x"82",
           499 => x"82",
           500 => x"81",
           501 => x"82",
           502 => x"82",
           503 => x"82",
           504 => x"81",
           505 => x"82",
           506 => x"82",
           507 => x"82",
           508 => x"81",
           509 => x"82",
           510 => x"82",
           511 => x"82",
           512 => x"81",
           513 => x"82",
           514 => x"82",
           515 => x"82",
           516 => x"81",
           517 => x"82",
           518 => x"82",
           519 => x"82",
           520 => x"81",
           521 => x"82",
           522 => x"82",
           523 => x"82",
           524 => x"81",
           525 => x"82",
           526 => x"82",
           527 => x"82",
           528 => x"81",
           529 => x"82",
           530 => x"82",
           531 => x"82",
           532 => x"82",
           533 => x"82",
           534 => x"82",
           535 => x"82",
           536 => x"82",
           537 => x"82",
           538 => x"82",
           539 => x"82",
           540 => x"81",
           541 => x"82",
           542 => x"82",
           543 => x"82",
           544 => x"82",
           545 => x"82",
           546 => x"82",
           547 => x"82",
           548 => x"82",
           549 => x"82",
           550 => x"82",
           551 => x"82",
           552 => x"82",
           553 => x"82",
           554 => x"82",
           555 => x"82",
           556 => x"81",
           557 => x"82",
           558 => x"82",
           559 => x"82",
           560 => x"81",
           561 => x"82",
           562 => x"82",
           563 => x"82",
           564 => x"81",
           565 => x"82",
           566 => x"82",
           567 => x"82",
           568 => x"80",
           569 => x"82",
           570 => x"82",
           571 => x"82",
           572 => x"80",
           573 => x"82",
           574 => x"82",
           575 => x"82",
           576 => x"80",
           577 => x"82",
           578 => x"82",
           579 => x"82",
           580 => x"80",
           581 => x"82",
           582 => x"82",
           583 => x"82",
           584 => x"81",
           585 => x"82",
           586 => x"82",
           587 => x"82",
           588 => x"81",
           589 => x"82",
           590 => x"82",
           591 => x"82",
           592 => x"81",
           593 => x"82",
           594 => x"82",
           595 => x"82",
           596 => x"81",
           597 => x"82",
           598 => x"82",
           599 => x"3c",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"51",
           609 => x"73",
           610 => x"73",
           611 => x"81",
           612 => x"10",
           613 => x"07",
           614 => x"0c",
           615 => x"72",
           616 => x"81",
           617 => x"09",
           618 => x"71",
           619 => x"0a",
           620 => x"72",
           621 => x"51",
           622 => x"82",
           623 => x"82",
           624 => x"8e",
           625 => x"70",
           626 => x"0c",
           627 => x"93",
           628 => x"81",
           629 => x"e2",
           630 => x"b5",
           631 => x"82",
           632 => x"fb",
           633 => x"b5",
           634 => x"05",
           635 => x"d4",
           636 => x"0c",
           637 => x"08",
           638 => x"54",
           639 => x"08",
           640 => x"53",
           641 => x"08",
           642 => x"9a",
           643 => x"c8",
           644 => x"b5",
           645 => x"05",
           646 => x"d4",
           647 => x"08",
           648 => x"c8",
           649 => x"87",
           650 => x"b5",
           651 => x"82",
           652 => x"02",
           653 => x"0c",
           654 => x"82",
           655 => x"90",
           656 => x"11",
           657 => x"32",
           658 => x"51",
           659 => x"71",
           660 => x"0b",
           661 => x"08",
           662 => x"25",
           663 => x"39",
           664 => x"b5",
           665 => x"05",
           666 => x"39",
           667 => x"08",
           668 => x"ff",
           669 => x"d4",
           670 => x"0c",
           671 => x"b5",
           672 => x"05",
           673 => x"d4",
           674 => x"08",
           675 => x"08",
           676 => x"82",
           677 => x"f8",
           678 => x"2e",
           679 => x"80",
           680 => x"d4",
           681 => x"08",
           682 => x"38",
           683 => x"08",
           684 => x"51",
           685 => x"82",
           686 => x"70",
           687 => x"08",
           688 => x"52",
           689 => x"08",
           690 => x"ff",
           691 => x"06",
           692 => x"0b",
           693 => x"08",
           694 => x"80",
           695 => x"b5",
           696 => x"05",
           697 => x"d4",
           698 => x"08",
           699 => x"73",
           700 => x"d4",
           701 => x"08",
           702 => x"b5",
           703 => x"05",
           704 => x"d4",
           705 => x"08",
           706 => x"b5",
           707 => x"05",
           708 => x"39",
           709 => x"08",
           710 => x"52",
           711 => x"82",
           712 => x"88",
           713 => x"82",
           714 => x"f4",
           715 => x"82",
           716 => x"f4",
           717 => x"b5",
           718 => x"3d",
           719 => x"d4",
           720 => x"b5",
           721 => x"82",
           722 => x"f4",
           723 => x"0b",
           724 => x"08",
           725 => x"82",
           726 => x"88",
           727 => x"b5",
           728 => x"05",
           729 => x"0b",
           730 => x"08",
           731 => x"82",
           732 => x"90",
           733 => x"b5",
           734 => x"05",
           735 => x"d4",
           736 => x"08",
           737 => x"d4",
           738 => x"08",
           739 => x"d4",
           740 => x"70",
           741 => x"81",
           742 => x"b5",
           743 => x"82",
           744 => x"dc",
           745 => x"b5",
           746 => x"05",
           747 => x"d4",
           748 => x"08",
           749 => x"80",
           750 => x"b5",
           751 => x"05",
           752 => x"b5",
           753 => x"8e",
           754 => x"b5",
           755 => x"82",
           756 => x"02",
           757 => x"0c",
           758 => x"82",
           759 => x"90",
           760 => x"b5",
           761 => x"05",
           762 => x"d4",
           763 => x"08",
           764 => x"d4",
           765 => x"08",
           766 => x"d4",
           767 => x"08",
           768 => x"3f",
           769 => x"08",
           770 => x"d4",
           771 => x"0c",
           772 => x"08",
           773 => x"70",
           774 => x"0c",
           775 => x"3d",
           776 => x"d4",
           777 => x"b5",
           778 => x"82",
           779 => x"ed",
           780 => x"0b",
           781 => x"08",
           782 => x"82",
           783 => x"88",
           784 => x"80",
           785 => x"0c",
           786 => x"08",
           787 => x"85",
           788 => x"81",
           789 => x"32",
           790 => x"51",
           791 => x"53",
           792 => x"8d",
           793 => x"82",
           794 => x"e0",
           795 => x"ac",
           796 => x"d4",
           797 => x"08",
           798 => x"53",
           799 => x"d4",
           800 => x"34",
           801 => x"06",
           802 => x"2e",
           803 => x"82",
           804 => x"8c",
           805 => x"05",
           806 => x"08",
           807 => x"82",
           808 => x"e4",
           809 => x"81",
           810 => x"72",
           811 => x"8b",
           812 => x"d4",
           813 => x"33",
           814 => x"27",
           815 => x"82",
           816 => x"f8",
           817 => x"72",
           818 => x"ee",
           819 => x"d4",
           820 => x"33",
           821 => x"2e",
           822 => x"80",
           823 => x"b5",
           824 => x"05",
           825 => x"2b",
           826 => x"51",
           827 => x"b2",
           828 => x"d4",
           829 => x"22",
           830 => x"70",
           831 => x"81",
           832 => x"51",
           833 => x"2e",
           834 => x"b5",
           835 => x"05",
           836 => x"80",
           837 => x"72",
           838 => x"08",
           839 => x"fe",
           840 => x"b5",
           841 => x"05",
           842 => x"2b",
           843 => x"70",
           844 => x"72",
           845 => x"51",
           846 => x"51",
           847 => x"82",
           848 => x"e8",
           849 => x"b5",
           850 => x"05",
           851 => x"b5",
           852 => x"05",
           853 => x"d0",
           854 => x"53",
           855 => x"d4",
           856 => x"34",
           857 => x"08",
           858 => x"70",
           859 => x"98",
           860 => x"53",
           861 => x"8b",
           862 => x"0b",
           863 => x"08",
           864 => x"82",
           865 => x"e4",
           866 => x"83",
           867 => x"06",
           868 => x"72",
           869 => x"82",
           870 => x"e8",
           871 => x"88",
           872 => x"2b",
           873 => x"70",
           874 => x"51",
           875 => x"72",
           876 => x"08",
           877 => x"fd",
           878 => x"b5",
           879 => x"05",
           880 => x"2a",
           881 => x"51",
           882 => x"80",
           883 => x"82",
           884 => x"e8",
           885 => x"98",
           886 => x"2c",
           887 => x"72",
           888 => x"0b",
           889 => x"08",
           890 => x"82",
           891 => x"f8",
           892 => x"11",
           893 => x"08",
           894 => x"53",
           895 => x"08",
           896 => x"80",
           897 => x"94",
           898 => x"d4",
           899 => x"08",
           900 => x"82",
           901 => x"70",
           902 => x"51",
           903 => x"82",
           904 => x"e4",
           905 => x"90",
           906 => x"72",
           907 => x"08",
           908 => x"82",
           909 => x"e4",
           910 => x"a0",
           911 => x"72",
           912 => x"08",
           913 => x"fc",
           914 => x"b5",
           915 => x"05",
           916 => x"80",
           917 => x"72",
           918 => x"08",
           919 => x"fc",
           920 => x"b5",
           921 => x"05",
           922 => x"c0",
           923 => x"72",
           924 => x"08",
           925 => x"fb",
           926 => x"b5",
           927 => x"05",
           928 => x"07",
           929 => x"82",
           930 => x"e4",
           931 => x"0b",
           932 => x"08",
           933 => x"fb",
           934 => x"b5",
           935 => x"05",
           936 => x"07",
           937 => x"82",
           938 => x"e4",
           939 => x"c1",
           940 => x"82",
           941 => x"fc",
           942 => x"b5",
           943 => x"05",
           944 => x"51",
           945 => x"b5",
           946 => x"05",
           947 => x"0b",
           948 => x"08",
           949 => x"8d",
           950 => x"b5",
           951 => x"05",
           952 => x"d4",
           953 => x"08",
           954 => x"b5",
           955 => x"05",
           956 => x"51",
           957 => x"b5",
           958 => x"05",
           959 => x"d4",
           960 => x"22",
           961 => x"53",
           962 => x"d4",
           963 => x"23",
           964 => x"82",
           965 => x"90",
           966 => x"b5",
           967 => x"05",
           968 => x"82",
           969 => x"90",
           970 => x"08",
           971 => x"08",
           972 => x"82",
           973 => x"e4",
           974 => x"83",
           975 => x"06",
           976 => x"53",
           977 => x"ab",
           978 => x"d4",
           979 => x"33",
           980 => x"53",
           981 => x"53",
           982 => x"08",
           983 => x"52",
           984 => x"3f",
           985 => x"08",
           986 => x"b5",
           987 => x"05",
           988 => x"82",
           989 => x"fc",
           990 => x"9d",
           991 => x"b5",
           992 => x"72",
           993 => x"08",
           994 => x"82",
           995 => x"ec",
           996 => x"82",
           997 => x"f4",
           998 => x"71",
           999 => x"72",
          1000 => x"08",
          1001 => x"8b",
          1002 => x"b5",
          1003 => x"05",
          1004 => x"d4",
          1005 => x"08",
          1006 => x"b5",
          1007 => x"05",
          1008 => x"82",
          1009 => x"fc",
          1010 => x"b5",
          1011 => x"05",
          1012 => x"2a",
          1013 => x"51",
          1014 => x"72",
          1015 => x"38",
          1016 => x"08",
          1017 => x"70",
          1018 => x"72",
          1019 => x"82",
          1020 => x"fc",
          1021 => x"53",
          1022 => x"82",
          1023 => x"53",
          1024 => x"d4",
          1025 => x"23",
          1026 => x"b5",
          1027 => x"05",
          1028 => x"f3",
          1029 => x"c8",
          1030 => x"82",
          1031 => x"f4",
          1032 => x"b5",
          1033 => x"05",
          1034 => x"b5",
          1035 => x"05",
          1036 => x"31",
          1037 => x"82",
          1038 => x"ec",
          1039 => x"c1",
          1040 => x"d4",
          1041 => x"22",
          1042 => x"70",
          1043 => x"51",
          1044 => x"2e",
          1045 => x"b5",
          1046 => x"05",
          1047 => x"d4",
          1048 => x"08",
          1049 => x"b5",
          1050 => x"05",
          1051 => x"82",
          1052 => x"dc",
          1053 => x"a2",
          1054 => x"d4",
          1055 => x"08",
          1056 => x"08",
          1057 => x"84",
          1058 => x"d4",
          1059 => x"0c",
          1060 => x"b5",
          1061 => x"05",
          1062 => x"b5",
          1063 => x"05",
          1064 => x"d4",
          1065 => x"0c",
          1066 => x"08",
          1067 => x"80",
          1068 => x"82",
          1069 => x"e4",
          1070 => x"82",
          1071 => x"72",
          1072 => x"08",
          1073 => x"82",
          1074 => x"fc",
          1075 => x"82",
          1076 => x"fc",
          1077 => x"b5",
          1078 => x"05",
          1079 => x"bf",
          1080 => x"72",
          1081 => x"08",
          1082 => x"81",
          1083 => x"0b",
          1084 => x"08",
          1085 => x"a9",
          1086 => x"d4",
          1087 => x"22",
          1088 => x"07",
          1089 => x"82",
          1090 => x"e4",
          1091 => x"f8",
          1092 => x"d4",
          1093 => x"34",
          1094 => x"b5",
          1095 => x"05",
          1096 => x"d4",
          1097 => x"22",
          1098 => x"70",
          1099 => x"51",
          1100 => x"2e",
          1101 => x"b5",
          1102 => x"05",
          1103 => x"d4",
          1104 => x"08",
          1105 => x"b5",
          1106 => x"05",
          1107 => x"82",
          1108 => x"d8",
          1109 => x"a2",
          1110 => x"d4",
          1111 => x"08",
          1112 => x"08",
          1113 => x"84",
          1114 => x"d4",
          1115 => x"0c",
          1116 => x"b5",
          1117 => x"05",
          1118 => x"b5",
          1119 => x"05",
          1120 => x"d4",
          1121 => x"0c",
          1122 => x"08",
          1123 => x"70",
          1124 => x"53",
          1125 => x"d4",
          1126 => x"23",
          1127 => x"0b",
          1128 => x"08",
          1129 => x"82",
          1130 => x"f0",
          1131 => x"b5",
          1132 => x"05",
          1133 => x"d4",
          1134 => x"08",
          1135 => x"54",
          1136 => x"a3",
          1137 => x"b5",
          1138 => x"72",
          1139 => x"b5",
          1140 => x"05",
          1141 => x"d4",
          1142 => x"0c",
          1143 => x"08",
          1144 => x"70",
          1145 => x"89",
          1146 => x"38",
          1147 => x"08",
          1148 => x"53",
          1149 => x"82",
          1150 => x"f8",
          1151 => x"15",
          1152 => x"51",
          1153 => x"b5",
          1154 => x"05",
          1155 => x"82",
          1156 => x"f0",
          1157 => x"72",
          1158 => x"51",
          1159 => x"b5",
          1160 => x"05",
          1161 => x"d4",
          1162 => x"08",
          1163 => x"d4",
          1164 => x"33",
          1165 => x"b5",
          1166 => x"05",
          1167 => x"82",
          1168 => x"f0",
          1169 => x"b5",
          1170 => x"05",
          1171 => x"82",
          1172 => x"fc",
          1173 => x"53",
          1174 => x"82",
          1175 => x"70",
          1176 => x"08",
          1177 => x"53",
          1178 => x"08",
          1179 => x"80",
          1180 => x"fe",
          1181 => x"b5",
          1182 => x"05",
          1183 => x"d8",
          1184 => x"54",
          1185 => x"31",
          1186 => x"82",
          1187 => x"fc",
          1188 => x"b5",
          1189 => x"05",
          1190 => x"06",
          1191 => x"80",
          1192 => x"82",
          1193 => x"ec",
          1194 => x"11",
          1195 => x"82",
          1196 => x"ec",
          1197 => x"b5",
          1198 => x"05",
          1199 => x"2a",
          1200 => x"51",
          1201 => x"80",
          1202 => x"38",
          1203 => x"08",
          1204 => x"70",
          1205 => x"b5",
          1206 => x"05",
          1207 => x"d4",
          1208 => x"08",
          1209 => x"b5",
          1210 => x"05",
          1211 => x"d4",
          1212 => x"22",
          1213 => x"90",
          1214 => x"06",
          1215 => x"b5",
          1216 => x"05",
          1217 => x"53",
          1218 => x"d4",
          1219 => x"23",
          1220 => x"b5",
          1221 => x"05",
          1222 => x"53",
          1223 => x"d4",
          1224 => x"23",
          1225 => x"08",
          1226 => x"82",
          1227 => x"ec",
          1228 => x"b5",
          1229 => x"05",
          1230 => x"2a",
          1231 => x"51",
          1232 => x"80",
          1233 => x"38",
          1234 => x"08",
          1235 => x"70",
          1236 => x"98",
          1237 => x"d4",
          1238 => x"33",
          1239 => x"53",
          1240 => x"97",
          1241 => x"d4",
          1242 => x"22",
          1243 => x"51",
          1244 => x"b5",
          1245 => x"05",
          1246 => x"82",
          1247 => x"e8",
          1248 => x"82",
          1249 => x"fc",
          1250 => x"71",
          1251 => x"72",
          1252 => x"08",
          1253 => x"82",
          1254 => x"e4",
          1255 => x"83",
          1256 => x"06",
          1257 => x"72",
          1258 => x"38",
          1259 => x"08",
          1260 => x"70",
          1261 => x"90",
          1262 => x"2c",
          1263 => x"51",
          1264 => x"53",
          1265 => x"b5",
          1266 => x"05",
          1267 => x"31",
          1268 => x"82",
          1269 => x"ec",
          1270 => x"39",
          1271 => x"08",
          1272 => x"70",
          1273 => x"90",
          1274 => x"2c",
          1275 => x"51",
          1276 => x"53",
          1277 => x"b5",
          1278 => x"05",
          1279 => x"31",
          1280 => x"82",
          1281 => x"ec",
          1282 => x"b5",
          1283 => x"05",
          1284 => x"80",
          1285 => x"72",
          1286 => x"b5",
          1287 => x"05",
          1288 => x"54",
          1289 => x"b5",
          1290 => x"05",
          1291 => x"2b",
          1292 => x"51",
          1293 => x"25",
          1294 => x"b5",
          1295 => x"05",
          1296 => x"51",
          1297 => x"d2",
          1298 => x"d4",
          1299 => x"22",
          1300 => x"70",
          1301 => x"51",
          1302 => x"2e",
          1303 => x"b5",
          1304 => x"05",
          1305 => x"51",
          1306 => x"80",
          1307 => x"b5",
          1308 => x"05",
          1309 => x"2a",
          1310 => x"51",
          1311 => x"80",
          1312 => x"82",
          1313 => x"88",
          1314 => x"ab",
          1315 => x"3f",
          1316 => x"b5",
          1317 => x"05",
          1318 => x"2a",
          1319 => x"51",
          1320 => x"80",
          1321 => x"82",
          1322 => x"88",
          1323 => x"a0",
          1324 => x"3f",
          1325 => x"08",
          1326 => x"70",
          1327 => x"81",
          1328 => x"53",
          1329 => x"b1",
          1330 => x"d4",
          1331 => x"08",
          1332 => x"89",
          1333 => x"b5",
          1334 => x"05",
          1335 => x"90",
          1336 => x"06",
          1337 => x"b5",
          1338 => x"05",
          1339 => x"b5",
          1340 => x"05",
          1341 => x"bc",
          1342 => x"d4",
          1343 => x"22",
          1344 => x"70",
          1345 => x"51",
          1346 => x"2e",
          1347 => x"b5",
          1348 => x"05",
          1349 => x"54",
          1350 => x"b5",
          1351 => x"05",
          1352 => x"2b",
          1353 => x"51",
          1354 => x"25",
          1355 => x"b5",
          1356 => x"05",
          1357 => x"51",
          1358 => x"d2",
          1359 => x"d4",
          1360 => x"22",
          1361 => x"70",
          1362 => x"51",
          1363 => x"2e",
          1364 => x"b5",
          1365 => x"05",
          1366 => x"54",
          1367 => x"b5",
          1368 => x"05",
          1369 => x"2b",
          1370 => x"51",
          1371 => x"25",
          1372 => x"b5",
          1373 => x"05",
          1374 => x"51",
          1375 => x"d2",
          1376 => x"d4",
          1377 => x"22",
          1378 => x"70",
          1379 => x"51",
          1380 => x"38",
          1381 => x"08",
          1382 => x"ff",
          1383 => x"72",
          1384 => x"08",
          1385 => x"73",
          1386 => x"90",
          1387 => x"80",
          1388 => x"38",
          1389 => x"08",
          1390 => x"52",
          1391 => x"f4",
          1392 => x"82",
          1393 => x"f8",
          1394 => x"72",
          1395 => x"09",
          1396 => x"38",
          1397 => x"08",
          1398 => x"52",
          1399 => x"08",
          1400 => x"51",
          1401 => x"81",
          1402 => x"b5",
          1403 => x"05",
          1404 => x"80",
          1405 => x"81",
          1406 => x"38",
          1407 => x"08",
          1408 => x"ff",
          1409 => x"72",
          1410 => x"08",
          1411 => x"72",
          1412 => x"06",
          1413 => x"ff",
          1414 => x"bb",
          1415 => x"d4",
          1416 => x"08",
          1417 => x"d4",
          1418 => x"08",
          1419 => x"82",
          1420 => x"fc",
          1421 => x"05",
          1422 => x"08",
          1423 => x"53",
          1424 => x"ff",
          1425 => x"b5",
          1426 => x"05",
          1427 => x"80",
          1428 => x"81",
          1429 => x"38",
          1430 => x"08",
          1431 => x"ff",
          1432 => x"72",
          1433 => x"08",
          1434 => x"72",
          1435 => x"06",
          1436 => x"ff",
          1437 => x"df",
          1438 => x"d4",
          1439 => x"08",
          1440 => x"d4",
          1441 => x"08",
          1442 => x"53",
          1443 => x"82",
          1444 => x"fc",
          1445 => x"05",
          1446 => x"08",
          1447 => x"ff",
          1448 => x"b5",
          1449 => x"05",
          1450 => x"d8",
          1451 => x"82",
          1452 => x"88",
          1453 => x"82",
          1454 => x"f0",
          1455 => x"05",
          1456 => x"08",
          1457 => x"82",
          1458 => x"f0",
          1459 => x"33",
          1460 => x"e0",
          1461 => x"82",
          1462 => x"e4",
          1463 => x"87",
          1464 => x"06",
          1465 => x"72",
          1466 => x"c3",
          1467 => x"d4",
          1468 => x"22",
          1469 => x"54",
          1470 => x"d4",
          1471 => x"23",
          1472 => x"70",
          1473 => x"53",
          1474 => x"a3",
          1475 => x"d4",
          1476 => x"08",
          1477 => x"85",
          1478 => x"39",
          1479 => x"08",
          1480 => x"52",
          1481 => x"08",
          1482 => x"51",
          1483 => x"80",
          1484 => x"d4",
          1485 => x"23",
          1486 => x"82",
          1487 => x"f8",
          1488 => x"72",
          1489 => x"81",
          1490 => x"81",
          1491 => x"d4",
          1492 => x"23",
          1493 => x"b5",
          1494 => x"05",
          1495 => x"82",
          1496 => x"e8",
          1497 => x"0b",
          1498 => x"08",
          1499 => x"ea",
          1500 => x"b5",
          1501 => x"05",
          1502 => x"b5",
          1503 => x"05",
          1504 => x"b0",
          1505 => x"39",
          1506 => x"08",
          1507 => x"8c",
          1508 => x"82",
          1509 => x"e0",
          1510 => x"53",
          1511 => x"08",
          1512 => x"82",
          1513 => x"95",
          1514 => x"b5",
          1515 => x"82",
          1516 => x"02",
          1517 => x"0c",
          1518 => x"82",
          1519 => x"53",
          1520 => x"08",
          1521 => x"52",
          1522 => x"08",
          1523 => x"51",
          1524 => x"82",
          1525 => x"70",
          1526 => x"0c",
          1527 => x"0d",
          1528 => x"0c",
          1529 => x"d4",
          1530 => x"b5",
          1531 => x"3d",
          1532 => x"82",
          1533 => x"f8",
          1534 => x"cd",
          1535 => x"11",
          1536 => x"2a",
          1537 => x"70",
          1538 => x"51",
          1539 => x"72",
          1540 => x"38",
          1541 => x"b5",
          1542 => x"05",
          1543 => x"39",
          1544 => x"08",
          1545 => x"53",
          1546 => x"b5",
          1547 => x"05",
          1548 => x"82",
          1549 => x"88",
          1550 => x"72",
          1551 => x"08",
          1552 => x"72",
          1553 => x"53",
          1554 => x"b0",
          1555 => x"9c",
          1556 => x"9c",
          1557 => x"b5",
          1558 => x"05",
          1559 => x"11",
          1560 => x"72",
          1561 => x"c8",
          1562 => x"80",
          1563 => x"38",
          1564 => x"b5",
          1565 => x"05",
          1566 => x"39",
          1567 => x"08",
          1568 => x"08",
          1569 => x"51",
          1570 => x"53",
          1571 => x"b5",
          1572 => x"72",
          1573 => x"38",
          1574 => x"b5",
          1575 => x"05",
          1576 => x"d4",
          1577 => x"08",
          1578 => x"d4",
          1579 => x"0c",
          1580 => x"d4",
          1581 => x"08",
          1582 => x"0c",
          1583 => x"82",
          1584 => x"04",
          1585 => x"08",
          1586 => x"d4",
          1587 => x"0d",
          1588 => x"b5",
          1589 => x"05",
          1590 => x"d4",
          1591 => x"08",
          1592 => x"70",
          1593 => x"81",
          1594 => x"06",
          1595 => x"51",
          1596 => x"2e",
          1597 => x"0b",
          1598 => x"08",
          1599 => x"80",
          1600 => x"b5",
          1601 => x"05",
          1602 => x"33",
          1603 => x"08",
          1604 => x"81",
          1605 => x"d4",
          1606 => x"0c",
          1607 => x"b5",
          1608 => x"05",
          1609 => x"ff",
          1610 => x"80",
          1611 => x"82",
          1612 => x"8c",
          1613 => x"b5",
          1614 => x"05",
          1615 => x"b5",
          1616 => x"05",
          1617 => x"11",
          1618 => x"72",
          1619 => x"c8",
          1620 => x"80",
          1621 => x"38",
          1622 => x"b5",
          1623 => x"05",
          1624 => x"39",
          1625 => x"08",
          1626 => x"70",
          1627 => x"08",
          1628 => x"53",
          1629 => x"08",
          1630 => x"82",
          1631 => x"87",
          1632 => x"b5",
          1633 => x"82",
          1634 => x"02",
          1635 => x"0c",
          1636 => x"82",
          1637 => x"52",
          1638 => x"08",
          1639 => x"51",
          1640 => x"b5",
          1641 => x"82",
          1642 => x"53",
          1643 => x"82",
          1644 => x"04",
          1645 => x"08",
          1646 => x"d4",
          1647 => x"0d",
          1648 => x"08",
          1649 => x"85",
          1650 => x"81",
          1651 => x"32",
          1652 => x"51",
          1653 => x"53",
          1654 => x"8d",
          1655 => x"82",
          1656 => x"fc",
          1657 => x"cb",
          1658 => x"d4",
          1659 => x"08",
          1660 => x"70",
          1661 => x"81",
          1662 => x"51",
          1663 => x"2e",
          1664 => x"82",
          1665 => x"8c",
          1666 => x"b5",
          1667 => x"05",
          1668 => x"8c",
          1669 => x"14",
          1670 => x"38",
          1671 => x"08",
          1672 => x"70",
          1673 => x"b5",
          1674 => x"05",
          1675 => x"54",
          1676 => x"34",
          1677 => x"05",
          1678 => x"b5",
          1679 => x"05",
          1680 => x"08",
          1681 => x"12",
          1682 => x"d4",
          1683 => x"08",
          1684 => x"d4",
          1685 => x"0c",
          1686 => x"d7",
          1687 => x"d4",
          1688 => x"08",
          1689 => x"08",
          1690 => x"53",
          1691 => x"08",
          1692 => x"70",
          1693 => x"53",
          1694 => x"51",
          1695 => x"2d",
          1696 => x"08",
          1697 => x"38",
          1698 => x"08",
          1699 => x"8c",
          1700 => x"05",
          1701 => x"82",
          1702 => x"88",
          1703 => x"82",
          1704 => x"fc",
          1705 => x"53",
          1706 => x"0b",
          1707 => x"08",
          1708 => x"82",
          1709 => x"fc",
          1710 => x"b5",
          1711 => x"3d",
          1712 => x"d4",
          1713 => x"b5",
          1714 => x"82",
          1715 => x"f9",
          1716 => x"b5",
          1717 => x"05",
          1718 => x"33",
          1719 => x"70",
          1720 => x"51",
          1721 => x"80",
          1722 => x"ff",
          1723 => x"d4",
          1724 => x"0c",
          1725 => x"82",
          1726 => x"88",
          1727 => x"11",
          1728 => x"2a",
          1729 => x"51",
          1730 => x"71",
          1731 => x"c5",
          1732 => x"d4",
          1733 => x"08",
          1734 => x"08",
          1735 => x"53",
          1736 => x"33",
          1737 => x"06",
          1738 => x"85",
          1739 => x"b5",
          1740 => x"05",
          1741 => x"08",
          1742 => x"12",
          1743 => x"d4",
          1744 => x"08",
          1745 => x"70",
          1746 => x"08",
          1747 => x"51",
          1748 => x"b6",
          1749 => x"d4",
          1750 => x"08",
          1751 => x"70",
          1752 => x"81",
          1753 => x"51",
          1754 => x"2e",
          1755 => x"82",
          1756 => x"88",
          1757 => x"08",
          1758 => x"b5",
          1759 => x"05",
          1760 => x"82",
          1761 => x"fc",
          1762 => x"38",
          1763 => x"08",
          1764 => x"82",
          1765 => x"88",
          1766 => x"53",
          1767 => x"70",
          1768 => x"52",
          1769 => x"34",
          1770 => x"b5",
          1771 => x"05",
          1772 => x"39",
          1773 => x"08",
          1774 => x"70",
          1775 => x"71",
          1776 => x"a1",
          1777 => x"d4",
          1778 => x"08",
          1779 => x"08",
          1780 => x"52",
          1781 => x"51",
          1782 => x"82",
          1783 => x"70",
          1784 => x"08",
          1785 => x"52",
          1786 => x"08",
          1787 => x"80",
          1788 => x"38",
          1789 => x"08",
          1790 => x"82",
          1791 => x"f4",
          1792 => x"b5",
          1793 => x"05",
          1794 => x"33",
          1795 => x"08",
          1796 => x"52",
          1797 => x"08",
          1798 => x"ff",
          1799 => x"06",
          1800 => x"b5",
          1801 => x"05",
          1802 => x"52",
          1803 => x"d4",
          1804 => x"34",
          1805 => x"b5",
          1806 => x"05",
          1807 => x"52",
          1808 => x"d4",
          1809 => x"34",
          1810 => x"08",
          1811 => x"52",
          1812 => x"08",
          1813 => x"85",
          1814 => x"0b",
          1815 => x"08",
          1816 => x"a6",
          1817 => x"d4",
          1818 => x"08",
          1819 => x"81",
          1820 => x"0c",
          1821 => x"08",
          1822 => x"70",
          1823 => x"70",
          1824 => x"08",
          1825 => x"51",
          1826 => x"b5",
          1827 => x"05",
          1828 => x"c8",
          1829 => x"0d",
          1830 => x"0c",
          1831 => x"d4",
          1832 => x"b5",
          1833 => x"3d",
          1834 => x"d4",
          1835 => x"08",
          1836 => x"08",
          1837 => x"82",
          1838 => x"8c",
          1839 => x"b5",
          1840 => x"05",
          1841 => x"d4",
          1842 => x"08",
          1843 => x"a2",
          1844 => x"d4",
          1845 => x"08",
          1846 => x"08",
          1847 => x"26",
          1848 => x"82",
          1849 => x"f8",
          1850 => x"b5",
          1851 => x"05",
          1852 => x"82",
          1853 => x"fc",
          1854 => x"27",
          1855 => x"82",
          1856 => x"fc",
          1857 => x"b5",
          1858 => x"05",
          1859 => x"b5",
          1860 => x"05",
          1861 => x"d4",
          1862 => x"08",
          1863 => x"08",
          1864 => x"05",
          1865 => x"08",
          1866 => x"82",
          1867 => x"90",
          1868 => x"05",
          1869 => x"08",
          1870 => x"82",
          1871 => x"90",
          1872 => x"05",
          1873 => x"08",
          1874 => x"82",
          1875 => x"90",
          1876 => x"2e",
          1877 => x"82",
          1878 => x"fc",
          1879 => x"05",
          1880 => x"08",
          1881 => x"82",
          1882 => x"f8",
          1883 => x"05",
          1884 => x"08",
          1885 => x"82",
          1886 => x"fc",
          1887 => x"b5",
          1888 => x"05",
          1889 => x"71",
          1890 => x"ff",
          1891 => x"b5",
          1892 => x"05",
          1893 => x"82",
          1894 => x"90",
          1895 => x"b5",
          1896 => x"05",
          1897 => x"82",
          1898 => x"90",
          1899 => x"b5",
          1900 => x"05",
          1901 => x"ba",
          1902 => x"d4",
          1903 => x"08",
          1904 => x"82",
          1905 => x"f8",
          1906 => x"05",
          1907 => x"08",
          1908 => x"82",
          1909 => x"fc",
          1910 => x"52",
          1911 => x"82",
          1912 => x"fc",
          1913 => x"05",
          1914 => x"08",
          1915 => x"ff",
          1916 => x"b5",
          1917 => x"05",
          1918 => x"b5",
          1919 => x"85",
          1920 => x"b5",
          1921 => x"82",
          1922 => x"02",
          1923 => x"0c",
          1924 => x"82",
          1925 => x"88",
          1926 => x"b5",
          1927 => x"05",
          1928 => x"d4",
          1929 => x"08",
          1930 => x"82",
          1931 => x"fc",
          1932 => x"05",
          1933 => x"08",
          1934 => x"70",
          1935 => x"51",
          1936 => x"2e",
          1937 => x"39",
          1938 => x"08",
          1939 => x"ff",
          1940 => x"d4",
          1941 => x"0c",
          1942 => x"08",
          1943 => x"82",
          1944 => x"88",
          1945 => x"70",
          1946 => x"0c",
          1947 => x"0d",
          1948 => x"0c",
          1949 => x"d4",
          1950 => x"b5",
          1951 => x"3d",
          1952 => x"d4",
          1953 => x"08",
          1954 => x"08",
          1955 => x"82",
          1956 => x"8c",
          1957 => x"71",
          1958 => x"d4",
          1959 => x"08",
          1960 => x"b5",
          1961 => x"05",
          1962 => x"d4",
          1963 => x"08",
          1964 => x"72",
          1965 => x"d4",
          1966 => x"08",
          1967 => x"b5",
          1968 => x"05",
          1969 => x"ff",
          1970 => x"80",
          1971 => x"ff",
          1972 => x"b5",
          1973 => x"05",
          1974 => x"b5",
          1975 => x"84",
          1976 => x"b5",
          1977 => x"82",
          1978 => x"02",
          1979 => x"0c",
          1980 => x"82",
          1981 => x"88",
          1982 => x"b5",
          1983 => x"05",
          1984 => x"d4",
          1985 => x"08",
          1986 => x"08",
          1987 => x"82",
          1988 => x"90",
          1989 => x"2e",
          1990 => x"82",
          1991 => x"90",
          1992 => x"05",
          1993 => x"08",
          1994 => x"82",
          1995 => x"90",
          1996 => x"05",
          1997 => x"08",
          1998 => x"82",
          1999 => x"90",
          2000 => x"2e",
          2001 => x"b5",
          2002 => x"05",
          2003 => x"33",
          2004 => x"08",
          2005 => x"81",
          2006 => x"d4",
          2007 => x"0c",
          2008 => x"08",
          2009 => x"52",
          2010 => x"34",
          2011 => x"08",
          2012 => x"81",
          2013 => x"d4",
          2014 => x"0c",
          2015 => x"82",
          2016 => x"88",
          2017 => x"82",
          2018 => x"51",
          2019 => x"82",
          2020 => x"04",
          2021 => x"08",
          2022 => x"d4",
          2023 => x"0d",
          2024 => x"08",
          2025 => x"80",
          2026 => x"38",
          2027 => x"08",
          2028 => x"52",
          2029 => x"b5",
          2030 => x"05",
          2031 => x"82",
          2032 => x"8c",
          2033 => x"b5",
          2034 => x"05",
          2035 => x"72",
          2036 => x"53",
          2037 => x"71",
          2038 => x"38",
          2039 => x"82",
          2040 => x"88",
          2041 => x"71",
          2042 => x"d4",
          2043 => x"08",
          2044 => x"b5",
          2045 => x"05",
          2046 => x"ff",
          2047 => x"70",
          2048 => x"0b",
          2049 => x"08",
          2050 => x"81",
          2051 => x"b5",
          2052 => x"05",
          2053 => x"82",
          2054 => x"90",
          2055 => x"b5",
          2056 => x"05",
          2057 => x"84",
          2058 => x"39",
          2059 => x"08",
          2060 => x"80",
          2061 => x"38",
          2062 => x"08",
          2063 => x"70",
          2064 => x"70",
          2065 => x"0b",
          2066 => x"08",
          2067 => x"80",
          2068 => x"b5",
          2069 => x"05",
          2070 => x"82",
          2071 => x"8c",
          2072 => x"b5",
          2073 => x"05",
          2074 => x"52",
          2075 => x"38",
          2076 => x"b5",
          2077 => x"05",
          2078 => x"82",
          2079 => x"88",
          2080 => x"33",
          2081 => x"08",
          2082 => x"70",
          2083 => x"31",
          2084 => x"d4",
          2085 => x"0c",
          2086 => x"52",
          2087 => x"80",
          2088 => x"d4",
          2089 => x"0c",
          2090 => x"08",
          2091 => x"82",
          2092 => x"85",
          2093 => x"b5",
          2094 => x"82",
          2095 => x"02",
          2096 => x"0c",
          2097 => x"82",
          2098 => x"88",
          2099 => x"b5",
          2100 => x"05",
          2101 => x"d4",
          2102 => x"08",
          2103 => x"0b",
          2104 => x"08",
          2105 => x"80",
          2106 => x"b5",
          2107 => x"05",
          2108 => x"33",
          2109 => x"08",
          2110 => x"81",
          2111 => x"d4",
          2112 => x"0c",
          2113 => x"06",
          2114 => x"80",
          2115 => x"82",
          2116 => x"8c",
          2117 => x"05",
          2118 => x"08",
          2119 => x"82",
          2120 => x"8c",
          2121 => x"2e",
          2122 => x"be",
          2123 => x"d4",
          2124 => x"08",
          2125 => x"b5",
          2126 => x"05",
          2127 => x"d4",
          2128 => x"08",
          2129 => x"08",
          2130 => x"31",
          2131 => x"d4",
          2132 => x"0c",
          2133 => x"d4",
          2134 => x"08",
          2135 => x"0c",
          2136 => x"82",
          2137 => x"04",
          2138 => x"08",
          2139 => x"d4",
          2140 => x"0d",
          2141 => x"08",
          2142 => x"82",
          2143 => x"fc",
          2144 => x"b5",
          2145 => x"05",
          2146 => x"80",
          2147 => x"b5",
          2148 => x"05",
          2149 => x"82",
          2150 => x"90",
          2151 => x"b5",
          2152 => x"05",
          2153 => x"82",
          2154 => x"90",
          2155 => x"b5",
          2156 => x"05",
          2157 => x"a9",
          2158 => x"d4",
          2159 => x"08",
          2160 => x"b5",
          2161 => x"05",
          2162 => x"71",
          2163 => x"b5",
          2164 => x"05",
          2165 => x"82",
          2166 => x"fc",
          2167 => x"be",
          2168 => x"d4",
          2169 => x"08",
          2170 => x"c8",
          2171 => x"3d",
          2172 => x"d4",
          2173 => x"b5",
          2174 => x"82",
          2175 => x"f9",
          2176 => x"0b",
          2177 => x"08",
          2178 => x"82",
          2179 => x"88",
          2180 => x"25",
          2181 => x"b5",
          2182 => x"05",
          2183 => x"b5",
          2184 => x"05",
          2185 => x"82",
          2186 => x"f4",
          2187 => x"b5",
          2188 => x"05",
          2189 => x"81",
          2190 => x"d4",
          2191 => x"0c",
          2192 => x"08",
          2193 => x"82",
          2194 => x"fc",
          2195 => x"b5",
          2196 => x"05",
          2197 => x"b9",
          2198 => x"d4",
          2199 => x"08",
          2200 => x"d4",
          2201 => x"0c",
          2202 => x"b5",
          2203 => x"05",
          2204 => x"d4",
          2205 => x"08",
          2206 => x"0b",
          2207 => x"08",
          2208 => x"82",
          2209 => x"f0",
          2210 => x"b5",
          2211 => x"05",
          2212 => x"82",
          2213 => x"8c",
          2214 => x"82",
          2215 => x"88",
          2216 => x"82",
          2217 => x"b5",
          2218 => x"82",
          2219 => x"f8",
          2220 => x"82",
          2221 => x"fc",
          2222 => x"2e",
          2223 => x"b5",
          2224 => x"05",
          2225 => x"b5",
          2226 => x"05",
          2227 => x"d4",
          2228 => x"08",
          2229 => x"c8",
          2230 => x"3d",
          2231 => x"d4",
          2232 => x"b5",
          2233 => x"82",
          2234 => x"fb",
          2235 => x"0b",
          2236 => x"08",
          2237 => x"82",
          2238 => x"88",
          2239 => x"25",
          2240 => x"b5",
          2241 => x"05",
          2242 => x"b5",
          2243 => x"05",
          2244 => x"82",
          2245 => x"fc",
          2246 => x"b5",
          2247 => x"05",
          2248 => x"90",
          2249 => x"d4",
          2250 => x"08",
          2251 => x"d4",
          2252 => x"0c",
          2253 => x"b5",
          2254 => x"05",
          2255 => x"b5",
          2256 => x"05",
          2257 => x"a2",
          2258 => x"c8",
          2259 => x"b5",
          2260 => x"05",
          2261 => x"b5",
          2262 => x"05",
          2263 => x"90",
          2264 => x"d4",
          2265 => x"08",
          2266 => x"d4",
          2267 => x"0c",
          2268 => x"08",
          2269 => x"70",
          2270 => x"0c",
          2271 => x"0d",
          2272 => x"0c",
          2273 => x"d4",
          2274 => x"b5",
          2275 => x"3d",
          2276 => x"82",
          2277 => x"8c",
          2278 => x"82",
          2279 => x"88",
          2280 => x"80",
          2281 => x"b5",
          2282 => x"82",
          2283 => x"54",
          2284 => x"82",
          2285 => x"04",
          2286 => x"08",
          2287 => x"d4",
          2288 => x"0d",
          2289 => x"b5",
          2290 => x"05",
          2291 => x"b5",
          2292 => x"05",
          2293 => x"3f",
          2294 => x"08",
          2295 => x"c8",
          2296 => x"3d",
          2297 => x"d4",
          2298 => x"b5",
          2299 => x"82",
          2300 => x"fd",
          2301 => x"0b",
          2302 => x"08",
          2303 => x"80",
          2304 => x"d4",
          2305 => x"0c",
          2306 => x"08",
          2307 => x"82",
          2308 => x"88",
          2309 => x"b9",
          2310 => x"d4",
          2311 => x"08",
          2312 => x"38",
          2313 => x"b5",
          2314 => x"05",
          2315 => x"38",
          2316 => x"08",
          2317 => x"10",
          2318 => x"08",
          2319 => x"82",
          2320 => x"fc",
          2321 => x"82",
          2322 => x"fc",
          2323 => x"b8",
          2324 => x"d4",
          2325 => x"08",
          2326 => x"e1",
          2327 => x"d4",
          2328 => x"08",
          2329 => x"08",
          2330 => x"26",
          2331 => x"b5",
          2332 => x"05",
          2333 => x"d4",
          2334 => x"08",
          2335 => x"d4",
          2336 => x"0c",
          2337 => x"08",
          2338 => x"82",
          2339 => x"fc",
          2340 => x"82",
          2341 => x"f8",
          2342 => x"b5",
          2343 => x"05",
          2344 => x"82",
          2345 => x"fc",
          2346 => x"b5",
          2347 => x"05",
          2348 => x"82",
          2349 => x"8c",
          2350 => x"95",
          2351 => x"d4",
          2352 => x"08",
          2353 => x"38",
          2354 => x"08",
          2355 => x"70",
          2356 => x"08",
          2357 => x"51",
          2358 => x"b5",
          2359 => x"05",
          2360 => x"b5",
          2361 => x"05",
          2362 => x"b5",
          2363 => x"05",
          2364 => x"c8",
          2365 => x"0d",
          2366 => x"0c",
          2367 => x"d4",
          2368 => x"b5",
          2369 => x"3d",
          2370 => x"82",
          2371 => x"f0",
          2372 => x"b5",
          2373 => x"05",
          2374 => x"73",
          2375 => x"d4",
          2376 => x"08",
          2377 => x"53",
          2378 => x"72",
          2379 => x"08",
          2380 => x"72",
          2381 => x"53",
          2382 => x"09",
          2383 => x"38",
          2384 => x"08",
          2385 => x"70",
          2386 => x"71",
          2387 => x"39",
          2388 => x"08",
          2389 => x"53",
          2390 => x"09",
          2391 => x"38",
          2392 => x"b5",
          2393 => x"05",
          2394 => x"d4",
          2395 => x"08",
          2396 => x"05",
          2397 => x"08",
          2398 => x"33",
          2399 => x"08",
          2400 => x"82",
          2401 => x"f8",
          2402 => x"72",
          2403 => x"81",
          2404 => x"38",
          2405 => x"08",
          2406 => x"70",
          2407 => x"71",
          2408 => x"51",
          2409 => x"82",
          2410 => x"f8",
          2411 => x"b5",
          2412 => x"05",
          2413 => x"d4",
          2414 => x"0c",
          2415 => x"08",
          2416 => x"80",
          2417 => x"38",
          2418 => x"08",
          2419 => x"80",
          2420 => x"38",
          2421 => x"90",
          2422 => x"d4",
          2423 => x"34",
          2424 => x"08",
          2425 => x"70",
          2426 => x"71",
          2427 => x"51",
          2428 => x"82",
          2429 => x"f8",
          2430 => x"a4",
          2431 => x"82",
          2432 => x"f4",
          2433 => x"b5",
          2434 => x"05",
          2435 => x"81",
          2436 => x"70",
          2437 => x"72",
          2438 => x"d4",
          2439 => x"34",
          2440 => x"82",
          2441 => x"f8",
          2442 => x"72",
          2443 => x"38",
          2444 => x"b5",
          2445 => x"05",
          2446 => x"39",
          2447 => x"08",
          2448 => x"53",
          2449 => x"90",
          2450 => x"d4",
          2451 => x"33",
          2452 => x"26",
          2453 => x"39",
          2454 => x"b5",
          2455 => x"05",
          2456 => x"39",
          2457 => x"b5",
          2458 => x"05",
          2459 => x"82",
          2460 => x"f8",
          2461 => x"af",
          2462 => x"38",
          2463 => x"08",
          2464 => x"53",
          2465 => x"83",
          2466 => x"80",
          2467 => x"d4",
          2468 => x"0c",
          2469 => x"8a",
          2470 => x"d4",
          2471 => x"34",
          2472 => x"b5",
          2473 => x"05",
          2474 => x"d4",
          2475 => x"33",
          2476 => x"27",
          2477 => x"82",
          2478 => x"f8",
          2479 => x"80",
          2480 => x"94",
          2481 => x"d4",
          2482 => x"33",
          2483 => x"53",
          2484 => x"d4",
          2485 => x"34",
          2486 => x"08",
          2487 => x"d0",
          2488 => x"72",
          2489 => x"08",
          2490 => x"82",
          2491 => x"f8",
          2492 => x"90",
          2493 => x"38",
          2494 => x"08",
          2495 => x"f9",
          2496 => x"72",
          2497 => x"08",
          2498 => x"82",
          2499 => x"f8",
          2500 => x"72",
          2501 => x"38",
          2502 => x"b5",
          2503 => x"05",
          2504 => x"39",
          2505 => x"08",
          2506 => x"82",
          2507 => x"f4",
          2508 => x"54",
          2509 => x"8d",
          2510 => x"82",
          2511 => x"ec",
          2512 => x"f7",
          2513 => x"d4",
          2514 => x"33",
          2515 => x"d4",
          2516 => x"08",
          2517 => x"d4",
          2518 => x"33",
          2519 => x"b5",
          2520 => x"05",
          2521 => x"d4",
          2522 => x"08",
          2523 => x"05",
          2524 => x"08",
          2525 => x"55",
          2526 => x"82",
          2527 => x"f8",
          2528 => x"a5",
          2529 => x"d4",
          2530 => x"33",
          2531 => x"2e",
          2532 => x"b5",
          2533 => x"05",
          2534 => x"b5",
          2535 => x"05",
          2536 => x"d4",
          2537 => x"08",
          2538 => x"08",
          2539 => x"71",
          2540 => x"0b",
          2541 => x"08",
          2542 => x"82",
          2543 => x"ec",
          2544 => x"b5",
          2545 => x"3d",
          2546 => x"d4",
          2547 => x"b5",
          2548 => x"82",
          2549 => x"f7",
          2550 => x"0b",
          2551 => x"08",
          2552 => x"82",
          2553 => x"8c",
          2554 => x"80",
          2555 => x"b5",
          2556 => x"05",
          2557 => x"51",
          2558 => x"53",
          2559 => x"d4",
          2560 => x"34",
          2561 => x"06",
          2562 => x"2e",
          2563 => x"91",
          2564 => x"d4",
          2565 => x"08",
          2566 => x"05",
          2567 => x"ce",
          2568 => x"d4",
          2569 => x"33",
          2570 => x"2e",
          2571 => x"a4",
          2572 => x"82",
          2573 => x"f0",
          2574 => x"b5",
          2575 => x"05",
          2576 => x"81",
          2577 => x"70",
          2578 => x"72",
          2579 => x"d4",
          2580 => x"34",
          2581 => x"08",
          2582 => x"53",
          2583 => x"09",
          2584 => x"dc",
          2585 => x"d4",
          2586 => x"08",
          2587 => x"05",
          2588 => x"08",
          2589 => x"33",
          2590 => x"08",
          2591 => x"82",
          2592 => x"f8",
          2593 => x"b5",
          2594 => x"05",
          2595 => x"d4",
          2596 => x"08",
          2597 => x"b6",
          2598 => x"d4",
          2599 => x"08",
          2600 => x"84",
          2601 => x"39",
          2602 => x"b5",
          2603 => x"05",
          2604 => x"d4",
          2605 => x"08",
          2606 => x"05",
          2607 => x"08",
          2608 => x"33",
          2609 => x"08",
          2610 => x"81",
          2611 => x"0b",
          2612 => x"08",
          2613 => x"82",
          2614 => x"88",
          2615 => x"08",
          2616 => x"0c",
          2617 => x"53",
          2618 => x"b5",
          2619 => x"05",
          2620 => x"39",
          2621 => x"08",
          2622 => x"53",
          2623 => x"8d",
          2624 => x"82",
          2625 => x"ec",
          2626 => x"80",
          2627 => x"d4",
          2628 => x"33",
          2629 => x"27",
          2630 => x"b5",
          2631 => x"05",
          2632 => x"b9",
          2633 => x"8d",
          2634 => x"82",
          2635 => x"ec",
          2636 => x"d8",
          2637 => x"82",
          2638 => x"f4",
          2639 => x"39",
          2640 => x"08",
          2641 => x"53",
          2642 => x"90",
          2643 => x"d4",
          2644 => x"33",
          2645 => x"26",
          2646 => x"39",
          2647 => x"b5",
          2648 => x"05",
          2649 => x"39",
          2650 => x"b5",
          2651 => x"05",
          2652 => x"82",
          2653 => x"fc",
          2654 => x"b5",
          2655 => x"05",
          2656 => x"73",
          2657 => x"38",
          2658 => x"08",
          2659 => x"53",
          2660 => x"27",
          2661 => x"b5",
          2662 => x"05",
          2663 => x"51",
          2664 => x"b5",
          2665 => x"05",
          2666 => x"d4",
          2667 => x"33",
          2668 => x"53",
          2669 => x"d4",
          2670 => x"34",
          2671 => x"08",
          2672 => x"53",
          2673 => x"ad",
          2674 => x"d4",
          2675 => x"33",
          2676 => x"53",
          2677 => x"d4",
          2678 => x"34",
          2679 => x"08",
          2680 => x"53",
          2681 => x"8d",
          2682 => x"82",
          2683 => x"ec",
          2684 => x"98",
          2685 => x"d4",
          2686 => x"33",
          2687 => x"08",
          2688 => x"54",
          2689 => x"26",
          2690 => x"0b",
          2691 => x"08",
          2692 => x"80",
          2693 => x"b5",
          2694 => x"05",
          2695 => x"b5",
          2696 => x"05",
          2697 => x"b5",
          2698 => x"05",
          2699 => x"82",
          2700 => x"fc",
          2701 => x"b5",
          2702 => x"05",
          2703 => x"81",
          2704 => x"70",
          2705 => x"52",
          2706 => x"33",
          2707 => x"08",
          2708 => x"fe",
          2709 => x"b5",
          2710 => x"05",
          2711 => x"80",
          2712 => x"82",
          2713 => x"fc",
          2714 => x"82",
          2715 => x"fc",
          2716 => x"b5",
          2717 => x"05",
          2718 => x"d4",
          2719 => x"08",
          2720 => x"81",
          2721 => x"d4",
          2722 => x"0c",
          2723 => x"08",
          2724 => x"82",
          2725 => x"8b",
          2726 => x"b5",
          2727 => x"f9",
          2728 => x"70",
          2729 => x"56",
          2730 => x"2e",
          2731 => x"95",
          2732 => x"51",
          2733 => x"82",
          2734 => x"15",
          2735 => x"16",
          2736 => x"cd",
          2737 => x"54",
          2738 => x"09",
          2739 => x"38",
          2740 => x"f1",
          2741 => x"76",
          2742 => x"b0",
          2743 => x"08",
          2744 => x"a3",
          2745 => x"c8",
          2746 => x"52",
          2747 => x"e9",
          2748 => x"b5",
          2749 => x"38",
          2750 => x"54",
          2751 => x"ff",
          2752 => x"17",
          2753 => x"06",
          2754 => x"77",
          2755 => x"ff",
          2756 => x"b5",
          2757 => x"3d",
          2758 => x"3d",
          2759 => x"71",
          2760 => x"8e",
          2761 => x"29",
          2762 => x"05",
          2763 => x"04",
          2764 => x"51",
          2765 => x"82",
          2766 => x"80",
          2767 => x"9b",
          2768 => x"f2",
          2769 => x"a0",
          2770 => x"39",
          2771 => x"51",
          2772 => x"82",
          2773 => x"80",
          2774 => x"9b",
          2775 => x"d6",
          2776 => x"e4",
          2777 => x"39",
          2778 => x"51",
          2779 => x"82",
          2780 => x"80",
          2781 => x"9c",
          2782 => x"39",
          2783 => x"51",
          2784 => x"9c",
          2785 => x"39",
          2786 => x"51",
          2787 => x"9d",
          2788 => x"39",
          2789 => x"51",
          2790 => x"9d",
          2791 => x"39",
          2792 => x"51",
          2793 => x"9d",
          2794 => x"39",
          2795 => x"51",
          2796 => x"9e",
          2797 => x"ad",
          2798 => x"0d",
          2799 => x"0d",
          2800 => x"56",
          2801 => x"26",
          2802 => x"52",
          2803 => x"29",
          2804 => x"87",
          2805 => x"51",
          2806 => x"82",
          2807 => x"52",
          2808 => x"a1",
          2809 => x"c8",
          2810 => x"53",
          2811 => x"9e",
          2812 => x"bb",
          2813 => x"3d",
          2814 => x"3d",
          2815 => x"84",
          2816 => x"05",
          2817 => x"80",
          2818 => x"70",
          2819 => x"25",
          2820 => x"59",
          2821 => x"87",
          2822 => x"38",
          2823 => x"76",
          2824 => x"ff",
          2825 => x"93",
          2826 => x"82",
          2827 => x"76",
          2828 => x"70",
          2829 => x"ff",
          2830 => x"b5",
          2831 => x"82",
          2832 => x"b9",
          2833 => x"c8",
          2834 => x"98",
          2835 => x"b5",
          2836 => x"96",
          2837 => x"54",
          2838 => x"77",
          2839 => x"81",
          2840 => x"82",
          2841 => x"57",
          2842 => x"08",
          2843 => x"55",
          2844 => x"89",
          2845 => x"75",
          2846 => x"d7",
          2847 => x"d8",
          2848 => x"8b",
          2849 => x"30",
          2850 => x"80",
          2851 => x"70",
          2852 => x"06",
          2853 => x"56",
          2854 => x"90",
          2855 => x"cc",
          2856 => x"98",
          2857 => x"78",
          2858 => x"3f",
          2859 => x"82",
          2860 => x"96",
          2861 => x"f8",
          2862 => x"02",
          2863 => x"05",
          2864 => x"ff",
          2865 => x"7b",
          2866 => x"fe",
          2867 => x"b5",
          2868 => x"38",
          2869 => x"88",
          2870 => x"2e",
          2871 => x"39",
          2872 => x"56",
          2873 => x"54",
          2874 => x"53",
          2875 => x"51",
          2876 => x"b5",
          2877 => x"83",
          2878 => x"77",
          2879 => x"0c",
          2880 => x"04",
          2881 => x"7f",
          2882 => x"8c",
          2883 => x"05",
          2884 => x"15",
          2885 => x"5c",
          2886 => x"5e",
          2887 => x"9e",
          2888 => x"b9",
          2889 => x"9e",
          2890 => x"b9",
          2891 => x"55",
          2892 => x"81",
          2893 => x"90",
          2894 => x"7b",
          2895 => x"38",
          2896 => x"74",
          2897 => x"7a",
          2898 => x"72",
          2899 => x"9e",
          2900 => x"b9",
          2901 => x"39",
          2902 => x"51",
          2903 => x"3f",
          2904 => x"80",
          2905 => x"18",
          2906 => x"27",
          2907 => x"08",
          2908 => x"d4",
          2909 => x"e2",
          2910 => x"82",
          2911 => x"ff",
          2912 => x"84",
          2913 => x"39",
          2914 => x"72",
          2915 => x"38",
          2916 => x"82",
          2917 => x"ff",
          2918 => x"89",
          2919 => x"fc",
          2920 => x"b6",
          2921 => x"55",
          2922 => x"08",
          2923 => x"d8",
          2924 => x"fc",
          2925 => x"80",
          2926 => x"9e",
          2927 => x"74",
          2928 => x"c6",
          2929 => x"70",
          2930 => x"80",
          2931 => x"27",
          2932 => x"56",
          2933 => x"74",
          2934 => x"81",
          2935 => x"06",
          2936 => x"06",
          2937 => x"80",
          2938 => x"73",
          2939 => x"8a",
          2940 => x"9c",
          2941 => x"51",
          2942 => x"cd",
          2943 => x"a0",
          2944 => x"3f",
          2945 => x"ff",
          2946 => x"9f",
          2947 => x"d5",
          2948 => x"79",
          2949 => x"9c",
          2950 => x"b5",
          2951 => x"2b",
          2952 => x"51",
          2953 => x"2e",
          2954 => x"aa",
          2955 => x"3f",
          2956 => x"08",
          2957 => x"98",
          2958 => x"32",
          2959 => x"9b",
          2960 => x"70",
          2961 => x"75",
          2962 => x"58",
          2963 => x"51",
          2964 => x"24",
          2965 => x"9b",
          2966 => x"06",
          2967 => x"53",
          2968 => x"1e",
          2969 => x"26",
          2970 => x"ff",
          2971 => x"b5",
          2972 => x"3d",
          2973 => x"3d",
          2974 => x"05",
          2975 => x"88",
          2976 => x"8c",
          2977 => x"b6",
          2978 => x"b4",
          2979 => x"a5",
          2980 => x"9f",
          2981 => x"9f",
          2982 => x"b4",
          2983 => x"82",
          2984 => x"ff",
          2985 => x"74",
          2986 => x"38",
          2987 => x"86",
          2988 => x"fe",
          2989 => x"c0",
          2990 => x"53",
          2991 => x"81",
          2992 => x"3f",
          2993 => x"51",
          2994 => x"80",
          2995 => x"3f",
          2996 => x"70",
          2997 => x"52",
          2998 => x"92",
          2999 => x"97",
          3000 => x"9f",
          3001 => x"85",
          3002 => x"97",
          3003 => x"82",
          3004 => x"06",
          3005 => x"80",
          3006 => x"81",
          3007 => x"3f",
          3008 => x"51",
          3009 => x"80",
          3010 => x"3f",
          3011 => x"70",
          3012 => x"52",
          3013 => x"92",
          3014 => x"97",
          3015 => x"a0",
          3016 => x"c9",
          3017 => x"97",
          3018 => x"84",
          3019 => x"06",
          3020 => x"80",
          3021 => x"81",
          3022 => x"3f",
          3023 => x"51",
          3024 => x"80",
          3025 => x"3f",
          3026 => x"70",
          3027 => x"52",
          3028 => x"92",
          3029 => x"96",
          3030 => x"a0",
          3031 => x"8d",
          3032 => x"96",
          3033 => x"86",
          3034 => x"06",
          3035 => x"80",
          3036 => x"81",
          3037 => x"3f",
          3038 => x"51",
          3039 => x"80",
          3040 => x"3f",
          3041 => x"70",
          3042 => x"52",
          3043 => x"92",
          3044 => x"96",
          3045 => x"a0",
          3046 => x"d1",
          3047 => x"96",
          3048 => x"88",
          3049 => x"06",
          3050 => x"80",
          3051 => x"81",
          3052 => x"3f",
          3053 => x"51",
          3054 => x"80",
          3055 => x"3f",
          3056 => x"84",
          3057 => x"fb",
          3058 => x"02",
          3059 => x"05",
          3060 => x"56",
          3061 => x"75",
          3062 => x"3f",
          3063 => x"b0",
          3064 => x"73",
          3065 => x"53",
          3066 => x"52",
          3067 => x"51",
          3068 => x"3f",
          3069 => x"08",
          3070 => x"b5",
          3071 => x"80",
          3072 => x"31",
          3073 => x"73",
          3074 => x"b0",
          3075 => x"0b",
          3076 => x"33",
          3077 => x"2e",
          3078 => x"af",
          3079 => x"c8",
          3080 => x"75",
          3081 => x"bc",
          3082 => x"c8",
          3083 => x"8b",
          3084 => x"c8",
          3085 => x"ad",
          3086 => x"82",
          3087 => x"81",
          3088 => x"82",
          3089 => x"82",
          3090 => x"0b",
          3091 => x"c4",
          3092 => x"82",
          3093 => x"06",
          3094 => x"a1",
          3095 => x"52",
          3096 => x"be",
          3097 => x"82",
          3098 => x"87",
          3099 => x"ce",
          3100 => x"70",
          3101 => x"c4",
          3102 => x"81",
          3103 => x"80",
          3104 => x"82",
          3105 => x"81",
          3106 => x"78",
          3107 => x"81",
          3108 => x"96",
          3109 => x"53",
          3110 => x"52",
          3111 => x"c7",
          3112 => x"78",
          3113 => x"f4",
          3114 => x"f1",
          3115 => x"c8",
          3116 => x"88",
          3117 => x"bc",
          3118 => x"39",
          3119 => x"5d",
          3120 => x"51",
          3121 => x"3f",
          3122 => x"46",
          3123 => x"52",
          3124 => x"f3",
          3125 => x"ff",
          3126 => x"f3",
          3127 => x"b5",
          3128 => x"2b",
          3129 => x"51",
          3130 => x"c2",
          3131 => x"38",
          3132 => x"24",
          3133 => x"bd",
          3134 => x"38",
          3135 => x"90",
          3136 => x"2e",
          3137 => x"78",
          3138 => x"da",
          3139 => x"39",
          3140 => x"2e",
          3141 => x"78",
          3142 => x"85",
          3143 => x"bf",
          3144 => x"38",
          3145 => x"78",
          3146 => x"89",
          3147 => x"80",
          3148 => x"38",
          3149 => x"2e",
          3150 => x"78",
          3151 => x"89",
          3152 => x"9f",
          3153 => x"83",
          3154 => x"38",
          3155 => x"24",
          3156 => x"81",
          3157 => x"eb",
          3158 => x"39",
          3159 => x"2e",
          3160 => x"89",
          3161 => x"3d",
          3162 => x"53",
          3163 => x"51",
          3164 => x"82",
          3165 => x"80",
          3166 => x"38",
          3167 => x"fc",
          3168 => x"84",
          3169 => x"c6",
          3170 => x"c8",
          3171 => x"fe",
          3172 => x"3d",
          3173 => x"53",
          3174 => x"51",
          3175 => x"82",
          3176 => x"86",
          3177 => x"c8",
          3178 => x"a1",
          3179 => x"b0",
          3180 => x"63",
          3181 => x"7b",
          3182 => x"38",
          3183 => x"7a",
          3184 => x"5c",
          3185 => x"26",
          3186 => x"db",
          3187 => x"ff",
          3188 => x"ff",
          3189 => x"eb",
          3190 => x"b5",
          3191 => x"2e",
          3192 => x"b4",
          3193 => x"11",
          3194 => x"05",
          3195 => x"3f",
          3196 => x"08",
          3197 => x"c8",
          3198 => x"fe",
          3199 => x"ff",
          3200 => x"eb",
          3201 => x"b5",
          3202 => x"2e",
          3203 => x"82",
          3204 => x"ff",
          3205 => x"63",
          3206 => x"27",
          3207 => x"61",
          3208 => x"81",
          3209 => x"79",
          3210 => x"05",
          3211 => x"b4",
          3212 => x"11",
          3213 => x"05",
          3214 => x"3f",
          3215 => x"08",
          3216 => x"fc",
          3217 => x"fe",
          3218 => x"ff",
          3219 => x"ea",
          3220 => x"b5",
          3221 => x"2e",
          3222 => x"b4",
          3223 => x"11",
          3224 => x"05",
          3225 => x"3f",
          3226 => x"08",
          3227 => x"d0",
          3228 => x"94",
          3229 => x"e2",
          3230 => x"79",
          3231 => x"38",
          3232 => x"7b",
          3233 => x"5b",
          3234 => x"92",
          3235 => x"7a",
          3236 => x"53",
          3237 => x"a2",
          3238 => x"ae",
          3239 => x"1a",
          3240 => x"43",
          3241 => x"8a",
          3242 => x"3f",
          3243 => x"b4",
          3244 => x"11",
          3245 => x"05",
          3246 => x"3f",
          3247 => x"08",
          3248 => x"82",
          3249 => x"59",
          3250 => x"89",
          3251 => x"ec",
          3252 => x"cd",
          3253 => x"b5",
          3254 => x"80",
          3255 => x"82",
          3256 => x"44",
          3257 => x"b4",
          3258 => x"78",
          3259 => x"38",
          3260 => x"08",
          3261 => x"82",
          3262 => x"59",
          3263 => x"88",
          3264 => x"84",
          3265 => x"39",
          3266 => x"33",
          3267 => x"2e",
          3268 => x"b4",
          3269 => x"89",
          3270 => x"9c",
          3271 => x"05",
          3272 => x"fe",
          3273 => x"ff",
          3274 => x"e9",
          3275 => x"b5",
          3276 => x"de",
          3277 => x"b4",
          3278 => x"80",
          3279 => x"82",
          3280 => x"43",
          3281 => x"82",
          3282 => x"59",
          3283 => x"88",
          3284 => x"f8",
          3285 => x"39",
          3286 => x"33",
          3287 => x"2e",
          3288 => x"b4",
          3289 => x"aa",
          3290 => x"b7",
          3291 => x"80",
          3292 => x"82",
          3293 => x"43",
          3294 => x"b4",
          3295 => x"78",
          3296 => x"38",
          3297 => x"08",
          3298 => x"82",
          3299 => x"88",
          3300 => x"3d",
          3301 => x"53",
          3302 => x"51",
          3303 => x"82",
          3304 => x"80",
          3305 => x"80",
          3306 => x"7a",
          3307 => x"38",
          3308 => x"90",
          3309 => x"70",
          3310 => x"2a",
          3311 => x"51",
          3312 => x"78",
          3313 => x"38",
          3314 => x"83",
          3315 => x"82",
          3316 => x"c8",
          3317 => x"55",
          3318 => x"53",
          3319 => x"51",
          3320 => x"82",
          3321 => x"86",
          3322 => x"3d",
          3323 => x"53",
          3324 => x"51",
          3325 => x"82",
          3326 => x"80",
          3327 => x"38",
          3328 => x"fc",
          3329 => x"84",
          3330 => x"c2",
          3331 => x"c8",
          3332 => x"a4",
          3333 => x"02",
          3334 => x"33",
          3335 => x"81",
          3336 => x"3d",
          3337 => x"53",
          3338 => x"51",
          3339 => x"82",
          3340 => x"e1",
          3341 => x"39",
          3342 => x"54",
          3343 => x"d8",
          3344 => x"96",
          3345 => x"98",
          3346 => x"f8",
          3347 => x"ff",
          3348 => x"79",
          3349 => x"59",
          3350 => x"f8",
          3351 => x"79",
          3352 => x"b4",
          3353 => x"11",
          3354 => x"05",
          3355 => x"3f",
          3356 => x"08",
          3357 => x"38",
          3358 => x"80",
          3359 => x"79",
          3360 => x"05",
          3361 => x"39",
          3362 => x"51",
          3363 => x"ff",
          3364 => x"3d",
          3365 => x"53",
          3366 => x"51",
          3367 => x"82",
          3368 => x"80",
          3369 => x"38",
          3370 => x"f0",
          3371 => x"84",
          3372 => x"c9",
          3373 => x"c8",
          3374 => x"a5",
          3375 => x"02",
          3376 => x"79",
          3377 => x"5b",
          3378 => x"b4",
          3379 => x"11",
          3380 => x"05",
          3381 => x"3f",
          3382 => x"08",
          3383 => x"e0",
          3384 => x"22",
          3385 => x"a2",
          3386 => x"a9",
          3387 => x"cd",
          3388 => x"80",
          3389 => x"51",
          3390 => x"3f",
          3391 => x"33",
          3392 => x"2e",
          3393 => x"78",
          3394 => x"38",
          3395 => x"41",
          3396 => x"3d",
          3397 => x"53",
          3398 => x"51",
          3399 => x"82",
          3400 => x"80",
          3401 => x"60",
          3402 => x"05",
          3403 => x"82",
          3404 => x"78",
          3405 => x"39",
          3406 => x"51",
          3407 => x"ff",
          3408 => x"3d",
          3409 => x"53",
          3410 => x"51",
          3411 => x"82",
          3412 => x"80",
          3413 => x"38",
          3414 => x"f0",
          3415 => x"84",
          3416 => x"99",
          3417 => x"c8",
          3418 => x"a0",
          3419 => x"71",
          3420 => x"84",
          3421 => x"3d",
          3422 => x"53",
          3423 => x"51",
          3424 => x"82",
          3425 => x"e5",
          3426 => x"39",
          3427 => x"54",
          3428 => x"f4",
          3429 => x"c2",
          3430 => x"98",
          3431 => x"f8",
          3432 => x"ff",
          3433 => x"79",
          3434 => x"59",
          3435 => x"f6",
          3436 => x"79",
          3437 => x"b4",
          3438 => x"11",
          3439 => x"05",
          3440 => x"3f",
          3441 => x"08",
          3442 => x"38",
          3443 => x"0c",
          3444 => x"05",
          3445 => x"39",
          3446 => x"51",
          3447 => x"ff",
          3448 => x"3d",
          3449 => x"53",
          3450 => x"51",
          3451 => x"82",
          3452 => x"80",
          3453 => x"38",
          3454 => x"a3",
          3455 => x"a7",
          3456 => x"59",
          3457 => x"3d",
          3458 => x"53",
          3459 => x"51",
          3460 => x"82",
          3461 => x"80",
          3462 => x"38",
          3463 => x"a3",
          3464 => x"a7",
          3465 => x"59",
          3466 => x"b5",
          3467 => x"2e",
          3468 => x"82",
          3469 => x"52",
          3470 => x"51",
          3471 => x"3f",
          3472 => x"82",
          3473 => x"c3",
          3474 => x"a6",
          3475 => x"f0",
          3476 => x"f4",
          3477 => x"3f",
          3478 => x"a8",
          3479 => x"3f",
          3480 => x"79",
          3481 => x"59",
          3482 => x"f4",
          3483 => x"7d",
          3484 => x"80",
          3485 => x"38",
          3486 => x"84",
          3487 => x"ca",
          3488 => x"c8",
          3489 => x"5b",
          3490 => x"b2",
          3491 => x"24",
          3492 => x"81",
          3493 => x"80",
          3494 => x"83",
          3495 => x"80",
          3496 => x"a4",
          3497 => x"55",
          3498 => x"54",
          3499 => x"a4",
          3500 => x"3d",
          3501 => x"51",
          3502 => x"3f",
          3503 => x"52",
          3504 => x"b0",
          3505 => x"ad",
          3506 => x"7b",
          3507 => x"8c",
          3508 => x"82",
          3509 => x"b4",
          3510 => x"05",
          3511 => x"e2",
          3512 => x"7b",
          3513 => x"82",
          3514 => x"b4",
          3515 => x"05",
          3516 => x"ce",
          3517 => x"ec",
          3518 => x"f8",
          3519 => x"64",
          3520 => x"82",
          3521 => x"82",
          3522 => x"b4",
          3523 => x"05",
          3524 => x"3f",
          3525 => x"08",
          3526 => x"08",
          3527 => x"70",
          3528 => x"25",
          3529 => x"5f",
          3530 => x"83",
          3531 => x"81",
          3532 => x"06",
          3533 => x"2e",
          3534 => x"1b",
          3535 => x"06",
          3536 => x"fe",
          3537 => x"81",
          3538 => x"32",
          3539 => x"8a",
          3540 => x"2e",
          3541 => x"f2",
          3542 => x"a4",
          3543 => x"85",
          3544 => x"39",
          3545 => x"80",
          3546 => x"f8",
          3547 => x"94",
          3548 => x"54",
          3549 => x"80",
          3550 => x"d8",
          3551 => x"b5",
          3552 => x"2b",
          3553 => x"53",
          3554 => x"52",
          3555 => x"f5",
          3556 => x"b5",
          3557 => x"75",
          3558 => x"94",
          3559 => x"54",
          3560 => x"80",
          3561 => x"d7",
          3562 => x"b5",
          3563 => x"2b",
          3564 => x"53",
          3565 => x"52",
          3566 => x"c9",
          3567 => x"b5",
          3568 => x"75",
          3569 => x"83",
          3570 => x"94",
          3571 => x"80",
          3572 => x"c0",
          3573 => x"80",
          3574 => x"80",
          3575 => x"83",
          3576 => x"99",
          3577 => x"5c",
          3578 => x"0b",
          3579 => x"88",
          3580 => x"72",
          3581 => x"9c",
          3582 => x"be",
          3583 => x"3f",
          3584 => x"51",
          3585 => x"3f",
          3586 => x"51",
          3587 => x"3f",
          3588 => x"51",
          3589 => x"81",
          3590 => x"3f",
          3591 => x"80",
          3592 => x"0d",
          3593 => x"53",
          3594 => x"52",
          3595 => x"82",
          3596 => x"81",
          3597 => x"07",
          3598 => x"52",
          3599 => x"e8",
          3600 => x"b5",
          3601 => x"3d",
          3602 => x"3d",
          3603 => x"08",
          3604 => x"73",
          3605 => x"74",
          3606 => x"38",
          3607 => x"70",
          3608 => x"81",
          3609 => x"81",
          3610 => x"39",
          3611 => x"70",
          3612 => x"81",
          3613 => x"81",
          3614 => x"54",
          3615 => x"81",
          3616 => x"06",
          3617 => x"39",
          3618 => x"80",
          3619 => x"54",
          3620 => x"83",
          3621 => x"70",
          3622 => x"38",
          3623 => x"98",
          3624 => x"52",
          3625 => x"52",
          3626 => x"2e",
          3627 => x"54",
          3628 => x"84",
          3629 => x"38",
          3630 => x"52",
          3631 => x"2e",
          3632 => x"83",
          3633 => x"70",
          3634 => x"30",
          3635 => x"76",
          3636 => x"51",
          3637 => x"88",
          3638 => x"70",
          3639 => x"34",
          3640 => x"72",
          3641 => x"b5",
          3642 => x"3d",
          3643 => x"3d",
          3644 => x"72",
          3645 => x"91",
          3646 => x"fc",
          3647 => x"51",
          3648 => x"82",
          3649 => x"85",
          3650 => x"83",
          3651 => x"72",
          3652 => x"0c",
          3653 => x"04",
          3654 => x"76",
          3655 => x"ff",
          3656 => x"81",
          3657 => x"26",
          3658 => x"83",
          3659 => x"05",
          3660 => x"70",
          3661 => x"8a",
          3662 => x"33",
          3663 => x"70",
          3664 => x"fe",
          3665 => x"33",
          3666 => x"70",
          3667 => x"f2",
          3668 => x"33",
          3669 => x"70",
          3670 => x"e6",
          3671 => x"22",
          3672 => x"74",
          3673 => x"80",
          3674 => x"13",
          3675 => x"52",
          3676 => x"26",
          3677 => x"81",
          3678 => x"98",
          3679 => x"22",
          3680 => x"bc",
          3681 => x"33",
          3682 => x"b8",
          3683 => x"33",
          3684 => x"b4",
          3685 => x"33",
          3686 => x"b0",
          3687 => x"33",
          3688 => x"ac",
          3689 => x"33",
          3690 => x"a8",
          3691 => x"c0",
          3692 => x"73",
          3693 => x"a0",
          3694 => x"87",
          3695 => x"0c",
          3696 => x"82",
          3697 => x"86",
          3698 => x"f3",
          3699 => x"5b",
          3700 => x"9c",
          3701 => x"0c",
          3702 => x"bc",
          3703 => x"7b",
          3704 => x"98",
          3705 => x"79",
          3706 => x"87",
          3707 => x"08",
          3708 => x"1c",
          3709 => x"98",
          3710 => x"79",
          3711 => x"87",
          3712 => x"08",
          3713 => x"1c",
          3714 => x"98",
          3715 => x"79",
          3716 => x"87",
          3717 => x"08",
          3718 => x"1c",
          3719 => x"98",
          3720 => x"79",
          3721 => x"80",
          3722 => x"83",
          3723 => x"59",
          3724 => x"ff",
          3725 => x"1b",
          3726 => x"1b",
          3727 => x"1b",
          3728 => x"1b",
          3729 => x"1b",
          3730 => x"83",
          3731 => x"52",
          3732 => x"51",
          3733 => x"3f",
          3734 => x"04",
          3735 => x"02",
          3736 => x"82",
          3737 => x"70",
          3738 => x"58",
          3739 => x"c0",
          3740 => x"75",
          3741 => x"38",
          3742 => x"94",
          3743 => x"70",
          3744 => x"81",
          3745 => x"52",
          3746 => x"8c",
          3747 => x"2a",
          3748 => x"51",
          3749 => x"38",
          3750 => x"70",
          3751 => x"51",
          3752 => x"8d",
          3753 => x"2a",
          3754 => x"51",
          3755 => x"be",
          3756 => x"ff",
          3757 => x"c0",
          3758 => x"70",
          3759 => x"38",
          3760 => x"90",
          3761 => x"0c",
          3762 => x"c8",
          3763 => x"0d",
          3764 => x"0d",
          3765 => x"33",
          3766 => x"9f",
          3767 => x"52",
          3768 => x"e8",
          3769 => x"0d",
          3770 => x"0d",
          3771 => x"33",
          3772 => x"2e",
          3773 => x"87",
          3774 => x"8d",
          3775 => x"82",
          3776 => x"70",
          3777 => x"58",
          3778 => x"94",
          3779 => x"80",
          3780 => x"87",
          3781 => x"53",
          3782 => x"96",
          3783 => x"06",
          3784 => x"72",
          3785 => x"38",
          3786 => x"70",
          3787 => x"53",
          3788 => x"74",
          3789 => x"81",
          3790 => x"72",
          3791 => x"38",
          3792 => x"70",
          3793 => x"53",
          3794 => x"38",
          3795 => x"06",
          3796 => x"94",
          3797 => x"80",
          3798 => x"87",
          3799 => x"54",
          3800 => x"80",
          3801 => x"c8",
          3802 => x"0d",
          3803 => x"0d",
          3804 => x"74",
          3805 => x"ff",
          3806 => x"57",
          3807 => x"80",
          3808 => x"81",
          3809 => x"15",
          3810 => x"33",
          3811 => x"06",
          3812 => x"58",
          3813 => x"84",
          3814 => x"2e",
          3815 => x"c0",
          3816 => x"70",
          3817 => x"2a",
          3818 => x"53",
          3819 => x"80",
          3820 => x"71",
          3821 => x"81",
          3822 => x"70",
          3823 => x"81",
          3824 => x"06",
          3825 => x"80",
          3826 => x"71",
          3827 => x"81",
          3828 => x"70",
          3829 => x"74",
          3830 => x"51",
          3831 => x"80",
          3832 => x"2e",
          3833 => x"c0",
          3834 => x"77",
          3835 => x"17",
          3836 => x"81",
          3837 => x"53",
          3838 => x"86",
          3839 => x"b5",
          3840 => x"3d",
          3841 => x"3d",
          3842 => x"e8",
          3843 => x"ff",
          3844 => x"87",
          3845 => x"51",
          3846 => x"86",
          3847 => x"94",
          3848 => x"08",
          3849 => x"70",
          3850 => x"51",
          3851 => x"2e",
          3852 => x"81",
          3853 => x"87",
          3854 => x"52",
          3855 => x"86",
          3856 => x"94",
          3857 => x"08",
          3858 => x"06",
          3859 => x"0c",
          3860 => x"0d",
          3861 => x"3f",
          3862 => x"08",
          3863 => x"82",
          3864 => x"04",
          3865 => x"82",
          3866 => x"70",
          3867 => x"52",
          3868 => x"94",
          3869 => x"80",
          3870 => x"87",
          3871 => x"52",
          3872 => x"82",
          3873 => x"06",
          3874 => x"ff",
          3875 => x"2e",
          3876 => x"81",
          3877 => x"87",
          3878 => x"52",
          3879 => x"86",
          3880 => x"94",
          3881 => x"08",
          3882 => x"70",
          3883 => x"53",
          3884 => x"b5",
          3885 => x"3d",
          3886 => x"3d",
          3887 => x"9e",
          3888 => x"9c",
          3889 => x"51",
          3890 => x"2e",
          3891 => x"87",
          3892 => x"08",
          3893 => x"0c",
          3894 => x"a8",
          3895 => x"f0",
          3896 => x"9e",
          3897 => x"b3",
          3898 => x"c0",
          3899 => x"82",
          3900 => x"87",
          3901 => x"08",
          3902 => x"0c",
          3903 => x"a0",
          3904 => x"80",
          3905 => x"9e",
          3906 => x"b4",
          3907 => x"c0",
          3908 => x"82",
          3909 => x"87",
          3910 => x"08",
          3911 => x"0c",
          3912 => x"b8",
          3913 => x"90",
          3914 => x"9e",
          3915 => x"b4",
          3916 => x"c0",
          3917 => x"82",
          3918 => x"87",
          3919 => x"08",
          3920 => x"0c",
          3921 => x"80",
          3922 => x"82",
          3923 => x"87",
          3924 => x"08",
          3925 => x"0c",
          3926 => x"88",
          3927 => x"a8",
          3928 => x"9e",
          3929 => x"b4",
          3930 => x"0b",
          3931 => x"34",
          3932 => x"c0",
          3933 => x"70",
          3934 => x"06",
          3935 => x"70",
          3936 => x"38",
          3937 => x"82",
          3938 => x"80",
          3939 => x"9e",
          3940 => x"88",
          3941 => x"51",
          3942 => x"80",
          3943 => x"81",
          3944 => x"b4",
          3945 => x"0b",
          3946 => x"90",
          3947 => x"80",
          3948 => x"52",
          3949 => x"2e",
          3950 => x"52",
          3951 => x"b3",
          3952 => x"87",
          3953 => x"08",
          3954 => x"80",
          3955 => x"52",
          3956 => x"83",
          3957 => x"71",
          3958 => x"34",
          3959 => x"c0",
          3960 => x"70",
          3961 => x"06",
          3962 => x"70",
          3963 => x"38",
          3964 => x"82",
          3965 => x"80",
          3966 => x"9e",
          3967 => x"90",
          3968 => x"51",
          3969 => x"80",
          3970 => x"81",
          3971 => x"b4",
          3972 => x"0b",
          3973 => x"90",
          3974 => x"80",
          3975 => x"52",
          3976 => x"2e",
          3977 => x"52",
          3978 => x"b7",
          3979 => x"87",
          3980 => x"08",
          3981 => x"80",
          3982 => x"52",
          3983 => x"83",
          3984 => x"71",
          3985 => x"34",
          3986 => x"c0",
          3987 => x"70",
          3988 => x"06",
          3989 => x"70",
          3990 => x"38",
          3991 => x"82",
          3992 => x"80",
          3993 => x"9e",
          3994 => x"80",
          3995 => x"51",
          3996 => x"80",
          3997 => x"81",
          3998 => x"b4",
          3999 => x"0b",
          4000 => x"90",
          4001 => x"80",
          4002 => x"52",
          4003 => x"83",
          4004 => x"71",
          4005 => x"34",
          4006 => x"90",
          4007 => x"80",
          4008 => x"2a",
          4009 => x"70",
          4010 => x"34",
          4011 => x"c0",
          4012 => x"70",
          4013 => x"51",
          4014 => x"80",
          4015 => x"81",
          4016 => x"b4",
          4017 => x"c0",
          4018 => x"70",
          4019 => x"70",
          4020 => x"51",
          4021 => x"b4",
          4022 => x"0b",
          4023 => x"90",
          4024 => x"06",
          4025 => x"70",
          4026 => x"38",
          4027 => x"82",
          4028 => x"87",
          4029 => x"08",
          4030 => x"51",
          4031 => x"b4",
          4032 => x"3d",
          4033 => x"3d",
          4034 => x"80",
          4035 => x"d5",
          4036 => x"b0",
          4037 => x"80",
          4038 => x"82",
          4039 => x"ff",
          4040 => x"82",
          4041 => x"ff",
          4042 => x"82",
          4043 => x"54",
          4044 => x"94",
          4045 => x"8c",
          4046 => x"90",
          4047 => x"52",
          4048 => x"51",
          4049 => x"3f",
          4050 => x"33",
          4051 => x"2e",
          4052 => x"b4",
          4053 => x"b4",
          4054 => x"54",
          4055 => x"dc",
          4056 => x"f6",
          4057 => x"b4",
          4058 => x"80",
          4059 => x"82",
          4060 => x"82",
          4061 => x"11",
          4062 => x"a5",
          4063 => x"94",
          4064 => x"b4",
          4065 => x"73",
          4066 => x"38",
          4067 => x"08",
          4068 => x"08",
          4069 => x"82",
          4070 => x"ff",
          4071 => x"82",
          4072 => x"54",
          4073 => x"94",
          4074 => x"fc",
          4075 => x"80",
          4076 => x"52",
          4077 => x"51",
          4078 => x"3f",
          4079 => x"33",
          4080 => x"2e",
          4081 => x"b4",
          4082 => x"82",
          4083 => x"ff",
          4084 => x"82",
          4085 => x"54",
          4086 => x"8e",
          4087 => x"c0",
          4088 => x"a6",
          4089 => x"93",
          4090 => x"b4",
          4091 => x"73",
          4092 => x"38",
          4093 => x"33",
          4094 => x"8c",
          4095 => x"da",
          4096 => x"b1",
          4097 => x"80",
          4098 => x"82",
          4099 => x"ff",
          4100 => x"82",
          4101 => x"54",
          4102 => x"89",
          4103 => x"c0",
          4104 => x"c1",
          4105 => x"b8",
          4106 => x"80",
          4107 => x"82",
          4108 => x"ff",
          4109 => x"82",
          4110 => x"54",
          4111 => x"89",
          4112 => x"d8",
          4113 => x"9d",
          4114 => x"ba",
          4115 => x"80",
          4116 => x"82",
          4117 => x"ff",
          4118 => x"82",
          4119 => x"ff",
          4120 => x"82",
          4121 => x"52",
          4122 => x"51",
          4123 => x"3f",
          4124 => x"08",
          4125 => x"a4",
          4126 => x"de",
          4127 => x"9c",
          4128 => x"a8",
          4129 => x"92",
          4130 => x"a8",
          4131 => x"ae",
          4132 => x"b4",
          4133 => x"82",
          4134 => x"ff",
          4135 => x"82",
          4136 => x"56",
          4137 => x"52",
          4138 => x"d9",
          4139 => x"c8",
          4140 => x"c0",
          4141 => x"31",
          4142 => x"b5",
          4143 => x"82",
          4144 => x"ff",
          4145 => x"82",
          4146 => x"54",
          4147 => x"a9",
          4148 => x"a8",
          4149 => x"84",
          4150 => x"51",
          4151 => x"82",
          4152 => x"bd",
          4153 => x"76",
          4154 => x"54",
          4155 => x"08",
          4156 => x"d0",
          4157 => x"e2",
          4158 => x"b2",
          4159 => x"80",
          4160 => x"82",
          4161 => x"56",
          4162 => x"52",
          4163 => x"f5",
          4164 => x"c8",
          4165 => x"c0",
          4166 => x"31",
          4167 => x"b5",
          4168 => x"82",
          4169 => x"ff",
          4170 => x"82",
          4171 => x"ff",
          4172 => x"87",
          4173 => x"fe",
          4174 => x"92",
          4175 => x"05",
          4176 => x"26",
          4177 => x"84",
          4178 => x"f8",
          4179 => x"08",
          4180 => x"a8",
          4181 => x"82",
          4182 => x"97",
          4183 => x"b8",
          4184 => x"82",
          4185 => x"8b",
          4186 => x"c4",
          4187 => x"82",
          4188 => x"ff",
          4189 => x"84",
          4190 => x"71",
          4191 => x"04",
          4192 => x"c0",
          4193 => x"04",
          4194 => x"08",
          4195 => x"84",
          4196 => x"3d",
          4197 => x"2b",
          4198 => x"79",
          4199 => x"98",
          4200 => x"13",
          4201 => x"51",
          4202 => x"51",
          4203 => x"82",
          4204 => x"33",
          4205 => x"74",
          4206 => x"82",
          4207 => x"08",
          4208 => x"05",
          4209 => x"71",
          4210 => x"52",
          4211 => x"09",
          4212 => x"38",
          4213 => x"82",
          4214 => x"85",
          4215 => x"fb",
          4216 => x"02",
          4217 => x"05",
          4218 => x"55",
          4219 => x"80",
          4220 => x"82",
          4221 => x"52",
          4222 => x"af",
          4223 => x"cd",
          4224 => x"a0",
          4225 => x"ac",
          4226 => x"9c",
          4227 => x"51",
          4228 => x"3f",
          4229 => x"05",
          4230 => x"34",
          4231 => x"06",
          4232 => x"77",
          4233 => x"b2",
          4234 => x"34",
          4235 => x"04",
          4236 => x"7c",
          4237 => x"b7",
          4238 => x"88",
          4239 => x"33",
          4240 => x"33",
          4241 => x"82",
          4242 => x"70",
          4243 => x"59",
          4244 => x"74",
          4245 => x"38",
          4246 => x"fa",
          4247 => x"a0",
          4248 => x"29",
          4249 => x"05",
          4250 => x"54",
          4251 => x"9d",
          4252 => x"b5",
          4253 => x"0c",
          4254 => x"33",
          4255 => x"82",
          4256 => x"70",
          4257 => x"5a",
          4258 => x"a7",
          4259 => x"78",
          4260 => x"ff",
          4261 => x"82",
          4262 => x"81",
          4263 => x"82",
          4264 => x"74",
          4265 => x"55",
          4266 => x"87",
          4267 => x"82",
          4268 => x"77",
          4269 => x"38",
          4270 => x"08",
          4271 => x"2e",
          4272 => x"b5",
          4273 => x"74",
          4274 => x"3d",
          4275 => x"76",
          4276 => x"75",
          4277 => x"88",
          4278 => x"9c",
          4279 => x"51",
          4280 => x"3f",
          4281 => x"08",
          4282 => x"e5",
          4283 => x"0d",
          4284 => x"0d",
          4285 => x"53",
          4286 => x"08",
          4287 => x"2e",
          4288 => x"51",
          4289 => x"80",
          4290 => x"14",
          4291 => x"54",
          4292 => x"e6",
          4293 => x"82",
          4294 => x"82",
          4295 => x"52",
          4296 => x"95",
          4297 => x"80",
          4298 => x"82",
          4299 => x"51",
          4300 => x"80",
          4301 => x"9c",
          4302 => x"0d",
          4303 => x"0d",
          4304 => x"52",
          4305 => x"08",
          4306 => x"b2",
          4307 => x"c8",
          4308 => x"38",
          4309 => x"08",
          4310 => x"52",
          4311 => x"52",
          4312 => x"80",
          4313 => x"c8",
          4314 => x"ba",
          4315 => x"ff",
          4316 => x"82",
          4317 => x"55",
          4318 => x"b5",
          4319 => x"9d",
          4320 => x"c8",
          4321 => x"70",
          4322 => x"80",
          4323 => x"53",
          4324 => x"17",
          4325 => x"52",
          4326 => x"be",
          4327 => x"2e",
          4328 => x"ff",
          4329 => x"3d",
          4330 => x"3d",
          4331 => x"08",
          4332 => x"5a",
          4333 => x"58",
          4334 => x"82",
          4335 => x"51",
          4336 => x"3f",
          4337 => x"08",
          4338 => x"ff",
          4339 => x"9c",
          4340 => x"80",
          4341 => x"3d",
          4342 => x"81",
          4343 => x"82",
          4344 => x"80",
          4345 => x"75",
          4346 => x"9b",
          4347 => x"c8",
          4348 => x"58",
          4349 => x"82",
          4350 => x"25",
          4351 => x"b5",
          4352 => x"05",
          4353 => x"55",
          4354 => x"74",
          4355 => x"70",
          4356 => x"2a",
          4357 => x"78",
          4358 => x"38",
          4359 => x"38",
          4360 => x"08",
          4361 => x"53",
          4362 => x"d2",
          4363 => x"c8",
          4364 => x"89",
          4365 => x"d4",
          4366 => x"9e",
          4367 => x"2e",
          4368 => x"9b",
          4369 => x"79",
          4370 => x"a9",
          4371 => x"ff",
          4372 => x"ab",
          4373 => x"82",
          4374 => x"74",
          4375 => x"77",
          4376 => x"0c",
          4377 => x"04",
          4378 => x"7c",
          4379 => x"71",
          4380 => x"59",
          4381 => x"a0",
          4382 => x"06",
          4383 => x"33",
          4384 => x"77",
          4385 => x"38",
          4386 => x"5b",
          4387 => x"56",
          4388 => x"a0",
          4389 => x"06",
          4390 => x"75",
          4391 => x"80",
          4392 => x"29",
          4393 => x"05",
          4394 => x"55",
          4395 => x"3f",
          4396 => x"08",
          4397 => x"74",
          4398 => x"b5",
          4399 => x"b5",
          4400 => x"c5",
          4401 => x"33",
          4402 => x"2e",
          4403 => x"82",
          4404 => x"b5",
          4405 => x"3f",
          4406 => x"1a",
          4407 => x"fc",
          4408 => x"05",
          4409 => x"3f",
          4410 => x"08",
          4411 => x"38",
          4412 => x"78",
          4413 => x"fd",
          4414 => x"b5",
          4415 => x"ff",
          4416 => x"85",
          4417 => x"91",
          4418 => x"70",
          4419 => x"51",
          4420 => x"27",
          4421 => x"80",
          4422 => x"b5",
          4423 => x"3d",
          4424 => x"3d",
          4425 => x"08",
          4426 => x"b4",
          4427 => x"5f",
          4428 => x"af",
          4429 => x"b5",
          4430 => x"b5",
          4431 => x"5b",
          4432 => x"38",
          4433 => x"98",
          4434 => x"73",
          4435 => x"55",
          4436 => x"81",
          4437 => x"70",
          4438 => x"56",
          4439 => x"81",
          4440 => x"51",
          4441 => x"82",
          4442 => x"82",
          4443 => x"82",
          4444 => x"80",
          4445 => x"38",
          4446 => x"52",
          4447 => x"08",
          4448 => x"fa",
          4449 => x"c8",
          4450 => x"8c",
          4451 => x"80",
          4452 => x"d1",
          4453 => x"39",
          4454 => x"08",
          4455 => x"9c",
          4456 => x"f8",
          4457 => x"70",
          4458 => x"87",
          4459 => x"b5",
          4460 => x"82",
          4461 => x"74",
          4462 => x"06",
          4463 => x"82",
          4464 => x"51",
          4465 => x"3f",
          4466 => x"08",
          4467 => x"82",
          4468 => x"25",
          4469 => x"b5",
          4470 => x"05",
          4471 => x"55",
          4472 => x"80",
          4473 => x"ff",
          4474 => x"51",
          4475 => x"81",
          4476 => x"ff",
          4477 => x"93",
          4478 => x"38",
          4479 => x"ff",
          4480 => x"06",
          4481 => x"86",
          4482 => x"b5",
          4483 => x"8c",
          4484 => x"9c",
          4485 => x"84",
          4486 => x"3f",
          4487 => x"ec",
          4488 => x"b5",
          4489 => x"2b",
          4490 => x"51",
          4491 => x"2e",
          4492 => x"81",
          4493 => x"cc",
          4494 => x"98",
          4495 => x"2c",
          4496 => x"33",
          4497 => x"70",
          4498 => x"98",
          4499 => x"84",
          4500 => x"d4",
          4501 => x"15",
          4502 => x"51",
          4503 => x"59",
          4504 => x"58",
          4505 => x"78",
          4506 => x"38",
          4507 => x"b4",
          4508 => x"80",
          4509 => x"ff",
          4510 => x"98",
          4511 => x"80",
          4512 => x"ce",
          4513 => x"74",
          4514 => x"f6",
          4515 => x"b5",
          4516 => x"ff",
          4517 => x"80",
          4518 => x"74",
          4519 => x"34",
          4520 => x"39",
          4521 => x"0a",
          4522 => x"0a",
          4523 => x"2c",
          4524 => x"06",
          4525 => x"73",
          4526 => x"38",
          4527 => x"52",
          4528 => x"ce",
          4529 => x"c8",
          4530 => x"06",
          4531 => x"38",
          4532 => x"56",
          4533 => x"80",
          4534 => x"1c",
          4535 => x"cc",
          4536 => x"98",
          4537 => x"2c",
          4538 => x"33",
          4539 => x"70",
          4540 => x"10",
          4541 => x"2b",
          4542 => x"11",
          4543 => x"51",
          4544 => x"51",
          4545 => x"2e",
          4546 => x"fe",
          4547 => x"aa",
          4548 => x"7d",
          4549 => x"82",
          4550 => x"80",
          4551 => x"f0",
          4552 => x"75",
          4553 => x"34",
          4554 => x"f0",
          4555 => x"3d",
          4556 => x"0c",
          4557 => x"95",
          4558 => x"38",
          4559 => x"82",
          4560 => x"54",
          4561 => x"82",
          4562 => x"54",
          4563 => x"fd",
          4564 => x"cc",
          4565 => x"73",
          4566 => x"38",
          4567 => x"70",
          4568 => x"55",
          4569 => x"9e",
          4570 => x"54",
          4571 => x"15",
          4572 => x"80",
          4573 => x"ff",
          4574 => x"98",
          4575 => x"fc",
          4576 => x"55",
          4577 => x"cc",
          4578 => x"11",
          4579 => x"82",
          4580 => x"73",
          4581 => x"3d",
          4582 => x"82",
          4583 => x"54",
          4584 => x"89",
          4585 => x"54",
          4586 => x"f8",
          4587 => x"fc",
          4588 => x"80",
          4589 => x"ff",
          4590 => x"98",
          4591 => x"f8",
          4592 => x"56",
          4593 => x"25",
          4594 => x"cd",
          4595 => x"74",
          4596 => x"52",
          4597 => x"dc",
          4598 => x"80",
          4599 => x"80",
          4600 => x"98",
          4601 => x"f8",
          4602 => x"55",
          4603 => x"da",
          4604 => x"fc",
          4605 => x"2b",
          4606 => x"82",
          4607 => x"5a",
          4608 => x"74",
          4609 => x"94",
          4610 => x"9c",
          4611 => x"51",
          4612 => x"3f",
          4613 => x"0a",
          4614 => x"0a",
          4615 => x"2c",
          4616 => x"33",
          4617 => x"73",
          4618 => x"38",
          4619 => x"83",
          4620 => x"0b",
          4621 => x"82",
          4622 => x"80",
          4623 => x"c8",
          4624 => x"3f",
          4625 => x"82",
          4626 => x"70",
          4627 => x"55",
          4628 => x"2e",
          4629 => x"82",
          4630 => x"ff",
          4631 => x"82",
          4632 => x"ff",
          4633 => x"82",
          4634 => x"82",
          4635 => x"52",
          4636 => x"a2",
          4637 => x"cc",
          4638 => x"98",
          4639 => x"2c",
          4640 => x"33",
          4641 => x"57",
          4642 => x"ad",
          4643 => x"54",
          4644 => x"74",
          4645 => x"9c",
          4646 => x"33",
          4647 => x"94",
          4648 => x"80",
          4649 => x"80",
          4650 => x"98",
          4651 => x"f8",
          4652 => x"55",
          4653 => x"d5",
          4654 => x"9c",
          4655 => x"51",
          4656 => x"3f",
          4657 => x"33",
          4658 => x"70",
          4659 => x"cc",
          4660 => x"51",
          4661 => x"74",
          4662 => x"38",
          4663 => x"08",
          4664 => x"ff",
          4665 => x"74",
          4666 => x"29",
          4667 => x"05",
          4668 => x"82",
          4669 => x"58",
          4670 => x"75",
          4671 => x"fa",
          4672 => x"cc",
          4673 => x"05",
          4674 => x"34",
          4675 => x"08",
          4676 => x"ff",
          4677 => x"82",
          4678 => x"79",
          4679 => x"3f",
          4680 => x"08",
          4681 => x"54",
          4682 => x"82",
          4683 => x"54",
          4684 => x"8f",
          4685 => x"73",
          4686 => x"f1",
          4687 => x"39",
          4688 => x"80",
          4689 => x"fc",
          4690 => x"82",
          4691 => x"79",
          4692 => x"0c",
          4693 => x"04",
          4694 => x"33",
          4695 => x"2e",
          4696 => x"82",
          4697 => x"52",
          4698 => x"a0",
          4699 => x"cc",
          4700 => x"05",
          4701 => x"cc",
          4702 => x"81",
          4703 => x"dd",
          4704 => x"fc",
          4705 => x"f8",
          4706 => x"73",
          4707 => x"8c",
          4708 => x"54",
          4709 => x"f8",
          4710 => x"2b",
          4711 => x"75",
          4712 => x"56",
          4713 => x"74",
          4714 => x"74",
          4715 => x"14",
          4716 => x"82",
          4717 => x"52",
          4718 => x"ff",
          4719 => x"74",
          4720 => x"29",
          4721 => x"05",
          4722 => x"82",
          4723 => x"58",
          4724 => x"75",
          4725 => x"82",
          4726 => x"52",
          4727 => x"9f",
          4728 => x"cc",
          4729 => x"98",
          4730 => x"2c",
          4731 => x"33",
          4732 => x"57",
          4733 => x"f8",
          4734 => x"cd",
          4735 => x"88",
          4736 => x"b0",
          4737 => x"80",
          4738 => x"80",
          4739 => x"98",
          4740 => x"f8",
          4741 => x"55",
          4742 => x"de",
          4743 => x"39",
          4744 => x"33",
          4745 => x"06",
          4746 => x"33",
          4747 => x"74",
          4748 => x"e8",
          4749 => x"9c",
          4750 => x"14",
          4751 => x"cc",
          4752 => x"1a",
          4753 => x"54",
          4754 => x"3f",
          4755 => x"33",
          4756 => x"06",
          4757 => x"33",
          4758 => x"75",
          4759 => x"38",
          4760 => x"82",
          4761 => x"80",
          4762 => x"c8",
          4763 => x"3f",
          4764 => x"cc",
          4765 => x"0b",
          4766 => x"34",
          4767 => x"7a",
          4768 => x"b5",
          4769 => x"74",
          4770 => x"38",
          4771 => x"a6",
          4772 => x"b5",
          4773 => x"cc",
          4774 => x"b5",
          4775 => x"ff",
          4776 => x"53",
          4777 => x"51",
          4778 => x"3f",
          4779 => x"c0",
          4780 => x"29",
          4781 => x"05",
          4782 => x"56",
          4783 => x"2e",
          4784 => x"51",
          4785 => x"3f",
          4786 => x"08",
          4787 => x"34",
          4788 => x"08",
          4789 => x"81",
          4790 => x"52",
          4791 => x"a8",
          4792 => x"1b",
          4793 => x"39",
          4794 => x"74",
          4795 => x"ac",
          4796 => x"ff",
          4797 => x"99",
          4798 => x"2e",
          4799 => x"ae",
          4800 => x"c8",
          4801 => x"80",
          4802 => x"74",
          4803 => x"f7",
          4804 => x"c8",
          4805 => x"f8",
          4806 => x"c8",
          4807 => x"06",
          4808 => x"74",
          4809 => x"ff",
          4810 => x"80",
          4811 => x"84",
          4812 => x"cc",
          4813 => x"56",
          4814 => x"2e",
          4815 => x"51",
          4816 => x"3f",
          4817 => x"08",
          4818 => x"34",
          4819 => x"08",
          4820 => x"81",
          4821 => x"52",
          4822 => x"a7",
          4823 => x"1b",
          4824 => x"ff",
          4825 => x"39",
          4826 => x"f8",
          4827 => x"34",
          4828 => x"53",
          4829 => x"33",
          4830 => x"ec",
          4831 => x"9c",
          4832 => x"fc",
          4833 => x"ff",
          4834 => x"f8",
          4835 => x"54",
          4836 => x"f5",
          4837 => x"cd",
          4838 => x"81",
          4839 => x"82",
          4840 => x"74",
          4841 => x"52",
          4842 => x"88",
          4843 => x"39",
          4844 => x"33",
          4845 => x"2e",
          4846 => x"82",
          4847 => x"52",
          4848 => x"9b",
          4849 => x"cc",
          4850 => x"05",
          4851 => x"cc",
          4852 => x"c8",
          4853 => x"0d",
          4854 => x"0b",
          4855 => x"0c",
          4856 => x"82",
          4857 => x"a0",
          4858 => x"52",
          4859 => x"51",
          4860 => x"3f",
          4861 => x"08",
          4862 => x"77",
          4863 => x"57",
          4864 => x"34",
          4865 => x"08",
          4866 => x"15",
          4867 => x"15",
          4868 => x"c0",
          4869 => x"86",
          4870 => x"87",
          4871 => x"b5",
          4872 => x"b5",
          4873 => x"05",
          4874 => x"07",
          4875 => x"ff",
          4876 => x"2a",
          4877 => x"56",
          4878 => x"34",
          4879 => x"34",
          4880 => x"22",
          4881 => x"82",
          4882 => x"05",
          4883 => x"55",
          4884 => x"15",
          4885 => x"15",
          4886 => x"0d",
          4887 => x"0d",
          4888 => x"51",
          4889 => x"8f",
          4890 => x"83",
          4891 => x"70",
          4892 => x"06",
          4893 => x"70",
          4894 => x"0c",
          4895 => x"04",
          4896 => x"02",
          4897 => x"02",
          4898 => x"05",
          4899 => x"82",
          4900 => x"71",
          4901 => x"11",
          4902 => x"73",
          4903 => x"81",
          4904 => x"88",
          4905 => x"a4",
          4906 => x"22",
          4907 => x"ff",
          4908 => x"88",
          4909 => x"52",
          4910 => x"5b",
          4911 => x"55",
          4912 => x"70",
          4913 => x"82",
          4914 => x"14",
          4915 => x"52",
          4916 => x"15",
          4917 => x"15",
          4918 => x"c0",
          4919 => x"70",
          4920 => x"33",
          4921 => x"07",
          4922 => x"8f",
          4923 => x"51",
          4924 => x"71",
          4925 => x"ff",
          4926 => x"88",
          4927 => x"51",
          4928 => x"34",
          4929 => x"06",
          4930 => x"12",
          4931 => x"c0",
          4932 => x"71",
          4933 => x"81",
          4934 => x"3d",
          4935 => x"3d",
          4936 => x"c0",
          4937 => x"05",
          4938 => x"70",
          4939 => x"11",
          4940 => x"87",
          4941 => x"8b",
          4942 => x"2b",
          4943 => x"59",
          4944 => x"72",
          4945 => x"33",
          4946 => x"71",
          4947 => x"70",
          4948 => x"56",
          4949 => x"84",
          4950 => x"85",
          4951 => x"b5",
          4952 => x"14",
          4953 => x"85",
          4954 => x"8b",
          4955 => x"2b",
          4956 => x"57",
          4957 => x"86",
          4958 => x"13",
          4959 => x"2b",
          4960 => x"2a",
          4961 => x"52",
          4962 => x"34",
          4963 => x"34",
          4964 => x"08",
          4965 => x"81",
          4966 => x"88",
          4967 => x"81",
          4968 => x"70",
          4969 => x"51",
          4970 => x"71",
          4971 => x"81",
          4972 => x"3d",
          4973 => x"3d",
          4974 => x"05",
          4975 => x"c0",
          4976 => x"2b",
          4977 => x"33",
          4978 => x"71",
          4979 => x"70",
          4980 => x"70",
          4981 => x"33",
          4982 => x"71",
          4983 => x"53",
          4984 => x"52",
          4985 => x"53",
          4986 => x"25",
          4987 => x"72",
          4988 => x"3f",
          4989 => x"08",
          4990 => x"33",
          4991 => x"71",
          4992 => x"83",
          4993 => x"11",
          4994 => x"12",
          4995 => x"2b",
          4996 => x"2b",
          4997 => x"06",
          4998 => x"51",
          4999 => x"53",
          5000 => x"88",
          5001 => x"72",
          5002 => x"73",
          5003 => x"82",
          5004 => x"70",
          5005 => x"81",
          5006 => x"8b",
          5007 => x"2b",
          5008 => x"57",
          5009 => x"70",
          5010 => x"33",
          5011 => x"07",
          5012 => x"ff",
          5013 => x"2a",
          5014 => x"58",
          5015 => x"34",
          5016 => x"34",
          5017 => x"04",
          5018 => x"82",
          5019 => x"02",
          5020 => x"05",
          5021 => x"2b",
          5022 => x"11",
          5023 => x"33",
          5024 => x"71",
          5025 => x"59",
          5026 => x"56",
          5027 => x"71",
          5028 => x"33",
          5029 => x"07",
          5030 => x"a2",
          5031 => x"07",
          5032 => x"53",
          5033 => x"53",
          5034 => x"70",
          5035 => x"82",
          5036 => x"70",
          5037 => x"81",
          5038 => x"8b",
          5039 => x"2b",
          5040 => x"57",
          5041 => x"82",
          5042 => x"13",
          5043 => x"2b",
          5044 => x"2a",
          5045 => x"52",
          5046 => x"34",
          5047 => x"34",
          5048 => x"08",
          5049 => x"33",
          5050 => x"71",
          5051 => x"82",
          5052 => x"52",
          5053 => x"0d",
          5054 => x"0d",
          5055 => x"c0",
          5056 => x"2a",
          5057 => x"ff",
          5058 => x"57",
          5059 => x"3f",
          5060 => x"08",
          5061 => x"71",
          5062 => x"33",
          5063 => x"71",
          5064 => x"83",
          5065 => x"11",
          5066 => x"12",
          5067 => x"2b",
          5068 => x"07",
          5069 => x"51",
          5070 => x"55",
          5071 => x"80",
          5072 => x"82",
          5073 => x"75",
          5074 => x"3f",
          5075 => x"84",
          5076 => x"15",
          5077 => x"2b",
          5078 => x"07",
          5079 => x"88",
          5080 => x"55",
          5081 => x"86",
          5082 => x"81",
          5083 => x"75",
          5084 => x"82",
          5085 => x"70",
          5086 => x"33",
          5087 => x"71",
          5088 => x"70",
          5089 => x"57",
          5090 => x"72",
          5091 => x"73",
          5092 => x"82",
          5093 => x"18",
          5094 => x"86",
          5095 => x"0b",
          5096 => x"82",
          5097 => x"53",
          5098 => x"34",
          5099 => x"34",
          5100 => x"08",
          5101 => x"81",
          5102 => x"88",
          5103 => x"82",
          5104 => x"70",
          5105 => x"51",
          5106 => x"74",
          5107 => x"81",
          5108 => x"3d",
          5109 => x"3d",
          5110 => x"82",
          5111 => x"84",
          5112 => x"3f",
          5113 => x"86",
          5114 => x"fe",
          5115 => x"3d",
          5116 => x"3d",
          5117 => x"52",
          5118 => x"3f",
          5119 => x"08",
          5120 => x"06",
          5121 => x"08",
          5122 => x"85",
          5123 => x"88",
          5124 => x"5f",
          5125 => x"5a",
          5126 => x"59",
          5127 => x"80",
          5128 => x"88",
          5129 => x"33",
          5130 => x"71",
          5131 => x"70",
          5132 => x"06",
          5133 => x"83",
          5134 => x"70",
          5135 => x"53",
          5136 => x"55",
          5137 => x"8a",
          5138 => x"2e",
          5139 => x"78",
          5140 => x"15",
          5141 => x"33",
          5142 => x"07",
          5143 => x"c2",
          5144 => x"ff",
          5145 => x"38",
          5146 => x"56",
          5147 => x"2b",
          5148 => x"08",
          5149 => x"81",
          5150 => x"88",
          5151 => x"81",
          5152 => x"51",
          5153 => x"5c",
          5154 => x"2e",
          5155 => x"55",
          5156 => x"78",
          5157 => x"38",
          5158 => x"80",
          5159 => x"38",
          5160 => x"09",
          5161 => x"38",
          5162 => x"f2",
          5163 => x"39",
          5164 => x"53",
          5165 => x"51",
          5166 => x"82",
          5167 => x"70",
          5168 => x"33",
          5169 => x"71",
          5170 => x"83",
          5171 => x"5a",
          5172 => x"05",
          5173 => x"83",
          5174 => x"70",
          5175 => x"59",
          5176 => x"84",
          5177 => x"81",
          5178 => x"76",
          5179 => x"82",
          5180 => x"75",
          5181 => x"11",
          5182 => x"11",
          5183 => x"33",
          5184 => x"07",
          5185 => x"53",
          5186 => x"5a",
          5187 => x"86",
          5188 => x"87",
          5189 => x"b5",
          5190 => x"1c",
          5191 => x"85",
          5192 => x"8b",
          5193 => x"2b",
          5194 => x"5a",
          5195 => x"54",
          5196 => x"34",
          5197 => x"34",
          5198 => x"08",
          5199 => x"1d",
          5200 => x"85",
          5201 => x"88",
          5202 => x"88",
          5203 => x"5f",
          5204 => x"73",
          5205 => x"75",
          5206 => x"82",
          5207 => x"1b",
          5208 => x"73",
          5209 => x"0c",
          5210 => x"04",
          5211 => x"74",
          5212 => x"c0",
          5213 => x"f4",
          5214 => x"53",
          5215 => x"8b",
          5216 => x"fc",
          5217 => x"b5",
          5218 => x"72",
          5219 => x"0c",
          5220 => x"04",
          5221 => x"64",
          5222 => x"80",
          5223 => x"82",
          5224 => x"60",
          5225 => x"06",
          5226 => x"a9",
          5227 => x"38",
          5228 => x"b8",
          5229 => x"c8",
          5230 => x"c7",
          5231 => x"38",
          5232 => x"92",
          5233 => x"83",
          5234 => x"51",
          5235 => x"82",
          5236 => x"83",
          5237 => x"82",
          5238 => x"7d",
          5239 => x"2a",
          5240 => x"ff",
          5241 => x"2b",
          5242 => x"33",
          5243 => x"71",
          5244 => x"70",
          5245 => x"83",
          5246 => x"70",
          5247 => x"05",
          5248 => x"1a",
          5249 => x"12",
          5250 => x"2b",
          5251 => x"2b",
          5252 => x"53",
          5253 => x"5c",
          5254 => x"5c",
          5255 => x"73",
          5256 => x"38",
          5257 => x"ff",
          5258 => x"70",
          5259 => x"06",
          5260 => x"16",
          5261 => x"33",
          5262 => x"07",
          5263 => x"1c",
          5264 => x"12",
          5265 => x"2b",
          5266 => x"07",
          5267 => x"52",
          5268 => x"80",
          5269 => x"78",
          5270 => x"83",
          5271 => x"41",
          5272 => x"27",
          5273 => x"60",
          5274 => x"7b",
          5275 => x"06",
          5276 => x"51",
          5277 => x"7a",
          5278 => x"06",
          5279 => x"39",
          5280 => x"7a",
          5281 => x"38",
          5282 => x"aa",
          5283 => x"39",
          5284 => x"7a",
          5285 => x"c8",
          5286 => x"82",
          5287 => x"12",
          5288 => x"2b",
          5289 => x"54",
          5290 => x"80",
          5291 => x"f7",
          5292 => x"b5",
          5293 => x"ff",
          5294 => x"54",
          5295 => x"83",
          5296 => x"c0",
          5297 => x"05",
          5298 => x"ff",
          5299 => x"82",
          5300 => x"14",
          5301 => x"83",
          5302 => x"59",
          5303 => x"39",
          5304 => x"7a",
          5305 => x"d4",
          5306 => x"f5",
          5307 => x"b5",
          5308 => x"82",
          5309 => x"12",
          5310 => x"2b",
          5311 => x"54",
          5312 => x"80",
          5313 => x"f6",
          5314 => x"b5",
          5315 => x"ff",
          5316 => x"54",
          5317 => x"83",
          5318 => x"c0",
          5319 => x"05",
          5320 => x"ff",
          5321 => x"82",
          5322 => x"14",
          5323 => x"62",
          5324 => x"5c",
          5325 => x"ff",
          5326 => x"39",
          5327 => x"54",
          5328 => x"82",
          5329 => x"5c",
          5330 => x"08",
          5331 => x"38",
          5332 => x"52",
          5333 => x"08",
          5334 => x"8b",
          5335 => x"f7",
          5336 => x"58",
          5337 => x"99",
          5338 => x"7a",
          5339 => x"f2",
          5340 => x"19",
          5341 => x"b5",
          5342 => x"84",
          5343 => x"f9",
          5344 => x"73",
          5345 => x"0c",
          5346 => x"04",
          5347 => x"77",
          5348 => x"52",
          5349 => x"3f",
          5350 => x"08",
          5351 => x"c8",
          5352 => x"8e",
          5353 => x"80",
          5354 => x"c8",
          5355 => x"9b",
          5356 => x"82",
          5357 => x"86",
          5358 => x"ff",
          5359 => x"8f",
          5360 => x"81",
          5361 => x"26",
          5362 => x"b5",
          5363 => x"52",
          5364 => x"c8",
          5365 => x"0d",
          5366 => x"0d",
          5367 => x"33",
          5368 => x"9f",
          5369 => x"53",
          5370 => x"81",
          5371 => x"38",
          5372 => x"87",
          5373 => x"11",
          5374 => x"54",
          5375 => x"84",
          5376 => x"54",
          5377 => x"87",
          5378 => x"11",
          5379 => x"0c",
          5380 => x"c0",
          5381 => x"70",
          5382 => x"70",
          5383 => x"51",
          5384 => x"8a",
          5385 => x"98",
          5386 => x"70",
          5387 => x"08",
          5388 => x"06",
          5389 => x"38",
          5390 => x"8c",
          5391 => x"80",
          5392 => x"71",
          5393 => x"14",
          5394 => x"c4",
          5395 => x"70",
          5396 => x"0c",
          5397 => x"04",
          5398 => x"60",
          5399 => x"8c",
          5400 => x"33",
          5401 => x"5b",
          5402 => x"5a",
          5403 => x"82",
          5404 => x"81",
          5405 => x"52",
          5406 => x"38",
          5407 => x"84",
          5408 => x"92",
          5409 => x"c0",
          5410 => x"87",
          5411 => x"13",
          5412 => x"57",
          5413 => x"0b",
          5414 => x"8c",
          5415 => x"0c",
          5416 => x"75",
          5417 => x"2a",
          5418 => x"51",
          5419 => x"80",
          5420 => x"7b",
          5421 => x"7b",
          5422 => x"5d",
          5423 => x"59",
          5424 => x"06",
          5425 => x"73",
          5426 => x"81",
          5427 => x"ff",
          5428 => x"72",
          5429 => x"38",
          5430 => x"8c",
          5431 => x"c3",
          5432 => x"98",
          5433 => x"71",
          5434 => x"38",
          5435 => x"2e",
          5436 => x"76",
          5437 => x"92",
          5438 => x"72",
          5439 => x"06",
          5440 => x"f7",
          5441 => x"5a",
          5442 => x"80",
          5443 => x"70",
          5444 => x"5a",
          5445 => x"80",
          5446 => x"73",
          5447 => x"06",
          5448 => x"38",
          5449 => x"fe",
          5450 => x"fc",
          5451 => x"52",
          5452 => x"83",
          5453 => x"71",
          5454 => x"b5",
          5455 => x"3d",
          5456 => x"3d",
          5457 => x"64",
          5458 => x"bf",
          5459 => x"40",
          5460 => x"59",
          5461 => x"58",
          5462 => x"82",
          5463 => x"81",
          5464 => x"52",
          5465 => x"09",
          5466 => x"b1",
          5467 => x"84",
          5468 => x"92",
          5469 => x"c0",
          5470 => x"87",
          5471 => x"13",
          5472 => x"56",
          5473 => x"87",
          5474 => x"0c",
          5475 => x"82",
          5476 => x"58",
          5477 => x"84",
          5478 => x"06",
          5479 => x"71",
          5480 => x"38",
          5481 => x"05",
          5482 => x"0c",
          5483 => x"73",
          5484 => x"81",
          5485 => x"71",
          5486 => x"38",
          5487 => x"8c",
          5488 => x"d0",
          5489 => x"98",
          5490 => x"71",
          5491 => x"38",
          5492 => x"2e",
          5493 => x"76",
          5494 => x"92",
          5495 => x"72",
          5496 => x"06",
          5497 => x"f7",
          5498 => x"59",
          5499 => x"1a",
          5500 => x"06",
          5501 => x"59",
          5502 => x"80",
          5503 => x"73",
          5504 => x"06",
          5505 => x"38",
          5506 => x"fe",
          5507 => x"fc",
          5508 => x"52",
          5509 => x"83",
          5510 => x"71",
          5511 => x"b5",
          5512 => x"3d",
          5513 => x"3d",
          5514 => x"84",
          5515 => x"33",
          5516 => x"a7",
          5517 => x"54",
          5518 => x"fa",
          5519 => x"b5",
          5520 => x"06",
          5521 => x"72",
          5522 => x"85",
          5523 => x"98",
          5524 => x"56",
          5525 => x"80",
          5526 => x"76",
          5527 => x"74",
          5528 => x"c0",
          5529 => x"54",
          5530 => x"2e",
          5531 => x"d4",
          5532 => x"2e",
          5533 => x"80",
          5534 => x"08",
          5535 => x"70",
          5536 => x"51",
          5537 => x"2e",
          5538 => x"c0",
          5539 => x"52",
          5540 => x"87",
          5541 => x"08",
          5542 => x"38",
          5543 => x"87",
          5544 => x"14",
          5545 => x"70",
          5546 => x"52",
          5547 => x"96",
          5548 => x"92",
          5549 => x"0a",
          5550 => x"39",
          5551 => x"0c",
          5552 => x"39",
          5553 => x"54",
          5554 => x"c8",
          5555 => x"0d",
          5556 => x"0d",
          5557 => x"33",
          5558 => x"88",
          5559 => x"b5",
          5560 => x"51",
          5561 => x"04",
          5562 => x"75",
          5563 => x"82",
          5564 => x"90",
          5565 => x"2b",
          5566 => x"33",
          5567 => x"88",
          5568 => x"71",
          5569 => x"c8",
          5570 => x"54",
          5571 => x"85",
          5572 => x"ff",
          5573 => x"02",
          5574 => x"05",
          5575 => x"70",
          5576 => x"05",
          5577 => x"88",
          5578 => x"72",
          5579 => x"0d",
          5580 => x"0d",
          5581 => x"52",
          5582 => x"81",
          5583 => x"70",
          5584 => x"70",
          5585 => x"05",
          5586 => x"88",
          5587 => x"72",
          5588 => x"54",
          5589 => x"2a",
          5590 => x"34",
          5591 => x"04",
          5592 => x"76",
          5593 => x"54",
          5594 => x"2e",
          5595 => x"70",
          5596 => x"33",
          5597 => x"05",
          5598 => x"11",
          5599 => x"84",
          5600 => x"fe",
          5601 => x"77",
          5602 => x"53",
          5603 => x"81",
          5604 => x"ff",
          5605 => x"f4",
          5606 => x"0d",
          5607 => x"0d",
          5608 => x"56",
          5609 => x"70",
          5610 => x"33",
          5611 => x"05",
          5612 => x"71",
          5613 => x"56",
          5614 => x"72",
          5615 => x"38",
          5616 => x"e2",
          5617 => x"b5",
          5618 => x"3d",
          5619 => x"3d",
          5620 => x"54",
          5621 => x"71",
          5622 => x"38",
          5623 => x"70",
          5624 => x"f3",
          5625 => x"82",
          5626 => x"84",
          5627 => x"80",
          5628 => x"c8",
          5629 => x"0b",
          5630 => x"0c",
          5631 => x"0d",
          5632 => x"0b",
          5633 => x"56",
          5634 => x"2e",
          5635 => x"81",
          5636 => x"08",
          5637 => x"70",
          5638 => x"33",
          5639 => x"a2",
          5640 => x"c8",
          5641 => x"09",
          5642 => x"38",
          5643 => x"08",
          5644 => x"b0",
          5645 => x"a4",
          5646 => x"9c",
          5647 => x"56",
          5648 => x"27",
          5649 => x"16",
          5650 => x"82",
          5651 => x"06",
          5652 => x"54",
          5653 => x"78",
          5654 => x"33",
          5655 => x"3f",
          5656 => x"5a",
          5657 => x"c8",
          5658 => x"0d",
          5659 => x"0d",
          5660 => x"56",
          5661 => x"b0",
          5662 => x"af",
          5663 => x"fe",
          5664 => x"b5",
          5665 => x"82",
          5666 => x"9f",
          5667 => x"74",
          5668 => x"52",
          5669 => x"51",
          5670 => x"82",
          5671 => x"80",
          5672 => x"ff",
          5673 => x"74",
          5674 => x"76",
          5675 => x"0c",
          5676 => x"04",
          5677 => x"7a",
          5678 => x"fe",
          5679 => x"b5",
          5680 => x"82",
          5681 => x"81",
          5682 => x"33",
          5683 => x"2e",
          5684 => x"80",
          5685 => x"17",
          5686 => x"81",
          5687 => x"06",
          5688 => x"84",
          5689 => x"b5",
          5690 => x"b4",
          5691 => x"56",
          5692 => x"82",
          5693 => x"84",
          5694 => x"fc",
          5695 => x"8b",
          5696 => x"52",
          5697 => x"a9",
          5698 => x"85",
          5699 => x"84",
          5700 => x"fc",
          5701 => x"17",
          5702 => x"9c",
          5703 => x"91",
          5704 => x"08",
          5705 => x"17",
          5706 => x"3f",
          5707 => x"81",
          5708 => x"19",
          5709 => x"53",
          5710 => x"17",
          5711 => x"82",
          5712 => x"18",
          5713 => x"80",
          5714 => x"33",
          5715 => x"3f",
          5716 => x"08",
          5717 => x"38",
          5718 => x"82",
          5719 => x"8a",
          5720 => x"fb",
          5721 => x"fe",
          5722 => x"08",
          5723 => x"56",
          5724 => x"74",
          5725 => x"38",
          5726 => x"75",
          5727 => x"16",
          5728 => x"53",
          5729 => x"c8",
          5730 => x"0d",
          5731 => x"0d",
          5732 => x"08",
          5733 => x"81",
          5734 => x"df",
          5735 => x"15",
          5736 => x"d7",
          5737 => x"33",
          5738 => x"82",
          5739 => x"38",
          5740 => x"89",
          5741 => x"2e",
          5742 => x"bf",
          5743 => x"2e",
          5744 => x"81",
          5745 => x"81",
          5746 => x"89",
          5747 => x"08",
          5748 => x"52",
          5749 => x"3f",
          5750 => x"08",
          5751 => x"74",
          5752 => x"14",
          5753 => x"81",
          5754 => x"2a",
          5755 => x"05",
          5756 => x"57",
          5757 => x"f5",
          5758 => x"c8",
          5759 => x"38",
          5760 => x"06",
          5761 => x"33",
          5762 => x"78",
          5763 => x"06",
          5764 => x"5c",
          5765 => x"53",
          5766 => x"38",
          5767 => x"06",
          5768 => x"39",
          5769 => x"a4",
          5770 => x"52",
          5771 => x"bd",
          5772 => x"c8",
          5773 => x"38",
          5774 => x"fe",
          5775 => x"b4",
          5776 => x"8d",
          5777 => x"c8",
          5778 => x"ff",
          5779 => x"39",
          5780 => x"a4",
          5781 => x"52",
          5782 => x"91",
          5783 => x"c8",
          5784 => x"76",
          5785 => x"fc",
          5786 => x"b4",
          5787 => x"f8",
          5788 => x"c8",
          5789 => x"06",
          5790 => x"81",
          5791 => x"b5",
          5792 => x"3d",
          5793 => x"3d",
          5794 => x"7e",
          5795 => x"82",
          5796 => x"27",
          5797 => x"76",
          5798 => x"27",
          5799 => x"75",
          5800 => x"79",
          5801 => x"38",
          5802 => x"89",
          5803 => x"2e",
          5804 => x"80",
          5805 => x"2e",
          5806 => x"81",
          5807 => x"81",
          5808 => x"89",
          5809 => x"08",
          5810 => x"52",
          5811 => x"3f",
          5812 => x"08",
          5813 => x"c8",
          5814 => x"38",
          5815 => x"06",
          5816 => x"81",
          5817 => x"06",
          5818 => x"77",
          5819 => x"2e",
          5820 => x"84",
          5821 => x"06",
          5822 => x"06",
          5823 => x"53",
          5824 => x"81",
          5825 => x"34",
          5826 => x"a4",
          5827 => x"52",
          5828 => x"d9",
          5829 => x"c8",
          5830 => x"b5",
          5831 => x"94",
          5832 => x"ff",
          5833 => x"05",
          5834 => x"54",
          5835 => x"38",
          5836 => x"74",
          5837 => x"06",
          5838 => x"07",
          5839 => x"74",
          5840 => x"39",
          5841 => x"a4",
          5842 => x"52",
          5843 => x"9d",
          5844 => x"c8",
          5845 => x"b5",
          5846 => x"d8",
          5847 => x"ff",
          5848 => x"76",
          5849 => x"06",
          5850 => x"05",
          5851 => x"3f",
          5852 => x"87",
          5853 => x"08",
          5854 => x"51",
          5855 => x"82",
          5856 => x"59",
          5857 => x"08",
          5858 => x"f0",
          5859 => x"82",
          5860 => x"06",
          5861 => x"05",
          5862 => x"54",
          5863 => x"3f",
          5864 => x"08",
          5865 => x"74",
          5866 => x"51",
          5867 => x"81",
          5868 => x"34",
          5869 => x"c8",
          5870 => x"0d",
          5871 => x"0d",
          5872 => x"72",
          5873 => x"56",
          5874 => x"27",
          5875 => x"98",
          5876 => x"9d",
          5877 => x"2e",
          5878 => x"53",
          5879 => x"51",
          5880 => x"82",
          5881 => x"54",
          5882 => x"08",
          5883 => x"93",
          5884 => x"80",
          5885 => x"54",
          5886 => x"82",
          5887 => x"54",
          5888 => x"74",
          5889 => x"fb",
          5890 => x"b5",
          5891 => x"82",
          5892 => x"80",
          5893 => x"38",
          5894 => x"08",
          5895 => x"38",
          5896 => x"08",
          5897 => x"38",
          5898 => x"52",
          5899 => x"d6",
          5900 => x"c8",
          5901 => x"98",
          5902 => x"11",
          5903 => x"57",
          5904 => x"74",
          5905 => x"81",
          5906 => x"0c",
          5907 => x"81",
          5908 => x"84",
          5909 => x"55",
          5910 => x"ff",
          5911 => x"54",
          5912 => x"c8",
          5913 => x"0d",
          5914 => x"0d",
          5915 => x"08",
          5916 => x"79",
          5917 => x"17",
          5918 => x"80",
          5919 => x"98",
          5920 => x"26",
          5921 => x"58",
          5922 => x"52",
          5923 => x"fd",
          5924 => x"74",
          5925 => x"08",
          5926 => x"38",
          5927 => x"08",
          5928 => x"c8",
          5929 => x"82",
          5930 => x"17",
          5931 => x"c8",
          5932 => x"c7",
          5933 => x"90",
          5934 => x"56",
          5935 => x"2e",
          5936 => x"77",
          5937 => x"81",
          5938 => x"38",
          5939 => x"98",
          5940 => x"26",
          5941 => x"56",
          5942 => x"51",
          5943 => x"80",
          5944 => x"c8",
          5945 => x"09",
          5946 => x"38",
          5947 => x"08",
          5948 => x"c8",
          5949 => x"30",
          5950 => x"80",
          5951 => x"07",
          5952 => x"08",
          5953 => x"55",
          5954 => x"ef",
          5955 => x"c8",
          5956 => x"95",
          5957 => x"08",
          5958 => x"27",
          5959 => x"98",
          5960 => x"89",
          5961 => x"85",
          5962 => x"db",
          5963 => x"81",
          5964 => x"17",
          5965 => x"89",
          5966 => x"75",
          5967 => x"ac",
          5968 => x"7a",
          5969 => x"3f",
          5970 => x"08",
          5971 => x"38",
          5972 => x"b5",
          5973 => x"2e",
          5974 => x"86",
          5975 => x"c8",
          5976 => x"b5",
          5977 => x"70",
          5978 => x"07",
          5979 => x"7c",
          5980 => x"55",
          5981 => x"f8",
          5982 => x"2e",
          5983 => x"ff",
          5984 => x"55",
          5985 => x"ff",
          5986 => x"76",
          5987 => x"3f",
          5988 => x"08",
          5989 => x"08",
          5990 => x"b5",
          5991 => x"80",
          5992 => x"55",
          5993 => x"94",
          5994 => x"2e",
          5995 => x"53",
          5996 => x"51",
          5997 => x"82",
          5998 => x"55",
          5999 => x"75",
          6000 => x"98",
          6001 => x"05",
          6002 => x"56",
          6003 => x"26",
          6004 => x"15",
          6005 => x"84",
          6006 => x"07",
          6007 => x"18",
          6008 => x"ff",
          6009 => x"2e",
          6010 => x"39",
          6011 => x"39",
          6012 => x"08",
          6013 => x"81",
          6014 => x"74",
          6015 => x"0c",
          6016 => x"04",
          6017 => x"7a",
          6018 => x"f3",
          6019 => x"b5",
          6020 => x"81",
          6021 => x"c8",
          6022 => x"38",
          6023 => x"51",
          6024 => x"82",
          6025 => x"82",
          6026 => x"b0",
          6027 => x"84",
          6028 => x"52",
          6029 => x"52",
          6030 => x"3f",
          6031 => x"39",
          6032 => x"8a",
          6033 => x"75",
          6034 => x"38",
          6035 => x"19",
          6036 => x"81",
          6037 => x"ed",
          6038 => x"b5",
          6039 => x"2e",
          6040 => x"15",
          6041 => x"70",
          6042 => x"07",
          6043 => x"53",
          6044 => x"75",
          6045 => x"0c",
          6046 => x"04",
          6047 => x"7a",
          6048 => x"58",
          6049 => x"f0",
          6050 => x"80",
          6051 => x"9f",
          6052 => x"80",
          6053 => x"90",
          6054 => x"17",
          6055 => x"aa",
          6056 => x"53",
          6057 => x"88",
          6058 => x"08",
          6059 => x"38",
          6060 => x"53",
          6061 => x"17",
          6062 => x"72",
          6063 => x"fe",
          6064 => x"08",
          6065 => x"80",
          6066 => x"16",
          6067 => x"2b",
          6068 => x"75",
          6069 => x"73",
          6070 => x"f5",
          6071 => x"b5",
          6072 => x"82",
          6073 => x"ff",
          6074 => x"81",
          6075 => x"c8",
          6076 => x"38",
          6077 => x"82",
          6078 => x"26",
          6079 => x"58",
          6080 => x"73",
          6081 => x"39",
          6082 => x"51",
          6083 => x"82",
          6084 => x"98",
          6085 => x"94",
          6086 => x"17",
          6087 => x"58",
          6088 => x"9a",
          6089 => x"81",
          6090 => x"74",
          6091 => x"98",
          6092 => x"83",
          6093 => x"b4",
          6094 => x"0c",
          6095 => x"82",
          6096 => x"8a",
          6097 => x"f8",
          6098 => x"70",
          6099 => x"08",
          6100 => x"57",
          6101 => x"0a",
          6102 => x"38",
          6103 => x"15",
          6104 => x"08",
          6105 => x"72",
          6106 => x"cb",
          6107 => x"ff",
          6108 => x"81",
          6109 => x"13",
          6110 => x"94",
          6111 => x"74",
          6112 => x"85",
          6113 => x"22",
          6114 => x"73",
          6115 => x"38",
          6116 => x"8a",
          6117 => x"05",
          6118 => x"06",
          6119 => x"8a",
          6120 => x"73",
          6121 => x"3f",
          6122 => x"08",
          6123 => x"81",
          6124 => x"c8",
          6125 => x"ff",
          6126 => x"82",
          6127 => x"ff",
          6128 => x"38",
          6129 => x"82",
          6130 => x"26",
          6131 => x"7b",
          6132 => x"98",
          6133 => x"55",
          6134 => x"94",
          6135 => x"73",
          6136 => x"3f",
          6137 => x"08",
          6138 => x"82",
          6139 => x"80",
          6140 => x"38",
          6141 => x"b5",
          6142 => x"2e",
          6143 => x"55",
          6144 => x"08",
          6145 => x"38",
          6146 => x"08",
          6147 => x"fb",
          6148 => x"b5",
          6149 => x"38",
          6150 => x"0c",
          6151 => x"51",
          6152 => x"82",
          6153 => x"98",
          6154 => x"90",
          6155 => x"16",
          6156 => x"15",
          6157 => x"74",
          6158 => x"0c",
          6159 => x"04",
          6160 => x"7b",
          6161 => x"5b",
          6162 => x"52",
          6163 => x"ac",
          6164 => x"c8",
          6165 => x"b5",
          6166 => x"ec",
          6167 => x"c8",
          6168 => x"17",
          6169 => x"51",
          6170 => x"82",
          6171 => x"54",
          6172 => x"08",
          6173 => x"82",
          6174 => x"9c",
          6175 => x"33",
          6176 => x"72",
          6177 => x"09",
          6178 => x"38",
          6179 => x"b5",
          6180 => x"72",
          6181 => x"55",
          6182 => x"53",
          6183 => x"8e",
          6184 => x"56",
          6185 => x"09",
          6186 => x"38",
          6187 => x"b5",
          6188 => x"81",
          6189 => x"fd",
          6190 => x"b5",
          6191 => x"82",
          6192 => x"80",
          6193 => x"38",
          6194 => x"09",
          6195 => x"38",
          6196 => x"82",
          6197 => x"8b",
          6198 => x"fd",
          6199 => x"9a",
          6200 => x"eb",
          6201 => x"b5",
          6202 => x"ff",
          6203 => x"70",
          6204 => x"53",
          6205 => x"09",
          6206 => x"38",
          6207 => x"eb",
          6208 => x"b5",
          6209 => x"2b",
          6210 => x"72",
          6211 => x"0c",
          6212 => x"04",
          6213 => x"77",
          6214 => x"ff",
          6215 => x"9a",
          6216 => x"55",
          6217 => x"76",
          6218 => x"53",
          6219 => x"09",
          6220 => x"38",
          6221 => x"52",
          6222 => x"eb",
          6223 => x"3d",
          6224 => x"3d",
          6225 => x"5b",
          6226 => x"08",
          6227 => x"15",
          6228 => x"81",
          6229 => x"15",
          6230 => x"51",
          6231 => x"82",
          6232 => x"58",
          6233 => x"08",
          6234 => x"9c",
          6235 => x"33",
          6236 => x"86",
          6237 => x"80",
          6238 => x"13",
          6239 => x"06",
          6240 => x"06",
          6241 => x"72",
          6242 => x"82",
          6243 => x"53",
          6244 => x"2e",
          6245 => x"53",
          6246 => x"a9",
          6247 => x"74",
          6248 => x"72",
          6249 => x"38",
          6250 => x"99",
          6251 => x"c8",
          6252 => x"06",
          6253 => x"88",
          6254 => x"06",
          6255 => x"54",
          6256 => x"a0",
          6257 => x"74",
          6258 => x"3f",
          6259 => x"08",
          6260 => x"c8",
          6261 => x"98",
          6262 => x"fa",
          6263 => x"80",
          6264 => x"0c",
          6265 => x"c8",
          6266 => x"0d",
          6267 => x"0d",
          6268 => x"57",
          6269 => x"73",
          6270 => x"3f",
          6271 => x"08",
          6272 => x"c8",
          6273 => x"98",
          6274 => x"75",
          6275 => x"3f",
          6276 => x"08",
          6277 => x"c8",
          6278 => x"a0",
          6279 => x"c8",
          6280 => x"14",
          6281 => x"db",
          6282 => x"a0",
          6283 => x"14",
          6284 => x"ac",
          6285 => x"83",
          6286 => x"82",
          6287 => x"87",
          6288 => x"fd",
          6289 => x"70",
          6290 => x"08",
          6291 => x"55",
          6292 => x"3f",
          6293 => x"08",
          6294 => x"13",
          6295 => x"73",
          6296 => x"83",
          6297 => x"3d",
          6298 => x"3d",
          6299 => x"57",
          6300 => x"89",
          6301 => x"17",
          6302 => x"81",
          6303 => x"70",
          6304 => x"55",
          6305 => x"08",
          6306 => x"81",
          6307 => x"52",
          6308 => x"a8",
          6309 => x"2e",
          6310 => x"84",
          6311 => x"52",
          6312 => x"09",
          6313 => x"38",
          6314 => x"81",
          6315 => x"81",
          6316 => x"73",
          6317 => x"55",
          6318 => x"55",
          6319 => x"c5",
          6320 => x"88",
          6321 => x"0b",
          6322 => x"9c",
          6323 => x"8b",
          6324 => x"17",
          6325 => x"08",
          6326 => x"52",
          6327 => x"82",
          6328 => x"76",
          6329 => x"51",
          6330 => x"82",
          6331 => x"86",
          6332 => x"12",
          6333 => x"3f",
          6334 => x"08",
          6335 => x"88",
          6336 => x"f3",
          6337 => x"70",
          6338 => x"80",
          6339 => x"51",
          6340 => x"af",
          6341 => x"81",
          6342 => x"dc",
          6343 => x"74",
          6344 => x"38",
          6345 => x"88",
          6346 => x"39",
          6347 => x"80",
          6348 => x"56",
          6349 => x"af",
          6350 => x"06",
          6351 => x"56",
          6352 => x"32",
          6353 => x"80",
          6354 => x"51",
          6355 => x"dc",
          6356 => x"1c",
          6357 => x"33",
          6358 => x"9f",
          6359 => x"ff",
          6360 => x"1c",
          6361 => x"7a",
          6362 => x"3f",
          6363 => x"08",
          6364 => x"39",
          6365 => x"a0",
          6366 => x"5e",
          6367 => x"52",
          6368 => x"ff",
          6369 => x"59",
          6370 => x"33",
          6371 => x"ae",
          6372 => x"06",
          6373 => x"78",
          6374 => x"81",
          6375 => x"32",
          6376 => x"9f",
          6377 => x"26",
          6378 => x"53",
          6379 => x"73",
          6380 => x"17",
          6381 => x"34",
          6382 => x"db",
          6383 => x"32",
          6384 => x"9f",
          6385 => x"54",
          6386 => x"2e",
          6387 => x"80",
          6388 => x"75",
          6389 => x"bd",
          6390 => x"7e",
          6391 => x"a0",
          6392 => x"bd",
          6393 => x"82",
          6394 => x"18",
          6395 => x"1a",
          6396 => x"a0",
          6397 => x"fc",
          6398 => x"32",
          6399 => x"80",
          6400 => x"30",
          6401 => x"71",
          6402 => x"51",
          6403 => x"55",
          6404 => x"ac",
          6405 => x"81",
          6406 => x"78",
          6407 => x"51",
          6408 => x"af",
          6409 => x"06",
          6410 => x"55",
          6411 => x"32",
          6412 => x"80",
          6413 => x"51",
          6414 => x"db",
          6415 => x"39",
          6416 => x"09",
          6417 => x"38",
          6418 => x"7c",
          6419 => x"54",
          6420 => x"a2",
          6421 => x"32",
          6422 => x"ae",
          6423 => x"72",
          6424 => x"9f",
          6425 => x"51",
          6426 => x"74",
          6427 => x"88",
          6428 => x"fe",
          6429 => x"98",
          6430 => x"80",
          6431 => x"75",
          6432 => x"82",
          6433 => x"33",
          6434 => x"51",
          6435 => x"82",
          6436 => x"80",
          6437 => x"78",
          6438 => x"81",
          6439 => x"5a",
          6440 => x"d2",
          6441 => x"c8",
          6442 => x"80",
          6443 => x"1c",
          6444 => x"27",
          6445 => x"79",
          6446 => x"74",
          6447 => x"7a",
          6448 => x"74",
          6449 => x"39",
          6450 => x"ae",
          6451 => x"fe",
          6452 => x"c8",
          6453 => x"ff",
          6454 => x"73",
          6455 => x"38",
          6456 => x"81",
          6457 => x"54",
          6458 => x"75",
          6459 => x"17",
          6460 => x"39",
          6461 => x"0c",
          6462 => x"99",
          6463 => x"54",
          6464 => x"2e",
          6465 => x"84",
          6466 => x"34",
          6467 => x"76",
          6468 => x"8b",
          6469 => x"81",
          6470 => x"56",
          6471 => x"80",
          6472 => x"1b",
          6473 => x"08",
          6474 => x"51",
          6475 => x"82",
          6476 => x"56",
          6477 => x"08",
          6478 => x"98",
          6479 => x"76",
          6480 => x"3f",
          6481 => x"08",
          6482 => x"c8",
          6483 => x"38",
          6484 => x"70",
          6485 => x"73",
          6486 => x"be",
          6487 => x"33",
          6488 => x"73",
          6489 => x"8b",
          6490 => x"83",
          6491 => x"06",
          6492 => x"73",
          6493 => x"53",
          6494 => x"51",
          6495 => x"82",
          6496 => x"80",
          6497 => x"75",
          6498 => x"f3",
          6499 => x"9f",
          6500 => x"1c",
          6501 => x"74",
          6502 => x"38",
          6503 => x"09",
          6504 => x"e7",
          6505 => x"2a",
          6506 => x"77",
          6507 => x"51",
          6508 => x"2e",
          6509 => x"81",
          6510 => x"80",
          6511 => x"38",
          6512 => x"ab",
          6513 => x"55",
          6514 => x"75",
          6515 => x"73",
          6516 => x"55",
          6517 => x"82",
          6518 => x"06",
          6519 => x"ab",
          6520 => x"33",
          6521 => x"70",
          6522 => x"55",
          6523 => x"2e",
          6524 => x"1b",
          6525 => x"06",
          6526 => x"52",
          6527 => x"db",
          6528 => x"c8",
          6529 => x"0c",
          6530 => x"74",
          6531 => x"0c",
          6532 => x"04",
          6533 => x"7c",
          6534 => x"08",
          6535 => x"55",
          6536 => x"59",
          6537 => x"81",
          6538 => x"70",
          6539 => x"33",
          6540 => x"52",
          6541 => x"2e",
          6542 => x"ee",
          6543 => x"2e",
          6544 => x"81",
          6545 => x"33",
          6546 => x"81",
          6547 => x"52",
          6548 => x"26",
          6549 => x"14",
          6550 => x"06",
          6551 => x"52",
          6552 => x"80",
          6553 => x"0b",
          6554 => x"59",
          6555 => x"7a",
          6556 => x"70",
          6557 => x"33",
          6558 => x"05",
          6559 => x"9f",
          6560 => x"53",
          6561 => x"89",
          6562 => x"70",
          6563 => x"54",
          6564 => x"12",
          6565 => x"26",
          6566 => x"12",
          6567 => x"06",
          6568 => x"30",
          6569 => x"51",
          6570 => x"2e",
          6571 => x"85",
          6572 => x"be",
          6573 => x"74",
          6574 => x"30",
          6575 => x"9f",
          6576 => x"2a",
          6577 => x"54",
          6578 => x"2e",
          6579 => x"15",
          6580 => x"55",
          6581 => x"ff",
          6582 => x"39",
          6583 => x"86",
          6584 => x"7c",
          6585 => x"51",
          6586 => x"cd",
          6587 => x"70",
          6588 => x"0c",
          6589 => x"04",
          6590 => x"78",
          6591 => x"83",
          6592 => x"0b",
          6593 => x"79",
          6594 => x"e2",
          6595 => x"55",
          6596 => x"08",
          6597 => x"84",
          6598 => x"df",
          6599 => x"b5",
          6600 => x"ff",
          6601 => x"83",
          6602 => x"d4",
          6603 => x"81",
          6604 => x"38",
          6605 => x"17",
          6606 => x"74",
          6607 => x"09",
          6608 => x"38",
          6609 => x"81",
          6610 => x"30",
          6611 => x"79",
          6612 => x"54",
          6613 => x"74",
          6614 => x"09",
          6615 => x"38",
          6616 => x"ae",
          6617 => x"ea",
          6618 => x"b1",
          6619 => x"c8",
          6620 => x"b5",
          6621 => x"2e",
          6622 => x"53",
          6623 => x"52",
          6624 => x"51",
          6625 => x"82",
          6626 => x"55",
          6627 => x"08",
          6628 => x"38",
          6629 => x"82",
          6630 => x"88",
          6631 => x"f2",
          6632 => x"02",
          6633 => x"cb",
          6634 => x"55",
          6635 => x"60",
          6636 => x"3f",
          6637 => x"08",
          6638 => x"80",
          6639 => x"c8",
          6640 => x"fc",
          6641 => x"c8",
          6642 => x"82",
          6643 => x"70",
          6644 => x"8c",
          6645 => x"2e",
          6646 => x"73",
          6647 => x"81",
          6648 => x"33",
          6649 => x"80",
          6650 => x"81",
          6651 => x"d7",
          6652 => x"b5",
          6653 => x"ff",
          6654 => x"06",
          6655 => x"98",
          6656 => x"2e",
          6657 => x"74",
          6658 => x"81",
          6659 => x"8a",
          6660 => x"ac",
          6661 => x"39",
          6662 => x"77",
          6663 => x"81",
          6664 => x"33",
          6665 => x"3f",
          6666 => x"08",
          6667 => x"70",
          6668 => x"55",
          6669 => x"86",
          6670 => x"80",
          6671 => x"74",
          6672 => x"81",
          6673 => x"8a",
          6674 => x"f4",
          6675 => x"53",
          6676 => x"fd",
          6677 => x"b5",
          6678 => x"ff",
          6679 => x"82",
          6680 => x"06",
          6681 => x"8c",
          6682 => x"58",
          6683 => x"f6",
          6684 => x"58",
          6685 => x"2e",
          6686 => x"fa",
          6687 => x"e8",
          6688 => x"c8",
          6689 => x"78",
          6690 => x"5a",
          6691 => x"90",
          6692 => x"75",
          6693 => x"38",
          6694 => x"3d",
          6695 => x"70",
          6696 => x"08",
          6697 => x"7a",
          6698 => x"38",
          6699 => x"51",
          6700 => x"82",
          6701 => x"81",
          6702 => x"81",
          6703 => x"38",
          6704 => x"83",
          6705 => x"38",
          6706 => x"84",
          6707 => x"38",
          6708 => x"81",
          6709 => x"38",
          6710 => x"db",
          6711 => x"b5",
          6712 => x"ff",
          6713 => x"72",
          6714 => x"09",
          6715 => x"d0",
          6716 => x"14",
          6717 => x"3f",
          6718 => x"08",
          6719 => x"06",
          6720 => x"38",
          6721 => x"51",
          6722 => x"82",
          6723 => x"58",
          6724 => x"0c",
          6725 => x"33",
          6726 => x"80",
          6727 => x"ff",
          6728 => x"ff",
          6729 => x"55",
          6730 => x"81",
          6731 => x"38",
          6732 => x"06",
          6733 => x"80",
          6734 => x"52",
          6735 => x"8a",
          6736 => x"80",
          6737 => x"ff",
          6738 => x"53",
          6739 => x"86",
          6740 => x"83",
          6741 => x"c5",
          6742 => x"f5",
          6743 => x"c8",
          6744 => x"b5",
          6745 => x"15",
          6746 => x"06",
          6747 => x"76",
          6748 => x"80",
          6749 => x"da",
          6750 => x"b5",
          6751 => x"ff",
          6752 => x"74",
          6753 => x"d4",
          6754 => x"dc",
          6755 => x"c8",
          6756 => x"c2",
          6757 => x"b9",
          6758 => x"c8",
          6759 => x"ff",
          6760 => x"56",
          6761 => x"83",
          6762 => x"14",
          6763 => x"71",
          6764 => x"5a",
          6765 => x"26",
          6766 => x"8a",
          6767 => x"74",
          6768 => x"fe",
          6769 => x"82",
          6770 => x"55",
          6771 => x"08",
          6772 => x"ec",
          6773 => x"c8",
          6774 => x"ff",
          6775 => x"83",
          6776 => x"74",
          6777 => x"26",
          6778 => x"57",
          6779 => x"26",
          6780 => x"57",
          6781 => x"56",
          6782 => x"82",
          6783 => x"15",
          6784 => x"0c",
          6785 => x"0c",
          6786 => x"a4",
          6787 => x"1d",
          6788 => x"54",
          6789 => x"2e",
          6790 => x"af",
          6791 => x"14",
          6792 => x"3f",
          6793 => x"08",
          6794 => x"06",
          6795 => x"72",
          6796 => x"79",
          6797 => x"80",
          6798 => x"d9",
          6799 => x"b5",
          6800 => x"15",
          6801 => x"2b",
          6802 => x"8d",
          6803 => x"2e",
          6804 => x"77",
          6805 => x"0c",
          6806 => x"76",
          6807 => x"38",
          6808 => x"70",
          6809 => x"81",
          6810 => x"53",
          6811 => x"89",
          6812 => x"56",
          6813 => x"08",
          6814 => x"38",
          6815 => x"15",
          6816 => x"8c",
          6817 => x"80",
          6818 => x"34",
          6819 => x"09",
          6820 => x"92",
          6821 => x"14",
          6822 => x"3f",
          6823 => x"08",
          6824 => x"06",
          6825 => x"2e",
          6826 => x"80",
          6827 => x"1b",
          6828 => x"db",
          6829 => x"b5",
          6830 => x"ea",
          6831 => x"c8",
          6832 => x"34",
          6833 => x"51",
          6834 => x"82",
          6835 => x"83",
          6836 => x"53",
          6837 => x"d5",
          6838 => x"06",
          6839 => x"b4",
          6840 => x"84",
          6841 => x"c8",
          6842 => x"85",
          6843 => x"09",
          6844 => x"38",
          6845 => x"51",
          6846 => x"82",
          6847 => x"86",
          6848 => x"f2",
          6849 => x"06",
          6850 => x"9c",
          6851 => x"d8",
          6852 => x"c8",
          6853 => x"0c",
          6854 => x"51",
          6855 => x"82",
          6856 => x"8c",
          6857 => x"74",
          6858 => x"90",
          6859 => x"53",
          6860 => x"90",
          6861 => x"15",
          6862 => x"94",
          6863 => x"56",
          6864 => x"c8",
          6865 => x"0d",
          6866 => x"0d",
          6867 => x"55",
          6868 => x"b9",
          6869 => x"53",
          6870 => x"b1",
          6871 => x"52",
          6872 => x"a9",
          6873 => x"22",
          6874 => x"57",
          6875 => x"2e",
          6876 => x"99",
          6877 => x"33",
          6878 => x"3f",
          6879 => x"08",
          6880 => x"71",
          6881 => x"74",
          6882 => x"83",
          6883 => x"78",
          6884 => x"52",
          6885 => x"c8",
          6886 => x"0d",
          6887 => x"0d",
          6888 => x"33",
          6889 => x"3d",
          6890 => x"56",
          6891 => x"8b",
          6892 => x"82",
          6893 => x"24",
          6894 => x"b5",
          6895 => x"29",
          6896 => x"05",
          6897 => x"55",
          6898 => x"84",
          6899 => x"34",
          6900 => x"80",
          6901 => x"80",
          6902 => x"75",
          6903 => x"75",
          6904 => x"38",
          6905 => x"3d",
          6906 => x"05",
          6907 => x"3f",
          6908 => x"08",
          6909 => x"b5",
          6910 => x"3d",
          6911 => x"3d",
          6912 => x"84",
          6913 => x"05",
          6914 => x"89",
          6915 => x"2e",
          6916 => x"77",
          6917 => x"54",
          6918 => x"05",
          6919 => x"84",
          6920 => x"f6",
          6921 => x"b5",
          6922 => x"82",
          6923 => x"84",
          6924 => x"5c",
          6925 => x"3d",
          6926 => x"ed",
          6927 => x"b5",
          6928 => x"82",
          6929 => x"92",
          6930 => x"d7",
          6931 => x"98",
          6932 => x"73",
          6933 => x"38",
          6934 => x"9c",
          6935 => x"80",
          6936 => x"38",
          6937 => x"95",
          6938 => x"2e",
          6939 => x"aa",
          6940 => x"ea",
          6941 => x"b5",
          6942 => x"9e",
          6943 => x"05",
          6944 => x"54",
          6945 => x"38",
          6946 => x"70",
          6947 => x"54",
          6948 => x"8e",
          6949 => x"83",
          6950 => x"88",
          6951 => x"83",
          6952 => x"83",
          6953 => x"06",
          6954 => x"80",
          6955 => x"38",
          6956 => x"51",
          6957 => x"82",
          6958 => x"56",
          6959 => x"0a",
          6960 => x"05",
          6961 => x"3f",
          6962 => x"0b",
          6963 => x"80",
          6964 => x"7a",
          6965 => x"3f",
          6966 => x"9c",
          6967 => x"d1",
          6968 => x"81",
          6969 => x"34",
          6970 => x"80",
          6971 => x"b0",
          6972 => x"54",
          6973 => x"52",
          6974 => x"05",
          6975 => x"3f",
          6976 => x"08",
          6977 => x"c8",
          6978 => x"38",
          6979 => x"82",
          6980 => x"b2",
          6981 => x"84",
          6982 => x"06",
          6983 => x"73",
          6984 => x"38",
          6985 => x"ad",
          6986 => x"2a",
          6987 => x"51",
          6988 => x"2e",
          6989 => x"81",
          6990 => x"80",
          6991 => x"87",
          6992 => x"39",
          6993 => x"51",
          6994 => x"82",
          6995 => x"7b",
          6996 => x"12",
          6997 => x"82",
          6998 => x"81",
          6999 => x"83",
          7000 => x"06",
          7001 => x"80",
          7002 => x"77",
          7003 => x"58",
          7004 => x"08",
          7005 => x"63",
          7006 => x"63",
          7007 => x"57",
          7008 => x"82",
          7009 => x"82",
          7010 => x"88",
          7011 => x"9c",
          7012 => x"d2",
          7013 => x"b5",
          7014 => x"b5",
          7015 => x"1b",
          7016 => x"0c",
          7017 => x"22",
          7018 => x"77",
          7019 => x"80",
          7020 => x"34",
          7021 => x"1a",
          7022 => x"94",
          7023 => x"85",
          7024 => x"06",
          7025 => x"80",
          7026 => x"38",
          7027 => x"08",
          7028 => x"84",
          7029 => x"c8",
          7030 => x"0c",
          7031 => x"70",
          7032 => x"52",
          7033 => x"39",
          7034 => x"51",
          7035 => x"82",
          7036 => x"57",
          7037 => x"08",
          7038 => x"38",
          7039 => x"b5",
          7040 => x"2e",
          7041 => x"83",
          7042 => x"75",
          7043 => x"74",
          7044 => x"07",
          7045 => x"54",
          7046 => x"8a",
          7047 => x"75",
          7048 => x"73",
          7049 => x"98",
          7050 => x"a9",
          7051 => x"ff",
          7052 => x"80",
          7053 => x"76",
          7054 => x"d6",
          7055 => x"b5",
          7056 => x"38",
          7057 => x"39",
          7058 => x"82",
          7059 => x"05",
          7060 => x"84",
          7061 => x"0c",
          7062 => x"82",
          7063 => x"97",
          7064 => x"f2",
          7065 => x"63",
          7066 => x"40",
          7067 => x"7e",
          7068 => x"fc",
          7069 => x"51",
          7070 => x"82",
          7071 => x"55",
          7072 => x"08",
          7073 => x"19",
          7074 => x"80",
          7075 => x"74",
          7076 => x"39",
          7077 => x"81",
          7078 => x"56",
          7079 => x"82",
          7080 => x"39",
          7081 => x"1a",
          7082 => x"82",
          7083 => x"0b",
          7084 => x"81",
          7085 => x"39",
          7086 => x"94",
          7087 => x"55",
          7088 => x"83",
          7089 => x"7b",
          7090 => x"89",
          7091 => x"08",
          7092 => x"06",
          7093 => x"81",
          7094 => x"8a",
          7095 => x"05",
          7096 => x"06",
          7097 => x"a8",
          7098 => x"38",
          7099 => x"55",
          7100 => x"19",
          7101 => x"51",
          7102 => x"82",
          7103 => x"55",
          7104 => x"ff",
          7105 => x"ff",
          7106 => x"38",
          7107 => x"0c",
          7108 => x"52",
          7109 => x"cb",
          7110 => x"c8",
          7111 => x"ff",
          7112 => x"b5",
          7113 => x"7c",
          7114 => x"57",
          7115 => x"80",
          7116 => x"1a",
          7117 => x"22",
          7118 => x"75",
          7119 => x"38",
          7120 => x"58",
          7121 => x"53",
          7122 => x"1b",
          7123 => x"88",
          7124 => x"c8",
          7125 => x"38",
          7126 => x"33",
          7127 => x"80",
          7128 => x"b0",
          7129 => x"31",
          7130 => x"27",
          7131 => x"80",
          7132 => x"52",
          7133 => x"77",
          7134 => x"7d",
          7135 => x"e0",
          7136 => x"2b",
          7137 => x"76",
          7138 => x"94",
          7139 => x"ff",
          7140 => x"71",
          7141 => x"7b",
          7142 => x"38",
          7143 => x"19",
          7144 => x"51",
          7145 => x"82",
          7146 => x"fe",
          7147 => x"53",
          7148 => x"83",
          7149 => x"b4",
          7150 => x"51",
          7151 => x"7b",
          7152 => x"08",
          7153 => x"76",
          7154 => x"08",
          7155 => x"0c",
          7156 => x"f3",
          7157 => x"75",
          7158 => x"0c",
          7159 => x"04",
          7160 => x"60",
          7161 => x"40",
          7162 => x"80",
          7163 => x"3d",
          7164 => x"77",
          7165 => x"3f",
          7166 => x"08",
          7167 => x"c8",
          7168 => x"91",
          7169 => x"74",
          7170 => x"38",
          7171 => x"b8",
          7172 => x"33",
          7173 => x"70",
          7174 => x"56",
          7175 => x"74",
          7176 => x"a4",
          7177 => x"82",
          7178 => x"34",
          7179 => x"98",
          7180 => x"91",
          7181 => x"56",
          7182 => x"94",
          7183 => x"11",
          7184 => x"76",
          7185 => x"75",
          7186 => x"80",
          7187 => x"38",
          7188 => x"70",
          7189 => x"56",
          7190 => x"fd",
          7191 => x"11",
          7192 => x"77",
          7193 => x"5c",
          7194 => x"38",
          7195 => x"88",
          7196 => x"74",
          7197 => x"52",
          7198 => x"18",
          7199 => x"51",
          7200 => x"82",
          7201 => x"55",
          7202 => x"08",
          7203 => x"ab",
          7204 => x"2e",
          7205 => x"74",
          7206 => x"95",
          7207 => x"19",
          7208 => x"08",
          7209 => x"88",
          7210 => x"55",
          7211 => x"9c",
          7212 => x"09",
          7213 => x"38",
          7214 => x"c1",
          7215 => x"c8",
          7216 => x"38",
          7217 => x"52",
          7218 => x"97",
          7219 => x"c8",
          7220 => x"fe",
          7221 => x"b5",
          7222 => x"7c",
          7223 => x"57",
          7224 => x"80",
          7225 => x"1b",
          7226 => x"22",
          7227 => x"75",
          7228 => x"38",
          7229 => x"59",
          7230 => x"53",
          7231 => x"1a",
          7232 => x"be",
          7233 => x"c8",
          7234 => x"38",
          7235 => x"08",
          7236 => x"56",
          7237 => x"9b",
          7238 => x"53",
          7239 => x"77",
          7240 => x"7d",
          7241 => x"16",
          7242 => x"3f",
          7243 => x"0b",
          7244 => x"78",
          7245 => x"80",
          7246 => x"18",
          7247 => x"08",
          7248 => x"7e",
          7249 => x"3f",
          7250 => x"08",
          7251 => x"7e",
          7252 => x"0c",
          7253 => x"19",
          7254 => x"08",
          7255 => x"84",
          7256 => x"57",
          7257 => x"27",
          7258 => x"56",
          7259 => x"52",
          7260 => x"f9",
          7261 => x"c8",
          7262 => x"38",
          7263 => x"52",
          7264 => x"83",
          7265 => x"b4",
          7266 => x"d4",
          7267 => x"81",
          7268 => x"34",
          7269 => x"7e",
          7270 => x"0c",
          7271 => x"1a",
          7272 => x"94",
          7273 => x"1b",
          7274 => x"5e",
          7275 => x"27",
          7276 => x"55",
          7277 => x"0c",
          7278 => x"90",
          7279 => x"c0",
          7280 => x"90",
          7281 => x"56",
          7282 => x"c8",
          7283 => x"0d",
          7284 => x"0d",
          7285 => x"fc",
          7286 => x"52",
          7287 => x"3f",
          7288 => x"08",
          7289 => x"c8",
          7290 => x"38",
          7291 => x"70",
          7292 => x"81",
          7293 => x"55",
          7294 => x"80",
          7295 => x"16",
          7296 => x"51",
          7297 => x"82",
          7298 => x"57",
          7299 => x"08",
          7300 => x"a4",
          7301 => x"11",
          7302 => x"55",
          7303 => x"16",
          7304 => x"08",
          7305 => x"75",
          7306 => x"e8",
          7307 => x"08",
          7308 => x"51",
          7309 => x"82",
          7310 => x"52",
          7311 => x"c9",
          7312 => x"52",
          7313 => x"c9",
          7314 => x"54",
          7315 => x"15",
          7316 => x"cc",
          7317 => x"b5",
          7318 => x"17",
          7319 => x"06",
          7320 => x"90",
          7321 => x"82",
          7322 => x"8a",
          7323 => x"fc",
          7324 => x"70",
          7325 => x"d9",
          7326 => x"c8",
          7327 => x"b5",
          7328 => x"38",
          7329 => x"05",
          7330 => x"f1",
          7331 => x"b5",
          7332 => x"82",
          7333 => x"87",
          7334 => x"c8",
          7335 => x"72",
          7336 => x"0c",
          7337 => x"04",
          7338 => x"84",
          7339 => x"e4",
          7340 => x"80",
          7341 => x"c8",
          7342 => x"38",
          7343 => x"08",
          7344 => x"34",
          7345 => x"82",
          7346 => x"83",
          7347 => x"ef",
          7348 => x"53",
          7349 => x"05",
          7350 => x"51",
          7351 => x"82",
          7352 => x"55",
          7353 => x"08",
          7354 => x"76",
          7355 => x"93",
          7356 => x"51",
          7357 => x"82",
          7358 => x"55",
          7359 => x"08",
          7360 => x"80",
          7361 => x"70",
          7362 => x"56",
          7363 => x"89",
          7364 => x"94",
          7365 => x"b2",
          7366 => x"05",
          7367 => x"2a",
          7368 => x"51",
          7369 => x"80",
          7370 => x"76",
          7371 => x"52",
          7372 => x"3f",
          7373 => x"08",
          7374 => x"8e",
          7375 => x"c8",
          7376 => x"09",
          7377 => x"38",
          7378 => x"82",
          7379 => x"93",
          7380 => x"e4",
          7381 => x"6f",
          7382 => x"7a",
          7383 => x"9e",
          7384 => x"05",
          7385 => x"51",
          7386 => x"82",
          7387 => x"57",
          7388 => x"08",
          7389 => x"7b",
          7390 => x"94",
          7391 => x"55",
          7392 => x"73",
          7393 => x"ed",
          7394 => x"93",
          7395 => x"55",
          7396 => x"82",
          7397 => x"57",
          7398 => x"08",
          7399 => x"68",
          7400 => x"c9",
          7401 => x"b5",
          7402 => x"82",
          7403 => x"82",
          7404 => x"52",
          7405 => x"a3",
          7406 => x"c8",
          7407 => x"52",
          7408 => x"b8",
          7409 => x"c8",
          7410 => x"b5",
          7411 => x"a2",
          7412 => x"74",
          7413 => x"3f",
          7414 => x"08",
          7415 => x"c8",
          7416 => x"69",
          7417 => x"d9",
          7418 => x"82",
          7419 => x"2e",
          7420 => x"52",
          7421 => x"cf",
          7422 => x"c8",
          7423 => x"b5",
          7424 => x"2e",
          7425 => x"84",
          7426 => x"06",
          7427 => x"57",
          7428 => x"76",
          7429 => x"9e",
          7430 => x"05",
          7431 => x"dc",
          7432 => x"90",
          7433 => x"81",
          7434 => x"56",
          7435 => x"80",
          7436 => x"02",
          7437 => x"81",
          7438 => x"70",
          7439 => x"56",
          7440 => x"81",
          7441 => x"78",
          7442 => x"38",
          7443 => x"99",
          7444 => x"81",
          7445 => x"18",
          7446 => x"18",
          7447 => x"58",
          7448 => x"33",
          7449 => x"ee",
          7450 => x"6f",
          7451 => x"af",
          7452 => x"8d",
          7453 => x"2e",
          7454 => x"8a",
          7455 => x"6f",
          7456 => x"af",
          7457 => x"0b",
          7458 => x"33",
          7459 => x"82",
          7460 => x"70",
          7461 => x"52",
          7462 => x"56",
          7463 => x"8d",
          7464 => x"70",
          7465 => x"51",
          7466 => x"f5",
          7467 => x"54",
          7468 => x"a7",
          7469 => x"74",
          7470 => x"38",
          7471 => x"73",
          7472 => x"81",
          7473 => x"81",
          7474 => x"39",
          7475 => x"81",
          7476 => x"74",
          7477 => x"81",
          7478 => x"91",
          7479 => x"6e",
          7480 => x"59",
          7481 => x"7a",
          7482 => x"5c",
          7483 => x"26",
          7484 => x"7a",
          7485 => x"b5",
          7486 => x"3d",
          7487 => x"3d",
          7488 => x"8d",
          7489 => x"54",
          7490 => x"55",
          7491 => x"82",
          7492 => x"53",
          7493 => x"08",
          7494 => x"91",
          7495 => x"72",
          7496 => x"8c",
          7497 => x"73",
          7498 => x"38",
          7499 => x"70",
          7500 => x"81",
          7501 => x"57",
          7502 => x"73",
          7503 => x"08",
          7504 => x"94",
          7505 => x"75",
          7506 => x"97",
          7507 => x"11",
          7508 => x"2b",
          7509 => x"73",
          7510 => x"38",
          7511 => x"16",
          7512 => x"a1",
          7513 => x"c8",
          7514 => x"78",
          7515 => x"55",
          7516 => x"91",
          7517 => x"c8",
          7518 => x"96",
          7519 => x"70",
          7520 => x"94",
          7521 => x"71",
          7522 => x"08",
          7523 => x"53",
          7524 => x"15",
          7525 => x"a6",
          7526 => x"74",
          7527 => x"3f",
          7528 => x"08",
          7529 => x"c8",
          7530 => x"81",
          7531 => x"b5",
          7532 => x"2e",
          7533 => x"82",
          7534 => x"88",
          7535 => x"98",
          7536 => x"80",
          7537 => x"38",
          7538 => x"80",
          7539 => x"77",
          7540 => x"08",
          7541 => x"0c",
          7542 => x"70",
          7543 => x"81",
          7544 => x"5a",
          7545 => x"2e",
          7546 => x"52",
          7547 => x"f9",
          7548 => x"c8",
          7549 => x"b5",
          7550 => x"38",
          7551 => x"08",
          7552 => x"73",
          7553 => x"c7",
          7554 => x"b5",
          7555 => x"73",
          7556 => x"38",
          7557 => x"af",
          7558 => x"73",
          7559 => x"27",
          7560 => x"98",
          7561 => x"a0",
          7562 => x"08",
          7563 => x"0c",
          7564 => x"06",
          7565 => x"2e",
          7566 => x"52",
          7567 => x"a3",
          7568 => x"c8",
          7569 => x"82",
          7570 => x"34",
          7571 => x"c4",
          7572 => x"91",
          7573 => x"53",
          7574 => x"89",
          7575 => x"c8",
          7576 => x"94",
          7577 => x"8c",
          7578 => x"27",
          7579 => x"8c",
          7580 => x"15",
          7581 => x"07",
          7582 => x"16",
          7583 => x"ff",
          7584 => x"80",
          7585 => x"77",
          7586 => x"2e",
          7587 => x"9c",
          7588 => x"53",
          7589 => x"c8",
          7590 => x"0d",
          7591 => x"0d",
          7592 => x"54",
          7593 => x"81",
          7594 => x"53",
          7595 => x"05",
          7596 => x"84",
          7597 => x"e7",
          7598 => x"c8",
          7599 => x"b5",
          7600 => x"ea",
          7601 => x"0c",
          7602 => x"51",
          7603 => x"82",
          7604 => x"55",
          7605 => x"08",
          7606 => x"ab",
          7607 => x"98",
          7608 => x"80",
          7609 => x"38",
          7610 => x"70",
          7611 => x"81",
          7612 => x"57",
          7613 => x"ad",
          7614 => x"08",
          7615 => x"d3",
          7616 => x"b5",
          7617 => x"17",
          7618 => x"86",
          7619 => x"17",
          7620 => x"75",
          7621 => x"3f",
          7622 => x"08",
          7623 => x"2e",
          7624 => x"85",
          7625 => x"86",
          7626 => x"2e",
          7627 => x"76",
          7628 => x"73",
          7629 => x"0c",
          7630 => x"04",
          7631 => x"76",
          7632 => x"05",
          7633 => x"53",
          7634 => x"82",
          7635 => x"87",
          7636 => x"c8",
          7637 => x"86",
          7638 => x"fb",
          7639 => x"79",
          7640 => x"05",
          7641 => x"56",
          7642 => x"3f",
          7643 => x"08",
          7644 => x"c8",
          7645 => x"38",
          7646 => x"82",
          7647 => x"52",
          7648 => x"f8",
          7649 => x"c8",
          7650 => x"ca",
          7651 => x"c8",
          7652 => x"51",
          7653 => x"82",
          7654 => x"53",
          7655 => x"08",
          7656 => x"81",
          7657 => x"80",
          7658 => x"82",
          7659 => x"a6",
          7660 => x"73",
          7661 => x"3f",
          7662 => x"51",
          7663 => x"82",
          7664 => x"84",
          7665 => x"70",
          7666 => x"2c",
          7667 => x"c8",
          7668 => x"51",
          7669 => x"82",
          7670 => x"87",
          7671 => x"ee",
          7672 => x"57",
          7673 => x"3d",
          7674 => x"3d",
          7675 => x"af",
          7676 => x"c8",
          7677 => x"b5",
          7678 => x"38",
          7679 => x"51",
          7680 => x"82",
          7681 => x"55",
          7682 => x"08",
          7683 => x"80",
          7684 => x"70",
          7685 => x"58",
          7686 => x"85",
          7687 => x"8d",
          7688 => x"2e",
          7689 => x"52",
          7690 => x"be",
          7691 => x"b5",
          7692 => x"3d",
          7693 => x"3d",
          7694 => x"55",
          7695 => x"92",
          7696 => x"52",
          7697 => x"de",
          7698 => x"b5",
          7699 => x"82",
          7700 => x"82",
          7701 => x"74",
          7702 => x"98",
          7703 => x"11",
          7704 => x"59",
          7705 => x"75",
          7706 => x"38",
          7707 => x"81",
          7708 => x"5b",
          7709 => x"82",
          7710 => x"39",
          7711 => x"08",
          7712 => x"59",
          7713 => x"09",
          7714 => x"38",
          7715 => x"57",
          7716 => x"3d",
          7717 => x"c1",
          7718 => x"b5",
          7719 => x"2e",
          7720 => x"b5",
          7721 => x"2e",
          7722 => x"b5",
          7723 => x"70",
          7724 => x"08",
          7725 => x"7a",
          7726 => x"7f",
          7727 => x"54",
          7728 => x"77",
          7729 => x"80",
          7730 => x"15",
          7731 => x"c8",
          7732 => x"75",
          7733 => x"52",
          7734 => x"52",
          7735 => x"8d",
          7736 => x"c8",
          7737 => x"b5",
          7738 => x"d6",
          7739 => x"33",
          7740 => x"1a",
          7741 => x"54",
          7742 => x"09",
          7743 => x"38",
          7744 => x"ff",
          7745 => x"82",
          7746 => x"83",
          7747 => x"70",
          7748 => x"25",
          7749 => x"59",
          7750 => x"9b",
          7751 => x"51",
          7752 => x"3f",
          7753 => x"08",
          7754 => x"70",
          7755 => x"25",
          7756 => x"59",
          7757 => x"75",
          7758 => x"7a",
          7759 => x"ff",
          7760 => x"7c",
          7761 => x"90",
          7762 => x"11",
          7763 => x"56",
          7764 => x"15",
          7765 => x"b5",
          7766 => x"3d",
          7767 => x"3d",
          7768 => x"3d",
          7769 => x"70",
          7770 => x"dd",
          7771 => x"c8",
          7772 => x"b5",
          7773 => x"a8",
          7774 => x"33",
          7775 => x"a0",
          7776 => x"33",
          7777 => x"70",
          7778 => x"55",
          7779 => x"73",
          7780 => x"8e",
          7781 => x"08",
          7782 => x"18",
          7783 => x"80",
          7784 => x"38",
          7785 => x"08",
          7786 => x"08",
          7787 => x"c4",
          7788 => x"b5",
          7789 => x"88",
          7790 => x"80",
          7791 => x"17",
          7792 => x"51",
          7793 => x"3f",
          7794 => x"08",
          7795 => x"81",
          7796 => x"81",
          7797 => x"c8",
          7798 => x"09",
          7799 => x"38",
          7800 => x"39",
          7801 => x"77",
          7802 => x"c8",
          7803 => x"08",
          7804 => x"98",
          7805 => x"82",
          7806 => x"52",
          7807 => x"bd",
          7808 => x"c8",
          7809 => x"17",
          7810 => x"0c",
          7811 => x"80",
          7812 => x"73",
          7813 => x"75",
          7814 => x"38",
          7815 => x"34",
          7816 => x"82",
          7817 => x"89",
          7818 => x"e2",
          7819 => x"53",
          7820 => x"a4",
          7821 => x"3d",
          7822 => x"3f",
          7823 => x"08",
          7824 => x"c8",
          7825 => x"38",
          7826 => x"3d",
          7827 => x"3d",
          7828 => x"d1",
          7829 => x"b5",
          7830 => x"82",
          7831 => x"81",
          7832 => x"80",
          7833 => x"70",
          7834 => x"81",
          7835 => x"56",
          7836 => x"81",
          7837 => x"98",
          7838 => x"74",
          7839 => x"38",
          7840 => x"05",
          7841 => x"06",
          7842 => x"55",
          7843 => x"38",
          7844 => x"51",
          7845 => x"82",
          7846 => x"74",
          7847 => x"81",
          7848 => x"56",
          7849 => x"80",
          7850 => x"54",
          7851 => x"08",
          7852 => x"2e",
          7853 => x"73",
          7854 => x"c8",
          7855 => x"52",
          7856 => x"52",
          7857 => x"3f",
          7858 => x"08",
          7859 => x"c8",
          7860 => x"38",
          7861 => x"08",
          7862 => x"cc",
          7863 => x"b5",
          7864 => x"82",
          7865 => x"86",
          7866 => x"80",
          7867 => x"b5",
          7868 => x"2e",
          7869 => x"b5",
          7870 => x"c0",
          7871 => x"ce",
          7872 => x"b5",
          7873 => x"b5",
          7874 => x"70",
          7875 => x"08",
          7876 => x"51",
          7877 => x"80",
          7878 => x"73",
          7879 => x"38",
          7880 => x"52",
          7881 => x"95",
          7882 => x"c8",
          7883 => x"8c",
          7884 => x"ff",
          7885 => x"82",
          7886 => x"55",
          7887 => x"c8",
          7888 => x"0d",
          7889 => x"0d",
          7890 => x"3d",
          7891 => x"9a",
          7892 => x"cb",
          7893 => x"c8",
          7894 => x"b5",
          7895 => x"b0",
          7896 => x"69",
          7897 => x"70",
          7898 => x"97",
          7899 => x"c8",
          7900 => x"b5",
          7901 => x"38",
          7902 => x"94",
          7903 => x"c8",
          7904 => x"09",
          7905 => x"88",
          7906 => x"df",
          7907 => x"85",
          7908 => x"51",
          7909 => x"74",
          7910 => x"78",
          7911 => x"8a",
          7912 => x"57",
          7913 => x"82",
          7914 => x"75",
          7915 => x"b5",
          7916 => x"38",
          7917 => x"b5",
          7918 => x"2e",
          7919 => x"83",
          7920 => x"82",
          7921 => x"ff",
          7922 => x"06",
          7923 => x"54",
          7924 => x"73",
          7925 => x"82",
          7926 => x"52",
          7927 => x"a4",
          7928 => x"c8",
          7929 => x"b5",
          7930 => x"9a",
          7931 => x"a0",
          7932 => x"51",
          7933 => x"3f",
          7934 => x"0b",
          7935 => x"78",
          7936 => x"bf",
          7937 => x"88",
          7938 => x"80",
          7939 => x"ff",
          7940 => x"75",
          7941 => x"11",
          7942 => x"f8",
          7943 => x"78",
          7944 => x"80",
          7945 => x"ff",
          7946 => x"78",
          7947 => x"80",
          7948 => x"7f",
          7949 => x"d4",
          7950 => x"c9",
          7951 => x"54",
          7952 => x"15",
          7953 => x"cb",
          7954 => x"b5",
          7955 => x"82",
          7956 => x"b2",
          7957 => x"b2",
          7958 => x"96",
          7959 => x"b5",
          7960 => x"53",
          7961 => x"51",
          7962 => x"64",
          7963 => x"8b",
          7964 => x"54",
          7965 => x"15",
          7966 => x"ff",
          7967 => x"82",
          7968 => x"54",
          7969 => x"53",
          7970 => x"51",
          7971 => x"3f",
          7972 => x"c8",
          7973 => x"0d",
          7974 => x"0d",
          7975 => x"05",
          7976 => x"3f",
          7977 => x"3d",
          7978 => x"52",
          7979 => x"d5",
          7980 => x"b5",
          7981 => x"82",
          7982 => x"82",
          7983 => x"4d",
          7984 => x"52",
          7985 => x"52",
          7986 => x"3f",
          7987 => x"08",
          7988 => x"c8",
          7989 => x"38",
          7990 => x"05",
          7991 => x"06",
          7992 => x"73",
          7993 => x"a0",
          7994 => x"08",
          7995 => x"ff",
          7996 => x"ff",
          7997 => x"ac",
          7998 => x"92",
          7999 => x"54",
          8000 => x"3f",
          8001 => x"52",
          8002 => x"f7",
          8003 => x"c8",
          8004 => x"b5",
          8005 => x"38",
          8006 => x"09",
          8007 => x"38",
          8008 => x"08",
          8009 => x"88",
          8010 => x"39",
          8011 => x"08",
          8012 => x"81",
          8013 => x"38",
          8014 => x"b1",
          8015 => x"c8",
          8016 => x"b5",
          8017 => x"c8",
          8018 => x"93",
          8019 => x"ff",
          8020 => x"8d",
          8021 => x"b4",
          8022 => x"af",
          8023 => x"17",
          8024 => x"33",
          8025 => x"70",
          8026 => x"55",
          8027 => x"38",
          8028 => x"54",
          8029 => x"34",
          8030 => x"0b",
          8031 => x"8b",
          8032 => x"84",
          8033 => x"06",
          8034 => x"73",
          8035 => x"e5",
          8036 => x"2e",
          8037 => x"75",
          8038 => x"c6",
          8039 => x"b5",
          8040 => x"78",
          8041 => x"bb",
          8042 => x"82",
          8043 => x"80",
          8044 => x"38",
          8045 => x"08",
          8046 => x"ff",
          8047 => x"82",
          8048 => x"79",
          8049 => x"58",
          8050 => x"b5",
          8051 => x"c0",
          8052 => x"33",
          8053 => x"2e",
          8054 => x"99",
          8055 => x"75",
          8056 => x"c6",
          8057 => x"54",
          8058 => x"15",
          8059 => x"82",
          8060 => x"9c",
          8061 => x"c8",
          8062 => x"b5",
          8063 => x"82",
          8064 => x"8c",
          8065 => x"ff",
          8066 => x"82",
          8067 => x"55",
          8068 => x"c8",
          8069 => x"0d",
          8070 => x"0d",
          8071 => x"05",
          8072 => x"05",
          8073 => x"33",
          8074 => x"53",
          8075 => x"05",
          8076 => x"51",
          8077 => x"82",
          8078 => x"55",
          8079 => x"08",
          8080 => x"78",
          8081 => x"95",
          8082 => x"51",
          8083 => x"82",
          8084 => x"55",
          8085 => x"08",
          8086 => x"80",
          8087 => x"81",
          8088 => x"86",
          8089 => x"38",
          8090 => x"61",
          8091 => x"12",
          8092 => x"7a",
          8093 => x"51",
          8094 => x"74",
          8095 => x"78",
          8096 => x"83",
          8097 => x"51",
          8098 => x"3f",
          8099 => x"08",
          8100 => x"b5",
          8101 => x"3d",
          8102 => x"3d",
          8103 => x"82",
          8104 => x"d0",
          8105 => x"3d",
          8106 => x"3f",
          8107 => x"08",
          8108 => x"c8",
          8109 => x"38",
          8110 => x"52",
          8111 => x"05",
          8112 => x"3f",
          8113 => x"08",
          8114 => x"c8",
          8115 => x"02",
          8116 => x"33",
          8117 => x"54",
          8118 => x"a6",
          8119 => x"22",
          8120 => x"71",
          8121 => x"53",
          8122 => x"51",
          8123 => x"3f",
          8124 => x"0b",
          8125 => x"76",
          8126 => x"b8",
          8127 => x"c8",
          8128 => x"82",
          8129 => x"93",
          8130 => x"ea",
          8131 => x"6b",
          8132 => x"53",
          8133 => x"05",
          8134 => x"51",
          8135 => x"82",
          8136 => x"82",
          8137 => x"30",
          8138 => x"c8",
          8139 => x"25",
          8140 => x"79",
          8141 => x"85",
          8142 => x"75",
          8143 => x"73",
          8144 => x"f9",
          8145 => x"80",
          8146 => x"8d",
          8147 => x"54",
          8148 => x"3f",
          8149 => x"08",
          8150 => x"c8",
          8151 => x"38",
          8152 => x"51",
          8153 => x"82",
          8154 => x"57",
          8155 => x"08",
          8156 => x"b5",
          8157 => x"b5",
          8158 => x"5b",
          8159 => x"18",
          8160 => x"18",
          8161 => x"74",
          8162 => x"81",
          8163 => x"78",
          8164 => x"8b",
          8165 => x"54",
          8166 => x"75",
          8167 => x"38",
          8168 => x"1b",
          8169 => x"55",
          8170 => x"2e",
          8171 => x"39",
          8172 => x"09",
          8173 => x"38",
          8174 => x"80",
          8175 => x"70",
          8176 => x"25",
          8177 => x"80",
          8178 => x"38",
          8179 => x"bc",
          8180 => x"11",
          8181 => x"ff",
          8182 => x"82",
          8183 => x"57",
          8184 => x"08",
          8185 => x"70",
          8186 => x"80",
          8187 => x"83",
          8188 => x"80",
          8189 => x"84",
          8190 => x"a7",
          8191 => x"b4",
          8192 => x"ad",
          8193 => x"b5",
          8194 => x"0c",
          8195 => x"c8",
          8196 => x"0d",
          8197 => x"0d",
          8198 => x"3d",
          8199 => x"52",
          8200 => x"ce",
          8201 => x"b5",
          8202 => x"b5",
          8203 => x"54",
          8204 => x"08",
          8205 => x"8b",
          8206 => x"8b",
          8207 => x"59",
          8208 => x"3f",
          8209 => x"33",
          8210 => x"06",
          8211 => x"57",
          8212 => x"81",
          8213 => x"58",
          8214 => x"06",
          8215 => x"4e",
          8216 => x"ff",
          8217 => x"82",
          8218 => x"80",
          8219 => x"6c",
          8220 => x"53",
          8221 => x"ae",
          8222 => x"b5",
          8223 => x"2e",
          8224 => x"88",
          8225 => x"6d",
          8226 => x"55",
          8227 => x"b5",
          8228 => x"ff",
          8229 => x"83",
          8230 => x"51",
          8231 => x"26",
          8232 => x"15",
          8233 => x"ff",
          8234 => x"80",
          8235 => x"87",
          8236 => x"90",
          8237 => x"74",
          8238 => x"38",
          8239 => x"b0",
          8240 => x"ae",
          8241 => x"b5",
          8242 => x"38",
          8243 => x"27",
          8244 => x"89",
          8245 => x"8b",
          8246 => x"27",
          8247 => x"55",
          8248 => x"81",
          8249 => x"8f",
          8250 => x"2a",
          8251 => x"70",
          8252 => x"34",
          8253 => x"74",
          8254 => x"05",
          8255 => x"17",
          8256 => x"70",
          8257 => x"52",
          8258 => x"73",
          8259 => x"c8",
          8260 => x"33",
          8261 => x"73",
          8262 => x"81",
          8263 => x"80",
          8264 => x"02",
          8265 => x"76",
          8266 => x"51",
          8267 => x"2e",
          8268 => x"87",
          8269 => x"57",
          8270 => x"79",
          8271 => x"80",
          8272 => x"70",
          8273 => x"ba",
          8274 => x"b5",
          8275 => x"82",
          8276 => x"80",
          8277 => x"52",
          8278 => x"bf",
          8279 => x"b5",
          8280 => x"82",
          8281 => x"8d",
          8282 => x"c4",
          8283 => x"e5",
          8284 => x"c6",
          8285 => x"c8",
          8286 => x"09",
          8287 => x"cc",
          8288 => x"76",
          8289 => x"c4",
          8290 => x"74",
          8291 => x"b0",
          8292 => x"c8",
          8293 => x"b5",
          8294 => x"38",
          8295 => x"b5",
          8296 => x"67",
          8297 => x"db",
          8298 => x"88",
          8299 => x"34",
          8300 => x"52",
          8301 => x"ab",
          8302 => x"54",
          8303 => x"15",
          8304 => x"ff",
          8305 => x"82",
          8306 => x"54",
          8307 => x"82",
          8308 => x"9c",
          8309 => x"f2",
          8310 => x"62",
          8311 => x"80",
          8312 => x"93",
          8313 => x"55",
          8314 => x"5e",
          8315 => x"3f",
          8316 => x"08",
          8317 => x"c8",
          8318 => x"38",
          8319 => x"58",
          8320 => x"38",
          8321 => x"97",
          8322 => x"08",
          8323 => x"38",
          8324 => x"70",
          8325 => x"81",
          8326 => x"55",
          8327 => x"87",
          8328 => x"39",
          8329 => x"90",
          8330 => x"82",
          8331 => x"8a",
          8332 => x"89",
          8333 => x"7f",
          8334 => x"56",
          8335 => x"3f",
          8336 => x"06",
          8337 => x"72",
          8338 => x"82",
          8339 => x"05",
          8340 => x"7c",
          8341 => x"55",
          8342 => x"27",
          8343 => x"16",
          8344 => x"83",
          8345 => x"76",
          8346 => x"80",
          8347 => x"79",
          8348 => x"99",
          8349 => x"7f",
          8350 => x"14",
          8351 => x"83",
          8352 => x"82",
          8353 => x"81",
          8354 => x"38",
          8355 => x"08",
          8356 => x"95",
          8357 => x"c8",
          8358 => x"81",
          8359 => x"7b",
          8360 => x"06",
          8361 => x"39",
          8362 => x"56",
          8363 => x"09",
          8364 => x"b9",
          8365 => x"80",
          8366 => x"80",
          8367 => x"78",
          8368 => x"7a",
          8369 => x"38",
          8370 => x"73",
          8371 => x"81",
          8372 => x"ff",
          8373 => x"74",
          8374 => x"ff",
          8375 => x"82",
          8376 => x"58",
          8377 => x"08",
          8378 => x"74",
          8379 => x"16",
          8380 => x"73",
          8381 => x"39",
          8382 => x"7e",
          8383 => x"0c",
          8384 => x"2e",
          8385 => x"88",
          8386 => x"8c",
          8387 => x"1a",
          8388 => x"07",
          8389 => x"1b",
          8390 => x"08",
          8391 => x"16",
          8392 => x"75",
          8393 => x"38",
          8394 => x"90",
          8395 => x"15",
          8396 => x"54",
          8397 => x"34",
          8398 => x"82",
          8399 => x"90",
          8400 => x"e9",
          8401 => x"6d",
          8402 => x"80",
          8403 => x"9d",
          8404 => x"5c",
          8405 => x"3f",
          8406 => x"0b",
          8407 => x"08",
          8408 => x"38",
          8409 => x"08",
          8410 => x"cd",
          8411 => x"08",
          8412 => x"80",
          8413 => x"80",
          8414 => x"b5",
          8415 => x"ff",
          8416 => x"52",
          8417 => x"a0",
          8418 => x"b5",
          8419 => x"ff",
          8420 => x"06",
          8421 => x"56",
          8422 => x"38",
          8423 => x"70",
          8424 => x"55",
          8425 => x"8b",
          8426 => x"3d",
          8427 => x"83",
          8428 => x"ff",
          8429 => x"82",
          8430 => x"99",
          8431 => x"74",
          8432 => x"38",
          8433 => x"80",
          8434 => x"ff",
          8435 => x"55",
          8436 => x"83",
          8437 => x"78",
          8438 => x"38",
          8439 => x"26",
          8440 => x"81",
          8441 => x"8b",
          8442 => x"79",
          8443 => x"80",
          8444 => x"93",
          8445 => x"39",
          8446 => x"6e",
          8447 => x"89",
          8448 => x"48",
          8449 => x"83",
          8450 => x"61",
          8451 => x"25",
          8452 => x"55",
          8453 => x"8a",
          8454 => x"3d",
          8455 => x"81",
          8456 => x"ff",
          8457 => x"81",
          8458 => x"c8",
          8459 => x"38",
          8460 => x"70",
          8461 => x"b5",
          8462 => x"56",
          8463 => x"38",
          8464 => x"55",
          8465 => x"75",
          8466 => x"38",
          8467 => x"70",
          8468 => x"ff",
          8469 => x"83",
          8470 => x"78",
          8471 => x"89",
          8472 => x"81",
          8473 => x"06",
          8474 => x"80",
          8475 => x"77",
          8476 => x"74",
          8477 => x"8d",
          8478 => x"06",
          8479 => x"2e",
          8480 => x"77",
          8481 => x"93",
          8482 => x"74",
          8483 => x"cb",
          8484 => x"7d",
          8485 => x"81",
          8486 => x"38",
          8487 => x"66",
          8488 => x"81",
          8489 => x"b4",
          8490 => x"74",
          8491 => x"38",
          8492 => x"98",
          8493 => x"b4",
          8494 => x"82",
          8495 => x"57",
          8496 => x"80",
          8497 => x"76",
          8498 => x"38",
          8499 => x"51",
          8500 => x"3f",
          8501 => x"08",
          8502 => x"87",
          8503 => x"2a",
          8504 => x"5c",
          8505 => x"b5",
          8506 => x"80",
          8507 => x"44",
          8508 => x"0a",
          8509 => x"ec",
          8510 => x"39",
          8511 => x"66",
          8512 => x"81",
          8513 => x"a4",
          8514 => x"74",
          8515 => x"38",
          8516 => x"98",
          8517 => x"a4",
          8518 => x"82",
          8519 => x"57",
          8520 => x"80",
          8521 => x"76",
          8522 => x"38",
          8523 => x"51",
          8524 => x"3f",
          8525 => x"08",
          8526 => x"57",
          8527 => x"08",
          8528 => x"96",
          8529 => x"82",
          8530 => x"10",
          8531 => x"08",
          8532 => x"72",
          8533 => x"59",
          8534 => x"ff",
          8535 => x"5d",
          8536 => x"44",
          8537 => x"11",
          8538 => x"70",
          8539 => x"71",
          8540 => x"06",
          8541 => x"52",
          8542 => x"40",
          8543 => x"09",
          8544 => x"38",
          8545 => x"18",
          8546 => x"39",
          8547 => x"79",
          8548 => x"70",
          8549 => x"58",
          8550 => x"76",
          8551 => x"38",
          8552 => x"7d",
          8553 => x"70",
          8554 => x"55",
          8555 => x"3f",
          8556 => x"08",
          8557 => x"2e",
          8558 => x"9b",
          8559 => x"c8",
          8560 => x"f5",
          8561 => x"38",
          8562 => x"38",
          8563 => x"59",
          8564 => x"38",
          8565 => x"7d",
          8566 => x"81",
          8567 => x"38",
          8568 => x"0b",
          8569 => x"08",
          8570 => x"78",
          8571 => x"1a",
          8572 => x"c0",
          8573 => x"74",
          8574 => x"39",
          8575 => x"55",
          8576 => x"8f",
          8577 => x"fd",
          8578 => x"b5",
          8579 => x"f5",
          8580 => x"78",
          8581 => x"79",
          8582 => x"80",
          8583 => x"f1",
          8584 => x"39",
          8585 => x"81",
          8586 => x"06",
          8587 => x"55",
          8588 => x"27",
          8589 => x"81",
          8590 => x"56",
          8591 => x"38",
          8592 => x"80",
          8593 => x"ff",
          8594 => x"8b",
          8595 => x"cc",
          8596 => x"ff",
          8597 => x"84",
          8598 => x"1b",
          8599 => x"b3",
          8600 => x"1c",
          8601 => x"ff",
          8602 => x"8e",
          8603 => x"a1",
          8604 => x"0b",
          8605 => x"7d",
          8606 => x"30",
          8607 => x"84",
          8608 => x"51",
          8609 => x"51",
          8610 => x"3f",
          8611 => x"83",
          8612 => x"90",
          8613 => x"ff",
          8614 => x"93",
          8615 => x"a0",
          8616 => x"39",
          8617 => x"1b",
          8618 => x"85",
          8619 => x"95",
          8620 => x"52",
          8621 => x"ff",
          8622 => x"81",
          8623 => x"1b",
          8624 => x"cf",
          8625 => x"9c",
          8626 => x"a0",
          8627 => x"83",
          8628 => x"06",
          8629 => x"82",
          8630 => x"52",
          8631 => x"51",
          8632 => x"3f",
          8633 => x"1b",
          8634 => x"c5",
          8635 => x"ac",
          8636 => x"a0",
          8637 => x"52",
          8638 => x"ff",
          8639 => x"86",
          8640 => x"51",
          8641 => x"3f",
          8642 => x"80",
          8643 => x"a9",
          8644 => x"1c",
          8645 => x"82",
          8646 => x"80",
          8647 => x"ae",
          8648 => x"b2",
          8649 => x"1b",
          8650 => x"85",
          8651 => x"ff",
          8652 => x"96",
          8653 => x"9f",
          8654 => x"80",
          8655 => x"34",
          8656 => x"1c",
          8657 => x"82",
          8658 => x"ab",
          8659 => x"a0",
          8660 => x"d4",
          8661 => x"fe",
          8662 => x"59",
          8663 => x"3f",
          8664 => x"53",
          8665 => x"51",
          8666 => x"3f",
          8667 => x"b5",
          8668 => x"e7",
          8669 => x"2e",
          8670 => x"80",
          8671 => x"54",
          8672 => x"53",
          8673 => x"51",
          8674 => x"3f",
          8675 => x"80",
          8676 => x"ff",
          8677 => x"84",
          8678 => x"d2",
          8679 => x"ff",
          8680 => x"86",
          8681 => x"f2",
          8682 => x"1b",
          8683 => x"81",
          8684 => x"52",
          8685 => x"51",
          8686 => x"3f",
          8687 => x"ec",
          8688 => x"9e",
          8689 => x"d4",
          8690 => x"51",
          8691 => x"3f",
          8692 => x"87",
          8693 => x"52",
          8694 => x"9a",
          8695 => x"54",
          8696 => x"7a",
          8697 => x"ff",
          8698 => x"65",
          8699 => x"7a",
          8700 => x"8f",
          8701 => x"80",
          8702 => x"2e",
          8703 => x"9a",
          8704 => x"7a",
          8705 => x"a9",
          8706 => x"84",
          8707 => x"9e",
          8708 => x"0a",
          8709 => x"51",
          8710 => x"ff",
          8711 => x"7d",
          8712 => x"38",
          8713 => x"52",
          8714 => x"9e",
          8715 => x"55",
          8716 => x"62",
          8717 => x"74",
          8718 => x"75",
          8719 => x"7e",
          8720 => x"fe",
          8721 => x"c8",
          8722 => x"38",
          8723 => x"82",
          8724 => x"52",
          8725 => x"9e",
          8726 => x"16",
          8727 => x"56",
          8728 => x"38",
          8729 => x"77",
          8730 => x"8d",
          8731 => x"7d",
          8732 => x"38",
          8733 => x"57",
          8734 => x"83",
          8735 => x"76",
          8736 => x"7a",
          8737 => x"ff",
          8738 => x"82",
          8739 => x"81",
          8740 => x"16",
          8741 => x"56",
          8742 => x"38",
          8743 => x"83",
          8744 => x"86",
          8745 => x"ff",
          8746 => x"38",
          8747 => x"82",
          8748 => x"81",
          8749 => x"06",
          8750 => x"fe",
          8751 => x"53",
          8752 => x"51",
          8753 => x"3f",
          8754 => x"52",
          8755 => x"9c",
          8756 => x"be",
          8757 => x"75",
          8758 => x"81",
          8759 => x"0b",
          8760 => x"77",
          8761 => x"75",
          8762 => x"60",
          8763 => x"80",
          8764 => x"75",
          8765 => x"8d",
          8766 => x"85",
          8767 => x"b5",
          8768 => x"2a",
          8769 => x"75",
          8770 => x"82",
          8771 => x"87",
          8772 => x"52",
          8773 => x"51",
          8774 => x"3f",
          8775 => x"ca",
          8776 => x"9c",
          8777 => x"54",
          8778 => x"52",
          8779 => x"98",
          8780 => x"56",
          8781 => x"08",
          8782 => x"53",
          8783 => x"51",
          8784 => x"3f",
          8785 => x"b5",
          8786 => x"38",
          8787 => x"56",
          8788 => x"56",
          8789 => x"b5",
          8790 => x"75",
          8791 => x"0c",
          8792 => x"04",
          8793 => x"7d",
          8794 => x"80",
          8795 => x"05",
          8796 => x"76",
          8797 => x"38",
          8798 => x"11",
          8799 => x"53",
          8800 => x"79",
          8801 => x"3f",
          8802 => x"09",
          8803 => x"38",
          8804 => x"55",
          8805 => x"db",
          8806 => x"70",
          8807 => x"34",
          8808 => x"74",
          8809 => x"81",
          8810 => x"80",
          8811 => x"55",
          8812 => x"76",
          8813 => x"b5",
          8814 => x"3d",
          8815 => x"3d",
          8816 => x"84",
          8817 => x"33",
          8818 => x"8a",
          8819 => x"06",
          8820 => x"52",
          8821 => x"3f",
          8822 => x"56",
          8823 => x"be",
          8824 => x"08",
          8825 => x"05",
          8826 => x"75",
          8827 => x"56",
          8828 => x"a1",
          8829 => x"fc",
          8830 => x"53",
          8831 => x"76",
          8832 => x"dc",
          8833 => x"32",
          8834 => x"72",
          8835 => x"70",
          8836 => x"56",
          8837 => x"18",
          8838 => x"88",
          8839 => x"3d",
          8840 => x"3d",
          8841 => x"11",
          8842 => x"80",
          8843 => x"38",
          8844 => x"05",
          8845 => x"8c",
          8846 => x"08",
          8847 => x"3f",
          8848 => x"08",
          8849 => x"16",
          8850 => x"09",
          8851 => x"38",
          8852 => x"55",
          8853 => x"55",
          8854 => x"c8",
          8855 => x"0d",
          8856 => x"0d",
          8857 => x"cc",
          8858 => x"73",
          8859 => x"93",
          8860 => x"0c",
          8861 => x"04",
          8862 => x"02",
          8863 => x"33",
          8864 => x"3d",
          8865 => x"54",
          8866 => x"52",
          8867 => x"ae",
          8868 => x"ff",
          8869 => x"3d",
          8870 => x"ff",
          8871 => x"00",
          8872 => x"ff",
          8873 => x"ff",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"69",
          9011 => x"00",
          9012 => x"69",
          9013 => x"6c",
          9014 => x"69",
          9015 => x"00",
          9016 => x"6c",
          9017 => x"00",
          9018 => x"65",
          9019 => x"00",
          9020 => x"63",
          9021 => x"72",
          9022 => x"63",
          9023 => x"00",
          9024 => x"64",
          9025 => x"00",
          9026 => x"64",
          9027 => x"00",
          9028 => x"65",
          9029 => x"65",
          9030 => x"65",
          9031 => x"69",
          9032 => x"69",
          9033 => x"66",
          9034 => x"66",
          9035 => x"61",
          9036 => x"00",
          9037 => x"6d",
          9038 => x"65",
          9039 => x"72",
          9040 => x"65",
          9041 => x"00",
          9042 => x"6e",
          9043 => x"00",
          9044 => x"65",
          9045 => x"00",
          9046 => x"62",
          9047 => x"63",
          9048 => x"62",
          9049 => x"63",
          9050 => x"69",
          9051 => x"00",
          9052 => x"64",
          9053 => x"69",
          9054 => x"45",
          9055 => x"72",
          9056 => x"6e",
          9057 => x"6e",
          9058 => x"65",
          9059 => x"72",
          9060 => x"69",
          9061 => x"6e",
          9062 => x"72",
          9063 => x"79",
          9064 => x"6f",
          9065 => x"6c",
          9066 => x"6f",
          9067 => x"2e",
          9068 => x"6f",
          9069 => x"74",
          9070 => x"6f",
          9071 => x"2e",
          9072 => x"6e",
          9073 => x"69",
          9074 => x"69",
          9075 => x"61",
          9076 => x"00",
          9077 => x"63",
          9078 => x"73",
          9079 => x"6e",
          9080 => x"2e",
          9081 => x"69",
          9082 => x"61",
          9083 => x"61",
          9084 => x"65",
          9085 => x"74",
          9086 => x"00",
          9087 => x"69",
          9088 => x"68",
          9089 => x"6c",
          9090 => x"6e",
          9091 => x"69",
          9092 => x"00",
          9093 => x"44",
          9094 => x"20",
          9095 => x"74",
          9096 => x"72",
          9097 => x"63",
          9098 => x"2e",
          9099 => x"72",
          9100 => x"20",
          9101 => x"62",
          9102 => x"69",
          9103 => x"6e",
          9104 => x"69",
          9105 => x"00",
          9106 => x"69",
          9107 => x"6e",
          9108 => x"65",
          9109 => x"6c",
          9110 => x"00",
          9111 => x"6f",
          9112 => x"6d",
          9113 => x"69",
          9114 => x"20",
          9115 => x"65",
          9116 => x"74",
          9117 => x"66",
          9118 => x"64",
          9119 => x"20",
          9120 => x"6b",
          9121 => x"6f",
          9122 => x"74",
          9123 => x"6f",
          9124 => x"64",
          9125 => x"69",
          9126 => x"75",
          9127 => x"6f",
          9128 => x"61",
          9129 => x"6e",
          9130 => x"6e",
          9131 => x"6c",
          9132 => x"00",
          9133 => x"69",
          9134 => x"69",
          9135 => x"6f",
          9136 => x"64",
          9137 => x"6e",
          9138 => x"66",
          9139 => x"65",
          9140 => x"6d",
          9141 => x"72",
          9142 => x"00",
          9143 => x"6f",
          9144 => x"61",
          9145 => x"6f",
          9146 => x"20",
          9147 => x"65",
          9148 => x"00",
          9149 => x"61",
          9150 => x"65",
          9151 => x"73",
          9152 => x"63",
          9153 => x"65",
          9154 => x"00",
          9155 => x"75",
          9156 => x"73",
          9157 => x"00",
          9158 => x"6e",
          9159 => x"77",
          9160 => x"72",
          9161 => x"2e",
          9162 => x"25",
          9163 => x"62",
          9164 => x"73",
          9165 => x"20",
          9166 => x"25",
          9167 => x"62",
          9168 => x"73",
          9169 => x"63",
          9170 => x"00",
          9171 => x"65",
          9172 => x"00",
          9173 => x"30",
          9174 => x"00",
          9175 => x"20",
          9176 => x"30",
          9177 => x"00",
          9178 => x"20",
          9179 => x"20",
          9180 => x"00",
          9181 => x"30",
          9182 => x"00",
          9183 => x"20",
          9184 => x"7c",
          9185 => x"00",
          9186 => x"4f",
          9187 => x"2a",
          9188 => x"73",
          9189 => x"00",
          9190 => x"32",
          9191 => x"2f",
          9192 => x"30",
          9193 => x"31",
          9194 => x"00",
          9195 => x"5a",
          9196 => x"20",
          9197 => x"20",
          9198 => x"78",
          9199 => x"73",
          9200 => x"20",
          9201 => x"0a",
          9202 => x"50",
          9203 => x"6e",
          9204 => x"72",
          9205 => x"20",
          9206 => x"64",
          9207 => x"00",
          9208 => x"69",
          9209 => x"20",
          9210 => x"65",
          9211 => x"70",
          9212 => x"53",
          9213 => x"6e",
          9214 => x"72",
          9215 => x"00",
          9216 => x"4f",
          9217 => x"20",
          9218 => x"69",
          9219 => x"72",
          9220 => x"74",
          9221 => x"4f",
          9222 => x"20",
          9223 => x"69",
          9224 => x"72",
          9225 => x"74",
          9226 => x"41",
          9227 => x"20",
          9228 => x"69",
          9229 => x"72",
          9230 => x"74",
          9231 => x"41",
          9232 => x"20",
          9233 => x"69",
          9234 => x"72",
          9235 => x"74",
          9236 => x"41",
          9237 => x"20",
          9238 => x"69",
          9239 => x"72",
          9240 => x"74",
          9241 => x"41",
          9242 => x"20",
          9243 => x"69",
          9244 => x"72",
          9245 => x"74",
          9246 => x"65",
          9247 => x"6e",
          9248 => x"70",
          9249 => x"6d",
          9250 => x"2e",
          9251 => x"6e",
          9252 => x"69",
          9253 => x"74",
          9254 => x"72",
          9255 => x"00",
          9256 => x"75",
          9257 => x"78",
          9258 => x"62",
          9259 => x"00",
          9260 => x"4f",
          9261 => x"73",
          9262 => x"3a",
          9263 => x"61",
          9264 => x"64",
          9265 => x"20",
          9266 => x"74",
          9267 => x"69",
          9268 => x"73",
          9269 => x"61",
          9270 => x"30",
          9271 => x"6c",
          9272 => x"65",
          9273 => x"69",
          9274 => x"61",
          9275 => x"6c",
          9276 => x"00",
          9277 => x"20",
          9278 => x"6c",
          9279 => x"69",
          9280 => x"2e",
          9281 => x"00",
          9282 => x"6f",
          9283 => x"6e",
          9284 => x"2e",
          9285 => x"6f",
          9286 => x"72",
          9287 => x"2e",
          9288 => x"00",
          9289 => x"30",
          9290 => x"28",
          9291 => x"78",
          9292 => x"25",
          9293 => x"78",
          9294 => x"38",
          9295 => x"00",
          9296 => x"75",
          9297 => x"4d",
          9298 => x"72",
          9299 => x"43",
          9300 => x"6c",
          9301 => x"2e",
          9302 => x"30",
          9303 => x"20",
          9304 => x"58",
          9305 => x"3f",
          9306 => x"30",
          9307 => x"20",
          9308 => x"58",
          9309 => x"30",
          9310 => x"20",
          9311 => x"6c",
          9312 => x"00",
          9313 => x"78",
          9314 => x"74",
          9315 => x"20",
          9316 => x"65",
          9317 => x"25",
          9318 => x"78",
          9319 => x"2e",
          9320 => x"61",
          9321 => x"6e",
          9322 => x"6f",
          9323 => x"40",
          9324 => x"38",
          9325 => x"2e",
          9326 => x"00",
          9327 => x"61",
          9328 => x"72",
          9329 => x"72",
          9330 => x"20",
          9331 => x"65",
          9332 => x"64",
          9333 => x"00",
          9334 => x"65",
          9335 => x"72",
          9336 => x"67",
          9337 => x"70",
          9338 => x"61",
          9339 => x"6e",
          9340 => x"00",
          9341 => x"6f",
          9342 => x"72",
          9343 => x"6f",
          9344 => x"67",
          9345 => x"00",
          9346 => x"50",
          9347 => x"69",
          9348 => x"64",
          9349 => x"73",
          9350 => x"2e",
          9351 => x"00",
          9352 => x"64",
          9353 => x"73",
          9354 => x"00",
          9355 => x"64",
          9356 => x"73",
          9357 => x"61",
          9358 => x"6f",
          9359 => x"6e",
          9360 => x"00",
          9361 => x"75",
          9362 => x"6e",
          9363 => x"2e",
          9364 => x"6e",
          9365 => x"69",
          9366 => x"69",
          9367 => x"72",
          9368 => x"74",
          9369 => x"2e",
          9370 => x"64",
          9371 => x"2f",
          9372 => x"25",
          9373 => x"64",
          9374 => x"2e",
          9375 => x"64",
          9376 => x"6f",
          9377 => x"6f",
          9378 => x"67",
          9379 => x"74",
          9380 => x"00",
          9381 => x"28",
          9382 => x"6d",
          9383 => x"43",
          9384 => x"6e",
          9385 => x"29",
          9386 => x"0a",
          9387 => x"69",
          9388 => x"20",
          9389 => x"6c",
          9390 => x"6e",
          9391 => x"3a",
          9392 => x"20",
          9393 => x"42",
          9394 => x"52",
          9395 => x"20",
          9396 => x"38",
          9397 => x"30",
          9398 => x"2e",
          9399 => x"20",
          9400 => x"44",
          9401 => x"20",
          9402 => x"20",
          9403 => x"38",
          9404 => x"30",
          9405 => x"2e",
          9406 => x"20",
          9407 => x"4e",
          9408 => x"42",
          9409 => x"20",
          9410 => x"38",
          9411 => x"30",
          9412 => x"2e",
          9413 => x"20",
          9414 => x"52",
          9415 => x"20",
          9416 => x"20",
          9417 => x"38",
          9418 => x"30",
          9419 => x"2e",
          9420 => x"20",
          9421 => x"41",
          9422 => x"20",
          9423 => x"20",
          9424 => x"38",
          9425 => x"30",
          9426 => x"2e",
          9427 => x"20",
          9428 => x"44",
          9429 => x"52",
          9430 => x"20",
          9431 => x"76",
          9432 => x"73",
          9433 => x"30",
          9434 => x"2e",
          9435 => x"20",
          9436 => x"49",
          9437 => x"31",
          9438 => x"20",
          9439 => x"6d",
          9440 => x"20",
          9441 => x"30",
          9442 => x"2e",
          9443 => x"20",
          9444 => x"4e",
          9445 => x"43",
          9446 => x"20",
          9447 => x"61",
          9448 => x"6c",
          9449 => x"30",
          9450 => x"2e",
          9451 => x"20",
          9452 => x"49",
          9453 => x"4f",
          9454 => x"42",
          9455 => x"00",
          9456 => x"20",
          9457 => x"42",
          9458 => x"43",
          9459 => x"20",
          9460 => x"4f",
          9461 => x"0a",
          9462 => x"20",
          9463 => x"53",
          9464 => x"00",
          9465 => x"20",
          9466 => x"50",
          9467 => x"00",
          9468 => x"64",
          9469 => x"73",
          9470 => x"3a",
          9471 => x"20",
          9472 => x"50",
          9473 => x"65",
          9474 => x"20",
          9475 => x"74",
          9476 => x"41",
          9477 => x"65",
          9478 => x"3d",
          9479 => x"38",
          9480 => x"00",
          9481 => x"20",
          9482 => x"50",
          9483 => x"65",
          9484 => x"79",
          9485 => x"61",
          9486 => x"41",
          9487 => x"65",
          9488 => x"3d",
          9489 => x"38",
          9490 => x"00",
          9491 => x"20",
          9492 => x"74",
          9493 => x"20",
          9494 => x"72",
          9495 => x"64",
          9496 => x"73",
          9497 => x"20",
          9498 => x"3d",
          9499 => x"38",
          9500 => x"00",
          9501 => x"69",
          9502 => x"0a",
          9503 => x"20",
          9504 => x"50",
          9505 => x"64",
          9506 => x"20",
          9507 => x"20",
          9508 => x"20",
          9509 => x"20",
          9510 => x"3d",
          9511 => x"34",
          9512 => x"00",
          9513 => x"20",
          9514 => x"79",
          9515 => x"6d",
          9516 => x"6f",
          9517 => x"46",
          9518 => x"20",
          9519 => x"20",
          9520 => x"3d",
          9521 => x"2e",
          9522 => x"64",
          9523 => x"0a",
          9524 => x"20",
          9525 => x"44",
          9526 => x"20",
          9527 => x"63",
          9528 => x"72",
          9529 => x"20",
          9530 => x"20",
          9531 => x"3d",
          9532 => x"2e",
          9533 => x"64",
          9534 => x"0a",
          9535 => x"20",
          9536 => x"69",
          9537 => x"6f",
          9538 => x"53",
          9539 => x"4d",
          9540 => x"6f",
          9541 => x"46",
          9542 => x"3d",
          9543 => x"2e",
          9544 => x"64",
          9545 => x"0a",
          9546 => x"6d",
          9547 => x"00",
          9548 => x"65",
          9549 => x"6d",
          9550 => x"6c",
          9551 => x"00",
          9552 => x"56",
          9553 => x"56",
          9554 => x"6e",
          9555 => x"6e",
          9556 => x"77",
          9557 => x"00",
          9558 => x"00",
          9559 => x"00",
          9560 => x"00",
          9561 => x"00",
          9562 => x"00",
          9563 => x"00",
          9564 => x"00",
          9565 => x"00",
          9566 => x"00",
          9567 => x"00",
          9568 => x"00",
          9569 => x"00",
          9570 => x"00",
          9571 => x"00",
          9572 => x"00",
          9573 => x"00",
          9574 => x"00",
          9575 => x"00",
          9576 => x"00",
          9577 => x"00",
          9578 => x"00",
          9579 => x"00",
          9580 => x"00",
          9581 => x"00",
          9582 => x"00",
          9583 => x"00",
          9584 => x"00",
          9585 => x"00",
          9586 => x"00",
          9587 => x"00",
          9588 => x"00",
          9589 => x"00",
          9590 => x"00",
          9591 => x"00",
          9592 => x"00",
          9593 => x"00",
          9594 => x"00",
          9595 => x"00",
          9596 => x"00",
          9597 => x"00",
          9598 => x"00",
          9599 => x"00",
          9600 => x"00",
          9601 => x"00",
          9602 => x"00",
          9603 => x"00",
          9604 => x"00",
          9605 => x"00",
          9606 => x"00",
          9607 => x"00",
          9608 => x"00",
          9609 => x"00",
          9610 => x"00",
          9611 => x"00",
          9612 => x"00",
          9613 => x"00",
          9614 => x"00",
          9615 => x"00",
          9616 => x"00",
          9617 => x"00",
          9618 => x"00",
          9619 => x"00",
          9620 => x"00",
          9621 => x"00",
          9622 => x"00",
          9623 => x"5b",
          9624 => x"5b",
          9625 => x"5b",
          9626 => x"5b",
          9627 => x"5b",
          9628 => x"5b",
          9629 => x"5b",
          9630 => x"30",
          9631 => x"5b",
          9632 => x"5b",
          9633 => x"5b",
          9634 => x"00",
          9635 => x"00",
          9636 => x"00",
          9637 => x"00",
          9638 => x"00",
          9639 => x"00",
          9640 => x"00",
          9641 => x"00",
          9642 => x"00",
          9643 => x"00",
          9644 => x"00",
          9645 => x"69",
          9646 => x"72",
          9647 => x"69",
          9648 => x"00",
          9649 => x"00",
          9650 => x"30",
          9651 => x"20",
          9652 => x"0a",
          9653 => x"61",
          9654 => x"64",
          9655 => x"20",
          9656 => x"65",
          9657 => x"68",
          9658 => x"69",
          9659 => x"72",
          9660 => x"69",
          9661 => x"74",
          9662 => x"4f",
          9663 => x"00",
          9664 => x"61",
          9665 => x"74",
          9666 => x"65",
          9667 => x"72",
          9668 => x"65",
          9669 => x"73",
          9670 => x"79",
          9671 => x"6c",
          9672 => x"64",
          9673 => x"62",
          9674 => x"67",
          9675 => x"44",
          9676 => x"2a",
          9677 => x"3b",
          9678 => x"3f",
          9679 => x"7f",
          9680 => x"41",
          9681 => x"41",
          9682 => x"00",
          9683 => x"fe",
          9684 => x"44",
          9685 => x"2e",
          9686 => x"4f",
          9687 => x"4d",
          9688 => x"20",
          9689 => x"54",
          9690 => x"20",
          9691 => x"4f",
          9692 => x"4d",
          9693 => x"20",
          9694 => x"54",
          9695 => x"20",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"9a",
          9701 => x"41",
          9702 => x"45",
          9703 => x"49",
          9704 => x"92",
          9705 => x"4f",
          9706 => x"99",
          9707 => x"9d",
          9708 => x"49",
          9709 => x"a5",
          9710 => x"a9",
          9711 => x"ad",
          9712 => x"b1",
          9713 => x"b5",
          9714 => x"b9",
          9715 => x"bd",
          9716 => x"c1",
          9717 => x"c5",
          9718 => x"c9",
          9719 => x"cd",
          9720 => x"d1",
          9721 => x"d5",
          9722 => x"d9",
          9723 => x"dd",
          9724 => x"e1",
          9725 => x"e5",
          9726 => x"e9",
          9727 => x"ed",
          9728 => x"f1",
          9729 => x"f5",
          9730 => x"f9",
          9731 => x"fd",
          9732 => x"2e",
          9733 => x"5b",
          9734 => x"22",
          9735 => x"3e",
          9736 => x"00",
          9737 => x"01",
          9738 => x"10",
          9739 => x"00",
          9740 => x"00",
          9741 => x"01",
          9742 => x"04",
          9743 => x"10",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"02",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"04",
          9752 => x"00",
          9753 => x"00",
          9754 => x"00",
          9755 => x"14",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"2b",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"30",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"3c",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"3d",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"3f",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"40",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"41",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"42",
          9788 => x"00",
          9789 => x"00",
          9790 => x"00",
          9791 => x"43",
          9792 => x"00",
          9793 => x"00",
          9794 => x"00",
          9795 => x"50",
          9796 => x"00",
          9797 => x"00",
          9798 => x"00",
          9799 => x"51",
          9800 => x"00",
          9801 => x"00",
          9802 => x"00",
          9803 => x"54",
          9804 => x"00",
          9805 => x"00",
          9806 => x"00",
          9807 => x"55",
          9808 => x"00",
          9809 => x"00",
          9810 => x"00",
          9811 => x"79",
          9812 => x"00",
          9813 => x"00",
          9814 => x"00",
          9815 => x"78",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"82",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"83",
          9824 => x"00",
          9825 => x"00",
          9826 => x"00",
          9827 => x"85",
          9828 => x"00",
          9829 => x"00",
          9830 => x"00",
          9831 => x"87",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"8c",
          9836 => x"00",
          9837 => x"00",
          9838 => x"00",
          9839 => x"8d",
          9840 => x"00",
          9841 => x"00",
          9842 => x"00",
          9843 => x"8e",
          9844 => x"00",
          9845 => x"00",
          9846 => x"00",
          9847 => x"8f",
          9848 => x"00",
          9849 => x"00",
          9850 => x"00",
          9851 => x"00",
          9852 => x"00",
          9853 => x"00",
          9854 => x"00",
          9855 => x"01",
          9856 => x"00",
          9857 => x"01",
          9858 => x"81",
          9859 => x"00",
          9860 => x"7f",
          9861 => x"00",
          9862 => x"00",
          9863 => x"00",
          9864 => x"00",
          9865 => x"f5",
          9866 => x"f5",
          9867 => x"f5",
          9868 => x"00",
          9869 => x"01",
          9870 => x"01",
          9871 => x"01",
          9872 => x"00",
          9873 => x"00",
          9874 => x"00",
          9875 => x"00",
          9876 => x"00",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"00",
          9881 => x"00",
          9882 => x"00",
          9883 => x"00",
          9884 => x"00",
          9885 => x"00",
          9886 => x"00",
          9887 => x"00",
          9888 => x"00",
          9889 => x"00",
          9890 => x"00",
          9891 => x"00",
          9892 => x"00",
          9893 => x"00",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"00",
          9898 => x"00",
          9899 => x"00",
          9900 => x"00",
          9901 => x"00",
          9902 => x"00",
          9903 => x"00",
          9904 => x"00",
          9905 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"9d",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"98",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"f4",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"e0",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"95",
           269 => x"0b",
           270 => x"0b",
           271 => x"b3",
           272 => x"0b",
           273 => x"0b",
           274 => x"d1",
           275 => x"0b",
           276 => x"0b",
           277 => x"f0",
           278 => x"0b",
           279 => x"0b",
           280 => x"8f",
           281 => x"0b",
           282 => x"0b",
           283 => x"ad",
           284 => x"0b",
           285 => x"0b",
           286 => x"cd",
           287 => x"0b",
           288 => x"0b",
           289 => x"ed",
           290 => x"0b",
           291 => x"0b",
           292 => x"8d",
           293 => x"0b",
           294 => x"0b",
           295 => x"ad",
           296 => x"0b",
           297 => x"0b",
           298 => x"cd",
           299 => x"0b",
           300 => x"0b",
           301 => x"ed",
           302 => x"0b",
           303 => x"0b",
           304 => x"8d",
           305 => x"0b",
           306 => x"0b",
           307 => x"ad",
           308 => x"0b",
           309 => x"0b",
           310 => x"cd",
           311 => x"0b",
           312 => x"0b",
           313 => x"ed",
           314 => x"0b",
           315 => x"0b",
           316 => x"8d",
           317 => x"0b",
           318 => x"0b",
           319 => x"ad",
           320 => x"0b",
           321 => x"0b",
           322 => x"cd",
           323 => x"0b",
           324 => x"0b",
           325 => x"ed",
           326 => x"0b",
           327 => x"0b",
           328 => x"8d",
           329 => x"0b",
           330 => x"0b",
           331 => x"ad",
           332 => x"0b",
           333 => x"0b",
           334 => x"cd",
           335 => x"0b",
           336 => x"0b",
           337 => x"ed",
           338 => x"0b",
           339 => x"0b",
           340 => x"8d",
           341 => x"0b",
           342 => x"0b",
           343 => x"ad",
           344 => x"0b",
           345 => x"0b",
           346 => x"cd",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"04",
           390 => x"0c",
           391 => x"82",
           392 => x"82",
           393 => x"82",
           394 => x"af",
           395 => x"b5",
           396 => x"d0",
           397 => x"b5",
           398 => x"ad",
           399 => x"d4",
           400 => x"90",
           401 => x"d4",
           402 => x"2d",
           403 => x"08",
           404 => x"04",
           405 => x"0c",
           406 => x"82",
           407 => x"82",
           408 => x"82",
           409 => x"80",
           410 => x"82",
           411 => x"82",
           412 => x"82",
           413 => x"80",
           414 => x"82",
           415 => x"82",
           416 => x"82",
           417 => x"93",
           418 => x"b5",
           419 => x"d0",
           420 => x"b5",
           421 => x"c0",
           422 => x"d4",
           423 => x"90",
           424 => x"d4",
           425 => x"2d",
           426 => x"08",
           427 => x"04",
           428 => x"0c",
           429 => x"2d",
           430 => x"08",
           431 => x"04",
           432 => x"0c",
           433 => x"2d",
           434 => x"08",
           435 => x"04",
           436 => x"0c",
           437 => x"2d",
           438 => x"08",
           439 => x"04",
           440 => x"0c",
           441 => x"2d",
           442 => x"08",
           443 => x"04",
           444 => x"0c",
           445 => x"2d",
           446 => x"08",
           447 => x"04",
           448 => x"0c",
           449 => x"2d",
           450 => x"08",
           451 => x"04",
           452 => x"0c",
           453 => x"2d",
           454 => x"08",
           455 => x"04",
           456 => x"0c",
           457 => x"2d",
           458 => x"08",
           459 => x"04",
           460 => x"0c",
           461 => x"2d",
           462 => x"08",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"04",
           468 => x"0c",
           469 => x"2d",
           470 => x"08",
           471 => x"04",
           472 => x"0c",
           473 => x"2d",
           474 => x"08",
           475 => x"04",
           476 => x"0c",
           477 => x"2d",
           478 => x"08",
           479 => x"04",
           480 => x"0c",
           481 => x"2d",
           482 => x"08",
           483 => x"04",
           484 => x"0c",
           485 => x"2d",
           486 => x"08",
           487 => x"04",
           488 => x"0c",
           489 => x"2d",
           490 => x"08",
           491 => x"04",
           492 => x"0c",
           493 => x"2d",
           494 => x"08",
           495 => x"04",
           496 => x"0c",
           497 => x"2d",
           498 => x"08",
           499 => x"04",
           500 => x"0c",
           501 => x"2d",
           502 => x"08",
           503 => x"04",
           504 => x"0c",
           505 => x"2d",
           506 => x"08",
           507 => x"04",
           508 => x"0c",
           509 => x"2d",
           510 => x"08",
           511 => x"04",
           512 => x"0c",
           513 => x"2d",
           514 => x"08",
           515 => x"04",
           516 => x"0c",
           517 => x"2d",
           518 => x"08",
           519 => x"04",
           520 => x"0c",
           521 => x"2d",
           522 => x"08",
           523 => x"04",
           524 => x"0c",
           525 => x"2d",
           526 => x"08",
           527 => x"04",
           528 => x"0c",
           529 => x"2d",
           530 => x"08",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"04",
           536 => x"0c",
           537 => x"2d",
           538 => x"08",
           539 => x"04",
           540 => x"0c",
           541 => x"2d",
           542 => x"08",
           543 => x"04",
           544 => x"0c",
           545 => x"2d",
           546 => x"08",
           547 => x"04",
           548 => x"0c",
           549 => x"2d",
           550 => x"08",
           551 => x"04",
           552 => x"0c",
           553 => x"2d",
           554 => x"08",
           555 => x"04",
           556 => x"0c",
           557 => x"2d",
           558 => x"08",
           559 => x"04",
           560 => x"0c",
           561 => x"2d",
           562 => x"08",
           563 => x"04",
           564 => x"0c",
           565 => x"2d",
           566 => x"08",
           567 => x"04",
           568 => x"0c",
           569 => x"2d",
           570 => x"08",
           571 => x"04",
           572 => x"0c",
           573 => x"2d",
           574 => x"08",
           575 => x"04",
           576 => x"0c",
           577 => x"2d",
           578 => x"08",
           579 => x"04",
           580 => x"0c",
           581 => x"2d",
           582 => x"08",
           583 => x"04",
           584 => x"0c",
           585 => x"2d",
           586 => x"08",
           587 => x"04",
           588 => x"0c",
           589 => x"2d",
           590 => x"08",
           591 => x"04",
           592 => x"0c",
           593 => x"2d",
           594 => x"08",
           595 => x"04",
           596 => x"0c",
           597 => x"2d",
           598 => x"08",
           599 => x"04",
           600 => x"00",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"53",
           609 => x"00",
           610 => x"06",
           611 => x"09",
           612 => x"05",
           613 => x"2b",
           614 => x"06",
           615 => x"04",
           616 => x"72",
           617 => x"05",
           618 => x"05",
           619 => x"72",
           620 => x"53",
           621 => x"51",
           622 => x"04",
           623 => x"70",
           624 => x"27",
           625 => x"71",
           626 => x"53",
           627 => x"0b",
           628 => x"8c",
           629 => x"ee",
           630 => x"82",
           631 => x"02",
           632 => x"0c",
           633 => x"82",
           634 => x"8c",
           635 => x"b5",
           636 => x"05",
           637 => x"d4",
           638 => x"08",
           639 => x"d4",
           640 => x"08",
           641 => x"9c",
           642 => x"84",
           643 => x"b5",
           644 => x"82",
           645 => x"f8",
           646 => x"b5",
           647 => x"05",
           648 => x"b5",
           649 => x"54",
           650 => x"82",
           651 => x"04",
           652 => x"08",
           653 => x"d4",
           654 => x"0d",
           655 => x"08",
           656 => x"85",
           657 => x"81",
           658 => x"06",
           659 => x"52",
           660 => x"80",
           661 => x"d4",
           662 => x"08",
           663 => x"8d",
           664 => x"82",
           665 => x"f4",
           666 => x"c4",
           667 => x"d4",
           668 => x"08",
           669 => x"b5",
           670 => x"05",
           671 => x"82",
           672 => x"f8",
           673 => x"b5",
           674 => x"05",
           675 => x"d4",
           676 => x"0c",
           677 => x"08",
           678 => x"8a",
           679 => x"38",
           680 => x"b5",
           681 => x"05",
           682 => x"e9",
           683 => x"d4",
           684 => x"08",
           685 => x"3f",
           686 => x"08",
           687 => x"d4",
           688 => x"0c",
           689 => x"d4",
           690 => x"08",
           691 => x"81",
           692 => x"80",
           693 => x"d4",
           694 => x"0c",
           695 => x"82",
           696 => x"fc",
           697 => x"b5",
           698 => x"05",
           699 => x"71",
           700 => x"b5",
           701 => x"05",
           702 => x"82",
           703 => x"8c",
           704 => x"b5",
           705 => x"05",
           706 => x"82",
           707 => x"fc",
           708 => x"80",
           709 => x"d4",
           710 => x"08",
           711 => x"34",
           712 => x"08",
           713 => x"70",
           714 => x"08",
           715 => x"52",
           716 => x"08",
           717 => x"82",
           718 => x"87",
           719 => x"b5",
           720 => x"82",
           721 => x"02",
           722 => x"0c",
           723 => x"86",
           724 => x"d4",
           725 => x"34",
           726 => x"08",
           727 => x"82",
           728 => x"e0",
           729 => x"0a",
           730 => x"d4",
           731 => x"0c",
           732 => x"08",
           733 => x"82",
           734 => x"fc",
           735 => x"b5",
           736 => x"05",
           737 => x"b5",
           738 => x"05",
           739 => x"b5",
           740 => x"05",
           741 => x"54",
           742 => x"82",
           743 => x"70",
           744 => x"08",
           745 => x"82",
           746 => x"ec",
           747 => x"b5",
           748 => x"05",
           749 => x"54",
           750 => x"82",
           751 => x"dc",
           752 => x"82",
           753 => x"54",
           754 => x"82",
           755 => x"04",
           756 => x"08",
           757 => x"d4",
           758 => x"0d",
           759 => x"08",
           760 => x"82",
           761 => x"fc",
           762 => x"b5",
           763 => x"05",
           764 => x"b5",
           765 => x"05",
           766 => x"b5",
           767 => x"05",
           768 => x"a3",
           769 => x"c8",
           770 => x"b5",
           771 => x"05",
           772 => x"d4",
           773 => x"08",
           774 => x"c8",
           775 => x"87",
           776 => x"b5",
           777 => x"82",
           778 => x"02",
           779 => x"0c",
           780 => x"80",
           781 => x"d4",
           782 => x"23",
           783 => x"08",
           784 => x"53",
           785 => x"14",
           786 => x"d4",
           787 => x"08",
           788 => x"70",
           789 => x"81",
           790 => x"06",
           791 => x"51",
           792 => x"2e",
           793 => x"0b",
           794 => x"08",
           795 => x"96",
           796 => x"b5",
           797 => x"05",
           798 => x"33",
           799 => x"b5",
           800 => x"05",
           801 => x"ff",
           802 => x"80",
           803 => x"38",
           804 => x"08",
           805 => x"81",
           806 => x"d4",
           807 => x"0c",
           808 => x"08",
           809 => x"70",
           810 => x"53",
           811 => x"95",
           812 => x"b5",
           813 => x"05",
           814 => x"73",
           815 => x"38",
           816 => x"08",
           817 => x"53",
           818 => x"81",
           819 => x"b5",
           820 => x"05",
           821 => x"b0",
           822 => x"06",
           823 => x"82",
           824 => x"e8",
           825 => x"98",
           826 => x"2c",
           827 => x"72",
           828 => x"b5",
           829 => x"05",
           830 => x"2a",
           831 => x"70",
           832 => x"51",
           833 => x"80",
           834 => x"82",
           835 => x"e4",
           836 => x"82",
           837 => x"53",
           838 => x"d4",
           839 => x"23",
           840 => x"82",
           841 => x"e8",
           842 => x"98",
           843 => x"2c",
           844 => x"2b",
           845 => x"11",
           846 => x"53",
           847 => x"72",
           848 => x"08",
           849 => x"82",
           850 => x"e8",
           851 => x"82",
           852 => x"f8",
           853 => x"15",
           854 => x"51",
           855 => x"b5",
           856 => x"05",
           857 => x"d4",
           858 => x"33",
           859 => x"70",
           860 => x"51",
           861 => x"25",
           862 => x"ff",
           863 => x"d4",
           864 => x"34",
           865 => x"08",
           866 => x"70",
           867 => x"81",
           868 => x"53",
           869 => x"38",
           870 => x"08",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"53",
           876 => x"d4",
           877 => x"23",
           878 => x"82",
           879 => x"e4",
           880 => x"83",
           881 => x"06",
           882 => x"72",
           883 => x"38",
           884 => x"08",
           885 => x"70",
           886 => x"98",
           887 => x"53",
           888 => x"81",
           889 => x"d4",
           890 => x"34",
           891 => x"08",
           892 => x"e0",
           893 => x"d4",
           894 => x"0c",
           895 => x"d4",
           896 => x"08",
           897 => x"92",
           898 => x"b5",
           899 => x"05",
           900 => x"2b",
           901 => x"11",
           902 => x"51",
           903 => x"04",
           904 => x"08",
           905 => x"70",
           906 => x"53",
           907 => x"d4",
           908 => x"23",
           909 => x"08",
           910 => x"70",
           911 => x"53",
           912 => x"d4",
           913 => x"23",
           914 => x"82",
           915 => x"e4",
           916 => x"81",
           917 => x"53",
           918 => x"d4",
           919 => x"23",
           920 => x"82",
           921 => x"e4",
           922 => x"80",
           923 => x"53",
           924 => x"d4",
           925 => x"23",
           926 => x"82",
           927 => x"e4",
           928 => x"88",
           929 => x"72",
           930 => x"08",
           931 => x"80",
           932 => x"d4",
           933 => x"34",
           934 => x"82",
           935 => x"e4",
           936 => x"84",
           937 => x"72",
           938 => x"08",
           939 => x"fb",
           940 => x"0b",
           941 => x"08",
           942 => x"82",
           943 => x"ec",
           944 => x"11",
           945 => x"82",
           946 => x"ec",
           947 => x"e3",
           948 => x"d4",
           949 => x"34",
           950 => x"82",
           951 => x"90",
           952 => x"b5",
           953 => x"05",
           954 => x"82",
           955 => x"90",
           956 => x"08",
           957 => x"82",
           958 => x"fc",
           959 => x"b5",
           960 => x"05",
           961 => x"51",
           962 => x"b5",
           963 => x"05",
           964 => x"39",
           965 => x"08",
           966 => x"82",
           967 => x"90",
           968 => x"05",
           969 => x"08",
           970 => x"70",
           971 => x"d4",
           972 => x"0c",
           973 => x"08",
           974 => x"70",
           975 => x"81",
           976 => x"51",
           977 => x"2e",
           978 => x"b5",
           979 => x"05",
           980 => x"2b",
           981 => x"2c",
           982 => x"d4",
           983 => x"08",
           984 => x"d8",
           985 => x"c8",
           986 => x"82",
           987 => x"f4",
           988 => x"39",
           989 => x"08",
           990 => x"51",
           991 => x"82",
           992 => x"53",
           993 => x"d4",
           994 => x"23",
           995 => x"08",
           996 => x"53",
           997 => x"08",
           998 => x"73",
           999 => x"54",
          1000 => x"d4",
          1001 => x"23",
          1002 => x"82",
          1003 => x"90",
          1004 => x"b5",
          1005 => x"05",
          1006 => x"82",
          1007 => x"90",
          1008 => x"08",
          1009 => x"08",
          1010 => x"82",
          1011 => x"e4",
          1012 => x"83",
          1013 => x"06",
          1014 => x"53",
          1015 => x"ab",
          1016 => x"d4",
          1017 => x"33",
          1018 => x"53",
          1019 => x"53",
          1020 => x"08",
          1021 => x"52",
          1022 => x"3f",
          1023 => x"08",
          1024 => x"b5",
          1025 => x"05",
          1026 => x"82",
          1027 => x"fc",
          1028 => x"9b",
          1029 => x"b5",
          1030 => x"72",
          1031 => x"08",
          1032 => x"82",
          1033 => x"ec",
          1034 => x"82",
          1035 => x"f4",
          1036 => x"71",
          1037 => x"72",
          1038 => x"08",
          1039 => x"8a",
          1040 => x"b5",
          1041 => x"05",
          1042 => x"2a",
          1043 => x"51",
          1044 => x"80",
          1045 => x"82",
          1046 => x"90",
          1047 => x"b5",
          1048 => x"05",
          1049 => x"82",
          1050 => x"90",
          1051 => x"08",
          1052 => x"08",
          1053 => x"53",
          1054 => x"b5",
          1055 => x"05",
          1056 => x"d4",
          1057 => x"08",
          1058 => x"b5",
          1059 => x"05",
          1060 => x"82",
          1061 => x"dc",
          1062 => x"82",
          1063 => x"dc",
          1064 => x"b5",
          1065 => x"05",
          1066 => x"d4",
          1067 => x"08",
          1068 => x"38",
          1069 => x"08",
          1070 => x"70",
          1071 => x"53",
          1072 => x"d4",
          1073 => x"23",
          1074 => x"08",
          1075 => x"30",
          1076 => x"08",
          1077 => x"82",
          1078 => x"e4",
          1079 => x"ff",
          1080 => x"53",
          1081 => x"d4",
          1082 => x"23",
          1083 => x"88",
          1084 => x"d4",
          1085 => x"23",
          1086 => x"b5",
          1087 => x"05",
          1088 => x"c0",
          1089 => x"72",
          1090 => x"08",
          1091 => x"80",
          1092 => x"b5",
          1093 => x"05",
          1094 => x"82",
          1095 => x"f4",
          1096 => x"b5",
          1097 => x"05",
          1098 => x"2a",
          1099 => x"51",
          1100 => x"80",
          1101 => x"82",
          1102 => x"90",
          1103 => x"b5",
          1104 => x"05",
          1105 => x"82",
          1106 => x"90",
          1107 => x"08",
          1108 => x"08",
          1109 => x"53",
          1110 => x"b5",
          1111 => x"05",
          1112 => x"d4",
          1113 => x"08",
          1114 => x"b5",
          1115 => x"05",
          1116 => x"82",
          1117 => x"d8",
          1118 => x"82",
          1119 => x"d8",
          1120 => x"b5",
          1121 => x"05",
          1122 => x"d4",
          1123 => x"22",
          1124 => x"51",
          1125 => x"b5",
          1126 => x"05",
          1127 => x"d8",
          1128 => x"d4",
          1129 => x"0c",
          1130 => x"08",
          1131 => x"82",
          1132 => x"f4",
          1133 => x"b5",
          1134 => x"05",
          1135 => x"70",
          1136 => x"55",
          1137 => x"82",
          1138 => x"53",
          1139 => x"82",
          1140 => x"f0",
          1141 => x"b5",
          1142 => x"05",
          1143 => x"d4",
          1144 => x"08",
          1145 => x"53",
          1146 => x"a4",
          1147 => x"d4",
          1148 => x"08",
          1149 => x"54",
          1150 => x"08",
          1151 => x"70",
          1152 => x"51",
          1153 => x"82",
          1154 => x"d0",
          1155 => x"39",
          1156 => x"08",
          1157 => x"53",
          1158 => x"11",
          1159 => x"82",
          1160 => x"d0",
          1161 => x"b5",
          1162 => x"05",
          1163 => x"b5",
          1164 => x"05",
          1165 => x"82",
          1166 => x"f0",
          1167 => x"05",
          1168 => x"08",
          1169 => x"82",
          1170 => x"f4",
          1171 => x"53",
          1172 => x"08",
          1173 => x"52",
          1174 => x"3f",
          1175 => x"08",
          1176 => x"d4",
          1177 => x"0c",
          1178 => x"d4",
          1179 => x"08",
          1180 => x"38",
          1181 => x"82",
          1182 => x"f0",
          1183 => x"b5",
          1184 => x"72",
          1185 => x"75",
          1186 => x"72",
          1187 => x"08",
          1188 => x"82",
          1189 => x"e4",
          1190 => x"b2",
          1191 => x"72",
          1192 => x"38",
          1193 => x"08",
          1194 => x"ff",
          1195 => x"72",
          1196 => x"08",
          1197 => x"82",
          1198 => x"e4",
          1199 => x"86",
          1200 => x"06",
          1201 => x"72",
          1202 => x"e7",
          1203 => x"d4",
          1204 => x"22",
          1205 => x"82",
          1206 => x"cc",
          1207 => x"b5",
          1208 => x"05",
          1209 => x"82",
          1210 => x"cc",
          1211 => x"b5",
          1212 => x"05",
          1213 => x"72",
          1214 => x"81",
          1215 => x"82",
          1216 => x"cc",
          1217 => x"05",
          1218 => x"b5",
          1219 => x"05",
          1220 => x"82",
          1221 => x"cc",
          1222 => x"05",
          1223 => x"b5",
          1224 => x"05",
          1225 => x"d4",
          1226 => x"22",
          1227 => x"08",
          1228 => x"82",
          1229 => x"e4",
          1230 => x"83",
          1231 => x"06",
          1232 => x"72",
          1233 => x"d0",
          1234 => x"d4",
          1235 => x"33",
          1236 => x"70",
          1237 => x"b5",
          1238 => x"05",
          1239 => x"51",
          1240 => x"24",
          1241 => x"b5",
          1242 => x"05",
          1243 => x"06",
          1244 => x"82",
          1245 => x"e4",
          1246 => x"39",
          1247 => x"08",
          1248 => x"53",
          1249 => x"08",
          1250 => x"73",
          1251 => x"54",
          1252 => x"d4",
          1253 => x"34",
          1254 => x"08",
          1255 => x"70",
          1256 => x"81",
          1257 => x"53",
          1258 => x"b1",
          1259 => x"d4",
          1260 => x"33",
          1261 => x"70",
          1262 => x"90",
          1263 => x"2c",
          1264 => x"51",
          1265 => x"82",
          1266 => x"ec",
          1267 => x"75",
          1268 => x"72",
          1269 => x"08",
          1270 => x"af",
          1271 => x"d4",
          1272 => x"33",
          1273 => x"70",
          1274 => x"90",
          1275 => x"2c",
          1276 => x"51",
          1277 => x"82",
          1278 => x"ec",
          1279 => x"75",
          1280 => x"72",
          1281 => x"08",
          1282 => x"82",
          1283 => x"e4",
          1284 => x"83",
          1285 => x"53",
          1286 => x"82",
          1287 => x"ec",
          1288 => x"11",
          1289 => x"82",
          1290 => x"ec",
          1291 => x"90",
          1292 => x"2c",
          1293 => x"73",
          1294 => x"82",
          1295 => x"88",
          1296 => x"a0",
          1297 => x"3f",
          1298 => x"b5",
          1299 => x"05",
          1300 => x"2a",
          1301 => x"51",
          1302 => x"80",
          1303 => x"82",
          1304 => x"88",
          1305 => x"ad",
          1306 => x"3f",
          1307 => x"82",
          1308 => x"e4",
          1309 => x"84",
          1310 => x"06",
          1311 => x"72",
          1312 => x"38",
          1313 => x"08",
          1314 => x"52",
          1315 => x"a5",
          1316 => x"82",
          1317 => x"e4",
          1318 => x"85",
          1319 => x"06",
          1320 => x"72",
          1321 => x"38",
          1322 => x"08",
          1323 => x"52",
          1324 => x"81",
          1325 => x"d4",
          1326 => x"22",
          1327 => x"70",
          1328 => x"51",
          1329 => x"2e",
          1330 => x"b5",
          1331 => x"05",
          1332 => x"51",
          1333 => x"82",
          1334 => x"f4",
          1335 => x"72",
          1336 => x"81",
          1337 => x"82",
          1338 => x"88",
          1339 => x"82",
          1340 => x"f8",
          1341 => x"89",
          1342 => x"b5",
          1343 => x"05",
          1344 => x"2a",
          1345 => x"51",
          1346 => x"80",
          1347 => x"82",
          1348 => x"ec",
          1349 => x"11",
          1350 => x"82",
          1351 => x"ec",
          1352 => x"90",
          1353 => x"2c",
          1354 => x"73",
          1355 => x"82",
          1356 => x"88",
          1357 => x"b0",
          1358 => x"3f",
          1359 => x"b5",
          1360 => x"05",
          1361 => x"2a",
          1362 => x"51",
          1363 => x"80",
          1364 => x"82",
          1365 => x"e8",
          1366 => x"11",
          1367 => x"82",
          1368 => x"e8",
          1369 => x"98",
          1370 => x"2c",
          1371 => x"73",
          1372 => x"82",
          1373 => x"88",
          1374 => x"b0",
          1375 => x"3f",
          1376 => x"b5",
          1377 => x"05",
          1378 => x"2a",
          1379 => x"51",
          1380 => x"b0",
          1381 => x"d4",
          1382 => x"22",
          1383 => x"54",
          1384 => x"d4",
          1385 => x"23",
          1386 => x"70",
          1387 => x"53",
          1388 => x"90",
          1389 => x"d4",
          1390 => x"08",
          1391 => x"87",
          1392 => x"39",
          1393 => x"08",
          1394 => x"53",
          1395 => x"2e",
          1396 => x"97",
          1397 => x"d4",
          1398 => x"08",
          1399 => x"d4",
          1400 => x"33",
          1401 => x"3f",
          1402 => x"82",
          1403 => x"f8",
          1404 => x"72",
          1405 => x"09",
          1406 => x"cb",
          1407 => x"d4",
          1408 => x"22",
          1409 => x"53",
          1410 => x"d4",
          1411 => x"23",
          1412 => x"ff",
          1413 => x"83",
          1414 => x"81",
          1415 => x"b5",
          1416 => x"05",
          1417 => x"b5",
          1418 => x"05",
          1419 => x"52",
          1420 => x"08",
          1421 => x"81",
          1422 => x"d4",
          1423 => x"0c",
          1424 => x"3f",
          1425 => x"82",
          1426 => x"f8",
          1427 => x"72",
          1428 => x"09",
          1429 => x"cb",
          1430 => x"d4",
          1431 => x"22",
          1432 => x"53",
          1433 => x"d4",
          1434 => x"23",
          1435 => x"ff",
          1436 => x"83",
          1437 => x"80",
          1438 => x"b5",
          1439 => x"05",
          1440 => x"b5",
          1441 => x"05",
          1442 => x"52",
          1443 => x"3f",
          1444 => x"08",
          1445 => x"81",
          1446 => x"d4",
          1447 => x"0c",
          1448 => x"82",
          1449 => x"f0",
          1450 => x"b5",
          1451 => x"38",
          1452 => x"08",
          1453 => x"52",
          1454 => x"08",
          1455 => x"ff",
          1456 => x"d4",
          1457 => x"0c",
          1458 => x"08",
          1459 => x"70",
          1460 => x"85",
          1461 => x"39",
          1462 => x"08",
          1463 => x"70",
          1464 => x"81",
          1465 => x"53",
          1466 => x"80",
          1467 => x"b5",
          1468 => x"05",
          1469 => x"54",
          1470 => x"b5",
          1471 => x"05",
          1472 => x"2b",
          1473 => x"51",
          1474 => x"25",
          1475 => x"b5",
          1476 => x"05",
          1477 => x"51",
          1478 => x"d2",
          1479 => x"d4",
          1480 => x"08",
          1481 => x"d4",
          1482 => x"33",
          1483 => x"3f",
          1484 => x"b5",
          1485 => x"05",
          1486 => x"39",
          1487 => x"08",
          1488 => x"53",
          1489 => x"09",
          1490 => x"38",
          1491 => x"b5",
          1492 => x"05",
          1493 => x"82",
          1494 => x"ec",
          1495 => x"0b",
          1496 => x"08",
          1497 => x"8a",
          1498 => x"d4",
          1499 => x"23",
          1500 => x"82",
          1501 => x"88",
          1502 => x"82",
          1503 => x"f8",
          1504 => x"84",
          1505 => x"ea",
          1506 => x"d4",
          1507 => x"08",
          1508 => x"70",
          1509 => x"08",
          1510 => x"51",
          1511 => x"d4",
          1512 => x"08",
          1513 => x"0c",
          1514 => x"82",
          1515 => x"04",
          1516 => x"08",
          1517 => x"d4",
          1518 => x"0d",
          1519 => x"08",
          1520 => x"d4",
          1521 => x"08",
          1522 => x"d4",
          1523 => x"08",
          1524 => x"3f",
          1525 => x"08",
          1526 => x"c8",
          1527 => x"3d",
          1528 => x"d4",
          1529 => x"b5",
          1530 => x"82",
          1531 => x"fb",
          1532 => x"0b",
          1533 => x"08",
          1534 => x"82",
          1535 => x"85",
          1536 => x"81",
          1537 => x"32",
          1538 => x"51",
          1539 => x"53",
          1540 => x"8d",
          1541 => x"82",
          1542 => x"f4",
          1543 => x"92",
          1544 => x"d4",
          1545 => x"08",
          1546 => x"82",
          1547 => x"88",
          1548 => x"05",
          1549 => x"08",
          1550 => x"53",
          1551 => x"d4",
          1552 => x"34",
          1553 => x"06",
          1554 => x"2e",
          1555 => x"cd",
          1556 => x"cd",
          1557 => x"82",
          1558 => x"fc",
          1559 => x"90",
          1560 => x"53",
          1561 => x"b5",
          1562 => x"72",
          1563 => x"b1",
          1564 => x"82",
          1565 => x"f8",
          1566 => x"a5",
          1567 => x"9c",
          1568 => x"9c",
          1569 => x"8a",
          1570 => x"08",
          1571 => x"82",
          1572 => x"53",
          1573 => x"8a",
          1574 => x"82",
          1575 => x"f8",
          1576 => x"b5",
          1577 => x"05",
          1578 => x"b5",
          1579 => x"05",
          1580 => x"b5",
          1581 => x"05",
          1582 => x"c8",
          1583 => x"0d",
          1584 => x"0c",
          1585 => x"d4",
          1586 => x"b5",
          1587 => x"3d",
          1588 => x"82",
          1589 => x"f8",
          1590 => x"b5",
          1591 => x"05",
          1592 => x"33",
          1593 => x"70",
          1594 => x"81",
          1595 => x"51",
          1596 => x"80",
          1597 => x"ff",
          1598 => x"d4",
          1599 => x"0c",
          1600 => x"82",
          1601 => x"88",
          1602 => x"72",
          1603 => x"d4",
          1604 => x"08",
          1605 => x"b5",
          1606 => x"05",
          1607 => x"82",
          1608 => x"fc",
          1609 => x"81",
          1610 => x"72",
          1611 => x"38",
          1612 => x"08",
          1613 => x"82",
          1614 => x"8c",
          1615 => x"82",
          1616 => x"fc",
          1617 => x"90",
          1618 => x"53",
          1619 => x"b5",
          1620 => x"72",
          1621 => x"ab",
          1622 => x"82",
          1623 => x"f8",
          1624 => x"9f",
          1625 => x"d4",
          1626 => x"08",
          1627 => x"d4",
          1628 => x"0c",
          1629 => x"d4",
          1630 => x"08",
          1631 => x"0c",
          1632 => x"82",
          1633 => x"04",
          1634 => x"08",
          1635 => x"d4",
          1636 => x"0d",
          1637 => x"08",
          1638 => x"d4",
          1639 => x"08",
          1640 => x"82",
          1641 => x"70",
          1642 => x"0c",
          1643 => x"0d",
          1644 => x"0c",
          1645 => x"d4",
          1646 => x"b5",
          1647 => x"3d",
          1648 => x"d4",
          1649 => x"08",
          1650 => x"70",
          1651 => x"81",
          1652 => x"06",
          1653 => x"51",
          1654 => x"2e",
          1655 => x"0b",
          1656 => x"08",
          1657 => x"81",
          1658 => x"b5",
          1659 => x"05",
          1660 => x"33",
          1661 => x"70",
          1662 => x"51",
          1663 => x"80",
          1664 => x"38",
          1665 => x"08",
          1666 => x"82",
          1667 => x"8c",
          1668 => x"54",
          1669 => x"88",
          1670 => x"9f",
          1671 => x"d4",
          1672 => x"08",
          1673 => x"82",
          1674 => x"88",
          1675 => x"57",
          1676 => x"75",
          1677 => x"81",
          1678 => x"82",
          1679 => x"8c",
          1680 => x"11",
          1681 => x"8c",
          1682 => x"b5",
          1683 => x"05",
          1684 => x"b5",
          1685 => x"05",
          1686 => x"80",
          1687 => x"b5",
          1688 => x"05",
          1689 => x"d4",
          1690 => x"08",
          1691 => x"d4",
          1692 => x"08",
          1693 => x"06",
          1694 => x"08",
          1695 => x"72",
          1696 => x"c8",
          1697 => x"a3",
          1698 => x"d4",
          1699 => x"08",
          1700 => x"81",
          1701 => x"0c",
          1702 => x"08",
          1703 => x"70",
          1704 => x"08",
          1705 => x"51",
          1706 => x"ff",
          1707 => x"d4",
          1708 => x"0c",
          1709 => x"08",
          1710 => x"82",
          1711 => x"87",
          1712 => x"b5",
          1713 => x"82",
          1714 => x"02",
          1715 => x"0c",
          1716 => x"82",
          1717 => x"88",
          1718 => x"11",
          1719 => x"32",
          1720 => x"51",
          1721 => x"71",
          1722 => x"38",
          1723 => x"b5",
          1724 => x"05",
          1725 => x"39",
          1726 => x"08",
          1727 => x"85",
          1728 => x"86",
          1729 => x"06",
          1730 => x"52",
          1731 => x"80",
          1732 => x"b5",
          1733 => x"05",
          1734 => x"d4",
          1735 => x"08",
          1736 => x"12",
          1737 => x"bf",
          1738 => x"71",
          1739 => x"82",
          1740 => x"88",
          1741 => x"11",
          1742 => x"8c",
          1743 => x"b5",
          1744 => x"05",
          1745 => x"33",
          1746 => x"d4",
          1747 => x"0c",
          1748 => x"82",
          1749 => x"b5",
          1750 => x"05",
          1751 => x"33",
          1752 => x"70",
          1753 => x"51",
          1754 => x"80",
          1755 => x"38",
          1756 => x"08",
          1757 => x"70",
          1758 => x"82",
          1759 => x"fc",
          1760 => x"52",
          1761 => x"08",
          1762 => x"a9",
          1763 => x"d4",
          1764 => x"08",
          1765 => x"08",
          1766 => x"53",
          1767 => x"33",
          1768 => x"51",
          1769 => x"14",
          1770 => x"82",
          1771 => x"f8",
          1772 => x"d7",
          1773 => x"d4",
          1774 => x"08",
          1775 => x"05",
          1776 => x"81",
          1777 => x"b5",
          1778 => x"05",
          1779 => x"d4",
          1780 => x"08",
          1781 => x"08",
          1782 => x"2d",
          1783 => x"08",
          1784 => x"d4",
          1785 => x"0c",
          1786 => x"d4",
          1787 => x"08",
          1788 => x"f2",
          1789 => x"d4",
          1790 => x"08",
          1791 => x"08",
          1792 => x"82",
          1793 => x"88",
          1794 => x"11",
          1795 => x"d4",
          1796 => x"0c",
          1797 => x"d4",
          1798 => x"08",
          1799 => x"81",
          1800 => x"82",
          1801 => x"f0",
          1802 => x"07",
          1803 => x"b5",
          1804 => x"05",
          1805 => x"82",
          1806 => x"f0",
          1807 => x"07",
          1808 => x"b5",
          1809 => x"05",
          1810 => x"d4",
          1811 => x"08",
          1812 => x"d4",
          1813 => x"33",
          1814 => x"ff",
          1815 => x"d4",
          1816 => x"0c",
          1817 => x"b5",
          1818 => x"05",
          1819 => x"08",
          1820 => x"12",
          1821 => x"d4",
          1822 => x"08",
          1823 => x"06",
          1824 => x"d4",
          1825 => x"0c",
          1826 => x"82",
          1827 => x"f8",
          1828 => x"b5",
          1829 => x"3d",
          1830 => x"d4",
          1831 => x"b5",
          1832 => x"82",
          1833 => x"fd",
          1834 => x"b5",
          1835 => x"05",
          1836 => x"d4",
          1837 => x"0c",
          1838 => x"08",
          1839 => x"82",
          1840 => x"f8",
          1841 => x"b5",
          1842 => x"05",
          1843 => x"82",
          1844 => x"b5",
          1845 => x"05",
          1846 => x"d4",
          1847 => x"08",
          1848 => x"38",
          1849 => x"08",
          1850 => x"82",
          1851 => x"90",
          1852 => x"51",
          1853 => x"08",
          1854 => x"71",
          1855 => x"38",
          1856 => x"08",
          1857 => x"82",
          1858 => x"90",
          1859 => x"82",
          1860 => x"fc",
          1861 => x"b5",
          1862 => x"05",
          1863 => x"d4",
          1864 => x"08",
          1865 => x"d4",
          1866 => x"0c",
          1867 => x"08",
          1868 => x"81",
          1869 => x"d4",
          1870 => x"0c",
          1871 => x"08",
          1872 => x"ff",
          1873 => x"d4",
          1874 => x"0c",
          1875 => x"08",
          1876 => x"80",
          1877 => x"38",
          1878 => x"08",
          1879 => x"ff",
          1880 => x"d4",
          1881 => x"0c",
          1882 => x"08",
          1883 => x"ff",
          1884 => x"d4",
          1885 => x"0c",
          1886 => x"08",
          1887 => x"82",
          1888 => x"f8",
          1889 => x"51",
          1890 => x"34",
          1891 => x"82",
          1892 => x"90",
          1893 => x"05",
          1894 => x"08",
          1895 => x"82",
          1896 => x"90",
          1897 => x"05",
          1898 => x"08",
          1899 => x"82",
          1900 => x"90",
          1901 => x"2e",
          1902 => x"b5",
          1903 => x"05",
          1904 => x"33",
          1905 => x"08",
          1906 => x"81",
          1907 => x"d4",
          1908 => x"0c",
          1909 => x"08",
          1910 => x"52",
          1911 => x"34",
          1912 => x"08",
          1913 => x"81",
          1914 => x"d4",
          1915 => x"0c",
          1916 => x"82",
          1917 => x"88",
          1918 => x"82",
          1919 => x"51",
          1920 => x"82",
          1921 => x"04",
          1922 => x"08",
          1923 => x"d4",
          1924 => x"0d",
          1925 => x"08",
          1926 => x"82",
          1927 => x"fc",
          1928 => x"b5",
          1929 => x"05",
          1930 => x"33",
          1931 => x"08",
          1932 => x"81",
          1933 => x"d4",
          1934 => x"0c",
          1935 => x"06",
          1936 => x"80",
          1937 => x"da",
          1938 => x"d4",
          1939 => x"08",
          1940 => x"b5",
          1941 => x"05",
          1942 => x"d4",
          1943 => x"08",
          1944 => x"08",
          1945 => x"31",
          1946 => x"c8",
          1947 => x"3d",
          1948 => x"d4",
          1949 => x"b5",
          1950 => x"82",
          1951 => x"fe",
          1952 => x"b5",
          1953 => x"05",
          1954 => x"d4",
          1955 => x"0c",
          1956 => x"08",
          1957 => x"52",
          1958 => x"b5",
          1959 => x"05",
          1960 => x"82",
          1961 => x"8c",
          1962 => x"b5",
          1963 => x"05",
          1964 => x"70",
          1965 => x"b5",
          1966 => x"05",
          1967 => x"82",
          1968 => x"fc",
          1969 => x"81",
          1970 => x"70",
          1971 => x"38",
          1972 => x"82",
          1973 => x"88",
          1974 => x"82",
          1975 => x"51",
          1976 => x"82",
          1977 => x"04",
          1978 => x"08",
          1979 => x"d4",
          1980 => x"0d",
          1981 => x"08",
          1982 => x"82",
          1983 => x"fc",
          1984 => x"b5",
          1985 => x"05",
          1986 => x"d4",
          1987 => x"0c",
          1988 => x"08",
          1989 => x"80",
          1990 => x"38",
          1991 => x"08",
          1992 => x"81",
          1993 => x"d4",
          1994 => x"0c",
          1995 => x"08",
          1996 => x"ff",
          1997 => x"d4",
          1998 => x"0c",
          1999 => x"08",
          2000 => x"80",
          2001 => x"82",
          2002 => x"f8",
          2003 => x"70",
          2004 => x"d4",
          2005 => x"08",
          2006 => x"b5",
          2007 => x"05",
          2008 => x"d4",
          2009 => x"08",
          2010 => x"71",
          2011 => x"d4",
          2012 => x"08",
          2013 => x"b5",
          2014 => x"05",
          2015 => x"39",
          2016 => x"08",
          2017 => x"70",
          2018 => x"0c",
          2019 => x"0d",
          2020 => x"0c",
          2021 => x"d4",
          2022 => x"b5",
          2023 => x"3d",
          2024 => x"d4",
          2025 => x"08",
          2026 => x"f4",
          2027 => x"d4",
          2028 => x"08",
          2029 => x"82",
          2030 => x"8c",
          2031 => x"05",
          2032 => x"08",
          2033 => x"82",
          2034 => x"88",
          2035 => x"33",
          2036 => x"06",
          2037 => x"51",
          2038 => x"84",
          2039 => x"39",
          2040 => x"08",
          2041 => x"52",
          2042 => x"b5",
          2043 => x"05",
          2044 => x"82",
          2045 => x"88",
          2046 => x"81",
          2047 => x"51",
          2048 => x"80",
          2049 => x"d4",
          2050 => x"0c",
          2051 => x"82",
          2052 => x"90",
          2053 => x"05",
          2054 => x"08",
          2055 => x"82",
          2056 => x"90",
          2057 => x"2e",
          2058 => x"81",
          2059 => x"d4",
          2060 => x"08",
          2061 => x"e8",
          2062 => x"d4",
          2063 => x"08",
          2064 => x"53",
          2065 => x"ff",
          2066 => x"d4",
          2067 => x"0c",
          2068 => x"82",
          2069 => x"8c",
          2070 => x"05",
          2071 => x"08",
          2072 => x"82",
          2073 => x"8c",
          2074 => x"33",
          2075 => x"8c",
          2076 => x"82",
          2077 => x"fc",
          2078 => x"39",
          2079 => x"08",
          2080 => x"70",
          2081 => x"d4",
          2082 => x"08",
          2083 => x"71",
          2084 => x"b5",
          2085 => x"05",
          2086 => x"52",
          2087 => x"39",
          2088 => x"b5",
          2089 => x"05",
          2090 => x"d4",
          2091 => x"08",
          2092 => x"0c",
          2093 => x"82",
          2094 => x"04",
          2095 => x"08",
          2096 => x"d4",
          2097 => x"0d",
          2098 => x"08",
          2099 => x"82",
          2100 => x"f8",
          2101 => x"b5",
          2102 => x"05",
          2103 => x"80",
          2104 => x"d4",
          2105 => x"0c",
          2106 => x"82",
          2107 => x"f8",
          2108 => x"71",
          2109 => x"d4",
          2110 => x"08",
          2111 => x"b5",
          2112 => x"05",
          2113 => x"ff",
          2114 => x"70",
          2115 => x"38",
          2116 => x"08",
          2117 => x"ff",
          2118 => x"d4",
          2119 => x"0c",
          2120 => x"08",
          2121 => x"ff",
          2122 => x"ff",
          2123 => x"b5",
          2124 => x"05",
          2125 => x"82",
          2126 => x"f8",
          2127 => x"b5",
          2128 => x"05",
          2129 => x"d4",
          2130 => x"08",
          2131 => x"b5",
          2132 => x"05",
          2133 => x"b5",
          2134 => x"05",
          2135 => x"c8",
          2136 => x"0d",
          2137 => x"0c",
          2138 => x"d4",
          2139 => x"b5",
          2140 => x"3d",
          2141 => x"d4",
          2142 => x"08",
          2143 => x"08",
          2144 => x"82",
          2145 => x"90",
          2146 => x"2e",
          2147 => x"82",
          2148 => x"90",
          2149 => x"05",
          2150 => x"08",
          2151 => x"82",
          2152 => x"90",
          2153 => x"05",
          2154 => x"08",
          2155 => x"82",
          2156 => x"90",
          2157 => x"2e",
          2158 => x"b5",
          2159 => x"05",
          2160 => x"82",
          2161 => x"fc",
          2162 => x"52",
          2163 => x"82",
          2164 => x"fc",
          2165 => x"05",
          2166 => x"08",
          2167 => x"ff",
          2168 => x"b5",
          2169 => x"05",
          2170 => x"b5",
          2171 => x"84",
          2172 => x"b5",
          2173 => x"82",
          2174 => x"02",
          2175 => x"0c",
          2176 => x"80",
          2177 => x"d4",
          2178 => x"0c",
          2179 => x"08",
          2180 => x"80",
          2181 => x"82",
          2182 => x"88",
          2183 => x"82",
          2184 => x"88",
          2185 => x"0b",
          2186 => x"08",
          2187 => x"82",
          2188 => x"fc",
          2189 => x"38",
          2190 => x"b5",
          2191 => x"05",
          2192 => x"d4",
          2193 => x"08",
          2194 => x"08",
          2195 => x"82",
          2196 => x"8c",
          2197 => x"25",
          2198 => x"b5",
          2199 => x"05",
          2200 => x"b5",
          2201 => x"05",
          2202 => x"82",
          2203 => x"f0",
          2204 => x"b5",
          2205 => x"05",
          2206 => x"81",
          2207 => x"d4",
          2208 => x"0c",
          2209 => x"08",
          2210 => x"82",
          2211 => x"fc",
          2212 => x"53",
          2213 => x"08",
          2214 => x"52",
          2215 => x"08",
          2216 => x"51",
          2217 => x"82",
          2218 => x"70",
          2219 => x"08",
          2220 => x"54",
          2221 => x"08",
          2222 => x"80",
          2223 => x"82",
          2224 => x"f8",
          2225 => x"82",
          2226 => x"f8",
          2227 => x"b5",
          2228 => x"05",
          2229 => x"b5",
          2230 => x"89",
          2231 => x"b5",
          2232 => x"82",
          2233 => x"02",
          2234 => x"0c",
          2235 => x"80",
          2236 => x"d4",
          2237 => x"0c",
          2238 => x"08",
          2239 => x"80",
          2240 => x"82",
          2241 => x"88",
          2242 => x"82",
          2243 => x"88",
          2244 => x"0b",
          2245 => x"08",
          2246 => x"82",
          2247 => x"8c",
          2248 => x"25",
          2249 => x"b5",
          2250 => x"05",
          2251 => x"b5",
          2252 => x"05",
          2253 => x"82",
          2254 => x"8c",
          2255 => x"82",
          2256 => x"88",
          2257 => x"81",
          2258 => x"b5",
          2259 => x"82",
          2260 => x"f8",
          2261 => x"82",
          2262 => x"fc",
          2263 => x"2e",
          2264 => x"b5",
          2265 => x"05",
          2266 => x"b5",
          2267 => x"05",
          2268 => x"d4",
          2269 => x"08",
          2270 => x"c8",
          2271 => x"3d",
          2272 => x"d4",
          2273 => x"b5",
          2274 => x"82",
          2275 => x"fd",
          2276 => x"53",
          2277 => x"08",
          2278 => x"52",
          2279 => x"08",
          2280 => x"51",
          2281 => x"82",
          2282 => x"70",
          2283 => x"0c",
          2284 => x"0d",
          2285 => x"0c",
          2286 => x"d4",
          2287 => x"b5",
          2288 => x"3d",
          2289 => x"82",
          2290 => x"8c",
          2291 => x"82",
          2292 => x"88",
          2293 => x"93",
          2294 => x"c8",
          2295 => x"b5",
          2296 => x"85",
          2297 => x"b5",
          2298 => x"82",
          2299 => x"02",
          2300 => x"0c",
          2301 => x"81",
          2302 => x"d4",
          2303 => x"0c",
          2304 => x"b5",
          2305 => x"05",
          2306 => x"d4",
          2307 => x"08",
          2308 => x"08",
          2309 => x"27",
          2310 => x"b5",
          2311 => x"05",
          2312 => x"ae",
          2313 => x"82",
          2314 => x"8c",
          2315 => x"a2",
          2316 => x"d4",
          2317 => x"08",
          2318 => x"d4",
          2319 => x"0c",
          2320 => x"08",
          2321 => x"10",
          2322 => x"08",
          2323 => x"ff",
          2324 => x"b5",
          2325 => x"05",
          2326 => x"80",
          2327 => x"b5",
          2328 => x"05",
          2329 => x"d4",
          2330 => x"08",
          2331 => x"82",
          2332 => x"88",
          2333 => x"b5",
          2334 => x"05",
          2335 => x"b5",
          2336 => x"05",
          2337 => x"d4",
          2338 => x"08",
          2339 => x"08",
          2340 => x"07",
          2341 => x"08",
          2342 => x"82",
          2343 => x"fc",
          2344 => x"2a",
          2345 => x"08",
          2346 => x"82",
          2347 => x"8c",
          2348 => x"2a",
          2349 => x"08",
          2350 => x"ff",
          2351 => x"b5",
          2352 => x"05",
          2353 => x"93",
          2354 => x"d4",
          2355 => x"08",
          2356 => x"d4",
          2357 => x"0c",
          2358 => x"82",
          2359 => x"f8",
          2360 => x"82",
          2361 => x"f4",
          2362 => x"82",
          2363 => x"f4",
          2364 => x"b5",
          2365 => x"3d",
          2366 => x"d4",
          2367 => x"b5",
          2368 => x"82",
          2369 => x"f7",
          2370 => x"0b",
          2371 => x"08",
          2372 => x"82",
          2373 => x"8c",
          2374 => x"80",
          2375 => x"b5",
          2376 => x"05",
          2377 => x"51",
          2378 => x"53",
          2379 => x"d4",
          2380 => x"34",
          2381 => x"06",
          2382 => x"2e",
          2383 => x"91",
          2384 => x"d4",
          2385 => x"08",
          2386 => x"05",
          2387 => x"ce",
          2388 => x"d4",
          2389 => x"33",
          2390 => x"2e",
          2391 => x"a4",
          2392 => x"82",
          2393 => x"f0",
          2394 => x"b5",
          2395 => x"05",
          2396 => x"81",
          2397 => x"70",
          2398 => x"72",
          2399 => x"d4",
          2400 => x"34",
          2401 => x"08",
          2402 => x"53",
          2403 => x"09",
          2404 => x"dc",
          2405 => x"d4",
          2406 => x"08",
          2407 => x"05",
          2408 => x"08",
          2409 => x"33",
          2410 => x"08",
          2411 => x"82",
          2412 => x"f8",
          2413 => x"b5",
          2414 => x"05",
          2415 => x"d4",
          2416 => x"08",
          2417 => x"b6",
          2418 => x"d4",
          2419 => x"08",
          2420 => x"84",
          2421 => x"39",
          2422 => x"b5",
          2423 => x"05",
          2424 => x"d4",
          2425 => x"08",
          2426 => x"05",
          2427 => x"08",
          2428 => x"33",
          2429 => x"08",
          2430 => x"81",
          2431 => x"0b",
          2432 => x"08",
          2433 => x"82",
          2434 => x"88",
          2435 => x"08",
          2436 => x"0c",
          2437 => x"53",
          2438 => x"b5",
          2439 => x"05",
          2440 => x"39",
          2441 => x"08",
          2442 => x"53",
          2443 => x"8d",
          2444 => x"82",
          2445 => x"ec",
          2446 => x"80",
          2447 => x"d4",
          2448 => x"33",
          2449 => x"27",
          2450 => x"b5",
          2451 => x"05",
          2452 => x"b9",
          2453 => x"8d",
          2454 => x"82",
          2455 => x"ec",
          2456 => x"d8",
          2457 => x"82",
          2458 => x"f4",
          2459 => x"39",
          2460 => x"08",
          2461 => x"53",
          2462 => x"90",
          2463 => x"d4",
          2464 => x"33",
          2465 => x"26",
          2466 => x"39",
          2467 => x"b5",
          2468 => x"05",
          2469 => x"39",
          2470 => x"b5",
          2471 => x"05",
          2472 => x"82",
          2473 => x"fc",
          2474 => x"b5",
          2475 => x"05",
          2476 => x"73",
          2477 => x"38",
          2478 => x"08",
          2479 => x"53",
          2480 => x"27",
          2481 => x"b5",
          2482 => x"05",
          2483 => x"51",
          2484 => x"b5",
          2485 => x"05",
          2486 => x"d4",
          2487 => x"33",
          2488 => x"53",
          2489 => x"d4",
          2490 => x"34",
          2491 => x"08",
          2492 => x"53",
          2493 => x"ad",
          2494 => x"d4",
          2495 => x"33",
          2496 => x"53",
          2497 => x"d4",
          2498 => x"34",
          2499 => x"08",
          2500 => x"53",
          2501 => x"8d",
          2502 => x"82",
          2503 => x"ec",
          2504 => x"98",
          2505 => x"d4",
          2506 => x"33",
          2507 => x"08",
          2508 => x"54",
          2509 => x"26",
          2510 => x"0b",
          2511 => x"08",
          2512 => x"80",
          2513 => x"b5",
          2514 => x"05",
          2515 => x"b5",
          2516 => x"05",
          2517 => x"b5",
          2518 => x"05",
          2519 => x"82",
          2520 => x"fc",
          2521 => x"b5",
          2522 => x"05",
          2523 => x"81",
          2524 => x"70",
          2525 => x"52",
          2526 => x"33",
          2527 => x"08",
          2528 => x"fe",
          2529 => x"b5",
          2530 => x"05",
          2531 => x"80",
          2532 => x"82",
          2533 => x"fc",
          2534 => x"82",
          2535 => x"fc",
          2536 => x"b5",
          2537 => x"05",
          2538 => x"d4",
          2539 => x"08",
          2540 => x"81",
          2541 => x"d4",
          2542 => x"0c",
          2543 => x"08",
          2544 => x"82",
          2545 => x"8b",
          2546 => x"b5",
          2547 => x"82",
          2548 => x"02",
          2549 => x"0c",
          2550 => x"80",
          2551 => x"d4",
          2552 => x"34",
          2553 => x"08",
          2554 => x"53",
          2555 => x"82",
          2556 => x"88",
          2557 => x"08",
          2558 => x"33",
          2559 => x"b5",
          2560 => x"05",
          2561 => x"ff",
          2562 => x"a0",
          2563 => x"06",
          2564 => x"b5",
          2565 => x"05",
          2566 => x"81",
          2567 => x"53",
          2568 => x"b5",
          2569 => x"05",
          2570 => x"ad",
          2571 => x"06",
          2572 => x"0b",
          2573 => x"08",
          2574 => x"82",
          2575 => x"88",
          2576 => x"08",
          2577 => x"0c",
          2578 => x"53",
          2579 => x"b5",
          2580 => x"05",
          2581 => x"d4",
          2582 => x"33",
          2583 => x"2e",
          2584 => x"81",
          2585 => x"b5",
          2586 => x"05",
          2587 => x"81",
          2588 => x"70",
          2589 => x"72",
          2590 => x"d4",
          2591 => x"34",
          2592 => x"08",
          2593 => x"82",
          2594 => x"e8",
          2595 => x"b5",
          2596 => x"05",
          2597 => x"2e",
          2598 => x"b5",
          2599 => x"05",
          2600 => x"2e",
          2601 => x"cd",
          2602 => x"82",
          2603 => x"f4",
          2604 => x"b5",
          2605 => x"05",
          2606 => x"81",
          2607 => x"70",
          2608 => x"72",
          2609 => x"d4",
          2610 => x"34",
          2611 => x"82",
          2612 => x"d4",
          2613 => x"34",
          2614 => x"08",
          2615 => x"70",
          2616 => x"71",
          2617 => x"51",
          2618 => x"82",
          2619 => x"f8",
          2620 => x"fe",
          2621 => x"d4",
          2622 => x"33",
          2623 => x"26",
          2624 => x"0b",
          2625 => x"08",
          2626 => x"83",
          2627 => x"b5",
          2628 => x"05",
          2629 => x"73",
          2630 => x"82",
          2631 => x"f8",
          2632 => x"72",
          2633 => x"38",
          2634 => x"0b",
          2635 => x"08",
          2636 => x"82",
          2637 => x"0b",
          2638 => x"08",
          2639 => x"b2",
          2640 => x"d4",
          2641 => x"33",
          2642 => x"27",
          2643 => x"b5",
          2644 => x"05",
          2645 => x"b9",
          2646 => x"8d",
          2647 => x"82",
          2648 => x"ec",
          2649 => x"a5",
          2650 => x"82",
          2651 => x"f4",
          2652 => x"0b",
          2653 => x"08",
          2654 => x"82",
          2655 => x"f8",
          2656 => x"a0",
          2657 => x"cf",
          2658 => x"d4",
          2659 => x"33",
          2660 => x"73",
          2661 => x"82",
          2662 => x"f8",
          2663 => x"11",
          2664 => x"82",
          2665 => x"f8",
          2666 => x"b5",
          2667 => x"05",
          2668 => x"51",
          2669 => x"b5",
          2670 => x"05",
          2671 => x"d4",
          2672 => x"33",
          2673 => x"27",
          2674 => x"b5",
          2675 => x"05",
          2676 => x"51",
          2677 => x"b5",
          2678 => x"05",
          2679 => x"d4",
          2680 => x"33",
          2681 => x"26",
          2682 => x"0b",
          2683 => x"08",
          2684 => x"81",
          2685 => x"b5",
          2686 => x"05",
          2687 => x"d4",
          2688 => x"33",
          2689 => x"74",
          2690 => x"80",
          2691 => x"d4",
          2692 => x"0c",
          2693 => x"82",
          2694 => x"f4",
          2695 => x"82",
          2696 => x"fc",
          2697 => x"82",
          2698 => x"f8",
          2699 => x"12",
          2700 => x"08",
          2701 => x"82",
          2702 => x"88",
          2703 => x"08",
          2704 => x"0c",
          2705 => x"51",
          2706 => x"72",
          2707 => x"d4",
          2708 => x"34",
          2709 => x"82",
          2710 => x"f0",
          2711 => x"72",
          2712 => x"38",
          2713 => x"08",
          2714 => x"30",
          2715 => x"08",
          2716 => x"82",
          2717 => x"8c",
          2718 => x"b5",
          2719 => x"05",
          2720 => x"53",
          2721 => x"b5",
          2722 => x"05",
          2723 => x"d4",
          2724 => x"08",
          2725 => x"0c",
          2726 => x"82",
          2727 => x"04",
          2728 => x"79",
          2729 => x"56",
          2730 => x"80",
          2731 => x"38",
          2732 => x"08",
          2733 => x"3f",
          2734 => x"08",
          2735 => x"85",
          2736 => x"80",
          2737 => x"33",
          2738 => x"2e",
          2739 => x"86",
          2740 => x"55",
          2741 => x"57",
          2742 => x"82",
          2743 => x"70",
          2744 => x"e6",
          2745 => x"b5",
          2746 => x"74",
          2747 => x"51",
          2748 => x"82",
          2749 => x"8b",
          2750 => x"33",
          2751 => x"2e",
          2752 => x"81",
          2753 => x"ff",
          2754 => x"99",
          2755 => x"38",
          2756 => x"82",
          2757 => x"89",
          2758 => x"ff",
          2759 => x"52",
          2760 => x"81",
          2761 => x"84",
          2762 => x"a8",
          2763 => x"08",
          2764 => x"f4",
          2765 => x"39",
          2766 => x"51",
          2767 => x"82",
          2768 => x"80",
          2769 => x"9b",
          2770 => x"eb",
          2771 => x"b0",
          2772 => x"39",
          2773 => x"51",
          2774 => x"82",
          2775 => x"80",
          2776 => x"9b",
          2777 => x"cf",
          2778 => x"fc",
          2779 => x"39",
          2780 => x"51",
          2781 => x"82",
          2782 => x"bb",
          2783 => x"c8",
          2784 => x"82",
          2785 => x"af",
          2786 => x"84",
          2787 => x"82",
          2788 => x"a3",
          2789 => x"b4",
          2790 => x"82",
          2791 => x"97",
          2792 => x"dc",
          2793 => x"82",
          2794 => x"8b",
          2795 => x"8c",
          2796 => x"82",
          2797 => x"d8",
          2798 => x"3d",
          2799 => x"3d",
          2800 => x"56",
          2801 => x"e7",
          2802 => x"74",
          2803 => x"e8",
          2804 => x"39",
          2805 => x"74",
          2806 => x"3f",
          2807 => x"08",
          2808 => x"ef",
          2809 => x"b5",
          2810 => x"79",
          2811 => x"82",
          2812 => x"ff",
          2813 => x"87",
          2814 => x"ec",
          2815 => x"02",
          2816 => x"e3",
          2817 => x"57",
          2818 => x"30",
          2819 => x"73",
          2820 => x"59",
          2821 => x"77",
          2822 => x"83",
          2823 => x"74",
          2824 => x"81",
          2825 => x"55",
          2826 => x"81",
          2827 => x"53",
          2828 => x"3d",
          2829 => x"80",
          2830 => x"82",
          2831 => x"57",
          2832 => x"08",
          2833 => x"b5",
          2834 => x"c0",
          2835 => x"82",
          2836 => x"59",
          2837 => x"05",
          2838 => x"53",
          2839 => x"51",
          2840 => x"3f",
          2841 => x"08",
          2842 => x"c8",
          2843 => x"7a",
          2844 => x"2e",
          2845 => x"19",
          2846 => x"59",
          2847 => x"3d",
          2848 => x"81",
          2849 => x"76",
          2850 => x"07",
          2851 => x"30",
          2852 => x"72",
          2853 => x"51",
          2854 => x"2e",
          2855 => x"9e",
          2856 => x"c0",
          2857 => x"52",
          2858 => x"92",
          2859 => x"75",
          2860 => x"0c",
          2861 => x"04",
          2862 => x"7c",
          2863 => x"b7",
          2864 => x"59",
          2865 => x"53",
          2866 => x"51",
          2867 => x"82",
          2868 => x"a8",
          2869 => x"2e",
          2870 => x"81",
          2871 => x"9c",
          2872 => x"98",
          2873 => x"60",
          2874 => x"c8",
          2875 => x"7e",
          2876 => x"82",
          2877 => x"58",
          2878 => x"04",
          2879 => x"c8",
          2880 => x"0d",
          2881 => x"0d",
          2882 => x"02",
          2883 => x"cf",
          2884 => x"73",
          2885 => x"5f",
          2886 => x"5e",
          2887 => x"82",
          2888 => x"ff",
          2889 => x"82",
          2890 => x"ff",
          2891 => x"80",
          2892 => x"27",
          2893 => x"7b",
          2894 => x"38",
          2895 => x"a7",
          2896 => x"39",
          2897 => x"72",
          2898 => x"38",
          2899 => x"82",
          2900 => x"ff",
          2901 => x"89",
          2902 => x"ec",
          2903 => x"fb",
          2904 => x"55",
          2905 => x"74",
          2906 => x"7a",
          2907 => x"72",
          2908 => x"9e",
          2909 => x"b8",
          2910 => x"39",
          2911 => x"51",
          2912 => x"3f",
          2913 => x"a1",
          2914 => x"53",
          2915 => x"8e",
          2916 => x"52",
          2917 => x"51",
          2918 => x"3f",
          2919 => x"9e",
          2920 => x"b8",
          2921 => x"15",
          2922 => x"9c",
          2923 => x"51",
          2924 => x"fe",
          2925 => x"9f",
          2926 => x"b8",
          2927 => x"55",
          2928 => x"80",
          2929 => x"18",
          2930 => x"53",
          2931 => x"7a",
          2932 => x"81",
          2933 => x"9f",
          2934 => x"38",
          2935 => x"73",
          2936 => x"ff",
          2937 => x"72",
          2938 => x"38",
          2939 => x"26",
          2940 => x"cd",
          2941 => x"73",
          2942 => x"82",
          2943 => x"52",
          2944 => x"b1",
          2945 => x"55",
          2946 => x"82",
          2947 => x"d3",
          2948 => x"18",
          2949 => x"58",
          2950 => x"82",
          2951 => x"98",
          2952 => x"2c",
          2953 => x"a0",
          2954 => x"06",
          2955 => x"b5",
          2956 => x"c8",
          2957 => x"70",
          2958 => x"a0",
          2959 => x"72",
          2960 => x"30",
          2961 => x"73",
          2962 => x"51",
          2963 => x"57",
          2964 => x"73",
          2965 => x"76",
          2966 => x"81",
          2967 => x"80",
          2968 => x"7c",
          2969 => x"78",
          2970 => x"38",
          2971 => x"82",
          2972 => x"8f",
          2973 => x"fc",
          2974 => x"9b",
          2975 => x"9f",
          2976 => x"9f",
          2977 => x"ff",
          2978 => x"82",
          2979 => x"51",
          2980 => x"82",
          2981 => x"82",
          2982 => x"82",
          2983 => x"52",
          2984 => x"51",
          2985 => x"3f",
          2986 => x"84",
          2987 => x"3f",
          2988 => x"04",
          2989 => x"87",
          2990 => x"08",
          2991 => x"3f",
          2992 => x"8e",
          2993 => x"c8",
          2994 => x"3f",
          2995 => x"82",
          2996 => x"2a",
          2997 => x"51",
          2998 => x"2e",
          2999 => x"51",
          3000 => x"82",
          3001 => x"99",
          3002 => x"51",
          3003 => x"72",
          3004 => x"81",
          3005 => x"71",
          3006 => x"38",
          3007 => x"d2",
          3008 => x"f0",
          3009 => x"3f",
          3010 => x"c6",
          3011 => x"2a",
          3012 => x"51",
          3013 => x"2e",
          3014 => x"51",
          3015 => x"82",
          3016 => x"98",
          3017 => x"51",
          3018 => x"72",
          3019 => x"81",
          3020 => x"71",
          3021 => x"38",
          3022 => x"96",
          3023 => x"94",
          3024 => x"3f",
          3025 => x"8a",
          3026 => x"2a",
          3027 => x"51",
          3028 => x"2e",
          3029 => x"51",
          3030 => x"82",
          3031 => x"98",
          3032 => x"51",
          3033 => x"72",
          3034 => x"81",
          3035 => x"71",
          3036 => x"38",
          3037 => x"da",
          3038 => x"bc",
          3039 => x"3f",
          3040 => x"ce",
          3041 => x"2a",
          3042 => x"51",
          3043 => x"2e",
          3044 => x"51",
          3045 => x"82",
          3046 => x"97",
          3047 => x"51",
          3048 => x"72",
          3049 => x"81",
          3050 => x"71",
          3051 => x"38",
          3052 => x"9e",
          3053 => x"e4",
          3054 => x"3f",
          3055 => x"92",
          3056 => x"3f",
          3057 => x"04",
          3058 => x"77",
          3059 => x"a3",
          3060 => x"55",
          3061 => x"52",
          3062 => x"8d",
          3063 => x"82",
          3064 => x"54",
          3065 => x"81",
          3066 => x"a0",
          3067 => x"c8",
          3068 => x"8b",
          3069 => x"c8",
          3070 => x"82",
          3071 => x"07",
          3072 => x"71",
          3073 => x"54",
          3074 => x"82",
          3075 => x"0b",
          3076 => x"c4",
          3077 => x"81",
          3078 => x"06",
          3079 => x"cc",
          3080 => x"52",
          3081 => x"b2",
          3082 => x"b5",
          3083 => x"2e",
          3084 => x"b5",
          3085 => x"cf",
          3086 => x"39",
          3087 => x"51",
          3088 => x"3f",
          3089 => x"0b",
          3090 => x"34",
          3091 => x"b0",
          3092 => x"73",
          3093 => x"81",
          3094 => x"82",
          3095 => x"74",
          3096 => x"a9",
          3097 => x"0b",
          3098 => x"0c",
          3099 => x"04",
          3100 => x"80",
          3101 => x"cc",
          3102 => x"5d",
          3103 => x"51",
          3104 => x"3f",
          3105 => x"08",
          3106 => x"59",
          3107 => x"09",
          3108 => x"38",
          3109 => x"83",
          3110 => x"b8",
          3111 => x"dc",
          3112 => x"53",
          3113 => x"b6",
          3114 => x"f5",
          3115 => x"b5",
          3116 => x"2e",
          3117 => x"a1",
          3118 => x"a3",
          3119 => x"5f",
          3120 => x"f4",
          3121 => x"93",
          3122 => x"70",
          3123 => x"f8",
          3124 => x"fd",
          3125 => x"3d",
          3126 => x"51",
          3127 => x"82",
          3128 => x"90",
          3129 => x"2c",
          3130 => x"80",
          3131 => x"a3",
          3132 => x"c2",
          3133 => x"78",
          3134 => x"d2",
          3135 => x"24",
          3136 => x"80",
          3137 => x"38",
          3138 => x"80",
          3139 => x"d4",
          3140 => x"c0",
          3141 => x"38",
          3142 => x"24",
          3143 => x"78",
          3144 => x"8c",
          3145 => x"39",
          3146 => x"2e",
          3147 => x"78",
          3148 => x"92",
          3149 => x"c3",
          3150 => x"38",
          3151 => x"2e",
          3152 => x"8a",
          3153 => x"81",
          3154 => x"86",
          3155 => x"83",
          3156 => x"78",
          3157 => x"89",
          3158 => x"88",
          3159 => x"85",
          3160 => x"38",
          3161 => x"b4",
          3162 => x"11",
          3163 => x"05",
          3164 => x"3f",
          3165 => x"08",
          3166 => x"c5",
          3167 => x"fe",
          3168 => x"ff",
          3169 => x"ec",
          3170 => x"b5",
          3171 => x"2e",
          3172 => x"b4",
          3173 => x"11",
          3174 => x"05",
          3175 => x"3f",
          3176 => x"08",
          3177 => x"b5",
          3178 => x"82",
          3179 => x"ff",
          3180 => x"63",
          3181 => x"79",
          3182 => x"ec",
          3183 => x"78",
          3184 => x"05",
          3185 => x"7a",
          3186 => x"81",
          3187 => x"3d",
          3188 => x"53",
          3189 => x"51",
          3190 => x"82",
          3191 => x"80",
          3192 => x"38",
          3193 => x"fc",
          3194 => x"84",
          3195 => x"df",
          3196 => x"c8",
          3197 => x"fd",
          3198 => x"3d",
          3199 => x"53",
          3200 => x"51",
          3201 => x"82",
          3202 => x"80",
          3203 => x"38",
          3204 => x"51",
          3205 => x"3f",
          3206 => x"63",
          3207 => x"38",
          3208 => x"70",
          3209 => x"33",
          3210 => x"81",
          3211 => x"39",
          3212 => x"80",
          3213 => x"84",
          3214 => x"93",
          3215 => x"c8",
          3216 => x"fc",
          3217 => x"3d",
          3218 => x"53",
          3219 => x"51",
          3220 => x"82",
          3221 => x"80",
          3222 => x"38",
          3223 => x"f8",
          3224 => x"84",
          3225 => x"e7",
          3226 => x"c8",
          3227 => x"fc",
          3228 => x"a2",
          3229 => x"ae",
          3230 => x"5a",
          3231 => x"a8",
          3232 => x"33",
          3233 => x"5a",
          3234 => x"2e",
          3235 => x"55",
          3236 => x"33",
          3237 => x"82",
          3238 => x"ff",
          3239 => x"81",
          3240 => x"05",
          3241 => x"39",
          3242 => x"dc",
          3243 => x"39",
          3244 => x"80",
          3245 => x"84",
          3246 => x"93",
          3247 => x"c8",
          3248 => x"38",
          3249 => x"33",
          3250 => x"2e",
          3251 => x"b3",
          3252 => x"80",
          3253 => x"b4",
          3254 => x"78",
          3255 => x"38",
          3256 => x"08",
          3257 => x"82",
          3258 => x"59",
          3259 => x"88",
          3260 => x"fc",
          3261 => x"39",
          3262 => x"33",
          3263 => x"2e",
          3264 => x"b4",
          3265 => x"9a",
          3266 => x"b2",
          3267 => x"80",
          3268 => x"82",
          3269 => x"44",
          3270 => x"b4",
          3271 => x"80",
          3272 => x"3d",
          3273 => x"53",
          3274 => x"51",
          3275 => x"82",
          3276 => x"80",
          3277 => x"b4",
          3278 => x"78",
          3279 => x"38",
          3280 => x"08",
          3281 => x"39",
          3282 => x"33",
          3283 => x"2e",
          3284 => x"b3",
          3285 => x"bb",
          3286 => x"b6",
          3287 => x"80",
          3288 => x"82",
          3289 => x"43",
          3290 => x"b4",
          3291 => x"78",
          3292 => x"38",
          3293 => x"08",
          3294 => x"82",
          3295 => x"59",
          3296 => x"88",
          3297 => x"90",
          3298 => x"39",
          3299 => x"08",
          3300 => x"b4",
          3301 => x"11",
          3302 => x"05",
          3303 => x"3f",
          3304 => x"08",
          3305 => x"38",
          3306 => x"5c",
          3307 => x"83",
          3308 => x"7a",
          3309 => x"30",
          3310 => x"9f",
          3311 => x"06",
          3312 => x"5a",
          3313 => x"88",
          3314 => x"2e",
          3315 => x"42",
          3316 => x"51",
          3317 => x"a0",
          3318 => x"61",
          3319 => x"63",
          3320 => x"3f",
          3321 => x"51",
          3322 => x"b4",
          3323 => x"11",
          3324 => x"05",
          3325 => x"3f",
          3326 => x"08",
          3327 => x"c1",
          3328 => x"fe",
          3329 => x"ff",
          3330 => x"e7",
          3331 => x"b5",
          3332 => x"2e",
          3333 => x"59",
          3334 => x"05",
          3335 => x"63",
          3336 => x"b4",
          3337 => x"11",
          3338 => x"05",
          3339 => x"3f",
          3340 => x"08",
          3341 => x"89",
          3342 => x"33",
          3343 => x"a2",
          3344 => x"ab",
          3345 => x"cd",
          3346 => x"80",
          3347 => x"51",
          3348 => x"3f",
          3349 => x"33",
          3350 => x"2e",
          3351 => x"9f",
          3352 => x"38",
          3353 => x"fc",
          3354 => x"84",
          3355 => x"df",
          3356 => x"c8",
          3357 => x"91",
          3358 => x"02",
          3359 => x"33",
          3360 => x"81",
          3361 => x"b1",
          3362 => x"e4",
          3363 => x"3f",
          3364 => x"b4",
          3365 => x"11",
          3366 => x"05",
          3367 => x"3f",
          3368 => x"08",
          3369 => x"99",
          3370 => x"fe",
          3371 => x"ff",
          3372 => x"e0",
          3373 => x"b5",
          3374 => x"2e",
          3375 => x"59",
          3376 => x"22",
          3377 => x"05",
          3378 => x"41",
          3379 => x"f0",
          3380 => x"84",
          3381 => x"a6",
          3382 => x"c8",
          3383 => x"f7",
          3384 => x"70",
          3385 => x"82",
          3386 => x"ff",
          3387 => x"82",
          3388 => x"53",
          3389 => x"79",
          3390 => x"b4",
          3391 => x"79",
          3392 => x"ae",
          3393 => x"38",
          3394 => x"87",
          3395 => x"05",
          3396 => x"b4",
          3397 => x"11",
          3398 => x"05",
          3399 => x"3f",
          3400 => x"08",
          3401 => x"38",
          3402 => x"be",
          3403 => x"70",
          3404 => x"23",
          3405 => x"aa",
          3406 => x"e4",
          3407 => x"3f",
          3408 => x"b4",
          3409 => x"11",
          3410 => x"05",
          3411 => x"3f",
          3412 => x"08",
          3413 => x"e9",
          3414 => x"fe",
          3415 => x"ff",
          3416 => x"df",
          3417 => x"b5",
          3418 => x"2e",
          3419 => x"60",
          3420 => x"60",
          3421 => x"b4",
          3422 => x"11",
          3423 => x"05",
          3424 => x"3f",
          3425 => x"08",
          3426 => x"b5",
          3427 => x"08",
          3428 => x"a2",
          3429 => x"a8",
          3430 => x"cd",
          3431 => x"80",
          3432 => x"51",
          3433 => x"3f",
          3434 => x"33",
          3435 => x"2e",
          3436 => x"9f",
          3437 => x"38",
          3438 => x"f0",
          3439 => x"84",
          3440 => x"ba",
          3441 => x"c8",
          3442 => x"8d",
          3443 => x"71",
          3444 => x"84",
          3445 => x"b5",
          3446 => x"e4",
          3447 => x"3f",
          3448 => x"b4",
          3449 => x"11",
          3450 => x"05",
          3451 => x"3f",
          3452 => x"08",
          3453 => x"c9",
          3454 => x"82",
          3455 => x"ff",
          3456 => x"63",
          3457 => x"b4",
          3458 => x"11",
          3459 => x"05",
          3460 => x"3f",
          3461 => x"08",
          3462 => x"a5",
          3463 => x"82",
          3464 => x"ff",
          3465 => x"63",
          3466 => x"82",
          3467 => x"80",
          3468 => x"38",
          3469 => x"08",
          3470 => x"bc",
          3471 => x"9b",
          3472 => x"39",
          3473 => x"51",
          3474 => x"ff",
          3475 => x"f4",
          3476 => x"a3",
          3477 => x"8e",
          3478 => x"ff",
          3479 => x"a7",
          3480 => x"39",
          3481 => x"33",
          3482 => x"2e",
          3483 => x"7d",
          3484 => x"78",
          3485 => x"cf",
          3486 => x"ff",
          3487 => x"83",
          3488 => x"b5",
          3489 => x"81",
          3490 => x"2e",
          3491 => x"82",
          3492 => x"7a",
          3493 => x"38",
          3494 => x"7a",
          3495 => x"38",
          3496 => x"82",
          3497 => x"7b",
          3498 => x"8c",
          3499 => x"82",
          3500 => x"b4",
          3501 => x"05",
          3502 => x"87",
          3503 => x"7b",
          3504 => x"ff",
          3505 => x"cf",
          3506 => x"39",
          3507 => x"a4",
          3508 => x"53",
          3509 => x"52",
          3510 => x"b0",
          3511 => x"a8",
          3512 => x"39",
          3513 => x"53",
          3514 => x"52",
          3515 => x"b0",
          3516 => x"a8",
          3517 => x"b3",
          3518 => x"b5",
          3519 => x"56",
          3520 => x"54",
          3521 => x"53",
          3522 => x"52",
          3523 => x"b0",
          3524 => x"a4",
          3525 => x"c8",
          3526 => x"c8",
          3527 => x"30",
          3528 => x"80",
          3529 => x"5b",
          3530 => x"7a",
          3531 => x"38",
          3532 => x"7a",
          3533 => x"80",
          3534 => x"81",
          3535 => x"ff",
          3536 => x"7a",
          3537 => x"7d",
          3538 => x"81",
          3539 => x"78",
          3540 => x"ff",
          3541 => x"06",
          3542 => x"82",
          3543 => x"c1",
          3544 => x"dd",
          3545 => x"0d",
          3546 => x"b5",
          3547 => x"c0",
          3548 => x"08",
          3549 => x"84",
          3550 => x"51",
          3551 => x"82",
          3552 => x"90",
          3553 => x"55",
          3554 => x"80",
          3555 => x"d7",
          3556 => x"82",
          3557 => x"07",
          3558 => x"c0",
          3559 => x"08",
          3560 => x"84",
          3561 => x"51",
          3562 => x"82",
          3563 => x"90",
          3564 => x"55",
          3565 => x"80",
          3566 => x"d7",
          3567 => x"82",
          3568 => x"07",
          3569 => x"80",
          3570 => x"c0",
          3571 => x"8c",
          3572 => x"87",
          3573 => x"0c",
          3574 => x"5a",
          3575 => x"5b",
          3576 => x"05",
          3577 => x"80",
          3578 => x"98",
          3579 => x"70",
          3580 => x"70",
          3581 => x"cd",
          3582 => x"89",
          3583 => x"81",
          3584 => x"c4",
          3585 => x"de",
          3586 => x"d0",
          3587 => x"d6",
          3588 => x"b1",
          3589 => x"3f",
          3590 => x"db",
          3591 => x"3f",
          3592 => x"3d",
          3593 => x"83",
          3594 => x"2b",
          3595 => x"3f",
          3596 => x"08",
          3597 => x"72",
          3598 => x"54",
          3599 => x"25",
          3600 => x"82",
          3601 => x"84",
          3602 => x"fc",
          3603 => x"70",
          3604 => x"80",
          3605 => x"72",
          3606 => x"8a",
          3607 => x"51",
          3608 => x"09",
          3609 => x"38",
          3610 => x"f1",
          3611 => x"51",
          3612 => x"09",
          3613 => x"38",
          3614 => x"81",
          3615 => x"73",
          3616 => x"81",
          3617 => x"84",
          3618 => x"52",
          3619 => x"52",
          3620 => x"2e",
          3621 => x"54",
          3622 => x"9d",
          3623 => x"38",
          3624 => x"12",
          3625 => x"33",
          3626 => x"a0",
          3627 => x"81",
          3628 => x"2e",
          3629 => x"ea",
          3630 => x"33",
          3631 => x"a0",
          3632 => x"06",
          3633 => x"54",
          3634 => x"70",
          3635 => x"25",
          3636 => x"51",
          3637 => x"2e",
          3638 => x"72",
          3639 => x"54",
          3640 => x"0c",
          3641 => x"82",
          3642 => x"86",
          3643 => x"fc",
          3644 => x"53",
          3645 => x"2e",
          3646 => x"3d",
          3647 => x"72",
          3648 => x"3f",
          3649 => x"08",
          3650 => x"53",
          3651 => x"53",
          3652 => x"c8",
          3653 => x"0d",
          3654 => x"0d",
          3655 => x"33",
          3656 => x"53",
          3657 => x"8b",
          3658 => x"38",
          3659 => x"ff",
          3660 => x"52",
          3661 => x"81",
          3662 => x"13",
          3663 => x"52",
          3664 => x"80",
          3665 => x"13",
          3666 => x"52",
          3667 => x"80",
          3668 => x"13",
          3669 => x"52",
          3670 => x"80",
          3671 => x"13",
          3672 => x"52",
          3673 => x"26",
          3674 => x"8a",
          3675 => x"87",
          3676 => x"e7",
          3677 => x"38",
          3678 => x"c0",
          3679 => x"72",
          3680 => x"98",
          3681 => x"13",
          3682 => x"98",
          3683 => x"13",
          3684 => x"98",
          3685 => x"13",
          3686 => x"98",
          3687 => x"13",
          3688 => x"98",
          3689 => x"13",
          3690 => x"98",
          3691 => x"87",
          3692 => x"0c",
          3693 => x"98",
          3694 => x"0b",
          3695 => x"9c",
          3696 => x"71",
          3697 => x"0c",
          3698 => x"04",
          3699 => x"7f",
          3700 => x"98",
          3701 => x"7d",
          3702 => x"98",
          3703 => x"7d",
          3704 => x"c0",
          3705 => x"5a",
          3706 => x"34",
          3707 => x"b4",
          3708 => x"83",
          3709 => x"c0",
          3710 => x"5a",
          3711 => x"34",
          3712 => x"ac",
          3713 => x"85",
          3714 => x"c0",
          3715 => x"5a",
          3716 => x"34",
          3717 => x"a4",
          3718 => x"88",
          3719 => x"c0",
          3720 => x"5a",
          3721 => x"23",
          3722 => x"79",
          3723 => x"06",
          3724 => x"ff",
          3725 => x"86",
          3726 => x"85",
          3727 => x"84",
          3728 => x"83",
          3729 => x"82",
          3730 => x"7d",
          3731 => x"06",
          3732 => x"e8",
          3733 => x"83",
          3734 => x"0d",
          3735 => x"0d",
          3736 => x"33",
          3737 => x"33",
          3738 => x"06",
          3739 => x"87",
          3740 => x"51",
          3741 => x"86",
          3742 => x"94",
          3743 => x"08",
          3744 => x"70",
          3745 => x"54",
          3746 => x"2e",
          3747 => x"91",
          3748 => x"06",
          3749 => x"d7",
          3750 => x"32",
          3751 => x"51",
          3752 => x"2e",
          3753 => x"93",
          3754 => x"06",
          3755 => x"ff",
          3756 => x"81",
          3757 => x"87",
          3758 => x"52",
          3759 => x"86",
          3760 => x"94",
          3761 => x"72",
          3762 => x"b5",
          3763 => x"3d",
          3764 => x"3d",
          3765 => x"05",
          3766 => x"70",
          3767 => x"52",
          3768 => x"b3",
          3769 => x"3d",
          3770 => x"3d",
          3771 => x"05",
          3772 => x"8a",
          3773 => x"06",
          3774 => x"52",
          3775 => x"3f",
          3776 => x"33",
          3777 => x"06",
          3778 => x"c0",
          3779 => x"76",
          3780 => x"38",
          3781 => x"94",
          3782 => x"70",
          3783 => x"81",
          3784 => x"54",
          3785 => x"8c",
          3786 => x"2a",
          3787 => x"51",
          3788 => x"38",
          3789 => x"70",
          3790 => x"53",
          3791 => x"8d",
          3792 => x"2a",
          3793 => x"51",
          3794 => x"be",
          3795 => x"ff",
          3796 => x"c0",
          3797 => x"72",
          3798 => x"38",
          3799 => x"90",
          3800 => x"0c",
          3801 => x"b5",
          3802 => x"3d",
          3803 => x"3d",
          3804 => x"80",
          3805 => x"81",
          3806 => x"53",
          3807 => x"2e",
          3808 => x"71",
          3809 => x"81",
          3810 => x"e8",
          3811 => x"ff",
          3812 => x"55",
          3813 => x"94",
          3814 => x"80",
          3815 => x"87",
          3816 => x"51",
          3817 => x"96",
          3818 => x"06",
          3819 => x"70",
          3820 => x"38",
          3821 => x"70",
          3822 => x"51",
          3823 => x"72",
          3824 => x"81",
          3825 => x"70",
          3826 => x"38",
          3827 => x"70",
          3828 => x"51",
          3829 => x"38",
          3830 => x"06",
          3831 => x"94",
          3832 => x"80",
          3833 => x"87",
          3834 => x"52",
          3835 => x"81",
          3836 => x"70",
          3837 => x"53",
          3838 => x"ff",
          3839 => x"82",
          3840 => x"89",
          3841 => x"fe",
          3842 => x"b3",
          3843 => x"81",
          3844 => x"52",
          3845 => x"84",
          3846 => x"2e",
          3847 => x"c0",
          3848 => x"70",
          3849 => x"2a",
          3850 => x"51",
          3851 => x"80",
          3852 => x"71",
          3853 => x"51",
          3854 => x"80",
          3855 => x"2e",
          3856 => x"c0",
          3857 => x"71",
          3858 => x"ff",
          3859 => x"c8",
          3860 => x"3d",
          3861 => x"af",
          3862 => x"c8",
          3863 => x"06",
          3864 => x"0c",
          3865 => x"0d",
          3866 => x"33",
          3867 => x"06",
          3868 => x"c0",
          3869 => x"70",
          3870 => x"38",
          3871 => x"94",
          3872 => x"70",
          3873 => x"81",
          3874 => x"51",
          3875 => x"80",
          3876 => x"72",
          3877 => x"51",
          3878 => x"80",
          3879 => x"2e",
          3880 => x"c0",
          3881 => x"71",
          3882 => x"2b",
          3883 => x"51",
          3884 => x"82",
          3885 => x"84",
          3886 => x"ff",
          3887 => x"c0",
          3888 => x"70",
          3889 => x"06",
          3890 => x"80",
          3891 => x"38",
          3892 => x"a4",
          3893 => x"ec",
          3894 => x"9e",
          3895 => x"b3",
          3896 => x"c0",
          3897 => x"82",
          3898 => x"87",
          3899 => x"08",
          3900 => x"0c",
          3901 => x"9c",
          3902 => x"fc",
          3903 => x"9e",
          3904 => x"b4",
          3905 => x"c0",
          3906 => x"82",
          3907 => x"87",
          3908 => x"08",
          3909 => x"0c",
          3910 => x"b4",
          3911 => x"8c",
          3912 => x"9e",
          3913 => x"b4",
          3914 => x"c0",
          3915 => x"82",
          3916 => x"87",
          3917 => x"08",
          3918 => x"0c",
          3919 => x"c4",
          3920 => x"9c",
          3921 => x"9e",
          3922 => x"70",
          3923 => x"23",
          3924 => x"84",
          3925 => x"a4",
          3926 => x"9e",
          3927 => x"b4",
          3928 => x"c0",
          3929 => x"82",
          3930 => x"81",
          3931 => x"b0",
          3932 => x"87",
          3933 => x"08",
          3934 => x"0a",
          3935 => x"52",
          3936 => x"83",
          3937 => x"71",
          3938 => x"34",
          3939 => x"c0",
          3940 => x"70",
          3941 => x"06",
          3942 => x"70",
          3943 => x"38",
          3944 => x"82",
          3945 => x"80",
          3946 => x"9e",
          3947 => x"90",
          3948 => x"51",
          3949 => x"80",
          3950 => x"81",
          3951 => x"b4",
          3952 => x"0b",
          3953 => x"90",
          3954 => x"80",
          3955 => x"52",
          3956 => x"2e",
          3957 => x"52",
          3958 => x"b4",
          3959 => x"87",
          3960 => x"08",
          3961 => x"80",
          3962 => x"52",
          3963 => x"83",
          3964 => x"71",
          3965 => x"34",
          3966 => x"c0",
          3967 => x"70",
          3968 => x"06",
          3969 => x"70",
          3970 => x"38",
          3971 => x"82",
          3972 => x"80",
          3973 => x"9e",
          3974 => x"84",
          3975 => x"51",
          3976 => x"80",
          3977 => x"81",
          3978 => x"b4",
          3979 => x"0b",
          3980 => x"90",
          3981 => x"80",
          3982 => x"52",
          3983 => x"2e",
          3984 => x"52",
          3985 => x"b8",
          3986 => x"87",
          3987 => x"08",
          3988 => x"80",
          3989 => x"52",
          3990 => x"83",
          3991 => x"71",
          3992 => x"34",
          3993 => x"c0",
          3994 => x"70",
          3995 => x"06",
          3996 => x"70",
          3997 => x"38",
          3998 => x"82",
          3999 => x"80",
          4000 => x"9e",
          4001 => x"a0",
          4002 => x"52",
          4003 => x"2e",
          4004 => x"52",
          4005 => x"bb",
          4006 => x"9e",
          4007 => x"98",
          4008 => x"8a",
          4009 => x"51",
          4010 => x"bc",
          4011 => x"87",
          4012 => x"08",
          4013 => x"06",
          4014 => x"70",
          4015 => x"38",
          4016 => x"82",
          4017 => x"87",
          4018 => x"08",
          4019 => x"06",
          4020 => x"51",
          4021 => x"82",
          4022 => x"80",
          4023 => x"9e",
          4024 => x"88",
          4025 => x"52",
          4026 => x"83",
          4027 => x"71",
          4028 => x"34",
          4029 => x"90",
          4030 => x"06",
          4031 => x"82",
          4032 => x"83",
          4033 => x"fb",
          4034 => x"a5",
          4035 => x"b1",
          4036 => x"b4",
          4037 => x"73",
          4038 => x"38",
          4039 => x"51",
          4040 => x"3f",
          4041 => x"51",
          4042 => x"3f",
          4043 => x"33",
          4044 => x"2e",
          4045 => x"b4",
          4046 => x"b4",
          4047 => x"54",
          4048 => x"c0",
          4049 => x"93",
          4050 => x"b7",
          4051 => x"80",
          4052 => x"82",
          4053 => x"82",
          4054 => x"11",
          4055 => x"a5",
          4056 => x"94",
          4057 => x"b4",
          4058 => x"73",
          4059 => x"38",
          4060 => x"08",
          4061 => x"08",
          4062 => x"82",
          4063 => x"ff",
          4064 => x"82",
          4065 => x"54",
          4066 => x"94",
          4067 => x"f4",
          4068 => x"f8",
          4069 => x"52",
          4070 => x"51",
          4071 => x"3f",
          4072 => x"33",
          4073 => x"2e",
          4074 => x"b3",
          4075 => x"b4",
          4076 => x"54",
          4077 => x"b0",
          4078 => x"9f",
          4079 => x"bb",
          4080 => x"80",
          4081 => x"82",
          4082 => x"52",
          4083 => x"51",
          4084 => x"3f",
          4085 => x"33",
          4086 => x"2e",
          4087 => x"b4",
          4088 => x"82",
          4089 => x"ff",
          4090 => x"82",
          4091 => x"54",
          4092 => x"8e",
          4093 => x"be",
          4094 => x"a7",
          4095 => x"93",
          4096 => x"b4",
          4097 => x"73",
          4098 => x"38",
          4099 => x"51",
          4100 => x"3f",
          4101 => x"33",
          4102 => x"2e",
          4103 => x"a7",
          4104 => x"af",
          4105 => x"b4",
          4106 => x"73",
          4107 => x"38",
          4108 => x"51",
          4109 => x"3f",
          4110 => x"33",
          4111 => x"2e",
          4112 => x"a7",
          4113 => x"af",
          4114 => x"b4",
          4115 => x"73",
          4116 => x"38",
          4117 => x"51",
          4118 => x"3f",
          4119 => x"51",
          4120 => x"3f",
          4121 => x"08",
          4122 => x"fc",
          4123 => x"eb",
          4124 => x"98",
          4125 => x"a8",
          4126 => x"92",
          4127 => x"b4",
          4128 => x"82",
          4129 => x"ff",
          4130 => x"82",
          4131 => x"ff",
          4132 => x"82",
          4133 => x"52",
          4134 => x"51",
          4135 => x"3f",
          4136 => x"08",
          4137 => x"c0",
          4138 => x"c5",
          4139 => x"b5",
          4140 => x"84",
          4141 => x"71",
          4142 => x"82",
          4143 => x"52",
          4144 => x"51",
          4145 => x"3f",
          4146 => x"33",
          4147 => x"2e",
          4148 => x"b4",
          4149 => x"bd",
          4150 => x"75",
          4151 => x"3f",
          4152 => x"08",
          4153 => x"29",
          4154 => x"54",
          4155 => x"c8",
          4156 => x"a9",
          4157 => x"91",
          4158 => x"b4",
          4159 => x"73",
          4160 => x"38",
          4161 => x"08",
          4162 => x"c0",
          4163 => x"c4",
          4164 => x"b5",
          4165 => x"84",
          4166 => x"71",
          4167 => x"82",
          4168 => x"52",
          4169 => x"51",
          4170 => x"3f",
          4171 => x"51",
          4172 => x"3f",
          4173 => x"04",
          4174 => x"02",
          4175 => x"ff",
          4176 => x"84",
          4177 => x"71",
          4178 => x"95",
          4179 => x"71",
          4180 => x"aa",
          4181 => x"39",
          4182 => x"51",
          4183 => x"aa",
          4184 => x"39",
          4185 => x"51",
          4186 => x"aa",
          4187 => x"39",
          4188 => x"51",
          4189 => x"3f",
          4190 => x"04",
          4191 => x"0c",
          4192 => x"87",
          4193 => x"0c",
          4194 => x"c4",
          4195 => x"96",
          4196 => x"fd",
          4197 => x"98",
          4198 => x"2c",
          4199 => x"70",
          4200 => x"10",
          4201 => x"2b",
          4202 => x"54",
          4203 => x"0b",
          4204 => x"12",
          4205 => x"71",
          4206 => x"38",
          4207 => x"11",
          4208 => x"84",
          4209 => x"33",
          4210 => x"52",
          4211 => x"2e",
          4212 => x"83",
          4213 => x"72",
          4214 => x"0c",
          4215 => x"04",
          4216 => x"79",
          4217 => x"a3",
          4218 => x"33",
          4219 => x"72",
          4220 => x"38",
          4221 => x"08",
          4222 => x"ff",
          4223 => x"82",
          4224 => x"52",
          4225 => x"af",
          4226 => x"cd",
          4227 => x"88",
          4228 => x"a1",
          4229 => x"ff",
          4230 => x"74",
          4231 => x"ff",
          4232 => x"39",
          4233 => x"8f",
          4234 => x"74",
          4235 => x"0d",
          4236 => x"0d",
          4237 => x"05",
          4238 => x"02",
          4239 => x"05",
          4240 => x"a0",
          4241 => x"29",
          4242 => x"05",
          4243 => x"59",
          4244 => x"59",
          4245 => x"86",
          4246 => x"9a",
          4247 => x"b5",
          4248 => x"84",
          4249 => x"c8",
          4250 => x"70",
          4251 => x"5a",
          4252 => x"82",
          4253 => x"75",
          4254 => x"a0",
          4255 => x"29",
          4256 => x"05",
          4257 => x"56",
          4258 => x"2e",
          4259 => x"53",
          4260 => x"51",
          4261 => x"3f",
          4262 => x"33",
          4263 => x"74",
          4264 => x"34",
          4265 => x"06",
          4266 => x"27",
          4267 => x"0b",
          4268 => x"34",
          4269 => x"b6",
          4270 => x"9c",
          4271 => x"80",
          4272 => x"82",
          4273 => x"55",
          4274 => x"8c",
          4275 => x"54",
          4276 => x"52",
          4277 => x"da",
          4278 => x"b5",
          4279 => x"8a",
          4280 => x"95",
          4281 => x"9c",
          4282 => x"dd",
          4283 => x"3d",
          4284 => x"3d",
          4285 => x"c8",
          4286 => x"72",
          4287 => x"80",
          4288 => x"71",
          4289 => x"3f",
          4290 => x"ff",
          4291 => x"54",
          4292 => x"25",
          4293 => x"0b",
          4294 => x"34",
          4295 => x"08",
          4296 => x"2e",
          4297 => x"51",
          4298 => x"3f",
          4299 => x"08",
          4300 => x"3f",
          4301 => x"b5",
          4302 => x"3d",
          4303 => x"3d",
          4304 => x"80",
          4305 => x"9c",
          4306 => x"e3",
          4307 => x"b5",
          4308 => x"d3",
          4309 => x"9c",
          4310 => x"f8",
          4311 => x"70",
          4312 => x"8c",
          4313 => x"b5",
          4314 => x"2e",
          4315 => x"51",
          4316 => x"3f",
          4317 => x"08",
          4318 => x"82",
          4319 => x"25",
          4320 => x"b5",
          4321 => x"05",
          4322 => x"55",
          4323 => x"75",
          4324 => x"81",
          4325 => x"c8",
          4326 => x"8c",
          4327 => x"ff",
          4328 => x"06",
          4329 => x"a6",
          4330 => x"d9",
          4331 => x"3d",
          4332 => x"08",
          4333 => x"70",
          4334 => x"52",
          4335 => x"08",
          4336 => x"bb",
          4337 => x"c8",
          4338 => x"38",
          4339 => x"b5",
          4340 => x"55",
          4341 => x"8b",
          4342 => x"56",
          4343 => x"3f",
          4344 => x"08",
          4345 => x"38",
          4346 => x"b4",
          4347 => x"b5",
          4348 => x"18",
          4349 => x"0b",
          4350 => x"08",
          4351 => x"82",
          4352 => x"ff",
          4353 => x"55",
          4354 => x"34",
          4355 => x"30",
          4356 => x"9f",
          4357 => x"55",
          4358 => x"85",
          4359 => x"ac",
          4360 => x"9c",
          4361 => x"08",
          4362 => x"e1",
          4363 => x"b5",
          4364 => x"2e",
          4365 => x"ad",
          4366 => x"8b",
          4367 => x"77",
          4368 => x"06",
          4369 => x"52",
          4370 => x"b4",
          4371 => x"51",
          4372 => x"3f",
          4373 => x"54",
          4374 => x"08",
          4375 => x"58",
          4376 => x"c8",
          4377 => x"0d",
          4378 => x"0d",
          4379 => x"5c",
          4380 => x"57",
          4381 => x"73",
          4382 => x"81",
          4383 => x"78",
          4384 => x"56",
          4385 => x"98",
          4386 => x"70",
          4387 => x"33",
          4388 => x"73",
          4389 => x"81",
          4390 => x"75",
          4391 => x"38",
          4392 => x"88",
          4393 => x"a4",
          4394 => x"52",
          4395 => x"d8",
          4396 => x"c8",
          4397 => x"52",
          4398 => x"ff",
          4399 => x"82",
          4400 => x"80",
          4401 => x"15",
          4402 => x"81",
          4403 => x"74",
          4404 => x"38",
          4405 => x"e6",
          4406 => x"81",
          4407 => x"3d",
          4408 => x"f8",
          4409 => x"e7",
          4410 => x"c8",
          4411 => x"9a",
          4412 => x"53",
          4413 => x"51",
          4414 => x"82",
          4415 => x"81",
          4416 => x"74",
          4417 => x"54",
          4418 => x"14",
          4419 => x"06",
          4420 => x"74",
          4421 => x"38",
          4422 => x"82",
          4423 => x"8c",
          4424 => x"d3",
          4425 => x"3d",
          4426 => x"08",
          4427 => x"59",
          4428 => x"0b",
          4429 => x"82",
          4430 => x"82",
          4431 => x"55",
          4432 => x"cb",
          4433 => x"b5",
          4434 => x"55",
          4435 => x"81",
          4436 => x"2e",
          4437 => x"81",
          4438 => x"55",
          4439 => x"2e",
          4440 => x"a8",
          4441 => x"3f",
          4442 => x"08",
          4443 => x"0c",
          4444 => x"08",
          4445 => x"92",
          4446 => x"76",
          4447 => x"c8",
          4448 => x"cc",
          4449 => x"b5",
          4450 => x"2e",
          4451 => x"ae",
          4452 => x"a4",
          4453 => x"f7",
          4454 => x"c8",
          4455 => x"b5",
          4456 => x"80",
          4457 => x"3d",
          4458 => x"81",
          4459 => x"82",
          4460 => x"56",
          4461 => x"08",
          4462 => x"81",
          4463 => x"38",
          4464 => x"08",
          4465 => x"c0",
          4466 => x"c8",
          4467 => x"0b",
          4468 => x"08",
          4469 => x"82",
          4470 => x"ff",
          4471 => x"55",
          4472 => x"34",
          4473 => x"81",
          4474 => x"75",
          4475 => x"3f",
          4476 => x"81",
          4477 => x"54",
          4478 => x"83",
          4479 => x"74",
          4480 => x"81",
          4481 => x"38",
          4482 => x"82",
          4483 => x"76",
          4484 => x"b5",
          4485 => x"2e",
          4486 => x"d6",
          4487 => x"5d",
          4488 => x"82",
          4489 => x"98",
          4490 => x"2c",
          4491 => x"ff",
          4492 => x"78",
          4493 => x"82",
          4494 => x"70",
          4495 => x"98",
          4496 => x"f0",
          4497 => x"2b",
          4498 => x"71",
          4499 => x"70",
          4500 => x"aa",
          4501 => x"08",
          4502 => x"51",
          4503 => x"59",
          4504 => x"5d",
          4505 => x"73",
          4506 => x"e9",
          4507 => x"27",
          4508 => x"81",
          4509 => x"81",
          4510 => x"70",
          4511 => x"55",
          4512 => x"80",
          4513 => x"53",
          4514 => x"51",
          4515 => x"82",
          4516 => x"81",
          4517 => x"73",
          4518 => x"38",
          4519 => x"f0",
          4520 => x"b1",
          4521 => x"80",
          4522 => x"80",
          4523 => x"98",
          4524 => x"ff",
          4525 => x"55",
          4526 => x"97",
          4527 => x"74",
          4528 => x"f5",
          4529 => x"b5",
          4530 => x"ff",
          4531 => x"cc",
          4532 => x"80",
          4533 => x"2e",
          4534 => x"81",
          4535 => x"82",
          4536 => x"74",
          4537 => x"98",
          4538 => x"f0",
          4539 => x"2b",
          4540 => x"70",
          4541 => x"82",
          4542 => x"d8",
          4543 => x"51",
          4544 => x"58",
          4545 => x"77",
          4546 => x"06",
          4547 => x"82",
          4548 => x"08",
          4549 => x"0b",
          4550 => x"34",
          4551 => x"cc",
          4552 => x"39",
          4553 => x"f4",
          4554 => x"cc",
          4555 => x"af",
          4556 => x"7d",
          4557 => x"73",
          4558 => x"e1",
          4559 => x"29",
          4560 => x"05",
          4561 => x"04",
          4562 => x"33",
          4563 => x"2e",
          4564 => x"82",
          4565 => x"55",
          4566 => x"ab",
          4567 => x"2b",
          4568 => x"51",
          4569 => x"24",
          4570 => x"1a",
          4571 => x"81",
          4572 => x"81",
          4573 => x"81",
          4574 => x"70",
          4575 => x"cc",
          4576 => x"51",
          4577 => x"82",
          4578 => x"81",
          4579 => x"74",
          4580 => x"34",
          4581 => x"ae",
          4582 => x"34",
          4583 => x"33",
          4584 => x"25",
          4585 => x"14",
          4586 => x"cc",
          4587 => x"cc",
          4588 => x"81",
          4589 => x"81",
          4590 => x"70",
          4591 => x"cc",
          4592 => x"51",
          4593 => x"77",
          4594 => x"82",
          4595 => x"52",
          4596 => x"33",
          4597 => x"a3",
          4598 => x"81",
          4599 => x"81",
          4600 => x"70",
          4601 => x"cc",
          4602 => x"51",
          4603 => x"24",
          4604 => x"cc",
          4605 => x"98",
          4606 => x"2c",
          4607 => x"33",
          4608 => x"56",
          4609 => x"fc",
          4610 => x"cd",
          4611 => x"88",
          4612 => x"a1",
          4613 => x"80",
          4614 => x"80",
          4615 => x"98",
          4616 => x"f8",
          4617 => x"55",
          4618 => x"de",
          4619 => x"39",
          4620 => x"80",
          4621 => x"34",
          4622 => x"53",
          4623 => x"9e",
          4624 => x"9c",
          4625 => x"39",
          4626 => x"33",
          4627 => x"06",
          4628 => x"80",
          4629 => x"38",
          4630 => x"33",
          4631 => x"73",
          4632 => x"34",
          4633 => x"73",
          4634 => x"34",
          4635 => x"08",
          4636 => x"ff",
          4637 => x"82",
          4638 => x"70",
          4639 => x"98",
          4640 => x"f8",
          4641 => x"56",
          4642 => x"25",
          4643 => x"1a",
          4644 => x"33",
          4645 => x"cd",
          4646 => x"73",
          4647 => x"a2",
          4648 => x"81",
          4649 => x"81",
          4650 => x"70",
          4651 => x"cc",
          4652 => x"51",
          4653 => x"24",
          4654 => x"cd",
          4655 => x"a0",
          4656 => x"f1",
          4657 => x"fc",
          4658 => x"2b",
          4659 => x"82",
          4660 => x"57",
          4661 => x"74",
          4662 => x"c1",
          4663 => x"9c",
          4664 => x"51",
          4665 => x"3f",
          4666 => x"0a",
          4667 => x"0a",
          4668 => x"2c",
          4669 => x"33",
          4670 => x"75",
          4671 => x"38",
          4672 => x"82",
          4673 => x"7a",
          4674 => x"74",
          4675 => x"9c",
          4676 => x"51",
          4677 => x"3f",
          4678 => x"52",
          4679 => x"c9",
          4680 => x"c8",
          4681 => x"06",
          4682 => x"38",
          4683 => x"33",
          4684 => x"2e",
          4685 => x"53",
          4686 => x"51",
          4687 => x"84",
          4688 => x"34",
          4689 => x"cc",
          4690 => x"0b",
          4691 => x"34",
          4692 => x"c8",
          4693 => x"0d",
          4694 => x"fc",
          4695 => x"80",
          4696 => x"38",
          4697 => x"08",
          4698 => x"ff",
          4699 => x"82",
          4700 => x"ff",
          4701 => x"82",
          4702 => x"73",
          4703 => x"54",
          4704 => x"cc",
          4705 => x"cc",
          4706 => x"55",
          4707 => x"f9",
          4708 => x"14",
          4709 => x"cc",
          4710 => x"98",
          4711 => x"2c",
          4712 => x"06",
          4713 => x"74",
          4714 => x"38",
          4715 => x"81",
          4716 => x"34",
          4717 => x"08",
          4718 => x"51",
          4719 => x"3f",
          4720 => x"0a",
          4721 => x"0a",
          4722 => x"2c",
          4723 => x"33",
          4724 => x"75",
          4725 => x"38",
          4726 => x"08",
          4727 => x"ff",
          4728 => x"82",
          4729 => x"70",
          4730 => x"98",
          4731 => x"f8",
          4732 => x"56",
          4733 => x"24",
          4734 => x"82",
          4735 => x"52",
          4736 => x"9f",
          4737 => x"81",
          4738 => x"81",
          4739 => x"70",
          4740 => x"cc",
          4741 => x"51",
          4742 => x"25",
          4743 => x"fd",
          4744 => x"fc",
          4745 => x"ff",
          4746 => x"f8",
          4747 => x"54",
          4748 => x"f7",
          4749 => x"cd",
          4750 => x"81",
          4751 => x"82",
          4752 => x"74",
          4753 => x"52",
          4754 => x"e9",
          4755 => x"fc",
          4756 => x"ff",
          4757 => x"f8",
          4758 => x"54",
          4759 => x"d6",
          4760 => x"39",
          4761 => x"53",
          4762 => x"9e",
          4763 => x"f0",
          4764 => x"82",
          4765 => x"80",
          4766 => x"f8",
          4767 => x"39",
          4768 => x"82",
          4769 => x"55",
          4770 => x"a6",
          4771 => x"ff",
          4772 => x"82",
          4773 => x"82",
          4774 => x"82",
          4775 => x"81",
          4776 => x"05",
          4777 => x"79",
          4778 => x"bc",
          4779 => x"81",
          4780 => x"84",
          4781 => x"c8",
          4782 => x"08",
          4783 => x"80",
          4784 => x"74",
          4785 => x"c0",
          4786 => x"c8",
          4787 => x"f8",
          4788 => x"c8",
          4789 => x"06",
          4790 => x"74",
          4791 => x"ff",
          4792 => x"ff",
          4793 => x"fa",
          4794 => x"55",
          4795 => x"f6",
          4796 => x"51",
          4797 => x"3f",
          4798 => x"93",
          4799 => x"06",
          4800 => x"b4",
          4801 => x"74",
          4802 => x"38",
          4803 => x"a5",
          4804 => x"b5",
          4805 => x"cc",
          4806 => x"b5",
          4807 => x"ff",
          4808 => x"53",
          4809 => x"51",
          4810 => x"3f",
          4811 => x"7a",
          4812 => x"b4",
          4813 => x"08",
          4814 => x"80",
          4815 => x"74",
          4816 => x"c4",
          4817 => x"c8",
          4818 => x"f8",
          4819 => x"c8",
          4820 => x"06",
          4821 => x"74",
          4822 => x"ff",
          4823 => x"81",
          4824 => x"81",
          4825 => x"89",
          4826 => x"cc",
          4827 => x"7a",
          4828 => x"fc",
          4829 => x"f8",
          4830 => x"51",
          4831 => x"f5",
          4832 => x"cc",
          4833 => x"81",
          4834 => x"cc",
          4835 => x"56",
          4836 => x"27",
          4837 => x"82",
          4838 => x"52",
          4839 => x"73",
          4840 => x"34",
          4841 => x"33",
          4842 => x"9c",
          4843 => x"ed",
          4844 => x"fc",
          4845 => x"80",
          4846 => x"38",
          4847 => x"08",
          4848 => x"ff",
          4849 => x"82",
          4850 => x"ff",
          4851 => x"82",
          4852 => x"f4",
          4853 => x"3d",
          4854 => x"f4",
          4855 => x"c0",
          4856 => x"0b",
          4857 => x"23",
          4858 => x"80",
          4859 => x"f4",
          4860 => x"f5",
          4861 => x"c0",
          4862 => x"58",
          4863 => x"81",
          4864 => x"15",
          4865 => x"c0",
          4866 => x"84",
          4867 => x"85",
          4868 => x"b5",
          4869 => x"77",
          4870 => x"76",
          4871 => x"82",
          4872 => x"82",
          4873 => x"ff",
          4874 => x"80",
          4875 => x"ff",
          4876 => x"88",
          4877 => x"55",
          4878 => x"17",
          4879 => x"17",
          4880 => x"bc",
          4881 => x"29",
          4882 => x"08",
          4883 => x"51",
          4884 => x"82",
          4885 => x"83",
          4886 => x"3d",
          4887 => x"3d",
          4888 => x"81",
          4889 => x"27",
          4890 => x"12",
          4891 => x"11",
          4892 => x"ff",
          4893 => x"51",
          4894 => x"c8",
          4895 => x"0d",
          4896 => x"0d",
          4897 => x"22",
          4898 => x"aa",
          4899 => x"05",
          4900 => x"08",
          4901 => x"71",
          4902 => x"2b",
          4903 => x"33",
          4904 => x"71",
          4905 => x"02",
          4906 => x"05",
          4907 => x"ff",
          4908 => x"70",
          4909 => x"51",
          4910 => x"5b",
          4911 => x"54",
          4912 => x"34",
          4913 => x"34",
          4914 => x"08",
          4915 => x"2a",
          4916 => x"82",
          4917 => x"83",
          4918 => x"b5",
          4919 => x"17",
          4920 => x"12",
          4921 => x"2b",
          4922 => x"2b",
          4923 => x"06",
          4924 => x"52",
          4925 => x"83",
          4926 => x"70",
          4927 => x"54",
          4928 => x"12",
          4929 => x"ff",
          4930 => x"83",
          4931 => x"b5",
          4932 => x"56",
          4933 => x"72",
          4934 => x"89",
          4935 => x"fb",
          4936 => x"b5",
          4937 => x"84",
          4938 => x"22",
          4939 => x"72",
          4940 => x"33",
          4941 => x"71",
          4942 => x"83",
          4943 => x"5b",
          4944 => x"52",
          4945 => x"12",
          4946 => x"33",
          4947 => x"07",
          4948 => x"54",
          4949 => x"70",
          4950 => x"73",
          4951 => x"82",
          4952 => x"70",
          4953 => x"33",
          4954 => x"71",
          4955 => x"83",
          4956 => x"59",
          4957 => x"05",
          4958 => x"87",
          4959 => x"88",
          4960 => x"88",
          4961 => x"56",
          4962 => x"13",
          4963 => x"13",
          4964 => x"c0",
          4965 => x"33",
          4966 => x"71",
          4967 => x"70",
          4968 => x"06",
          4969 => x"53",
          4970 => x"53",
          4971 => x"70",
          4972 => x"87",
          4973 => x"fa",
          4974 => x"a2",
          4975 => x"b5",
          4976 => x"83",
          4977 => x"70",
          4978 => x"33",
          4979 => x"07",
          4980 => x"15",
          4981 => x"12",
          4982 => x"2b",
          4983 => x"07",
          4984 => x"55",
          4985 => x"57",
          4986 => x"80",
          4987 => x"38",
          4988 => x"ab",
          4989 => x"c0",
          4990 => x"70",
          4991 => x"33",
          4992 => x"71",
          4993 => x"74",
          4994 => x"81",
          4995 => x"88",
          4996 => x"83",
          4997 => x"f8",
          4998 => x"54",
          4999 => x"58",
          5000 => x"74",
          5001 => x"52",
          5002 => x"34",
          5003 => x"34",
          5004 => x"08",
          5005 => x"33",
          5006 => x"71",
          5007 => x"83",
          5008 => x"59",
          5009 => x"05",
          5010 => x"12",
          5011 => x"2b",
          5012 => x"ff",
          5013 => x"88",
          5014 => x"52",
          5015 => x"74",
          5016 => x"15",
          5017 => x"0d",
          5018 => x"0d",
          5019 => x"08",
          5020 => x"9e",
          5021 => x"83",
          5022 => x"82",
          5023 => x"12",
          5024 => x"2b",
          5025 => x"07",
          5026 => x"52",
          5027 => x"05",
          5028 => x"13",
          5029 => x"2b",
          5030 => x"05",
          5031 => x"71",
          5032 => x"2a",
          5033 => x"53",
          5034 => x"34",
          5035 => x"34",
          5036 => x"08",
          5037 => x"33",
          5038 => x"71",
          5039 => x"83",
          5040 => x"59",
          5041 => x"05",
          5042 => x"83",
          5043 => x"88",
          5044 => x"88",
          5045 => x"56",
          5046 => x"13",
          5047 => x"13",
          5048 => x"c0",
          5049 => x"11",
          5050 => x"33",
          5051 => x"07",
          5052 => x"0c",
          5053 => x"3d",
          5054 => x"3d",
          5055 => x"b5",
          5056 => x"83",
          5057 => x"ff",
          5058 => x"53",
          5059 => x"a7",
          5060 => x"c0",
          5061 => x"2b",
          5062 => x"11",
          5063 => x"33",
          5064 => x"71",
          5065 => x"75",
          5066 => x"81",
          5067 => x"98",
          5068 => x"2b",
          5069 => x"40",
          5070 => x"58",
          5071 => x"72",
          5072 => x"38",
          5073 => x"52",
          5074 => x"9d",
          5075 => x"39",
          5076 => x"85",
          5077 => x"8b",
          5078 => x"2b",
          5079 => x"79",
          5080 => x"51",
          5081 => x"76",
          5082 => x"75",
          5083 => x"56",
          5084 => x"34",
          5085 => x"08",
          5086 => x"12",
          5087 => x"33",
          5088 => x"07",
          5089 => x"54",
          5090 => x"53",
          5091 => x"34",
          5092 => x"34",
          5093 => x"08",
          5094 => x"0b",
          5095 => x"80",
          5096 => x"34",
          5097 => x"08",
          5098 => x"14",
          5099 => x"14",
          5100 => x"c0",
          5101 => x"33",
          5102 => x"71",
          5103 => x"70",
          5104 => x"07",
          5105 => x"53",
          5106 => x"54",
          5107 => x"72",
          5108 => x"8b",
          5109 => x"ff",
          5110 => x"52",
          5111 => x"08",
          5112 => x"f2",
          5113 => x"2e",
          5114 => x"51",
          5115 => x"83",
          5116 => x"f5",
          5117 => x"7e",
          5118 => x"e2",
          5119 => x"c8",
          5120 => x"ff",
          5121 => x"c0",
          5122 => x"33",
          5123 => x"71",
          5124 => x"70",
          5125 => x"58",
          5126 => x"ff",
          5127 => x"2e",
          5128 => x"75",
          5129 => x"70",
          5130 => x"33",
          5131 => x"07",
          5132 => x"ff",
          5133 => x"70",
          5134 => x"06",
          5135 => x"52",
          5136 => x"59",
          5137 => x"27",
          5138 => x"80",
          5139 => x"75",
          5140 => x"84",
          5141 => x"16",
          5142 => x"2b",
          5143 => x"75",
          5144 => x"81",
          5145 => x"85",
          5146 => x"59",
          5147 => x"83",
          5148 => x"c0",
          5149 => x"33",
          5150 => x"71",
          5151 => x"70",
          5152 => x"06",
          5153 => x"56",
          5154 => x"75",
          5155 => x"81",
          5156 => x"79",
          5157 => x"cc",
          5158 => x"74",
          5159 => x"c4",
          5160 => x"2e",
          5161 => x"89",
          5162 => x"f8",
          5163 => x"ac",
          5164 => x"80",
          5165 => x"75",
          5166 => x"3f",
          5167 => x"08",
          5168 => x"11",
          5169 => x"33",
          5170 => x"71",
          5171 => x"53",
          5172 => x"74",
          5173 => x"70",
          5174 => x"06",
          5175 => x"5c",
          5176 => x"78",
          5177 => x"76",
          5178 => x"57",
          5179 => x"34",
          5180 => x"08",
          5181 => x"71",
          5182 => x"86",
          5183 => x"12",
          5184 => x"2b",
          5185 => x"2a",
          5186 => x"53",
          5187 => x"73",
          5188 => x"75",
          5189 => x"82",
          5190 => x"70",
          5191 => x"33",
          5192 => x"71",
          5193 => x"83",
          5194 => x"5d",
          5195 => x"05",
          5196 => x"15",
          5197 => x"15",
          5198 => x"c0",
          5199 => x"71",
          5200 => x"33",
          5201 => x"71",
          5202 => x"70",
          5203 => x"5a",
          5204 => x"54",
          5205 => x"34",
          5206 => x"34",
          5207 => x"08",
          5208 => x"54",
          5209 => x"c8",
          5210 => x"0d",
          5211 => x"0d",
          5212 => x"b5",
          5213 => x"38",
          5214 => x"71",
          5215 => x"2e",
          5216 => x"51",
          5217 => x"82",
          5218 => x"53",
          5219 => x"c8",
          5220 => x"0d",
          5221 => x"0d",
          5222 => x"5c",
          5223 => x"40",
          5224 => x"08",
          5225 => x"81",
          5226 => x"f4",
          5227 => x"8e",
          5228 => x"ff",
          5229 => x"b5",
          5230 => x"83",
          5231 => x"8b",
          5232 => x"fc",
          5233 => x"54",
          5234 => x"7e",
          5235 => x"3f",
          5236 => x"08",
          5237 => x"06",
          5238 => x"08",
          5239 => x"83",
          5240 => x"ff",
          5241 => x"83",
          5242 => x"70",
          5243 => x"33",
          5244 => x"07",
          5245 => x"70",
          5246 => x"06",
          5247 => x"fc",
          5248 => x"29",
          5249 => x"81",
          5250 => x"88",
          5251 => x"90",
          5252 => x"4e",
          5253 => x"52",
          5254 => x"41",
          5255 => x"5b",
          5256 => x"8f",
          5257 => x"ff",
          5258 => x"31",
          5259 => x"ff",
          5260 => x"82",
          5261 => x"17",
          5262 => x"2b",
          5263 => x"29",
          5264 => x"81",
          5265 => x"98",
          5266 => x"2b",
          5267 => x"45",
          5268 => x"73",
          5269 => x"38",
          5270 => x"70",
          5271 => x"06",
          5272 => x"7b",
          5273 => x"38",
          5274 => x"73",
          5275 => x"81",
          5276 => x"78",
          5277 => x"3f",
          5278 => x"ff",
          5279 => x"e5",
          5280 => x"38",
          5281 => x"89",
          5282 => x"f6",
          5283 => x"a5",
          5284 => x"55",
          5285 => x"80",
          5286 => x"1d",
          5287 => x"83",
          5288 => x"88",
          5289 => x"57",
          5290 => x"3f",
          5291 => x"51",
          5292 => x"82",
          5293 => x"83",
          5294 => x"7e",
          5295 => x"70",
          5296 => x"b5",
          5297 => x"84",
          5298 => x"59",
          5299 => x"3f",
          5300 => x"08",
          5301 => x"75",
          5302 => x"06",
          5303 => x"85",
          5304 => x"54",
          5305 => x"80",
          5306 => x"51",
          5307 => x"82",
          5308 => x"1d",
          5309 => x"83",
          5310 => x"88",
          5311 => x"43",
          5312 => x"3f",
          5313 => x"51",
          5314 => x"82",
          5315 => x"83",
          5316 => x"7e",
          5317 => x"70",
          5318 => x"b5",
          5319 => x"84",
          5320 => x"59",
          5321 => x"3f",
          5322 => x"08",
          5323 => x"60",
          5324 => x"55",
          5325 => x"ff",
          5326 => x"a9",
          5327 => x"52",
          5328 => x"3f",
          5329 => x"08",
          5330 => x"c8",
          5331 => x"93",
          5332 => x"73",
          5333 => x"c8",
          5334 => x"97",
          5335 => x"51",
          5336 => x"7a",
          5337 => x"27",
          5338 => x"53",
          5339 => x"51",
          5340 => x"7a",
          5341 => x"82",
          5342 => x"05",
          5343 => x"f6",
          5344 => x"54",
          5345 => x"c8",
          5346 => x"0d",
          5347 => x"0d",
          5348 => x"70",
          5349 => x"d5",
          5350 => x"c8",
          5351 => x"b5",
          5352 => x"2e",
          5353 => x"53",
          5354 => x"b5",
          5355 => x"ff",
          5356 => x"74",
          5357 => x"0c",
          5358 => x"04",
          5359 => x"02",
          5360 => x"51",
          5361 => x"72",
          5362 => x"82",
          5363 => x"33",
          5364 => x"b5",
          5365 => x"3d",
          5366 => x"3d",
          5367 => x"05",
          5368 => x"05",
          5369 => x"56",
          5370 => x"72",
          5371 => x"e0",
          5372 => x"2b",
          5373 => x"8c",
          5374 => x"88",
          5375 => x"2e",
          5376 => x"88",
          5377 => x"0c",
          5378 => x"8c",
          5379 => x"71",
          5380 => x"87",
          5381 => x"0c",
          5382 => x"08",
          5383 => x"51",
          5384 => x"2e",
          5385 => x"c0",
          5386 => x"51",
          5387 => x"71",
          5388 => x"80",
          5389 => x"92",
          5390 => x"98",
          5391 => x"70",
          5392 => x"38",
          5393 => x"c4",
          5394 => x"b5",
          5395 => x"51",
          5396 => x"c8",
          5397 => x"0d",
          5398 => x"0d",
          5399 => x"02",
          5400 => x"05",
          5401 => x"58",
          5402 => x"52",
          5403 => x"3f",
          5404 => x"08",
          5405 => x"54",
          5406 => x"be",
          5407 => x"75",
          5408 => x"c0",
          5409 => x"87",
          5410 => x"12",
          5411 => x"84",
          5412 => x"40",
          5413 => x"85",
          5414 => x"98",
          5415 => x"7d",
          5416 => x"0c",
          5417 => x"85",
          5418 => x"06",
          5419 => x"71",
          5420 => x"38",
          5421 => x"71",
          5422 => x"05",
          5423 => x"19",
          5424 => x"a2",
          5425 => x"71",
          5426 => x"38",
          5427 => x"83",
          5428 => x"38",
          5429 => x"8a",
          5430 => x"98",
          5431 => x"71",
          5432 => x"c0",
          5433 => x"52",
          5434 => x"87",
          5435 => x"80",
          5436 => x"81",
          5437 => x"c0",
          5438 => x"53",
          5439 => x"82",
          5440 => x"71",
          5441 => x"1a",
          5442 => x"84",
          5443 => x"19",
          5444 => x"06",
          5445 => x"79",
          5446 => x"38",
          5447 => x"80",
          5448 => x"87",
          5449 => x"26",
          5450 => x"73",
          5451 => x"06",
          5452 => x"2e",
          5453 => x"52",
          5454 => x"82",
          5455 => x"8f",
          5456 => x"f3",
          5457 => x"62",
          5458 => x"05",
          5459 => x"57",
          5460 => x"83",
          5461 => x"52",
          5462 => x"3f",
          5463 => x"08",
          5464 => x"54",
          5465 => x"2e",
          5466 => x"81",
          5467 => x"74",
          5468 => x"c0",
          5469 => x"87",
          5470 => x"12",
          5471 => x"84",
          5472 => x"5f",
          5473 => x"0b",
          5474 => x"8c",
          5475 => x"0c",
          5476 => x"80",
          5477 => x"70",
          5478 => x"81",
          5479 => x"54",
          5480 => x"8c",
          5481 => x"81",
          5482 => x"7c",
          5483 => x"58",
          5484 => x"70",
          5485 => x"52",
          5486 => x"8a",
          5487 => x"98",
          5488 => x"71",
          5489 => x"c0",
          5490 => x"52",
          5491 => x"87",
          5492 => x"80",
          5493 => x"81",
          5494 => x"c0",
          5495 => x"53",
          5496 => x"82",
          5497 => x"71",
          5498 => x"19",
          5499 => x"81",
          5500 => x"ff",
          5501 => x"19",
          5502 => x"78",
          5503 => x"38",
          5504 => x"80",
          5505 => x"87",
          5506 => x"26",
          5507 => x"73",
          5508 => x"06",
          5509 => x"2e",
          5510 => x"52",
          5511 => x"82",
          5512 => x"8f",
          5513 => x"fa",
          5514 => x"02",
          5515 => x"05",
          5516 => x"05",
          5517 => x"71",
          5518 => x"57",
          5519 => x"82",
          5520 => x"81",
          5521 => x"54",
          5522 => x"38",
          5523 => x"c0",
          5524 => x"81",
          5525 => x"2e",
          5526 => x"71",
          5527 => x"38",
          5528 => x"87",
          5529 => x"11",
          5530 => x"80",
          5531 => x"80",
          5532 => x"83",
          5533 => x"38",
          5534 => x"72",
          5535 => x"2a",
          5536 => x"51",
          5537 => x"80",
          5538 => x"87",
          5539 => x"08",
          5540 => x"38",
          5541 => x"8c",
          5542 => x"96",
          5543 => x"0c",
          5544 => x"8c",
          5545 => x"08",
          5546 => x"51",
          5547 => x"38",
          5548 => x"56",
          5549 => x"80",
          5550 => x"85",
          5551 => x"77",
          5552 => x"83",
          5553 => x"75",
          5554 => x"b5",
          5555 => x"3d",
          5556 => x"3d",
          5557 => x"11",
          5558 => x"71",
          5559 => x"82",
          5560 => x"53",
          5561 => x"0d",
          5562 => x"0d",
          5563 => x"33",
          5564 => x"71",
          5565 => x"88",
          5566 => x"14",
          5567 => x"07",
          5568 => x"33",
          5569 => x"b5",
          5570 => x"53",
          5571 => x"52",
          5572 => x"04",
          5573 => x"73",
          5574 => x"92",
          5575 => x"52",
          5576 => x"81",
          5577 => x"70",
          5578 => x"70",
          5579 => x"3d",
          5580 => x"3d",
          5581 => x"52",
          5582 => x"70",
          5583 => x"34",
          5584 => x"51",
          5585 => x"81",
          5586 => x"70",
          5587 => x"70",
          5588 => x"05",
          5589 => x"88",
          5590 => x"72",
          5591 => x"0d",
          5592 => x"0d",
          5593 => x"54",
          5594 => x"80",
          5595 => x"71",
          5596 => x"53",
          5597 => x"81",
          5598 => x"ff",
          5599 => x"39",
          5600 => x"04",
          5601 => x"75",
          5602 => x"52",
          5603 => x"70",
          5604 => x"34",
          5605 => x"70",
          5606 => x"3d",
          5607 => x"3d",
          5608 => x"79",
          5609 => x"74",
          5610 => x"56",
          5611 => x"81",
          5612 => x"71",
          5613 => x"16",
          5614 => x"52",
          5615 => x"86",
          5616 => x"2e",
          5617 => x"82",
          5618 => x"86",
          5619 => x"fe",
          5620 => x"76",
          5621 => x"39",
          5622 => x"8a",
          5623 => x"51",
          5624 => x"71",
          5625 => x"33",
          5626 => x"0c",
          5627 => x"04",
          5628 => x"b5",
          5629 => x"80",
          5630 => x"c8",
          5631 => x"3d",
          5632 => x"80",
          5633 => x"33",
          5634 => x"7a",
          5635 => x"38",
          5636 => x"16",
          5637 => x"16",
          5638 => x"17",
          5639 => x"fa",
          5640 => x"b5",
          5641 => x"2e",
          5642 => x"b7",
          5643 => x"c8",
          5644 => x"34",
          5645 => x"70",
          5646 => x"31",
          5647 => x"59",
          5648 => x"77",
          5649 => x"82",
          5650 => x"74",
          5651 => x"81",
          5652 => x"81",
          5653 => x"53",
          5654 => x"16",
          5655 => x"e3",
          5656 => x"81",
          5657 => x"b5",
          5658 => x"3d",
          5659 => x"3d",
          5660 => x"56",
          5661 => x"74",
          5662 => x"2e",
          5663 => x"51",
          5664 => x"82",
          5665 => x"57",
          5666 => x"08",
          5667 => x"54",
          5668 => x"16",
          5669 => x"33",
          5670 => x"3f",
          5671 => x"08",
          5672 => x"38",
          5673 => x"57",
          5674 => x"0c",
          5675 => x"c8",
          5676 => x"0d",
          5677 => x"0d",
          5678 => x"57",
          5679 => x"82",
          5680 => x"58",
          5681 => x"08",
          5682 => x"76",
          5683 => x"83",
          5684 => x"06",
          5685 => x"84",
          5686 => x"78",
          5687 => x"81",
          5688 => x"38",
          5689 => x"82",
          5690 => x"52",
          5691 => x"52",
          5692 => x"3f",
          5693 => x"52",
          5694 => x"51",
          5695 => x"84",
          5696 => x"d2",
          5697 => x"fc",
          5698 => x"8a",
          5699 => x"52",
          5700 => x"51",
          5701 => x"90",
          5702 => x"84",
          5703 => x"fc",
          5704 => x"17",
          5705 => x"a0",
          5706 => x"86",
          5707 => x"08",
          5708 => x"b0",
          5709 => x"55",
          5710 => x"81",
          5711 => x"f8",
          5712 => x"84",
          5713 => x"53",
          5714 => x"17",
          5715 => x"d7",
          5716 => x"c8",
          5717 => x"83",
          5718 => x"77",
          5719 => x"0c",
          5720 => x"04",
          5721 => x"77",
          5722 => x"12",
          5723 => x"55",
          5724 => x"56",
          5725 => x"8d",
          5726 => x"22",
          5727 => x"ac",
          5728 => x"57",
          5729 => x"b5",
          5730 => x"3d",
          5731 => x"3d",
          5732 => x"70",
          5733 => x"57",
          5734 => x"81",
          5735 => x"98",
          5736 => x"81",
          5737 => x"74",
          5738 => x"72",
          5739 => x"f5",
          5740 => x"24",
          5741 => x"81",
          5742 => x"81",
          5743 => x"83",
          5744 => x"38",
          5745 => x"76",
          5746 => x"70",
          5747 => x"16",
          5748 => x"74",
          5749 => x"96",
          5750 => x"c8",
          5751 => x"38",
          5752 => x"06",
          5753 => x"33",
          5754 => x"89",
          5755 => x"08",
          5756 => x"54",
          5757 => x"fc",
          5758 => x"b5",
          5759 => x"fe",
          5760 => x"ff",
          5761 => x"11",
          5762 => x"2b",
          5763 => x"81",
          5764 => x"2a",
          5765 => x"51",
          5766 => x"e2",
          5767 => x"ff",
          5768 => x"da",
          5769 => x"2a",
          5770 => x"05",
          5771 => x"fc",
          5772 => x"b5",
          5773 => x"c6",
          5774 => x"83",
          5775 => x"05",
          5776 => x"f9",
          5777 => x"b5",
          5778 => x"ff",
          5779 => x"ae",
          5780 => x"2a",
          5781 => x"05",
          5782 => x"fc",
          5783 => x"b5",
          5784 => x"38",
          5785 => x"83",
          5786 => x"05",
          5787 => x"f8",
          5788 => x"b5",
          5789 => x"0a",
          5790 => x"39",
          5791 => x"82",
          5792 => x"89",
          5793 => x"f8",
          5794 => x"7c",
          5795 => x"56",
          5796 => x"77",
          5797 => x"38",
          5798 => x"08",
          5799 => x"38",
          5800 => x"72",
          5801 => x"9d",
          5802 => x"24",
          5803 => x"81",
          5804 => x"82",
          5805 => x"83",
          5806 => x"38",
          5807 => x"76",
          5808 => x"70",
          5809 => x"18",
          5810 => x"76",
          5811 => x"9e",
          5812 => x"c8",
          5813 => x"b5",
          5814 => x"d9",
          5815 => x"ff",
          5816 => x"05",
          5817 => x"81",
          5818 => x"54",
          5819 => x"80",
          5820 => x"77",
          5821 => x"f0",
          5822 => x"8f",
          5823 => x"51",
          5824 => x"34",
          5825 => x"17",
          5826 => x"2a",
          5827 => x"05",
          5828 => x"fa",
          5829 => x"b5",
          5830 => x"82",
          5831 => x"81",
          5832 => x"83",
          5833 => x"b4",
          5834 => x"2a",
          5835 => x"8f",
          5836 => x"2a",
          5837 => x"f0",
          5838 => x"06",
          5839 => x"72",
          5840 => x"ec",
          5841 => x"2a",
          5842 => x"05",
          5843 => x"fa",
          5844 => x"b5",
          5845 => x"82",
          5846 => x"80",
          5847 => x"83",
          5848 => x"52",
          5849 => x"fe",
          5850 => x"b4",
          5851 => x"a4",
          5852 => x"76",
          5853 => x"17",
          5854 => x"75",
          5855 => x"3f",
          5856 => x"08",
          5857 => x"c8",
          5858 => x"77",
          5859 => x"77",
          5860 => x"fc",
          5861 => x"b4",
          5862 => x"51",
          5863 => x"c9",
          5864 => x"c8",
          5865 => x"06",
          5866 => x"72",
          5867 => x"3f",
          5868 => x"17",
          5869 => x"b5",
          5870 => x"3d",
          5871 => x"3d",
          5872 => x"7e",
          5873 => x"56",
          5874 => x"75",
          5875 => x"74",
          5876 => x"27",
          5877 => x"80",
          5878 => x"ff",
          5879 => x"75",
          5880 => x"3f",
          5881 => x"08",
          5882 => x"c8",
          5883 => x"38",
          5884 => x"54",
          5885 => x"81",
          5886 => x"39",
          5887 => x"08",
          5888 => x"39",
          5889 => x"51",
          5890 => x"82",
          5891 => x"58",
          5892 => x"08",
          5893 => x"c7",
          5894 => x"c8",
          5895 => x"d2",
          5896 => x"c8",
          5897 => x"cf",
          5898 => x"74",
          5899 => x"fc",
          5900 => x"b5",
          5901 => x"38",
          5902 => x"fe",
          5903 => x"08",
          5904 => x"74",
          5905 => x"38",
          5906 => x"17",
          5907 => x"33",
          5908 => x"73",
          5909 => x"77",
          5910 => x"26",
          5911 => x"80",
          5912 => x"b5",
          5913 => x"3d",
          5914 => x"3d",
          5915 => x"71",
          5916 => x"5b",
          5917 => x"8c",
          5918 => x"77",
          5919 => x"38",
          5920 => x"78",
          5921 => x"81",
          5922 => x"79",
          5923 => x"f9",
          5924 => x"55",
          5925 => x"c8",
          5926 => x"e0",
          5927 => x"c8",
          5928 => x"b5",
          5929 => x"2e",
          5930 => x"98",
          5931 => x"b5",
          5932 => x"82",
          5933 => x"58",
          5934 => x"70",
          5935 => x"80",
          5936 => x"38",
          5937 => x"09",
          5938 => x"e2",
          5939 => x"56",
          5940 => x"76",
          5941 => x"82",
          5942 => x"7a",
          5943 => x"3f",
          5944 => x"b5",
          5945 => x"2e",
          5946 => x"86",
          5947 => x"c8",
          5948 => x"b5",
          5949 => x"70",
          5950 => x"07",
          5951 => x"7c",
          5952 => x"c8",
          5953 => x"51",
          5954 => x"81",
          5955 => x"b5",
          5956 => x"2e",
          5957 => x"17",
          5958 => x"74",
          5959 => x"73",
          5960 => x"27",
          5961 => x"58",
          5962 => x"80",
          5963 => x"56",
          5964 => x"98",
          5965 => x"26",
          5966 => x"56",
          5967 => x"81",
          5968 => x"52",
          5969 => x"c6",
          5970 => x"c8",
          5971 => x"b8",
          5972 => x"82",
          5973 => x"81",
          5974 => x"06",
          5975 => x"b5",
          5976 => x"82",
          5977 => x"09",
          5978 => x"72",
          5979 => x"70",
          5980 => x"51",
          5981 => x"80",
          5982 => x"78",
          5983 => x"06",
          5984 => x"73",
          5985 => x"39",
          5986 => x"52",
          5987 => x"f7",
          5988 => x"c8",
          5989 => x"c8",
          5990 => x"82",
          5991 => x"07",
          5992 => x"55",
          5993 => x"2e",
          5994 => x"80",
          5995 => x"75",
          5996 => x"76",
          5997 => x"3f",
          5998 => x"08",
          5999 => x"38",
          6000 => x"0c",
          6001 => x"fe",
          6002 => x"08",
          6003 => x"74",
          6004 => x"ff",
          6005 => x"0c",
          6006 => x"81",
          6007 => x"84",
          6008 => x"39",
          6009 => x"81",
          6010 => x"8c",
          6011 => x"8c",
          6012 => x"c8",
          6013 => x"39",
          6014 => x"55",
          6015 => x"c8",
          6016 => x"0d",
          6017 => x"0d",
          6018 => x"55",
          6019 => x"82",
          6020 => x"58",
          6021 => x"b5",
          6022 => x"d8",
          6023 => x"74",
          6024 => x"3f",
          6025 => x"08",
          6026 => x"08",
          6027 => x"59",
          6028 => x"77",
          6029 => x"70",
          6030 => x"c8",
          6031 => x"84",
          6032 => x"56",
          6033 => x"58",
          6034 => x"97",
          6035 => x"75",
          6036 => x"52",
          6037 => x"51",
          6038 => x"82",
          6039 => x"80",
          6040 => x"8a",
          6041 => x"32",
          6042 => x"72",
          6043 => x"2a",
          6044 => x"56",
          6045 => x"c8",
          6046 => x"0d",
          6047 => x"0d",
          6048 => x"08",
          6049 => x"74",
          6050 => x"26",
          6051 => x"74",
          6052 => x"72",
          6053 => x"74",
          6054 => x"88",
          6055 => x"73",
          6056 => x"33",
          6057 => x"27",
          6058 => x"16",
          6059 => x"9b",
          6060 => x"2a",
          6061 => x"88",
          6062 => x"58",
          6063 => x"80",
          6064 => x"16",
          6065 => x"0c",
          6066 => x"8a",
          6067 => x"89",
          6068 => x"72",
          6069 => x"38",
          6070 => x"51",
          6071 => x"82",
          6072 => x"54",
          6073 => x"08",
          6074 => x"38",
          6075 => x"b5",
          6076 => x"8b",
          6077 => x"08",
          6078 => x"08",
          6079 => x"82",
          6080 => x"74",
          6081 => x"cb",
          6082 => x"75",
          6083 => x"3f",
          6084 => x"08",
          6085 => x"73",
          6086 => x"98",
          6087 => x"82",
          6088 => x"2e",
          6089 => x"39",
          6090 => x"39",
          6091 => x"13",
          6092 => x"74",
          6093 => x"16",
          6094 => x"18",
          6095 => x"77",
          6096 => x"0c",
          6097 => x"04",
          6098 => x"7a",
          6099 => x"12",
          6100 => x"59",
          6101 => x"80",
          6102 => x"86",
          6103 => x"98",
          6104 => x"14",
          6105 => x"55",
          6106 => x"81",
          6107 => x"83",
          6108 => x"77",
          6109 => x"81",
          6110 => x"0c",
          6111 => x"55",
          6112 => x"76",
          6113 => x"17",
          6114 => x"74",
          6115 => x"9b",
          6116 => x"39",
          6117 => x"ff",
          6118 => x"2a",
          6119 => x"81",
          6120 => x"52",
          6121 => x"e6",
          6122 => x"c8",
          6123 => x"55",
          6124 => x"b5",
          6125 => x"80",
          6126 => x"55",
          6127 => x"08",
          6128 => x"f4",
          6129 => x"08",
          6130 => x"08",
          6131 => x"38",
          6132 => x"77",
          6133 => x"84",
          6134 => x"39",
          6135 => x"52",
          6136 => x"86",
          6137 => x"c8",
          6138 => x"55",
          6139 => x"08",
          6140 => x"c4",
          6141 => x"82",
          6142 => x"81",
          6143 => x"81",
          6144 => x"c8",
          6145 => x"b0",
          6146 => x"c8",
          6147 => x"51",
          6148 => x"82",
          6149 => x"a0",
          6150 => x"15",
          6151 => x"75",
          6152 => x"3f",
          6153 => x"08",
          6154 => x"76",
          6155 => x"77",
          6156 => x"9c",
          6157 => x"55",
          6158 => x"c8",
          6159 => x"0d",
          6160 => x"0d",
          6161 => x"08",
          6162 => x"80",
          6163 => x"fc",
          6164 => x"b5",
          6165 => x"82",
          6166 => x"80",
          6167 => x"b5",
          6168 => x"98",
          6169 => x"78",
          6170 => x"3f",
          6171 => x"08",
          6172 => x"c8",
          6173 => x"38",
          6174 => x"08",
          6175 => x"70",
          6176 => x"58",
          6177 => x"2e",
          6178 => x"83",
          6179 => x"82",
          6180 => x"55",
          6181 => x"81",
          6182 => x"07",
          6183 => x"2e",
          6184 => x"16",
          6185 => x"2e",
          6186 => x"88",
          6187 => x"82",
          6188 => x"56",
          6189 => x"51",
          6190 => x"82",
          6191 => x"54",
          6192 => x"08",
          6193 => x"9b",
          6194 => x"2e",
          6195 => x"83",
          6196 => x"73",
          6197 => x"0c",
          6198 => x"04",
          6199 => x"76",
          6200 => x"54",
          6201 => x"82",
          6202 => x"83",
          6203 => x"76",
          6204 => x"53",
          6205 => x"2e",
          6206 => x"90",
          6207 => x"51",
          6208 => x"82",
          6209 => x"90",
          6210 => x"53",
          6211 => x"c8",
          6212 => x"0d",
          6213 => x"0d",
          6214 => x"83",
          6215 => x"54",
          6216 => x"55",
          6217 => x"3f",
          6218 => x"51",
          6219 => x"2e",
          6220 => x"8b",
          6221 => x"2a",
          6222 => x"51",
          6223 => x"86",
          6224 => x"f7",
          6225 => x"7d",
          6226 => x"75",
          6227 => x"98",
          6228 => x"2e",
          6229 => x"98",
          6230 => x"78",
          6231 => x"3f",
          6232 => x"08",
          6233 => x"c8",
          6234 => x"38",
          6235 => x"70",
          6236 => x"73",
          6237 => x"58",
          6238 => x"8b",
          6239 => x"bf",
          6240 => x"ff",
          6241 => x"53",
          6242 => x"34",
          6243 => x"08",
          6244 => x"e5",
          6245 => x"81",
          6246 => x"2e",
          6247 => x"70",
          6248 => x"57",
          6249 => x"9e",
          6250 => x"2e",
          6251 => x"b5",
          6252 => x"df",
          6253 => x"72",
          6254 => x"81",
          6255 => x"76",
          6256 => x"2e",
          6257 => x"52",
          6258 => x"fc",
          6259 => x"c8",
          6260 => x"b5",
          6261 => x"38",
          6262 => x"fe",
          6263 => x"39",
          6264 => x"16",
          6265 => x"b5",
          6266 => x"3d",
          6267 => x"3d",
          6268 => x"08",
          6269 => x"52",
          6270 => x"c5",
          6271 => x"c8",
          6272 => x"b5",
          6273 => x"38",
          6274 => x"52",
          6275 => x"de",
          6276 => x"c8",
          6277 => x"b5",
          6278 => x"38",
          6279 => x"b5",
          6280 => x"9c",
          6281 => x"ea",
          6282 => x"53",
          6283 => x"9c",
          6284 => x"ea",
          6285 => x"0b",
          6286 => x"74",
          6287 => x"0c",
          6288 => x"04",
          6289 => x"75",
          6290 => x"12",
          6291 => x"53",
          6292 => x"9a",
          6293 => x"c8",
          6294 => x"9c",
          6295 => x"e5",
          6296 => x"0b",
          6297 => x"85",
          6298 => x"fa",
          6299 => x"7a",
          6300 => x"0b",
          6301 => x"98",
          6302 => x"2e",
          6303 => x"80",
          6304 => x"55",
          6305 => x"17",
          6306 => x"33",
          6307 => x"51",
          6308 => x"2e",
          6309 => x"85",
          6310 => x"06",
          6311 => x"e5",
          6312 => x"2e",
          6313 => x"8b",
          6314 => x"70",
          6315 => x"34",
          6316 => x"71",
          6317 => x"05",
          6318 => x"15",
          6319 => x"27",
          6320 => x"15",
          6321 => x"80",
          6322 => x"34",
          6323 => x"52",
          6324 => x"88",
          6325 => x"17",
          6326 => x"52",
          6327 => x"3f",
          6328 => x"08",
          6329 => x"12",
          6330 => x"3f",
          6331 => x"08",
          6332 => x"98",
          6333 => x"da",
          6334 => x"c8",
          6335 => x"23",
          6336 => x"04",
          6337 => x"7f",
          6338 => x"5b",
          6339 => x"33",
          6340 => x"73",
          6341 => x"38",
          6342 => x"80",
          6343 => x"38",
          6344 => x"8c",
          6345 => x"08",
          6346 => x"aa",
          6347 => x"41",
          6348 => x"33",
          6349 => x"73",
          6350 => x"81",
          6351 => x"81",
          6352 => x"dc",
          6353 => x"70",
          6354 => x"07",
          6355 => x"73",
          6356 => x"88",
          6357 => x"70",
          6358 => x"73",
          6359 => x"38",
          6360 => x"ab",
          6361 => x"52",
          6362 => x"91",
          6363 => x"c8",
          6364 => x"98",
          6365 => x"61",
          6366 => x"5a",
          6367 => x"a0",
          6368 => x"e7",
          6369 => x"70",
          6370 => x"79",
          6371 => x"73",
          6372 => x"81",
          6373 => x"38",
          6374 => x"33",
          6375 => x"ae",
          6376 => x"70",
          6377 => x"82",
          6378 => x"51",
          6379 => x"54",
          6380 => x"79",
          6381 => x"74",
          6382 => x"57",
          6383 => x"af",
          6384 => x"70",
          6385 => x"51",
          6386 => x"dc",
          6387 => x"73",
          6388 => x"38",
          6389 => x"82",
          6390 => x"19",
          6391 => x"54",
          6392 => x"82",
          6393 => x"54",
          6394 => x"78",
          6395 => x"81",
          6396 => x"54",
          6397 => x"81",
          6398 => x"af",
          6399 => x"77",
          6400 => x"70",
          6401 => x"25",
          6402 => x"07",
          6403 => x"51",
          6404 => x"2e",
          6405 => x"39",
          6406 => x"80",
          6407 => x"33",
          6408 => x"73",
          6409 => x"81",
          6410 => x"81",
          6411 => x"dc",
          6412 => x"70",
          6413 => x"07",
          6414 => x"73",
          6415 => x"b5",
          6416 => x"2e",
          6417 => x"83",
          6418 => x"76",
          6419 => x"07",
          6420 => x"2e",
          6421 => x"8b",
          6422 => x"77",
          6423 => x"30",
          6424 => x"71",
          6425 => x"53",
          6426 => x"55",
          6427 => x"38",
          6428 => x"5c",
          6429 => x"75",
          6430 => x"73",
          6431 => x"38",
          6432 => x"06",
          6433 => x"11",
          6434 => x"75",
          6435 => x"3f",
          6436 => x"08",
          6437 => x"38",
          6438 => x"33",
          6439 => x"54",
          6440 => x"e6",
          6441 => x"b5",
          6442 => x"2e",
          6443 => x"ff",
          6444 => x"74",
          6445 => x"38",
          6446 => x"75",
          6447 => x"17",
          6448 => x"57",
          6449 => x"a7",
          6450 => x"82",
          6451 => x"e5",
          6452 => x"b5",
          6453 => x"38",
          6454 => x"54",
          6455 => x"89",
          6456 => x"70",
          6457 => x"57",
          6458 => x"54",
          6459 => x"81",
          6460 => x"f7",
          6461 => x"7e",
          6462 => x"2e",
          6463 => x"33",
          6464 => x"e5",
          6465 => x"06",
          6466 => x"7a",
          6467 => x"a0",
          6468 => x"38",
          6469 => x"55",
          6470 => x"84",
          6471 => x"39",
          6472 => x"8b",
          6473 => x"7b",
          6474 => x"7a",
          6475 => x"3f",
          6476 => x"08",
          6477 => x"c8",
          6478 => x"38",
          6479 => x"52",
          6480 => x"aa",
          6481 => x"c8",
          6482 => x"b5",
          6483 => x"c2",
          6484 => x"08",
          6485 => x"55",
          6486 => x"ff",
          6487 => x"15",
          6488 => x"54",
          6489 => x"34",
          6490 => x"70",
          6491 => x"81",
          6492 => x"58",
          6493 => x"8b",
          6494 => x"74",
          6495 => x"3f",
          6496 => x"08",
          6497 => x"38",
          6498 => x"51",
          6499 => x"ff",
          6500 => x"ab",
          6501 => x"55",
          6502 => x"bb",
          6503 => x"2e",
          6504 => x"80",
          6505 => x"85",
          6506 => x"06",
          6507 => x"58",
          6508 => x"80",
          6509 => x"75",
          6510 => x"73",
          6511 => x"b5",
          6512 => x"0b",
          6513 => x"80",
          6514 => x"39",
          6515 => x"54",
          6516 => x"85",
          6517 => x"75",
          6518 => x"81",
          6519 => x"73",
          6520 => x"1b",
          6521 => x"2a",
          6522 => x"51",
          6523 => x"80",
          6524 => x"90",
          6525 => x"ff",
          6526 => x"05",
          6527 => x"f5",
          6528 => x"b5",
          6529 => x"1c",
          6530 => x"39",
          6531 => x"c8",
          6532 => x"0d",
          6533 => x"0d",
          6534 => x"7b",
          6535 => x"73",
          6536 => x"55",
          6537 => x"2e",
          6538 => x"75",
          6539 => x"57",
          6540 => x"26",
          6541 => x"ba",
          6542 => x"70",
          6543 => x"ba",
          6544 => x"06",
          6545 => x"73",
          6546 => x"70",
          6547 => x"51",
          6548 => x"89",
          6549 => x"82",
          6550 => x"ff",
          6551 => x"56",
          6552 => x"2e",
          6553 => x"80",
          6554 => x"80",
          6555 => x"08",
          6556 => x"76",
          6557 => x"58",
          6558 => x"81",
          6559 => x"ff",
          6560 => x"53",
          6561 => x"26",
          6562 => x"13",
          6563 => x"06",
          6564 => x"9f",
          6565 => x"99",
          6566 => x"e0",
          6567 => x"ff",
          6568 => x"72",
          6569 => x"2a",
          6570 => x"72",
          6571 => x"06",
          6572 => x"ff",
          6573 => x"30",
          6574 => x"70",
          6575 => x"07",
          6576 => x"9f",
          6577 => x"54",
          6578 => x"80",
          6579 => x"81",
          6580 => x"59",
          6581 => x"25",
          6582 => x"8b",
          6583 => x"24",
          6584 => x"76",
          6585 => x"78",
          6586 => x"82",
          6587 => x"51",
          6588 => x"c8",
          6589 => x"0d",
          6590 => x"0d",
          6591 => x"0b",
          6592 => x"ff",
          6593 => x"0c",
          6594 => x"51",
          6595 => x"84",
          6596 => x"c8",
          6597 => x"38",
          6598 => x"51",
          6599 => x"82",
          6600 => x"83",
          6601 => x"54",
          6602 => x"82",
          6603 => x"09",
          6604 => x"e3",
          6605 => x"b4",
          6606 => x"57",
          6607 => x"2e",
          6608 => x"83",
          6609 => x"74",
          6610 => x"70",
          6611 => x"25",
          6612 => x"51",
          6613 => x"38",
          6614 => x"2e",
          6615 => x"b5",
          6616 => x"82",
          6617 => x"80",
          6618 => x"e0",
          6619 => x"b5",
          6620 => x"82",
          6621 => x"80",
          6622 => x"85",
          6623 => x"c4",
          6624 => x"16",
          6625 => x"3f",
          6626 => x"08",
          6627 => x"c8",
          6628 => x"83",
          6629 => x"74",
          6630 => x"0c",
          6631 => x"04",
          6632 => x"61",
          6633 => x"80",
          6634 => x"58",
          6635 => x"0c",
          6636 => x"e1",
          6637 => x"c8",
          6638 => x"56",
          6639 => x"b5",
          6640 => x"86",
          6641 => x"b5",
          6642 => x"29",
          6643 => x"05",
          6644 => x"53",
          6645 => x"80",
          6646 => x"38",
          6647 => x"76",
          6648 => x"74",
          6649 => x"72",
          6650 => x"38",
          6651 => x"51",
          6652 => x"82",
          6653 => x"81",
          6654 => x"81",
          6655 => x"72",
          6656 => x"80",
          6657 => x"38",
          6658 => x"70",
          6659 => x"53",
          6660 => x"86",
          6661 => x"a7",
          6662 => x"34",
          6663 => x"34",
          6664 => x"14",
          6665 => x"b2",
          6666 => x"c8",
          6667 => x"06",
          6668 => x"54",
          6669 => x"72",
          6670 => x"76",
          6671 => x"38",
          6672 => x"70",
          6673 => x"53",
          6674 => x"85",
          6675 => x"70",
          6676 => x"5b",
          6677 => x"82",
          6678 => x"81",
          6679 => x"76",
          6680 => x"81",
          6681 => x"38",
          6682 => x"56",
          6683 => x"83",
          6684 => x"70",
          6685 => x"80",
          6686 => x"83",
          6687 => x"dc",
          6688 => x"b5",
          6689 => x"76",
          6690 => x"05",
          6691 => x"16",
          6692 => x"56",
          6693 => x"d7",
          6694 => x"8d",
          6695 => x"72",
          6696 => x"54",
          6697 => x"57",
          6698 => x"95",
          6699 => x"73",
          6700 => x"3f",
          6701 => x"08",
          6702 => x"57",
          6703 => x"89",
          6704 => x"56",
          6705 => x"d7",
          6706 => x"76",
          6707 => x"f1",
          6708 => x"76",
          6709 => x"e9",
          6710 => x"51",
          6711 => x"82",
          6712 => x"83",
          6713 => x"53",
          6714 => x"2e",
          6715 => x"84",
          6716 => x"ca",
          6717 => x"da",
          6718 => x"c8",
          6719 => x"ff",
          6720 => x"8d",
          6721 => x"14",
          6722 => x"3f",
          6723 => x"08",
          6724 => x"15",
          6725 => x"14",
          6726 => x"34",
          6727 => x"33",
          6728 => x"81",
          6729 => x"54",
          6730 => x"72",
          6731 => x"91",
          6732 => x"ff",
          6733 => x"29",
          6734 => x"33",
          6735 => x"72",
          6736 => x"72",
          6737 => x"38",
          6738 => x"06",
          6739 => x"2e",
          6740 => x"56",
          6741 => x"80",
          6742 => x"da",
          6743 => x"b5",
          6744 => x"82",
          6745 => x"88",
          6746 => x"8f",
          6747 => x"56",
          6748 => x"38",
          6749 => x"51",
          6750 => x"82",
          6751 => x"83",
          6752 => x"55",
          6753 => x"80",
          6754 => x"da",
          6755 => x"b5",
          6756 => x"80",
          6757 => x"da",
          6758 => x"b5",
          6759 => x"ff",
          6760 => x"8d",
          6761 => x"2e",
          6762 => x"88",
          6763 => x"14",
          6764 => x"05",
          6765 => x"75",
          6766 => x"38",
          6767 => x"52",
          6768 => x"51",
          6769 => x"3f",
          6770 => x"08",
          6771 => x"c8",
          6772 => x"82",
          6773 => x"b5",
          6774 => x"ff",
          6775 => x"26",
          6776 => x"57",
          6777 => x"f5",
          6778 => x"82",
          6779 => x"f5",
          6780 => x"81",
          6781 => x"8d",
          6782 => x"2e",
          6783 => x"82",
          6784 => x"16",
          6785 => x"16",
          6786 => x"70",
          6787 => x"7a",
          6788 => x"0c",
          6789 => x"83",
          6790 => x"06",
          6791 => x"de",
          6792 => x"ae",
          6793 => x"c8",
          6794 => x"ff",
          6795 => x"56",
          6796 => x"38",
          6797 => x"38",
          6798 => x"51",
          6799 => x"82",
          6800 => x"a8",
          6801 => x"82",
          6802 => x"39",
          6803 => x"80",
          6804 => x"38",
          6805 => x"15",
          6806 => x"53",
          6807 => x"8d",
          6808 => x"15",
          6809 => x"76",
          6810 => x"51",
          6811 => x"13",
          6812 => x"8d",
          6813 => x"15",
          6814 => x"c5",
          6815 => x"90",
          6816 => x"0b",
          6817 => x"ff",
          6818 => x"15",
          6819 => x"2e",
          6820 => x"81",
          6821 => x"e4",
          6822 => x"b6",
          6823 => x"c8",
          6824 => x"ff",
          6825 => x"81",
          6826 => x"06",
          6827 => x"81",
          6828 => x"51",
          6829 => x"82",
          6830 => x"80",
          6831 => x"b5",
          6832 => x"15",
          6833 => x"14",
          6834 => x"3f",
          6835 => x"08",
          6836 => x"06",
          6837 => x"d4",
          6838 => x"81",
          6839 => x"38",
          6840 => x"d8",
          6841 => x"b5",
          6842 => x"8b",
          6843 => x"2e",
          6844 => x"b3",
          6845 => x"14",
          6846 => x"3f",
          6847 => x"08",
          6848 => x"e4",
          6849 => x"81",
          6850 => x"84",
          6851 => x"d7",
          6852 => x"b5",
          6853 => x"15",
          6854 => x"14",
          6855 => x"3f",
          6856 => x"08",
          6857 => x"76",
          6858 => x"cd",
          6859 => x"05",
          6860 => x"cd",
          6861 => x"86",
          6862 => x"0b",
          6863 => x"80",
          6864 => x"b5",
          6865 => x"3d",
          6866 => x"3d",
          6867 => x"89",
          6868 => x"2e",
          6869 => x"08",
          6870 => x"2e",
          6871 => x"33",
          6872 => x"2e",
          6873 => x"13",
          6874 => x"22",
          6875 => x"76",
          6876 => x"06",
          6877 => x"13",
          6878 => x"c0",
          6879 => x"c8",
          6880 => x"52",
          6881 => x"71",
          6882 => x"55",
          6883 => x"53",
          6884 => x"0c",
          6885 => x"b5",
          6886 => x"3d",
          6887 => x"3d",
          6888 => x"05",
          6889 => x"89",
          6890 => x"52",
          6891 => x"3f",
          6892 => x"0b",
          6893 => x"08",
          6894 => x"82",
          6895 => x"84",
          6896 => x"80",
          6897 => x"55",
          6898 => x"2e",
          6899 => x"74",
          6900 => x"73",
          6901 => x"38",
          6902 => x"78",
          6903 => x"54",
          6904 => x"92",
          6905 => x"89",
          6906 => x"84",
          6907 => x"b0",
          6908 => x"c8",
          6909 => x"82",
          6910 => x"88",
          6911 => x"eb",
          6912 => x"02",
          6913 => x"e7",
          6914 => x"59",
          6915 => x"80",
          6916 => x"38",
          6917 => x"70",
          6918 => x"d0",
          6919 => x"3d",
          6920 => x"58",
          6921 => x"82",
          6922 => x"55",
          6923 => x"08",
          6924 => x"7a",
          6925 => x"8c",
          6926 => x"56",
          6927 => x"82",
          6928 => x"55",
          6929 => x"08",
          6930 => x"80",
          6931 => x"70",
          6932 => x"57",
          6933 => x"83",
          6934 => x"77",
          6935 => x"73",
          6936 => x"ab",
          6937 => x"2e",
          6938 => x"84",
          6939 => x"06",
          6940 => x"51",
          6941 => x"82",
          6942 => x"55",
          6943 => x"b2",
          6944 => x"06",
          6945 => x"b8",
          6946 => x"2a",
          6947 => x"51",
          6948 => x"2e",
          6949 => x"55",
          6950 => x"77",
          6951 => x"74",
          6952 => x"77",
          6953 => x"81",
          6954 => x"73",
          6955 => x"af",
          6956 => x"7a",
          6957 => x"3f",
          6958 => x"08",
          6959 => x"b2",
          6960 => x"8e",
          6961 => x"ea",
          6962 => x"a0",
          6963 => x"34",
          6964 => x"52",
          6965 => x"bd",
          6966 => x"62",
          6967 => x"d4",
          6968 => x"54",
          6969 => x"15",
          6970 => x"2e",
          6971 => x"7a",
          6972 => x"51",
          6973 => x"75",
          6974 => x"d4",
          6975 => x"be",
          6976 => x"c8",
          6977 => x"b5",
          6978 => x"ca",
          6979 => x"74",
          6980 => x"02",
          6981 => x"70",
          6982 => x"81",
          6983 => x"56",
          6984 => x"86",
          6985 => x"82",
          6986 => x"81",
          6987 => x"06",
          6988 => x"80",
          6989 => x"75",
          6990 => x"73",
          6991 => x"38",
          6992 => x"92",
          6993 => x"7a",
          6994 => x"3f",
          6995 => x"08",
          6996 => x"8c",
          6997 => x"55",
          6998 => x"08",
          6999 => x"77",
          7000 => x"81",
          7001 => x"73",
          7002 => x"38",
          7003 => x"07",
          7004 => x"11",
          7005 => x"0c",
          7006 => x"0c",
          7007 => x"52",
          7008 => x"3f",
          7009 => x"08",
          7010 => x"08",
          7011 => x"63",
          7012 => x"5a",
          7013 => x"82",
          7014 => x"82",
          7015 => x"8c",
          7016 => x"7a",
          7017 => x"17",
          7018 => x"23",
          7019 => x"34",
          7020 => x"1a",
          7021 => x"9c",
          7022 => x"0b",
          7023 => x"77",
          7024 => x"81",
          7025 => x"73",
          7026 => x"8d",
          7027 => x"c8",
          7028 => x"81",
          7029 => x"b5",
          7030 => x"1a",
          7031 => x"22",
          7032 => x"7b",
          7033 => x"a8",
          7034 => x"78",
          7035 => x"3f",
          7036 => x"08",
          7037 => x"c8",
          7038 => x"83",
          7039 => x"82",
          7040 => x"ff",
          7041 => x"06",
          7042 => x"55",
          7043 => x"56",
          7044 => x"76",
          7045 => x"51",
          7046 => x"27",
          7047 => x"70",
          7048 => x"5a",
          7049 => x"76",
          7050 => x"74",
          7051 => x"83",
          7052 => x"73",
          7053 => x"38",
          7054 => x"51",
          7055 => x"82",
          7056 => x"85",
          7057 => x"8e",
          7058 => x"2a",
          7059 => x"08",
          7060 => x"0c",
          7061 => x"79",
          7062 => x"73",
          7063 => x"0c",
          7064 => x"04",
          7065 => x"60",
          7066 => x"40",
          7067 => x"80",
          7068 => x"3d",
          7069 => x"78",
          7070 => x"3f",
          7071 => x"08",
          7072 => x"c8",
          7073 => x"91",
          7074 => x"74",
          7075 => x"38",
          7076 => x"c4",
          7077 => x"33",
          7078 => x"87",
          7079 => x"2e",
          7080 => x"95",
          7081 => x"91",
          7082 => x"56",
          7083 => x"81",
          7084 => x"34",
          7085 => x"a0",
          7086 => x"08",
          7087 => x"31",
          7088 => x"27",
          7089 => x"5c",
          7090 => x"82",
          7091 => x"19",
          7092 => x"ff",
          7093 => x"74",
          7094 => x"7e",
          7095 => x"ff",
          7096 => x"2a",
          7097 => x"79",
          7098 => x"87",
          7099 => x"08",
          7100 => x"98",
          7101 => x"78",
          7102 => x"3f",
          7103 => x"08",
          7104 => x"27",
          7105 => x"74",
          7106 => x"a3",
          7107 => x"1a",
          7108 => x"08",
          7109 => x"d4",
          7110 => x"b5",
          7111 => x"2e",
          7112 => x"82",
          7113 => x"1a",
          7114 => x"59",
          7115 => x"2e",
          7116 => x"77",
          7117 => x"11",
          7118 => x"55",
          7119 => x"85",
          7120 => x"31",
          7121 => x"76",
          7122 => x"81",
          7123 => x"ca",
          7124 => x"b5",
          7125 => x"d7",
          7126 => x"11",
          7127 => x"74",
          7128 => x"38",
          7129 => x"77",
          7130 => x"78",
          7131 => x"84",
          7132 => x"16",
          7133 => x"08",
          7134 => x"2b",
          7135 => x"cf",
          7136 => x"89",
          7137 => x"39",
          7138 => x"0c",
          7139 => x"83",
          7140 => x"80",
          7141 => x"55",
          7142 => x"83",
          7143 => x"9c",
          7144 => x"7e",
          7145 => x"3f",
          7146 => x"08",
          7147 => x"75",
          7148 => x"08",
          7149 => x"1f",
          7150 => x"7c",
          7151 => x"3f",
          7152 => x"7e",
          7153 => x"0c",
          7154 => x"1b",
          7155 => x"1c",
          7156 => x"fd",
          7157 => x"56",
          7158 => x"c8",
          7159 => x"0d",
          7160 => x"0d",
          7161 => x"64",
          7162 => x"58",
          7163 => x"90",
          7164 => x"52",
          7165 => x"d2",
          7166 => x"c8",
          7167 => x"b5",
          7168 => x"38",
          7169 => x"55",
          7170 => x"86",
          7171 => x"83",
          7172 => x"18",
          7173 => x"2a",
          7174 => x"51",
          7175 => x"56",
          7176 => x"83",
          7177 => x"39",
          7178 => x"19",
          7179 => x"83",
          7180 => x"0b",
          7181 => x"81",
          7182 => x"39",
          7183 => x"7c",
          7184 => x"74",
          7185 => x"38",
          7186 => x"7b",
          7187 => x"ec",
          7188 => x"08",
          7189 => x"06",
          7190 => x"81",
          7191 => x"8a",
          7192 => x"05",
          7193 => x"06",
          7194 => x"bf",
          7195 => x"38",
          7196 => x"55",
          7197 => x"7a",
          7198 => x"98",
          7199 => x"77",
          7200 => x"3f",
          7201 => x"08",
          7202 => x"c8",
          7203 => x"82",
          7204 => x"81",
          7205 => x"38",
          7206 => x"ff",
          7207 => x"98",
          7208 => x"18",
          7209 => x"74",
          7210 => x"7e",
          7211 => x"08",
          7212 => x"2e",
          7213 => x"8d",
          7214 => x"ce",
          7215 => x"b5",
          7216 => x"ee",
          7217 => x"08",
          7218 => x"d1",
          7219 => x"b5",
          7220 => x"2e",
          7221 => x"82",
          7222 => x"1b",
          7223 => x"5a",
          7224 => x"2e",
          7225 => x"78",
          7226 => x"11",
          7227 => x"55",
          7228 => x"85",
          7229 => x"31",
          7230 => x"76",
          7231 => x"81",
          7232 => x"c8",
          7233 => x"b5",
          7234 => x"a6",
          7235 => x"11",
          7236 => x"56",
          7237 => x"27",
          7238 => x"80",
          7239 => x"08",
          7240 => x"2b",
          7241 => x"b4",
          7242 => x"b5",
          7243 => x"80",
          7244 => x"34",
          7245 => x"56",
          7246 => x"8c",
          7247 => x"19",
          7248 => x"38",
          7249 => x"b6",
          7250 => x"c8",
          7251 => x"38",
          7252 => x"12",
          7253 => x"9c",
          7254 => x"18",
          7255 => x"06",
          7256 => x"31",
          7257 => x"76",
          7258 => x"7b",
          7259 => x"08",
          7260 => x"cd",
          7261 => x"b5",
          7262 => x"b6",
          7263 => x"7c",
          7264 => x"08",
          7265 => x"1f",
          7266 => x"cb",
          7267 => x"55",
          7268 => x"16",
          7269 => x"31",
          7270 => x"7f",
          7271 => x"94",
          7272 => x"70",
          7273 => x"8c",
          7274 => x"58",
          7275 => x"76",
          7276 => x"75",
          7277 => x"19",
          7278 => x"39",
          7279 => x"80",
          7280 => x"74",
          7281 => x"80",
          7282 => x"b5",
          7283 => x"3d",
          7284 => x"3d",
          7285 => x"3d",
          7286 => x"70",
          7287 => x"ea",
          7288 => x"c8",
          7289 => x"b5",
          7290 => x"fb",
          7291 => x"33",
          7292 => x"70",
          7293 => x"55",
          7294 => x"2e",
          7295 => x"a0",
          7296 => x"78",
          7297 => x"3f",
          7298 => x"08",
          7299 => x"c8",
          7300 => x"38",
          7301 => x"8b",
          7302 => x"07",
          7303 => x"8b",
          7304 => x"16",
          7305 => x"52",
          7306 => x"dd",
          7307 => x"16",
          7308 => x"15",
          7309 => x"3f",
          7310 => x"0a",
          7311 => x"51",
          7312 => x"76",
          7313 => x"51",
          7314 => x"78",
          7315 => x"83",
          7316 => x"51",
          7317 => x"82",
          7318 => x"90",
          7319 => x"bf",
          7320 => x"73",
          7321 => x"76",
          7322 => x"0c",
          7323 => x"04",
          7324 => x"76",
          7325 => x"fe",
          7326 => x"b5",
          7327 => x"82",
          7328 => x"9c",
          7329 => x"fc",
          7330 => x"51",
          7331 => x"82",
          7332 => x"53",
          7333 => x"08",
          7334 => x"b5",
          7335 => x"0c",
          7336 => x"c8",
          7337 => x"0d",
          7338 => x"0d",
          7339 => x"e6",
          7340 => x"52",
          7341 => x"b5",
          7342 => x"8b",
          7343 => x"c8",
          7344 => x"94",
          7345 => x"71",
          7346 => x"0c",
          7347 => x"04",
          7348 => x"80",
          7349 => x"d0",
          7350 => x"3d",
          7351 => x"3f",
          7352 => x"08",
          7353 => x"c8",
          7354 => x"38",
          7355 => x"52",
          7356 => x"05",
          7357 => x"3f",
          7358 => x"08",
          7359 => x"c8",
          7360 => x"02",
          7361 => x"33",
          7362 => x"55",
          7363 => x"25",
          7364 => x"7a",
          7365 => x"54",
          7366 => x"a2",
          7367 => x"84",
          7368 => x"06",
          7369 => x"73",
          7370 => x"38",
          7371 => x"70",
          7372 => x"a8",
          7373 => x"c8",
          7374 => x"0c",
          7375 => x"b5",
          7376 => x"2e",
          7377 => x"83",
          7378 => x"74",
          7379 => x"0c",
          7380 => x"04",
          7381 => x"6f",
          7382 => x"80",
          7383 => x"53",
          7384 => x"b8",
          7385 => x"3d",
          7386 => x"3f",
          7387 => x"08",
          7388 => x"c8",
          7389 => x"38",
          7390 => x"7c",
          7391 => x"47",
          7392 => x"54",
          7393 => x"81",
          7394 => x"52",
          7395 => x"52",
          7396 => x"3f",
          7397 => x"08",
          7398 => x"c8",
          7399 => x"38",
          7400 => x"51",
          7401 => x"82",
          7402 => x"57",
          7403 => x"08",
          7404 => x"69",
          7405 => x"da",
          7406 => x"b5",
          7407 => x"76",
          7408 => x"d5",
          7409 => x"b5",
          7410 => x"82",
          7411 => x"82",
          7412 => x"52",
          7413 => x"eb",
          7414 => x"c8",
          7415 => x"b5",
          7416 => x"38",
          7417 => x"51",
          7418 => x"73",
          7419 => x"08",
          7420 => x"76",
          7421 => x"d6",
          7422 => x"b5",
          7423 => x"82",
          7424 => x"80",
          7425 => x"76",
          7426 => x"81",
          7427 => x"82",
          7428 => x"39",
          7429 => x"38",
          7430 => x"bc",
          7431 => x"51",
          7432 => x"76",
          7433 => x"11",
          7434 => x"51",
          7435 => x"73",
          7436 => x"38",
          7437 => x"55",
          7438 => x"16",
          7439 => x"56",
          7440 => x"38",
          7441 => x"73",
          7442 => x"90",
          7443 => x"2e",
          7444 => x"16",
          7445 => x"ff",
          7446 => x"ff",
          7447 => x"58",
          7448 => x"74",
          7449 => x"75",
          7450 => x"18",
          7451 => x"58",
          7452 => x"fe",
          7453 => x"7b",
          7454 => x"06",
          7455 => x"18",
          7456 => x"58",
          7457 => x"80",
          7458 => x"94",
          7459 => x"29",
          7460 => x"05",
          7461 => x"33",
          7462 => x"56",
          7463 => x"2e",
          7464 => x"16",
          7465 => x"33",
          7466 => x"73",
          7467 => x"16",
          7468 => x"26",
          7469 => x"55",
          7470 => x"91",
          7471 => x"54",
          7472 => x"70",
          7473 => x"34",
          7474 => x"ec",
          7475 => x"70",
          7476 => x"34",
          7477 => x"09",
          7478 => x"38",
          7479 => x"39",
          7480 => x"19",
          7481 => x"33",
          7482 => x"05",
          7483 => x"78",
          7484 => x"80",
          7485 => x"82",
          7486 => x"9e",
          7487 => x"f7",
          7488 => x"7d",
          7489 => x"05",
          7490 => x"57",
          7491 => x"3f",
          7492 => x"08",
          7493 => x"c8",
          7494 => x"38",
          7495 => x"53",
          7496 => x"38",
          7497 => x"54",
          7498 => x"92",
          7499 => x"33",
          7500 => x"70",
          7501 => x"54",
          7502 => x"38",
          7503 => x"15",
          7504 => x"70",
          7505 => x"58",
          7506 => x"82",
          7507 => x"8a",
          7508 => x"89",
          7509 => x"53",
          7510 => x"b7",
          7511 => x"ff",
          7512 => x"dc",
          7513 => x"b5",
          7514 => x"15",
          7515 => x"53",
          7516 => x"dc",
          7517 => x"b5",
          7518 => x"26",
          7519 => x"30",
          7520 => x"70",
          7521 => x"77",
          7522 => x"18",
          7523 => x"51",
          7524 => x"88",
          7525 => x"73",
          7526 => x"52",
          7527 => x"ca",
          7528 => x"c8",
          7529 => x"b5",
          7530 => x"2e",
          7531 => x"82",
          7532 => x"ff",
          7533 => x"38",
          7534 => x"08",
          7535 => x"73",
          7536 => x"73",
          7537 => x"9c",
          7538 => x"27",
          7539 => x"75",
          7540 => x"16",
          7541 => x"17",
          7542 => x"33",
          7543 => x"70",
          7544 => x"55",
          7545 => x"80",
          7546 => x"73",
          7547 => x"cc",
          7548 => x"b5",
          7549 => x"82",
          7550 => x"94",
          7551 => x"c8",
          7552 => x"39",
          7553 => x"51",
          7554 => x"82",
          7555 => x"54",
          7556 => x"be",
          7557 => x"27",
          7558 => x"53",
          7559 => x"08",
          7560 => x"73",
          7561 => x"ff",
          7562 => x"15",
          7563 => x"16",
          7564 => x"ff",
          7565 => x"80",
          7566 => x"73",
          7567 => x"c6",
          7568 => x"b5",
          7569 => x"38",
          7570 => x"16",
          7571 => x"80",
          7572 => x"0b",
          7573 => x"81",
          7574 => x"75",
          7575 => x"b5",
          7576 => x"58",
          7577 => x"54",
          7578 => x"74",
          7579 => x"73",
          7580 => x"90",
          7581 => x"c0",
          7582 => x"90",
          7583 => x"83",
          7584 => x"72",
          7585 => x"38",
          7586 => x"08",
          7587 => x"77",
          7588 => x"80",
          7589 => x"b5",
          7590 => x"3d",
          7591 => x"3d",
          7592 => x"89",
          7593 => x"2e",
          7594 => x"80",
          7595 => x"fc",
          7596 => x"3d",
          7597 => x"e1",
          7598 => x"b5",
          7599 => x"82",
          7600 => x"80",
          7601 => x"76",
          7602 => x"75",
          7603 => x"3f",
          7604 => x"08",
          7605 => x"c8",
          7606 => x"38",
          7607 => x"70",
          7608 => x"57",
          7609 => x"a2",
          7610 => x"33",
          7611 => x"70",
          7612 => x"55",
          7613 => x"2e",
          7614 => x"16",
          7615 => x"51",
          7616 => x"82",
          7617 => x"88",
          7618 => x"54",
          7619 => x"84",
          7620 => x"52",
          7621 => x"e5",
          7622 => x"c8",
          7623 => x"84",
          7624 => x"06",
          7625 => x"55",
          7626 => x"80",
          7627 => x"80",
          7628 => x"54",
          7629 => x"c8",
          7630 => x"0d",
          7631 => x"0d",
          7632 => x"fc",
          7633 => x"52",
          7634 => x"3f",
          7635 => x"08",
          7636 => x"b5",
          7637 => x"0c",
          7638 => x"04",
          7639 => x"77",
          7640 => x"fc",
          7641 => x"53",
          7642 => x"de",
          7643 => x"c8",
          7644 => x"b5",
          7645 => x"df",
          7646 => x"38",
          7647 => x"08",
          7648 => x"cd",
          7649 => x"b5",
          7650 => x"80",
          7651 => x"b5",
          7652 => x"73",
          7653 => x"3f",
          7654 => x"08",
          7655 => x"c8",
          7656 => x"09",
          7657 => x"38",
          7658 => x"39",
          7659 => x"08",
          7660 => x"52",
          7661 => x"b3",
          7662 => x"73",
          7663 => x"3f",
          7664 => x"08",
          7665 => x"30",
          7666 => x"9f",
          7667 => x"b5",
          7668 => x"51",
          7669 => x"72",
          7670 => x"0c",
          7671 => x"04",
          7672 => x"65",
          7673 => x"89",
          7674 => x"96",
          7675 => x"df",
          7676 => x"b5",
          7677 => x"82",
          7678 => x"b2",
          7679 => x"75",
          7680 => x"3f",
          7681 => x"08",
          7682 => x"c8",
          7683 => x"02",
          7684 => x"33",
          7685 => x"55",
          7686 => x"25",
          7687 => x"55",
          7688 => x"80",
          7689 => x"76",
          7690 => x"d4",
          7691 => x"82",
          7692 => x"94",
          7693 => x"f0",
          7694 => x"65",
          7695 => x"53",
          7696 => x"05",
          7697 => x"51",
          7698 => x"82",
          7699 => x"5b",
          7700 => x"08",
          7701 => x"7c",
          7702 => x"08",
          7703 => x"fe",
          7704 => x"08",
          7705 => x"55",
          7706 => x"91",
          7707 => x"0c",
          7708 => x"81",
          7709 => x"39",
          7710 => x"c7",
          7711 => x"c8",
          7712 => x"55",
          7713 => x"2e",
          7714 => x"bf",
          7715 => x"5f",
          7716 => x"92",
          7717 => x"51",
          7718 => x"82",
          7719 => x"ff",
          7720 => x"82",
          7721 => x"81",
          7722 => x"82",
          7723 => x"30",
          7724 => x"c8",
          7725 => x"25",
          7726 => x"19",
          7727 => x"5a",
          7728 => x"08",
          7729 => x"38",
          7730 => x"a4",
          7731 => x"b5",
          7732 => x"58",
          7733 => x"77",
          7734 => x"7d",
          7735 => x"bf",
          7736 => x"b5",
          7737 => x"82",
          7738 => x"80",
          7739 => x"70",
          7740 => x"ff",
          7741 => x"56",
          7742 => x"2e",
          7743 => x"9e",
          7744 => x"51",
          7745 => x"3f",
          7746 => x"08",
          7747 => x"06",
          7748 => x"80",
          7749 => x"19",
          7750 => x"54",
          7751 => x"14",
          7752 => x"c5",
          7753 => x"c8",
          7754 => x"06",
          7755 => x"80",
          7756 => x"19",
          7757 => x"54",
          7758 => x"06",
          7759 => x"79",
          7760 => x"78",
          7761 => x"79",
          7762 => x"84",
          7763 => x"07",
          7764 => x"84",
          7765 => x"82",
          7766 => x"92",
          7767 => x"f9",
          7768 => x"8a",
          7769 => x"53",
          7770 => x"e3",
          7771 => x"b5",
          7772 => x"82",
          7773 => x"81",
          7774 => x"17",
          7775 => x"81",
          7776 => x"17",
          7777 => x"2a",
          7778 => x"51",
          7779 => x"55",
          7780 => x"81",
          7781 => x"17",
          7782 => x"8c",
          7783 => x"81",
          7784 => x"9b",
          7785 => x"c8",
          7786 => x"17",
          7787 => x"51",
          7788 => x"82",
          7789 => x"74",
          7790 => x"56",
          7791 => x"98",
          7792 => x"76",
          7793 => x"c6",
          7794 => x"c8",
          7795 => x"09",
          7796 => x"38",
          7797 => x"b5",
          7798 => x"2e",
          7799 => x"85",
          7800 => x"a3",
          7801 => x"38",
          7802 => x"b5",
          7803 => x"15",
          7804 => x"38",
          7805 => x"53",
          7806 => x"08",
          7807 => x"c3",
          7808 => x"b5",
          7809 => x"94",
          7810 => x"18",
          7811 => x"33",
          7812 => x"54",
          7813 => x"34",
          7814 => x"85",
          7815 => x"18",
          7816 => x"74",
          7817 => x"0c",
          7818 => x"04",
          7819 => x"82",
          7820 => x"ff",
          7821 => x"a1",
          7822 => x"e4",
          7823 => x"c8",
          7824 => x"b5",
          7825 => x"f5",
          7826 => x"a1",
          7827 => x"95",
          7828 => x"58",
          7829 => x"82",
          7830 => x"55",
          7831 => x"08",
          7832 => x"02",
          7833 => x"33",
          7834 => x"70",
          7835 => x"55",
          7836 => x"73",
          7837 => x"75",
          7838 => x"80",
          7839 => x"bd",
          7840 => x"d6",
          7841 => x"81",
          7842 => x"87",
          7843 => x"ad",
          7844 => x"78",
          7845 => x"3f",
          7846 => x"08",
          7847 => x"70",
          7848 => x"55",
          7849 => x"2e",
          7850 => x"78",
          7851 => x"c8",
          7852 => x"08",
          7853 => x"38",
          7854 => x"b5",
          7855 => x"76",
          7856 => x"70",
          7857 => x"b5",
          7858 => x"c8",
          7859 => x"b5",
          7860 => x"e9",
          7861 => x"c8",
          7862 => x"51",
          7863 => x"82",
          7864 => x"55",
          7865 => x"08",
          7866 => x"55",
          7867 => x"82",
          7868 => x"84",
          7869 => x"82",
          7870 => x"80",
          7871 => x"51",
          7872 => x"82",
          7873 => x"82",
          7874 => x"30",
          7875 => x"c8",
          7876 => x"25",
          7877 => x"75",
          7878 => x"38",
          7879 => x"8f",
          7880 => x"75",
          7881 => x"c1",
          7882 => x"b5",
          7883 => x"74",
          7884 => x"51",
          7885 => x"3f",
          7886 => x"08",
          7887 => x"b5",
          7888 => x"3d",
          7889 => x"3d",
          7890 => x"99",
          7891 => x"52",
          7892 => x"d8",
          7893 => x"b5",
          7894 => x"82",
          7895 => x"82",
          7896 => x"5e",
          7897 => x"3d",
          7898 => x"cf",
          7899 => x"b5",
          7900 => x"82",
          7901 => x"86",
          7902 => x"82",
          7903 => x"b5",
          7904 => x"2e",
          7905 => x"82",
          7906 => x"80",
          7907 => x"70",
          7908 => x"06",
          7909 => x"54",
          7910 => x"38",
          7911 => x"52",
          7912 => x"52",
          7913 => x"3f",
          7914 => x"08",
          7915 => x"82",
          7916 => x"83",
          7917 => x"82",
          7918 => x"81",
          7919 => x"06",
          7920 => x"54",
          7921 => x"08",
          7922 => x"81",
          7923 => x"81",
          7924 => x"39",
          7925 => x"38",
          7926 => x"08",
          7927 => x"c4",
          7928 => x"b5",
          7929 => x"82",
          7930 => x"81",
          7931 => x"53",
          7932 => x"19",
          7933 => x"8c",
          7934 => x"ae",
          7935 => x"34",
          7936 => x"0b",
          7937 => x"82",
          7938 => x"52",
          7939 => x"51",
          7940 => x"3f",
          7941 => x"b4",
          7942 => x"c9",
          7943 => x"53",
          7944 => x"53",
          7945 => x"51",
          7946 => x"3f",
          7947 => x"0b",
          7948 => x"34",
          7949 => x"80",
          7950 => x"51",
          7951 => x"78",
          7952 => x"83",
          7953 => x"51",
          7954 => x"82",
          7955 => x"54",
          7956 => x"08",
          7957 => x"88",
          7958 => x"64",
          7959 => x"ff",
          7960 => x"75",
          7961 => x"78",
          7962 => x"3f",
          7963 => x"0b",
          7964 => x"78",
          7965 => x"83",
          7966 => x"51",
          7967 => x"3f",
          7968 => x"08",
          7969 => x"80",
          7970 => x"76",
          7971 => x"ae",
          7972 => x"b5",
          7973 => x"3d",
          7974 => x"3d",
          7975 => x"84",
          7976 => x"f1",
          7977 => x"a8",
          7978 => x"05",
          7979 => x"51",
          7980 => x"82",
          7981 => x"55",
          7982 => x"08",
          7983 => x"78",
          7984 => x"08",
          7985 => x"70",
          7986 => x"b8",
          7987 => x"c8",
          7988 => x"b5",
          7989 => x"b9",
          7990 => x"9b",
          7991 => x"a0",
          7992 => x"55",
          7993 => x"38",
          7994 => x"3d",
          7995 => x"3d",
          7996 => x"51",
          7997 => x"3f",
          7998 => x"52",
          7999 => x"52",
          8000 => x"dd",
          8001 => x"08",
          8002 => x"cb",
          8003 => x"b5",
          8004 => x"82",
          8005 => x"95",
          8006 => x"2e",
          8007 => x"88",
          8008 => x"3d",
          8009 => x"38",
          8010 => x"e5",
          8011 => x"c8",
          8012 => x"09",
          8013 => x"b8",
          8014 => x"c9",
          8015 => x"b5",
          8016 => x"82",
          8017 => x"81",
          8018 => x"56",
          8019 => x"3d",
          8020 => x"52",
          8021 => x"ff",
          8022 => x"02",
          8023 => x"8b",
          8024 => x"16",
          8025 => x"2a",
          8026 => x"51",
          8027 => x"89",
          8028 => x"07",
          8029 => x"17",
          8030 => x"81",
          8031 => x"34",
          8032 => x"70",
          8033 => x"81",
          8034 => x"55",
          8035 => x"80",
          8036 => x"64",
          8037 => x"38",
          8038 => x"51",
          8039 => x"82",
          8040 => x"52",
          8041 => x"b7",
          8042 => x"55",
          8043 => x"08",
          8044 => x"dd",
          8045 => x"c8",
          8046 => x"51",
          8047 => x"3f",
          8048 => x"08",
          8049 => x"11",
          8050 => x"82",
          8051 => x"80",
          8052 => x"16",
          8053 => x"ae",
          8054 => x"06",
          8055 => x"53",
          8056 => x"51",
          8057 => x"78",
          8058 => x"83",
          8059 => x"39",
          8060 => x"08",
          8061 => x"51",
          8062 => x"82",
          8063 => x"55",
          8064 => x"08",
          8065 => x"51",
          8066 => x"3f",
          8067 => x"08",
          8068 => x"b5",
          8069 => x"3d",
          8070 => x"3d",
          8071 => x"db",
          8072 => x"84",
          8073 => x"05",
          8074 => x"82",
          8075 => x"d0",
          8076 => x"3d",
          8077 => x"3f",
          8078 => x"08",
          8079 => x"c8",
          8080 => x"38",
          8081 => x"52",
          8082 => x"05",
          8083 => x"3f",
          8084 => x"08",
          8085 => x"c8",
          8086 => x"02",
          8087 => x"33",
          8088 => x"54",
          8089 => x"aa",
          8090 => x"06",
          8091 => x"8b",
          8092 => x"06",
          8093 => x"07",
          8094 => x"56",
          8095 => x"34",
          8096 => x"0b",
          8097 => x"78",
          8098 => x"a9",
          8099 => x"c8",
          8100 => x"82",
          8101 => x"95",
          8102 => x"ef",
          8103 => x"56",
          8104 => x"3d",
          8105 => x"94",
          8106 => x"f4",
          8107 => x"c8",
          8108 => x"b5",
          8109 => x"cb",
          8110 => x"63",
          8111 => x"d4",
          8112 => x"c0",
          8113 => x"c8",
          8114 => x"b5",
          8115 => x"38",
          8116 => x"05",
          8117 => x"06",
          8118 => x"73",
          8119 => x"16",
          8120 => x"22",
          8121 => x"07",
          8122 => x"1f",
          8123 => x"c2",
          8124 => x"81",
          8125 => x"34",
          8126 => x"b3",
          8127 => x"b5",
          8128 => x"74",
          8129 => x"0c",
          8130 => x"04",
          8131 => x"69",
          8132 => x"80",
          8133 => x"d0",
          8134 => x"3d",
          8135 => x"3f",
          8136 => x"08",
          8137 => x"08",
          8138 => x"b5",
          8139 => x"80",
          8140 => x"57",
          8141 => x"81",
          8142 => x"70",
          8143 => x"55",
          8144 => x"80",
          8145 => x"5d",
          8146 => x"52",
          8147 => x"52",
          8148 => x"a9",
          8149 => x"c8",
          8150 => x"b5",
          8151 => x"d1",
          8152 => x"73",
          8153 => x"3f",
          8154 => x"08",
          8155 => x"c8",
          8156 => x"82",
          8157 => x"82",
          8158 => x"65",
          8159 => x"78",
          8160 => x"7b",
          8161 => x"55",
          8162 => x"34",
          8163 => x"8a",
          8164 => x"38",
          8165 => x"1a",
          8166 => x"34",
          8167 => x"9e",
          8168 => x"70",
          8169 => x"51",
          8170 => x"a0",
          8171 => x"8e",
          8172 => x"2e",
          8173 => x"86",
          8174 => x"34",
          8175 => x"30",
          8176 => x"80",
          8177 => x"7a",
          8178 => x"c1",
          8179 => x"2e",
          8180 => x"a0",
          8181 => x"51",
          8182 => x"3f",
          8183 => x"08",
          8184 => x"c8",
          8185 => x"7b",
          8186 => x"55",
          8187 => x"73",
          8188 => x"38",
          8189 => x"73",
          8190 => x"38",
          8191 => x"15",
          8192 => x"ff",
          8193 => x"82",
          8194 => x"7b",
          8195 => x"b5",
          8196 => x"3d",
          8197 => x"3d",
          8198 => x"9c",
          8199 => x"05",
          8200 => x"51",
          8201 => x"82",
          8202 => x"82",
          8203 => x"56",
          8204 => x"c8",
          8205 => x"38",
          8206 => x"52",
          8207 => x"52",
          8208 => x"c0",
          8209 => x"70",
          8210 => x"ff",
          8211 => x"55",
          8212 => x"27",
          8213 => x"78",
          8214 => x"ff",
          8215 => x"05",
          8216 => x"55",
          8217 => x"3f",
          8218 => x"08",
          8219 => x"38",
          8220 => x"70",
          8221 => x"ff",
          8222 => x"82",
          8223 => x"80",
          8224 => x"74",
          8225 => x"07",
          8226 => x"4e",
          8227 => x"82",
          8228 => x"55",
          8229 => x"70",
          8230 => x"06",
          8231 => x"99",
          8232 => x"e0",
          8233 => x"ff",
          8234 => x"54",
          8235 => x"27",
          8236 => x"ae",
          8237 => x"55",
          8238 => x"a3",
          8239 => x"82",
          8240 => x"ff",
          8241 => x"82",
          8242 => x"93",
          8243 => x"75",
          8244 => x"76",
          8245 => x"38",
          8246 => x"77",
          8247 => x"86",
          8248 => x"39",
          8249 => x"27",
          8250 => x"88",
          8251 => x"78",
          8252 => x"5a",
          8253 => x"57",
          8254 => x"81",
          8255 => x"81",
          8256 => x"33",
          8257 => x"06",
          8258 => x"57",
          8259 => x"fe",
          8260 => x"3d",
          8261 => x"55",
          8262 => x"2e",
          8263 => x"76",
          8264 => x"38",
          8265 => x"55",
          8266 => x"33",
          8267 => x"a0",
          8268 => x"06",
          8269 => x"17",
          8270 => x"38",
          8271 => x"43",
          8272 => x"3d",
          8273 => x"ff",
          8274 => x"82",
          8275 => x"54",
          8276 => x"08",
          8277 => x"81",
          8278 => x"ff",
          8279 => x"82",
          8280 => x"54",
          8281 => x"08",
          8282 => x"80",
          8283 => x"54",
          8284 => x"80",
          8285 => x"b5",
          8286 => x"2e",
          8287 => x"80",
          8288 => x"54",
          8289 => x"80",
          8290 => x"52",
          8291 => x"bd",
          8292 => x"b5",
          8293 => x"82",
          8294 => x"b1",
          8295 => x"82",
          8296 => x"52",
          8297 => x"ab",
          8298 => x"54",
          8299 => x"15",
          8300 => x"78",
          8301 => x"ff",
          8302 => x"79",
          8303 => x"83",
          8304 => x"51",
          8305 => x"3f",
          8306 => x"08",
          8307 => x"74",
          8308 => x"0c",
          8309 => x"04",
          8310 => x"60",
          8311 => x"05",
          8312 => x"33",
          8313 => x"05",
          8314 => x"40",
          8315 => x"da",
          8316 => x"c8",
          8317 => x"b5",
          8318 => x"bd",
          8319 => x"33",
          8320 => x"b5",
          8321 => x"2e",
          8322 => x"1a",
          8323 => x"90",
          8324 => x"33",
          8325 => x"70",
          8326 => x"55",
          8327 => x"38",
          8328 => x"97",
          8329 => x"82",
          8330 => x"58",
          8331 => x"7e",
          8332 => x"70",
          8333 => x"55",
          8334 => x"56",
          8335 => x"c6",
          8336 => x"7d",
          8337 => x"70",
          8338 => x"2a",
          8339 => x"08",
          8340 => x"08",
          8341 => x"5d",
          8342 => x"77",
          8343 => x"98",
          8344 => x"26",
          8345 => x"57",
          8346 => x"59",
          8347 => x"52",
          8348 => x"ae",
          8349 => x"15",
          8350 => x"98",
          8351 => x"26",
          8352 => x"55",
          8353 => x"08",
          8354 => x"99",
          8355 => x"c8",
          8356 => x"ff",
          8357 => x"b5",
          8358 => x"38",
          8359 => x"75",
          8360 => x"81",
          8361 => x"93",
          8362 => x"80",
          8363 => x"2e",
          8364 => x"ff",
          8365 => x"58",
          8366 => x"7d",
          8367 => x"38",
          8368 => x"55",
          8369 => x"b4",
          8370 => x"56",
          8371 => x"09",
          8372 => x"38",
          8373 => x"53",
          8374 => x"51",
          8375 => x"3f",
          8376 => x"08",
          8377 => x"c8",
          8378 => x"38",
          8379 => x"ff",
          8380 => x"5c",
          8381 => x"84",
          8382 => x"5c",
          8383 => x"12",
          8384 => x"80",
          8385 => x"78",
          8386 => x"7c",
          8387 => x"90",
          8388 => x"c0",
          8389 => x"90",
          8390 => x"15",
          8391 => x"90",
          8392 => x"54",
          8393 => x"91",
          8394 => x"31",
          8395 => x"84",
          8396 => x"07",
          8397 => x"16",
          8398 => x"73",
          8399 => x"0c",
          8400 => x"04",
          8401 => x"6b",
          8402 => x"05",
          8403 => x"33",
          8404 => x"5a",
          8405 => x"bd",
          8406 => x"80",
          8407 => x"c8",
          8408 => x"f8",
          8409 => x"c8",
          8410 => x"82",
          8411 => x"70",
          8412 => x"74",
          8413 => x"38",
          8414 => x"82",
          8415 => x"81",
          8416 => x"81",
          8417 => x"ff",
          8418 => x"82",
          8419 => x"81",
          8420 => x"81",
          8421 => x"83",
          8422 => x"c0",
          8423 => x"2a",
          8424 => x"51",
          8425 => x"74",
          8426 => x"99",
          8427 => x"53",
          8428 => x"51",
          8429 => x"3f",
          8430 => x"08",
          8431 => x"55",
          8432 => x"92",
          8433 => x"80",
          8434 => x"38",
          8435 => x"06",
          8436 => x"2e",
          8437 => x"48",
          8438 => x"87",
          8439 => x"79",
          8440 => x"78",
          8441 => x"26",
          8442 => x"19",
          8443 => x"74",
          8444 => x"38",
          8445 => x"e4",
          8446 => x"2a",
          8447 => x"70",
          8448 => x"59",
          8449 => x"7a",
          8450 => x"56",
          8451 => x"80",
          8452 => x"51",
          8453 => x"74",
          8454 => x"99",
          8455 => x"53",
          8456 => x"51",
          8457 => x"3f",
          8458 => x"b5",
          8459 => x"ac",
          8460 => x"2a",
          8461 => x"82",
          8462 => x"43",
          8463 => x"83",
          8464 => x"66",
          8465 => x"60",
          8466 => x"90",
          8467 => x"31",
          8468 => x"80",
          8469 => x"8a",
          8470 => x"56",
          8471 => x"26",
          8472 => x"77",
          8473 => x"81",
          8474 => x"74",
          8475 => x"38",
          8476 => x"55",
          8477 => x"83",
          8478 => x"81",
          8479 => x"80",
          8480 => x"38",
          8481 => x"55",
          8482 => x"5e",
          8483 => x"89",
          8484 => x"5a",
          8485 => x"09",
          8486 => x"e1",
          8487 => x"38",
          8488 => x"57",
          8489 => x"b0",
          8490 => x"5a",
          8491 => x"9d",
          8492 => x"26",
          8493 => x"b0",
          8494 => x"10",
          8495 => x"22",
          8496 => x"74",
          8497 => x"38",
          8498 => x"ee",
          8499 => x"66",
          8500 => x"b2",
          8501 => x"c8",
          8502 => x"84",
          8503 => x"89",
          8504 => x"a0",
          8505 => x"82",
          8506 => x"fc",
          8507 => x"56",
          8508 => x"f0",
          8509 => x"80",
          8510 => x"d3",
          8511 => x"38",
          8512 => x"57",
          8513 => x"b0",
          8514 => x"5a",
          8515 => x"9d",
          8516 => x"26",
          8517 => x"b0",
          8518 => x"10",
          8519 => x"22",
          8520 => x"74",
          8521 => x"38",
          8522 => x"ee",
          8523 => x"66",
          8524 => x"d2",
          8525 => x"c8",
          8526 => x"05",
          8527 => x"c8",
          8528 => x"26",
          8529 => x"0b",
          8530 => x"08",
          8531 => x"c8",
          8532 => x"11",
          8533 => x"05",
          8534 => x"83",
          8535 => x"2a",
          8536 => x"a0",
          8537 => x"7d",
          8538 => x"69",
          8539 => x"05",
          8540 => x"72",
          8541 => x"5c",
          8542 => x"59",
          8543 => x"2e",
          8544 => x"89",
          8545 => x"60",
          8546 => x"84",
          8547 => x"5d",
          8548 => x"18",
          8549 => x"68",
          8550 => x"74",
          8551 => x"af",
          8552 => x"31",
          8553 => x"53",
          8554 => x"52",
          8555 => x"d6",
          8556 => x"c8",
          8557 => x"83",
          8558 => x"06",
          8559 => x"b5",
          8560 => x"ff",
          8561 => x"dd",
          8562 => x"83",
          8563 => x"2a",
          8564 => x"be",
          8565 => x"39",
          8566 => x"09",
          8567 => x"c5",
          8568 => x"f5",
          8569 => x"c8",
          8570 => x"38",
          8571 => x"79",
          8572 => x"80",
          8573 => x"38",
          8574 => x"96",
          8575 => x"06",
          8576 => x"2e",
          8577 => x"5e",
          8578 => x"82",
          8579 => x"9f",
          8580 => x"38",
          8581 => x"38",
          8582 => x"81",
          8583 => x"fc",
          8584 => x"ab",
          8585 => x"7d",
          8586 => x"81",
          8587 => x"7d",
          8588 => x"78",
          8589 => x"74",
          8590 => x"8e",
          8591 => x"9c",
          8592 => x"53",
          8593 => x"51",
          8594 => x"3f",
          8595 => x"ae",
          8596 => x"51",
          8597 => x"3f",
          8598 => x"8b",
          8599 => x"a1",
          8600 => x"8d",
          8601 => x"83",
          8602 => x"52",
          8603 => x"ff",
          8604 => x"81",
          8605 => x"34",
          8606 => x"70",
          8607 => x"2a",
          8608 => x"54",
          8609 => x"1b",
          8610 => x"88",
          8611 => x"74",
          8612 => x"26",
          8613 => x"83",
          8614 => x"52",
          8615 => x"ff",
          8616 => x"8a",
          8617 => x"a0",
          8618 => x"a1",
          8619 => x"0b",
          8620 => x"bf",
          8621 => x"51",
          8622 => x"3f",
          8623 => x"9a",
          8624 => x"a0",
          8625 => x"52",
          8626 => x"ff",
          8627 => x"7d",
          8628 => x"81",
          8629 => x"38",
          8630 => x"0a",
          8631 => x"1b",
          8632 => x"ce",
          8633 => x"a4",
          8634 => x"a0",
          8635 => x"52",
          8636 => x"ff",
          8637 => x"81",
          8638 => x"51",
          8639 => x"3f",
          8640 => x"1b",
          8641 => x"8c",
          8642 => x"0b",
          8643 => x"34",
          8644 => x"c2",
          8645 => x"53",
          8646 => x"52",
          8647 => x"51",
          8648 => x"88",
          8649 => x"a7",
          8650 => x"a0",
          8651 => x"83",
          8652 => x"52",
          8653 => x"ff",
          8654 => x"ff",
          8655 => x"1c",
          8656 => x"a6",
          8657 => x"53",
          8658 => x"52",
          8659 => x"ff",
          8660 => x"82",
          8661 => x"83",
          8662 => x"52",
          8663 => x"b4",
          8664 => x"60",
          8665 => x"7e",
          8666 => x"d7",
          8667 => x"82",
          8668 => x"83",
          8669 => x"83",
          8670 => x"06",
          8671 => x"75",
          8672 => x"05",
          8673 => x"7e",
          8674 => x"b7",
          8675 => x"53",
          8676 => x"51",
          8677 => x"3f",
          8678 => x"a4",
          8679 => x"51",
          8680 => x"3f",
          8681 => x"e4",
          8682 => x"e4",
          8683 => x"9f",
          8684 => x"18",
          8685 => x"1b",
          8686 => x"f6",
          8687 => x"83",
          8688 => x"ff",
          8689 => x"82",
          8690 => x"78",
          8691 => x"c4",
          8692 => x"60",
          8693 => x"7a",
          8694 => x"ff",
          8695 => x"75",
          8696 => x"53",
          8697 => x"51",
          8698 => x"3f",
          8699 => x"52",
          8700 => x"9f",
          8701 => x"56",
          8702 => x"83",
          8703 => x"06",
          8704 => x"52",
          8705 => x"9e",
          8706 => x"52",
          8707 => x"ff",
          8708 => x"f0",
          8709 => x"1b",
          8710 => x"87",
          8711 => x"55",
          8712 => x"83",
          8713 => x"74",
          8714 => x"ff",
          8715 => x"7c",
          8716 => x"74",
          8717 => x"38",
          8718 => x"54",
          8719 => x"52",
          8720 => x"99",
          8721 => x"b5",
          8722 => x"87",
          8723 => x"53",
          8724 => x"08",
          8725 => x"ff",
          8726 => x"76",
          8727 => x"31",
          8728 => x"cd",
          8729 => x"58",
          8730 => x"ff",
          8731 => x"55",
          8732 => x"83",
          8733 => x"61",
          8734 => x"26",
          8735 => x"57",
          8736 => x"53",
          8737 => x"51",
          8738 => x"3f",
          8739 => x"08",
          8740 => x"76",
          8741 => x"31",
          8742 => x"db",
          8743 => x"7d",
          8744 => x"38",
          8745 => x"83",
          8746 => x"8a",
          8747 => x"7d",
          8748 => x"38",
          8749 => x"81",
          8750 => x"80",
          8751 => x"80",
          8752 => x"7a",
          8753 => x"bc",
          8754 => x"d5",
          8755 => x"ff",
          8756 => x"83",
          8757 => x"77",
          8758 => x"0b",
          8759 => x"81",
          8760 => x"34",
          8761 => x"34",
          8762 => x"34",
          8763 => x"56",
          8764 => x"52",
          8765 => x"b5",
          8766 => x"0b",
          8767 => x"82",
          8768 => x"82",
          8769 => x"56",
          8770 => x"34",
          8771 => x"08",
          8772 => x"60",
          8773 => x"1b",
          8774 => x"96",
          8775 => x"83",
          8776 => x"ff",
          8777 => x"81",
          8778 => x"7a",
          8779 => x"ff",
          8780 => x"81",
          8781 => x"c8",
          8782 => x"80",
          8783 => x"7e",
          8784 => x"e3",
          8785 => x"82",
          8786 => x"90",
          8787 => x"8e",
          8788 => x"81",
          8789 => x"82",
          8790 => x"56",
          8791 => x"c8",
          8792 => x"0d",
          8793 => x"0d",
          8794 => x"59",
          8795 => x"ff",
          8796 => x"57",
          8797 => x"b4",
          8798 => x"f8",
          8799 => x"81",
          8800 => x"52",
          8801 => x"dc",
          8802 => x"2e",
          8803 => x"9c",
          8804 => x"33",
          8805 => x"2e",
          8806 => x"76",
          8807 => x"58",
          8808 => x"57",
          8809 => x"09",
          8810 => x"38",
          8811 => x"78",
          8812 => x"38",
          8813 => x"82",
          8814 => x"8d",
          8815 => x"f7",
          8816 => x"02",
          8817 => x"05",
          8818 => x"77",
          8819 => x"81",
          8820 => x"8d",
          8821 => x"e7",
          8822 => x"08",
          8823 => x"24",
          8824 => x"17",
          8825 => x"8c",
          8826 => x"77",
          8827 => x"16",
          8828 => x"25",
          8829 => x"3d",
          8830 => x"75",
          8831 => x"52",
          8832 => x"cb",
          8833 => x"76",
          8834 => x"70",
          8835 => x"2a",
          8836 => x"51",
          8837 => x"84",
          8838 => x"19",
          8839 => x"8b",
          8840 => x"f9",
          8841 => x"84",
          8842 => x"56",
          8843 => x"a7",
          8844 => x"fc",
          8845 => x"53",
          8846 => x"75",
          8847 => x"a1",
          8848 => x"c8",
          8849 => x"84",
          8850 => x"2e",
          8851 => x"87",
          8852 => x"08",
          8853 => x"ff",
          8854 => x"b5",
          8855 => x"3d",
          8856 => x"3d",
          8857 => x"80",
          8858 => x"52",
          8859 => x"9a",
          8860 => x"74",
          8861 => x"0d",
          8862 => x"0d",
          8863 => x"05",
          8864 => x"86",
          8865 => x"54",
          8866 => x"73",
          8867 => x"fe",
          8868 => x"51",
          8869 => x"98",
          8870 => x"00",
          8871 => x"ff",
          8872 => x"ff",
          8873 => x"ff",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"64",
          9011 => x"74",
          9012 => x"64",
          9013 => x"74",
          9014 => x"66",
          9015 => x"74",
          9016 => x"66",
          9017 => x"64",
          9018 => x"66",
          9019 => x"63",
          9020 => x"6d",
          9021 => x"61",
          9022 => x"6d",
          9023 => x"79",
          9024 => x"6d",
          9025 => x"66",
          9026 => x"6d",
          9027 => x"70",
          9028 => x"6d",
          9029 => x"6d",
          9030 => x"6d",
          9031 => x"68",
          9032 => x"68",
          9033 => x"68",
          9034 => x"68",
          9035 => x"63",
          9036 => x"00",
          9037 => x"6a",
          9038 => x"72",
          9039 => x"61",
          9040 => x"72",
          9041 => x"74",
          9042 => x"69",
          9043 => x"00",
          9044 => x"74",
          9045 => x"00",
          9046 => x"74",
          9047 => x"69",
          9048 => x"6d",
          9049 => x"69",
          9050 => x"6b",
          9051 => x"00",
          9052 => x"65",
          9053 => x"44",
          9054 => x"20",
          9055 => x"6f",
          9056 => x"49",
          9057 => x"72",
          9058 => x"20",
          9059 => x"6f",
          9060 => x"44",
          9061 => x"20",
          9062 => x"20",
          9063 => x"64",
          9064 => x"4e",
          9065 => x"69",
          9066 => x"66",
          9067 => x"64",
          9068 => x"4e",
          9069 => x"61",
          9070 => x"66",
          9071 => x"64",
          9072 => x"49",
          9073 => x"6c",
          9074 => x"66",
          9075 => x"6e",
          9076 => x"2e",
          9077 => x"41",
          9078 => x"73",
          9079 => x"65",
          9080 => x"64",
          9081 => x"46",
          9082 => x"20",
          9083 => x"65",
          9084 => x"20",
          9085 => x"73",
          9086 => x"00",
          9087 => x"46",
          9088 => x"20",
          9089 => x"64",
          9090 => x"69",
          9091 => x"6c",
          9092 => x"00",
          9093 => x"53",
          9094 => x"73",
          9095 => x"69",
          9096 => x"70",
          9097 => x"65",
          9098 => x"64",
          9099 => x"44",
          9100 => x"65",
          9101 => x"6d",
          9102 => x"20",
          9103 => x"69",
          9104 => x"6c",
          9105 => x"00",
          9106 => x"44",
          9107 => x"20",
          9108 => x"20",
          9109 => x"62",
          9110 => x"2e",
          9111 => x"4e",
          9112 => x"6f",
          9113 => x"74",
          9114 => x"65",
          9115 => x"6c",
          9116 => x"73",
          9117 => x"20",
          9118 => x"6e",
          9119 => x"6e",
          9120 => x"73",
          9121 => x"46",
          9122 => x"61",
          9123 => x"62",
          9124 => x"65",
          9125 => x"54",
          9126 => x"6f",
          9127 => x"20",
          9128 => x"72",
          9129 => x"6f",
          9130 => x"61",
          9131 => x"6c",
          9132 => x"2e",
          9133 => x"46",
          9134 => x"20",
          9135 => x"6c",
          9136 => x"65",
          9137 => x"49",
          9138 => x"66",
          9139 => x"69",
          9140 => x"20",
          9141 => x"6f",
          9142 => x"00",
          9143 => x"54",
          9144 => x"6d",
          9145 => x"20",
          9146 => x"6e",
          9147 => x"6c",
          9148 => x"00",
          9149 => x"50",
          9150 => x"6d",
          9151 => x"72",
          9152 => x"6e",
          9153 => x"72",
          9154 => x"2e",
          9155 => x"53",
          9156 => x"65",
          9157 => x"00",
          9158 => x"55",
          9159 => x"6f",
          9160 => x"65",
          9161 => x"72",
          9162 => x"0a",
          9163 => x"20",
          9164 => x"65",
          9165 => x"73",
          9166 => x"20",
          9167 => x"20",
          9168 => x"65",
          9169 => x"65",
          9170 => x"00",
          9171 => x"72",
          9172 => x"00",
          9173 => x"25",
          9174 => x"58",
          9175 => x"3a",
          9176 => x"25",
          9177 => x"00",
          9178 => x"20",
          9179 => x"20",
          9180 => x"00",
          9181 => x"25",
          9182 => x"00",
          9183 => x"20",
          9184 => x"20",
          9185 => x"7c",
          9186 => x"7a",
          9187 => x"0a",
          9188 => x"25",
          9189 => x"00",
          9190 => x"30",
          9191 => x"35",
          9192 => x"32",
          9193 => x"76",
          9194 => x"32",
          9195 => x"20",
          9196 => x"2c",
          9197 => x"76",
          9198 => x"32",
          9199 => x"25",
          9200 => x"73",
          9201 => x"0a",
          9202 => x"5a",
          9203 => x"49",
          9204 => x"72",
          9205 => x"74",
          9206 => x"6e",
          9207 => x"72",
          9208 => x"54",
          9209 => x"72",
          9210 => x"74",
          9211 => x"75",
          9212 => x"50",
          9213 => x"69",
          9214 => x"72",
          9215 => x"74",
          9216 => x"49",
          9217 => x"4c",
          9218 => x"20",
          9219 => x"65",
          9220 => x"70",
          9221 => x"49",
          9222 => x"4c",
          9223 => x"20",
          9224 => x"65",
          9225 => x"70",
          9226 => x"55",
          9227 => x"30",
          9228 => x"20",
          9229 => x"65",
          9230 => x"70",
          9231 => x"55",
          9232 => x"30",
          9233 => x"20",
          9234 => x"65",
          9235 => x"70",
          9236 => x"55",
          9237 => x"31",
          9238 => x"20",
          9239 => x"65",
          9240 => x"70",
          9241 => x"55",
          9242 => x"31",
          9243 => x"20",
          9244 => x"65",
          9245 => x"70",
          9246 => x"53",
          9247 => x"69",
          9248 => x"75",
          9249 => x"69",
          9250 => x"2e",
          9251 => x"45",
          9252 => x"6c",
          9253 => x"20",
          9254 => x"65",
          9255 => x"2e",
          9256 => x"61",
          9257 => x"65",
          9258 => x"2e",
          9259 => x"00",
          9260 => x"7a",
          9261 => x"68",
          9262 => x"30",
          9263 => x"46",
          9264 => x"65",
          9265 => x"6f",
          9266 => x"69",
          9267 => x"6c",
          9268 => x"20",
          9269 => x"63",
          9270 => x"20",
          9271 => x"70",
          9272 => x"73",
          9273 => x"6e",
          9274 => x"6d",
          9275 => x"61",
          9276 => x"2e",
          9277 => x"2a",
          9278 => x"43",
          9279 => x"72",
          9280 => x"2e",
          9281 => x"00",
          9282 => x"43",
          9283 => x"69",
          9284 => x"2e",
          9285 => x"43",
          9286 => x"61",
          9287 => x"67",
          9288 => x"00",
          9289 => x"25",
          9290 => x"78",
          9291 => x"38",
          9292 => x"3e",
          9293 => x"6c",
          9294 => x"30",
          9295 => x"0a",
          9296 => x"44",
          9297 => x"20",
          9298 => x"6f",
          9299 => x"0a",
          9300 => x"70",
          9301 => x"65",
          9302 => x"25",
          9303 => x"58",
          9304 => x"32",
          9305 => x"3f",
          9306 => x"25",
          9307 => x"58",
          9308 => x"34",
          9309 => x"25",
          9310 => x"58",
          9311 => x"38",
          9312 => x"00",
          9313 => x"45",
          9314 => x"75",
          9315 => x"67",
          9316 => x"64",
          9317 => x"20",
          9318 => x"6c",
          9319 => x"2e",
          9320 => x"43",
          9321 => x"69",
          9322 => x"63",
          9323 => x"20",
          9324 => x"30",
          9325 => x"20",
          9326 => x"0a",
          9327 => x"43",
          9328 => x"20",
          9329 => x"75",
          9330 => x"64",
          9331 => x"64",
          9332 => x"25",
          9333 => x"0a",
          9334 => x"52",
          9335 => x"61",
          9336 => x"6e",
          9337 => x"70",
          9338 => x"63",
          9339 => x"6f",
          9340 => x"2e",
          9341 => x"43",
          9342 => x"20",
          9343 => x"6f",
          9344 => x"6e",
          9345 => x"2e",
          9346 => x"5a",
          9347 => x"62",
          9348 => x"25",
          9349 => x"25",
          9350 => x"73",
          9351 => x"00",
          9352 => x"25",
          9353 => x"25",
          9354 => x"73",
          9355 => x"25",
          9356 => x"25",
          9357 => x"42",
          9358 => x"63",
          9359 => x"61",
          9360 => x"00",
          9361 => x"52",
          9362 => x"69",
          9363 => x"2e",
          9364 => x"45",
          9365 => x"6c",
          9366 => x"20",
          9367 => x"65",
          9368 => x"70",
          9369 => x"2e",
          9370 => x"25",
          9371 => x"64",
          9372 => x"20",
          9373 => x"25",
          9374 => x"64",
          9375 => x"25",
          9376 => x"53",
          9377 => x"43",
          9378 => x"69",
          9379 => x"61",
          9380 => x"6e",
          9381 => x"20",
          9382 => x"6f",
          9383 => x"6f",
          9384 => x"6f",
          9385 => x"67",
          9386 => x"3a",
          9387 => x"76",
          9388 => x"73",
          9389 => x"70",
          9390 => x"65",
          9391 => x"64",
          9392 => x"20",
          9393 => x"57",
          9394 => x"44",
          9395 => x"20",
          9396 => x"30",
          9397 => x"25",
          9398 => x"29",
          9399 => x"20",
          9400 => x"53",
          9401 => x"4d",
          9402 => x"20",
          9403 => x"30",
          9404 => x"25",
          9405 => x"29",
          9406 => x"20",
          9407 => x"49",
          9408 => x"20",
          9409 => x"4d",
          9410 => x"30",
          9411 => x"25",
          9412 => x"29",
          9413 => x"20",
          9414 => x"42",
          9415 => x"20",
          9416 => x"20",
          9417 => x"30",
          9418 => x"25",
          9419 => x"29",
          9420 => x"20",
          9421 => x"52",
          9422 => x"20",
          9423 => x"20",
          9424 => x"30",
          9425 => x"25",
          9426 => x"29",
          9427 => x"20",
          9428 => x"53",
          9429 => x"41",
          9430 => x"20",
          9431 => x"65",
          9432 => x"65",
          9433 => x"25",
          9434 => x"29",
          9435 => x"20",
          9436 => x"54",
          9437 => x"52",
          9438 => x"20",
          9439 => x"69",
          9440 => x"73",
          9441 => x"25",
          9442 => x"29",
          9443 => x"20",
          9444 => x"49",
          9445 => x"20",
          9446 => x"4c",
          9447 => x"68",
          9448 => x"65",
          9449 => x"25",
          9450 => x"29",
          9451 => x"20",
          9452 => x"57",
          9453 => x"42",
          9454 => x"20",
          9455 => x"0a",
          9456 => x"20",
          9457 => x"57",
          9458 => x"32",
          9459 => x"20",
          9460 => x"49",
          9461 => x"4c",
          9462 => x"20",
          9463 => x"50",
          9464 => x"00",
          9465 => x"20",
          9466 => x"53",
          9467 => x"00",
          9468 => x"41",
          9469 => x"65",
          9470 => x"73",
          9471 => x"20",
          9472 => x"43",
          9473 => x"52",
          9474 => x"74",
          9475 => x"63",
          9476 => x"20",
          9477 => x"72",
          9478 => x"20",
          9479 => x"30",
          9480 => x"00",
          9481 => x"20",
          9482 => x"43",
          9483 => x"4d",
          9484 => x"72",
          9485 => x"74",
          9486 => x"20",
          9487 => x"72",
          9488 => x"20",
          9489 => x"30",
          9490 => x"00",
          9491 => x"20",
          9492 => x"53",
          9493 => x"6b",
          9494 => x"61",
          9495 => x"41",
          9496 => x"65",
          9497 => x"20",
          9498 => x"20",
          9499 => x"30",
          9500 => x"00",
          9501 => x"4d",
          9502 => x"3a",
          9503 => x"20",
          9504 => x"5a",
          9505 => x"49",
          9506 => x"20",
          9507 => x"20",
          9508 => x"20",
          9509 => x"20",
          9510 => x"20",
          9511 => x"30",
          9512 => x"00",
          9513 => x"20",
          9514 => x"53",
          9515 => x"65",
          9516 => x"6c",
          9517 => x"20",
          9518 => x"71",
          9519 => x"20",
          9520 => x"20",
          9521 => x"64",
          9522 => x"34",
          9523 => x"7a",
          9524 => x"20",
          9525 => x"53",
          9526 => x"4d",
          9527 => x"6f",
          9528 => x"46",
          9529 => x"20",
          9530 => x"20",
          9531 => x"20",
          9532 => x"64",
          9533 => x"34",
          9534 => x"7a",
          9535 => x"20",
          9536 => x"57",
          9537 => x"62",
          9538 => x"20",
          9539 => x"41",
          9540 => x"6c",
          9541 => x"20",
          9542 => x"71",
          9543 => x"64",
          9544 => x"34",
          9545 => x"7a",
          9546 => x"53",
          9547 => x"6c",
          9548 => x"4d",
          9549 => x"75",
          9550 => x"46",
          9551 => x"00",
          9552 => x"45",
          9553 => x"45",
          9554 => x"69",
          9555 => x"55",
          9556 => x"6f",
          9557 => x"00",
          9558 => x"01",
          9559 => x"00",
          9560 => x"00",
          9561 => x"01",
          9562 => x"00",
          9563 => x"00",
          9564 => x"01",
          9565 => x"00",
          9566 => x"00",
          9567 => x"01",
          9568 => x"00",
          9569 => x"00",
          9570 => x"01",
          9571 => x"00",
          9572 => x"00",
          9573 => x"01",
          9574 => x"00",
          9575 => x"00",
          9576 => x"01",
          9577 => x"00",
          9578 => x"00",
          9579 => x"01",
          9580 => x"00",
          9581 => x"00",
          9582 => x"01",
          9583 => x"00",
          9584 => x"00",
          9585 => x"01",
          9586 => x"00",
          9587 => x"00",
          9588 => x"01",
          9589 => x"00",
          9590 => x"00",
          9591 => x"04",
          9592 => x"00",
          9593 => x"00",
          9594 => x"04",
          9595 => x"00",
          9596 => x"00",
          9597 => x"04",
          9598 => x"00",
          9599 => x"00",
          9600 => x"03",
          9601 => x"00",
          9602 => x"00",
          9603 => x"04",
          9604 => x"00",
          9605 => x"00",
          9606 => x"04",
          9607 => x"00",
          9608 => x"00",
          9609 => x"04",
          9610 => x"00",
          9611 => x"00",
          9612 => x"03",
          9613 => x"00",
          9614 => x"00",
          9615 => x"03",
          9616 => x"00",
          9617 => x"00",
          9618 => x"03",
          9619 => x"00",
          9620 => x"00",
          9621 => x"03",
          9622 => x"00",
          9623 => x"1b",
          9624 => x"1b",
          9625 => x"1b",
          9626 => x"1b",
          9627 => x"1b",
          9628 => x"1b",
          9629 => x"1b",
          9630 => x"1b",
          9631 => x"1b",
          9632 => x"1b",
          9633 => x"1b",
          9634 => x"10",
          9635 => x"0e",
          9636 => x"0d",
          9637 => x"0b",
          9638 => x"08",
          9639 => x"06",
          9640 => x"05",
          9641 => x"04",
          9642 => x"03",
          9643 => x"02",
          9644 => x"01",
          9645 => x"68",
          9646 => x"6f",
          9647 => x"68",
          9648 => x"00",
          9649 => x"21",
          9650 => x"25",
          9651 => x"75",
          9652 => x"73",
          9653 => x"46",
          9654 => x"65",
          9655 => x"6f",
          9656 => x"73",
          9657 => x"74",
          9658 => x"68",
          9659 => x"6f",
          9660 => x"66",
          9661 => x"20",
          9662 => x"45",
          9663 => x"00",
          9664 => x"43",
          9665 => x"6f",
          9666 => x"70",
          9667 => x"63",
          9668 => x"74",
          9669 => x"69",
          9670 => x"72",
          9671 => x"69",
          9672 => x"20",
          9673 => x"61",
          9674 => x"6e",
          9675 => x"53",
          9676 => x"22",
          9677 => x"3a",
          9678 => x"3e",
          9679 => x"7c",
          9680 => x"46",
          9681 => x"46",
          9682 => x"32",
          9683 => x"eb",
          9684 => x"53",
          9685 => x"35",
          9686 => x"4e",
          9687 => x"41",
          9688 => x"20",
          9689 => x"41",
          9690 => x"20",
          9691 => x"4e",
          9692 => x"41",
          9693 => x"20",
          9694 => x"41",
          9695 => x"20",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"80",
          9701 => x"8e",
          9702 => x"45",
          9703 => x"49",
          9704 => x"90",
          9705 => x"99",
          9706 => x"59",
          9707 => x"9c",
          9708 => x"41",
          9709 => x"a5",
          9710 => x"a8",
          9711 => x"ac",
          9712 => x"b0",
          9713 => x"b4",
          9714 => x"b8",
          9715 => x"bc",
          9716 => x"c0",
          9717 => x"c4",
          9718 => x"c8",
          9719 => x"cc",
          9720 => x"d0",
          9721 => x"d4",
          9722 => x"d8",
          9723 => x"dc",
          9724 => x"e0",
          9725 => x"e4",
          9726 => x"e8",
          9727 => x"ec",
          9728 => x"f0",
          9729 => x"f4",
          9730 => x"f8",
          9731 => x"fc",
          9732 => x"2b",
          9733 => x"3d",
          9734 => x"5c",
          9735 => x"3c",
          9736 => x"7f",
          9737 => x"00",
          9738 => x"00",
          9739 => x"01",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"01",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"01",
          9752 => x"00",
          9753 => x"00",
          9754 => x"00",
          9755 => x"01",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"01",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"01",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"01",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"01",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"01",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"01",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"01",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"01",
          9788 => x"00",
          9789 => x"00",
          9790 => x"00",
          9791 => x"01",
          9792 => x"00",
          9793 => x"00",
          9794 => x"00",
          9795 => x"01",
          9796 => x"00",
          9797 => x"00",
          9798 => x"00",
          9799 => x"01",
          9800 => x"00",
          9801 => x"00",
          9802 => x"00",
          9803 => x"01",
          9804 => x"00",
          9805 => x"00",
          9806 => x"00",
          9807 => x"01",
          9808 => x"00",
          9809 => x"00",
          9810 => x"00",
          9811 => x"01",
          9812 => x"00",
          9813 => x"00",
          9814 => x"00",
          9815 => x"01",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"01",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"01",
          9824 => x"00",
          9825 => x"00",
          9826 => x"00",
          9827 => x"01",
          9828 => x"00",
          9829 => x"00",
          9830 => x"00",
          9831 => x"01",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"01",
          9836 => x"00",
          9837 => x"00",
          9838 => x"00",
          9839 => x"01",
          9840 => x"00",
          9841 => x"00",
          9842 => x"00",
          9843 => x"01",
          9844 => x"00",
          9845 => x"00",
          9846 => x"00",
          9847 => x"01",
          9848 => x"00",
          9849 => x"00",
          9850 => x"00",
          9851 => x"00",
          9852 => x"00",
          9853 => x"00",
          9854 => x"00",
          9855 => x"00",
          9856 => x"00",
          9857 => x"00",
          9858 => x"00",
          9859 => x"01",
          9860 => x"01",
          9861 => x"00",
          9862 => x"00",
          9863 => x"00",
          9864 => x"00",
          9865 => x"05",
          9866 => x"05",
          9867 => x"05",
          9868 => x"00",
          9869 => x"01",
          9870 => x"01",
          9871 => x"01",
          9872 => x"01",
          9873 => x"00",
          9874 => x"00",
          9875 => x"00",
          9876 => x"00",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"00",
          9881 => x"00",
          9882 => x"00",
          9883 => x"00",
          9884 => x"00",
          9885 => x"00",
          9886 => x"00",
          9887 => x"00",
          9888 => x"00",
          9889 => x"00",
          9890 => x"00",
          9891 => x"00",
          9892 => x"00",
          9893 => x"00",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"00",
          9898 => x"01",
          9899 => x"00",
          9900 => x"01",
          9901 => x"00",
          9902 => x"02",
          9903 => x"00",
          9904 => x"00",
          9905 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
