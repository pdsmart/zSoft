-- Byte Addressed 32bit/64bit BRAM module for the ZPU Evo implementation.
--
-- This template provides a 32bit wide bus on port A and a 64bit bus
-- on port B. This is typically used for the ZPU Boot BRAM where port B
-- is used exclusively for instruction storage.
--
-- Copyright 2018-2021 - Philip Smart for the ZPU Evo implementation.
-- History:
--   20190618  - Initial 32 bit dual port BRAM described by inference rather than
--               using an IP Megacore. This was to make it more portable but also
--               to allow 8/16/32 bit writes to the memory.
--   20210108  - Updated to 64bit on Port B to allow for the 64bit decoder on the ZPU.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.softZPU_pkg.all;

entity DualPort3264BootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 3);
        memBWrite            : in  std_logic_vector(WORD_64BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_64BIT_RANGE)
    );
end DualPort3264BootBRAM;

architecture arch of DualPort3264BootBRAM is

    -- Declare 8 byte wide arrays for byte level addressing.
    type ramArray is array(natural range 0 to (2**(addrbits-3))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"fa",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"05",
            10 => x"52",
            11 => x"00",
            12 => x"08",
            13 => x"81",
            14 => x"06",
            15 => x"0b",
            16 => x"05",
            17 => x"06",
            18 => x"06",
            19 => x"00",
            20 => x"73",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"09",
            25 => x"72",
            26 => x"31",
            27 => x"51",
            28 => x"73",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"93",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"2b",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"06",
            45 => x"b0",
            46 => x"00",
            47 => x"00",
            48 => x"ff",
            49 => x"0a",
            50 => x"51",
            51 => x"00",
            52 => x"51",
            53 => x"05",
            54 => x"72",
            55 => x"00",
            56 => x"05",
            57 => x"06",
            58 => x"00",
            59 => x"00",
            60 => x"05",
            61 => x"06",
            62 => x"00",
            63 => x"00",
            64 => x"05",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"81",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"06",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"08",
            77 => x"05",
            78 => x"52",
            79 => x"00",
            80 => x"08",
            81 => x"06",
            82 => x"0b",
            83 => x"00",
            84 => x"08",
            85 => x"ac",
            86 => x"90",
            87 => x"00",
            88 => x"08",
            89 => x"ab",
            90 => x"90",
            91 => x"00",
            92 => x"81",
            93 => x"05",
            94 => x"74",
            95 => x"51",
            96 => x"81",
            97 => x"ff",
            98 => x"72",
            99 => x"51",
           100 => x"04",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"52",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"72",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"ff",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"8c",
           133 => x"04",
           134 => x"0b",
           135 => x"8c",
           136 => x"04",
           137 => x"0b",
           138 => x"8c",
           139 => x"04",
           140 => x"0b",
           141 => x"8d",
           142 => x"04",
           143 => x"0b",
           144 => x"8d",
           145 => x"04",
           146 => x"0b",
           147 => x"8e",
           148 => x"04",
           149 => x"0b",
           150 => x"8f",
           151 => x"04",
           152 => x"0b",
           153 => x"8f",
           154 => x"04",
           155 => x"0b",
           156 => x"90",
           157 => x"04",
           158 => x"0b",
           159 => x"90",
           160 => x"04",
           161 => x"0b",
           162 => x"91",
           163 => x"04",
           164 => x"0b",
           165 => x"91",
           166 => x"04",
           167 => x"0b",
           168 => x"92",
           169 => x"04",
           170 => x"0b",
           171 => x"92",
           172 => x"04",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"81",
           193 => x"87",
           194 => x"80",
           195 => x"ee",
           196 => x"80",
           197 => x"f3",
           198 => x"80",
           199 => x"e0",
           200 => x"80",
           201 => x"a3",
           202 => x"80",
           203 => x"f6",
           204 => x"80",
           205 => x"86",
           206 => x"80",
           207 => x"82",
           208 => x"80",
           209 => x"88",
           210 => x"80",
           211 => x"a8",
           212 => x"80",
           213 => x"d1",
           214 => x"80",
           215 => x"8a",
           216 => x"80",
           217 => x"d4",
           218 => x"c0",
           219 => x"80",
           220 => x"80",
           221 => x"0c",
           222 => x"08",
           223 => x"d4",
           224 => x"d4",
           225 => x"b9",
           226 => x"b9",
           227 => x"84",
           228 => x"84",
           229 => x"04",
           230 => x"2d",
           231 => x"90",
           232 => x"c0",
           233 => x"80",
           234 => x"ed",
           235 => x"c0",
           236 => x"82",
           237 => x"80",
           238 => x"0c",
           239 => x"08",
           240 => x"d4",
           241 => x"d4",
           242 => x"b9",
           243 => x"b9",
           244 => x"84",
           245 => x"84",
           246 => x"04",
           247 => x"2d",
           248 => x"90",
           249 => x"e7",
           250 => x"80",
           251 => x"8b",
           252 => x"c0",
           253 => x"82",
           254 => x"80",
           255 => x"0c",
           256 => x"08",
           257 => x"d4",
           258 => x"d4",
           259 => x"b9",
           260 => x"b9",
           261 => x"84",
           262 => x"84",
           263 => x"04",
           264 => x"2d",
           265 => x"90",
           266 => x"a7",
           267 => x"80",
           268 => x"96",
           269 => x"c0",
           270 => x"83",
           271 => x"80",
           272 => x"0c",
           273 => x"08",
           274 => x"d4",
           275 => x"d4",
           276 => x"b9",
           277 => x"b9",
           278 => x"84",
           279 => x"84",
           280 => x"04",
           281 => x"2d",
           282 => x"90",
           283 => x"e3",
           284 => x"80",
           285 => x"f4",
           286 => x"c0",
           287 => x"81",
           288 => x"80",
           289 => x"0c",
           290 => x"08",
           291 => x"d4",
           292 => x"d4",
           293 => x"b9",
           294 => x"b9",
           295 => x"84",
           296 => x"b9",
           297 => x"84",
           298 => x"84",
           299 => x"04",
           300 => x"2d",
           301 => x"90",
           302 => x"bd",
           303 => x"80",
           304 => x"d5",
           305 => x"c0",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"00",
           311 => x"06",
           312 => x"10",
           313 => x"51",
           314 => x"ff",
           315 => x"52",
           316 => x"38",
           317 => x"c8",
           318 => x"80",
           319 => x"0b",
           320 => x"80",
           321 => x"87",
           322 => x"56",
           323 => x"51",
           324 => x"fa",
           325 => x"33",
           326 => x"07",
           327 => x"72",
           328 => x"ff",
           329 => x"70",
           330 => x"56",
           331 => x"80",
           332 => x"3f",
           333 => x"c8",
           334 => x"c8",
           335 => x"ff",
           336 => x"72",
           337 => x"73",
           338 => x"76",
           339 => x"3d",
           340 => x"0c",
           341 => x"7d",
           342 => x"34",
           343 => x"88",
           344 => x"05",
           345 => x"74",
           346 => x"0d",
           347 => x"75",
           348 => x"f1",
           349 => x"5d",
           350 => x"33",
           351 => x"55",
           352 => x"09",
           353 => x"57",
           354 => x"1c",
           355 => x"2e",
           356 => x"89",
           357 => x"70",
           358 => x"78",
           359 => x"7a",
           360 => x"40",
           361 => x"82",
           362 => x"ff",
           363 => x"84",
           364 => x"7a",
           365 => x"79",
           366 => x"2c",
           367 => x"0a",
           368 => x"56",
           369 => x"73",
           370 => x"78",
           371 => x"38",
           372 => x"81",
           373 => x"5a",
           374 => x"fe",
           375 => x"76",
           376 => x"76",
           377 => x"83",
           378 => x"8a",
           379 => x"7e",
           380 => x"d8",
           381 => x"ca",
           382 => x"e0",
           383 => x"eb",
           384 => x"3f",
           385 => x"86",
           386 => x"fe",
           387 => x"05",
           388 => x"5e",
           389 => x"79",
           390 => x"b9",
           391 => x"c8",
           392 => x"89",
           393 => x"b0",
           394 => x"40",
           395 => x"3f",
           396 => x"c8",
           397 => x"31",
           398 => x"7e",
           399 => x"80",
           400 => x"2c",
           401 => x"06",
           402 => x"77",
           403 => x"05",
           404 => x"84",
           405 => x"53",
           406 => x"70",
           407 => x"9e",
           408 => x"06",
           409 => x"38",
           410 => x"2a",
           411 => x"81",
           412 => x"38",
           413 => x"2c",
           414 => x"73",
           415 => x"2a",
           416 => x"7a",
           417 => x"98",
           418 => x"73",
           419 => x"73",
           420 => x"06",
           421 => x"78",
           422 => x"05",
           423 => x"74",
           424 => x"88",
           425 => x"29",
           426 => x"5a",
           427 => x"74",
           428 => x"38",
           429 => x"ff",
           430 => x"55",
           431 => x"b0",
           432 => x"80",
           433 => x"98",
           434 => x"e5",
           435 => x"5c",
           436 => x"76",
           437 => x"80",
           438 => x"d3",
           439 => x"d8",
           440 => x"70",
           441 => x"84",
           442 => x"38",
           443 => x"fc",
           444 => x"29",
           445 => x"5a",
           446 => x"38",
           447 => x"e2",
           448 => x"07",
           449 => x"38",
           450 => x"5b",
           451 => x"05",
           452 => x"5f",
           453 => x"7f",
           454 => x"06",
           455 => x"07",
           456 => x"80",
           457 => x"56",
           458 => x"81",
           459 => x"77",
           460 => x"80",
           461 => x"80",
           462 => x"a0",
           463 => x"1a",
           464 => x"79",
           465 => x"7c",
           466 => x"51",
           467 => x"70",
           468 => x"83",
           469 => x"52",
           470 => x"85",
           471 => x"06",
           472 => x"80",
           473 => x"2c",
           474 => x"2a",
           475 => x"fd",
           476 => x"84",
           477 => x"56",
           478 => x"83",
           479 => x"5e",
           480 => x"33",
           481 => x"ca",
           482 => x"33",
           483 => x"ba",
           484 => x"77",
           485 => x"82",
           486 => x"84",
           487 => x"78",
           488 => x"90",
           489 => x"c0",
           490 => x"be",
           491 => x"05",
           492 => x"41",
           493 => x"87",
           494 => x"ff",
           495 => x"54",
           496 => x"7c",
           497 => x"f7",
           498 => x"29",
           499 => x"5a",
           500 => x"38",
           501 => x"e2",
           502 => x"3f",
           503 => x"e3",
           504 => x"3f",
           505 => x"80",
           506 => x"75",
           507 => x"70",
           508 => x"5a",
           509 => x"a2",
           510 => x"3f",
           511 => x"fa",
           512 => x"75",
           513 => x"81",
           514 => x"38",
           515 => x"2b",
           516 => x"39",
           517 => x"c8",
           518 => x"3f",
           519 => x"88",
           520 => x"ff",
           521 => x"54",
           522 => x"7e",
           523 => x"57",
           524 => x"84",
           525 => x"51",
           526 => x"fa",
           527 => x"d5",
           528 => x"2a",
           529 => x"58",
           530 => x"09",
           531 => x"81",
           532 => x"b0",
           533 => x"51",
           534 => x"b9",
           535 => x"57",
           536 => x"72",
           537 => x"08",
           538 => x"54",
           539 => x"90",
           540 => x"c8",
           541 => x"76",
           542 => x"3d",
           543 => x"56",
           544 => x"81",
           545 => x"55",
           546 => x"09",
           547 => x"05",
           548 => x"81",
           549 => x"b9",
           550 => x"70",
           551 => x"2e",
           552 => x"15",
           553 => x"08",
           554 => x"81",
           555 => x"38",
           556 => x"ac",
           557 => x"3d",
           558 => x"85",
           559 => x"81",
           560 => x"72",
           561 => x"54",
           562 => x"08",
           563 => x"38",
           564 => x"08",
           565 => x"53",
           566 => x"75",
           567 => x"04",
           568 => x"90",
           569 => x"84",
           570 => x"08",
           571 => x"d7",
           572 => x"33",
           573 => x"81",
           574 => x"71",
           575 => x"52",
           576 => x"06",
           577 => x"75",
           578 => x"2e",
           579 => x"8c",
           580 => x"71",
           581 => x"c8",
           582 => x"bf",
           583 => x"16",
           584 => x"16",
           585 => x"0d",
           586 => x"74",
           587 => x"b9",
           588 => x"85",
           589 => x"84",
           590 => x"71",
           591 => x"ff",
           592 => x"3d",
           593 => x"85",
           594 => x"3d",
           595 => x"71",
           596 => x"f7",
           597 => x"05",
           598 => x"05",
           599 => x"b9",
           600 => x"3d",
           601 => x"52",
           602 => x"72",
           603 => x"38",
           604 => x"70",
           605 => x"70",
           606 => x"86",
           607 => x"75",
           608 => x"53",
           609 => x"33",
           610 => x"2e",
           611 => x"53",
           612 => x"70",
           613 => x"74",
           614 => x"53",
           615 => x"70",
           616 => x"84",
           617 => x"77",
           618 => x"05",
           619 => x"05",
           620 => x"b9",
           621 => x"3d",
           622 => x"52",
           623 => x"70",
           624 => x"05",
           625 => x"38",
           626 => x"0d",
           627 => x"55",
           628 => x"73",
           629 => x"52",
           630 => x"9a",
           631 => x"b7",
           632 => x"80",
           633 => x"3d",
           634 => x"73",
           635 => x"e9",
           636 => x"71",
           637 => x"84",
           638 => x"71",
           639 => x"04",
           640 => x"52",
           641 => x"08",
           642 => x"55",
           643 => x"08",
           644 => x"9b",
           645 => x"80",
           646 => x"b9",
           647 => x"b9",
           648 => x"0c",
           649 => x"75",
           650 => x"71",
           651 => x"05",
           652 => x"38",
           653 => x"81",
           654 => x"31",
           655 => x"85",
           656 => x"77",
           657 => x"80",
           658 => x"05",
           659 => x"38",
           660 => x"0d",
           661 => x"54",
           662 => x"76",
           663 => x"08",
           664 => x"8d",
           665 => x"84",
           666 => x"72",
           667 => x"72",
           668 => x"74",
           669 => x"2b",
           670 => x"76",
           671 => x"2a",
           672 => x"31",
           673 => x"7b",
           674 => x"5c",
           675 => x"74",
           676 => x"71",
           677 => x"04",
           678 => x"80",
           679 => x"25",
           680 => x"71",
           681 => x"30",
           682 => x"31",
           683 => x"70",
           684 => x"71",
           685 => x"1b",
           686 => x"80",
           687 => x"2a",
           688 => x"06",
           689 => x"19",
           690 => x"54",
           691 => x"55",
           692 => x"58",
           693 => x"fd",
           694 => x"53",
           695 => x"c8",
           696 => x"b9",
           697 => x"fa",
           698 => x"53",
           699 => x"fe",
           700 => x"e0",
           701 => x"73",
           702 => x"c8",
           703 => x"26",
           704 => x"2e",
           705 => x"a0",
           706 => x"54",
           707 => x"38",
           708 => x"10",
           709 => x"9f",
           710 => x"75",
           711 => x"52",
           712 => x"72",
           713 => x"04",
           714 => x"9f",
           715 => x"9f",
           716 => x"74",
           717 => x"56",
           718 => x"b9",
           719 => x"b9",
           720 => x"3d",
           721 => x"7b",
           722 => x"59",
           723 => x"38",
           724 => x"55",
           725 => x"ad",
           726 => x"81",
           727 => x"77",
           728 => x"80",
           729 => x"80",
           730 => x"70",
           731 => x"70",
           732 => x"27",
           733 => x"06",
           734 => x"38",
           735 => x"76",
           736 => x"70",
           737 => x"ff",
           738 => x"75",
           739 => x"75",
           740 => x"04",
           741 => x"33",
           742 => x"81",
           743 => x"78",
           744 => x"e2",
           745 => x"f8",
           746 => x"27",
           747 => x"88",
           748 => x"75",
           749 => x"04",
           750 => x"70",
           751 => x"39",
           752 => x"3d",
           753 => x"5b",
           754 => x"70",
           755 => x"09",
           756 => x"78",
           757 => x"2e",
           758 => x"38",
           759 => x"14",
           760 => x"db",
           761 => x"27",
           762 => x"89",
           763 => x"55",
           764 => x"51",
           765 => x"13",
           766 => x"73",
           767 => x"81",
           768 => x"16",
           769 => x"56",
           770 => x"80",
           771 => x"7a",
           772 => x"0c",
           773 => x"70",
           774 => x"73",
           775 => x"38",
           776 => x"55",
           777 => x"90",
           778 => x"81",
           779 => x"14",
           780 => x"27",
           781 => x"0c",
           782 => x"15",
           783 => x"80",
           784 => x"b9",
           785 => x"d6",
           786 => x"ff",
           787 => x"3d",
           788 => x"38",
           789 => x"52",
           790 => x"ef",
           791 => x"ce",
           792 => x"0d",
           793 => x"3f",
           794 => x"51",
           795 => x"83",
           796 => x"3d",
           797 => x"87",
           798 => x"a4",
           799 => x"04",
           800 => x"83",
           801 => x"ee",
           802 => x"cf",
           803 => x"0d",
           804 => x"3f",
           805 => x"51",
           806 => x"83",
           807 => x"3d",
           808 => x"af",
           809 => x"e4",
           810 => x"04",
           811 => x"83",
           812 => x"ee",
           813 => x"d1",
           814 => x"0d",
           815 => x"3f",
           816 => x"51",
           817 => x"83",
           818 => x"3d",
           819 => x"84",
           820 => x"80",
           821 => x"25",
           822 => x"87",
           823 => x"77",
           824 => x"93",
           825 => x"77",
           826 => x"95",
           827 => x"84",
           828 => x"38",
           829 => x"30",
           830 => x"70",
           831 => x"58",
           832 => x"98",
           833 => x"80",
           834 => x"29",
           835 => x"08",
           836 => x"83",
           837 => x"84",
           838 => x"84",
           839 => x"0c",
           840 => x"d4",
           841 => x"77",
           842 => x"c8",
           843 => x"88",
           844 => x"80",
           845 => x"d5",
           846 => x"b1",
           847 => x"51",
           848 => x"54",
           849 => x"d1",
           850 => x"39",
           851 => x"b7",
           852 => x"53",
           853 => x"84",
           854 => x"2e",
           855 => x"77",
           856 => x"04",
           857 => x"55",
           858 => x"52",
           859 => x"08",
           860 => x"04",
           861 => x"8c",
           862 => x"15",
           863 => x"5e",
           864 => x"52",
           865 => x"83",
           866 => x"54",
           867 => x"2e",
           868 => x"a8",
           869 => x"81",
           870 => x"88",
           871 => x"d5",
           872 => x"aa",
           873 => x"d2",
           874 => x"75",
           875 => x"70",
           876 => x"27",
           877 => x"74",
           878 => x"06",
           879 => x"80",
           880 => x"81",
           881 => x"a0",
           882 => x"78",
           883 => x"51",
           884 => x"5c",
           885 => x"b9",
           886 => x"58",
           887 => x"76",
           888 => x"57",
           889 => x"0b",
           890 => x"04",
           891 => x"81",
           892 => x"a0",
           893 => x"fe",
           894 => x"a8",
           895 => x"d5",
           896 => x"ea",
           897 => x"73",
           898 => x"72",
           899 => x"ec",
           900 => x"53",
           901 => x"74",
           902 => x"d2",
           903 => x"84",
           904 => x"ea",
           905 => x"38",
           906 => x"38",
           907 => x"db",
           908 => x"08",
           909 => x"78",
           910 => x"84",
           911 => x"f2",
           912 => x"80",
           913 => x"81",
           914 => x"2e",
           915 => x"d0",
           916 => x"90",
           917 => x"c0",
           918 => x"70",
           919 => x"72",
           920 => x"73",
           921 => x"57",
           922 => x"38",
           923 => x"c8",
           924 => x"a0",
           925 => x"30",
           926 => x"51",
           927 => x"73",
           928 => x"80",
           929 => x"0d",
           930 => x"80",
           931 => x"9d",
           932 => x"99",
           933 => x"81",
           934 => x"82",
           935 => x"06",
           936 => x"83",
           937 => x"81",
           938 => x"06",
           939 => x"85",
           940 => x"80",
           941 => x"06",
           942 => x"87",
           943 => x"a9",
           944 => x"72",
           945 => x"0d",
           946 => x"d3",
           947 => x"9c",
           948 => x"0d",
           949 => x"d3",
           950 => x"9b",
           951 => x"53",
           952 => x"81",
           953 => x"51",
           954 => x"3f",
           955 => x"52",
           956 => x"39",
           957 => x"94",
           958 => x"b1",
           959 => x"51",
           960 => x"ff",
           961 => x"83",
           962 => x"51",
           963 => x"81",
           964 => x"c2",
           965 => x"f9",
           966 => x"3f",
           967 => x"2a",
           968 => x"2e",
           969 => x"51",
           970 => x"9a",
           971 => x"72",
           972 => x"71",
           973 => x"39",
           974 => x"e0",
           975 => x"a9",
           976 => x"51",
           977 => x"ff",
           978 => x"41",
           979 => x"42",
           980 => x"3f",
           981 => x"9b",
           982 => x"b1",
           983 => x"3f",
           984 => x"d6",
           985 => x"80",
           986 => x"0b",
           987 => x"06",
           988 => x"38",
           989 => x"81",
           990 => x"c1",
           991 => x"2e",
           992 => x"a0",
           993 => x"1a",
           994 => x"f6",
           995 => x"38",
           996 => x"70",
           997 => x"b9",
           998 => x"7a",
           999 => x"3f",
          1000 => x"1b",
          1001 => x"38",
          1002 => x"5b",
          1003 => x"33",
          1004 => x"80",
          1005 => x"84",
          1006 => x"08",
          1007 => x"c8",
          1008 => x"51",
          1009 => x"60",
          1010 => x"81",
          1011 => x"e7",
          1012 => x"26",
          1013 => x"5e",
          1014 => x"7a",
          1015 => x"2e",
          1016 => x"83",
          1017 => x"3f",
          1018 => x"57",
          1019 => x"80",
          1020 => x"51",
          1021 => x"84",
          1022 => x"72",
          1023 => x"80",
          1024 => x"5a",
          1025 => x"8d",
          1026 => x"5c",
          1027 => x"32",
          1028 => x"ee",
          1029 => x"7d",
          1030 => x"ec",
          1031 => x"f8",
          1032 => x"3f",
          1033 => x"81",
          1034 => x"38",
          1035 => x"d0",
          1036 => x"b9",
          1037 => x"0b",
          1038 => x"d8",
          1039 => x"f6",
          1040 => x"2e",
          1041 => x"df",
          1042 => x"33",
          1043 => x"82",
          1044 => x"91",
          1045 => x"d4",
          1046 => x"bc",
          1047 => x"52",
          1048 => x"5a",
          1049 => x"7c",
          1050 => x"78",
          1051 => x"10",
          1052 => x"08",
          1053 => x"7e",
          1054 => x"52",
          1055 => x"3f",
          1056 => x"81",
          1057 => x"3d",
          1058 => x"d5",
          1059 => x"81",
          1060 => x"d6",
          1061 => x"54",
          1062 => x"51",
          1063 => x"8c",
          1064 => x"3f",
          1065 => x"bf",
          1066 => x"d6",
          1067 => x"51",
          1068 => x"83",
          1069 => x"fd",
          1070 => x"84",
          1071 => x"8a",
          1072 => x"fa",
          1073 => x"51",
          1074 => x"84",
          1075 => x"38",
          1076 => x"f0",
          1077 => x"b8",
          1078 => x"05",
          1079 => x"08",
          1080 => x"83",
          1081 => x"59",
          1082 => x"53",
          1083 => x"84",
          1084 => x"38",
          1085 => x"80",
          1086 => x"c8",
          1087 => x"08",
          1088 => x"d0",
          1089 => x"80",
          1090 => x"7e",
          1091 => x"f9",
          1092 => x"38",
          1093 => x"39",
          1094 => x"80",
          1095 => x"c8",
          1096 => x"3d",
          1097 => x"51",
          1098 => x"86",
          1099 => x"78",
          1100 => x"3f",
          1101 => x"52",
          1102 => x"7e",
          1103 => x"38",
          1104 => x"82",
          1105 => x"3d",
          1106 => x"51",
          1107 => x"80",
          1108 => x"fc",
          1109 => x"da",
          1110 => x"f8",
          1111 => x"53",
          1112 => x"84",
          1113 => x"38",
          1114 => x"68",
          1115 => x"8d",
          1116 => x"5c",
          1117 => x"55",
          1118 => x"83",
          1119 => x"66",
          1120 => x"59",
          1121 => x"53",
          1122 => x"84",
          1123 => x"38",
          1124 => x"80",
          1125 => x"c8",
          1126 => x"3d",
          1127 => x"51",
          1128 => x"80",
          1129 => x"51",
          1130 => x"27",
          1131 => x"81",
          1132 => x"05",
          1133 => x"11",
          1134 => x"3f",
          1135 => x"c3",
          1136 => x"ff",
          1137 => x"b9",
          1138 => x"54",
          1139 => x"3f",
          1140 => x"52",
          1141 => x"7e",
          1142 => x"38",
          1143 => x"81",
          1144 => x"80",
          1145 => x"05",
          1146 => x"ff",
          1147 => x"b9",
          1148 => x"68",
          1149 => x"34",
          1150 => x"fc",
          1151 => x"8a",
          1152 => x"38",
          1153 => x"11",
          1154 => x"3f",
          1155 => x"a3",
          1156 => x"ff",
          1157 => x"b9",
          1158 => x"b8",
          1159 => x"05",
          1160 => x"08",
          1161 => x"83",
          1162 => x"67",
          1163 => x"65",
          1164 => x"0c",
          1165 => x"d9",
          1166 => x"ff",
          1167 => x"b9",
          1168 => x"52",
          1169 => x"b9",
          1170 => x"3f",
          1171 => x"a3",
          1172 => x"f6",
          1173 => x"84",
          1174 => x"d2",
          1175 => x"83",
          1176 => x"83",
          1177 => x"b8",
          1178 => x"05",
          1179 => x"08",
          1180 => x"79",
          1181 => x"88",
          1182 => x"53",
          1183 => x"84",
          1184 => x"80",
          1185 => x"38",
          1186 => x"70",
          1187 => x"5f",
          1188 => x"a0",
          1189 => x"98",
          1190 => x"54",
          1191 => x"a8",
          1192 => x"3f",
          1193 => x"59",
          1194 => x"f0",
          1195 => x"a6",
          1196 => x"f2",
          1197 => x"64",
          1198 => x"11",
          1199 => x"3f",
          1200 => x"bb",
          1201 => x"22",
          1202 => x"45",
          1203 => x"80",
          1204 => x"c8",
          1205 => x"5e",
          1206 => x"82",
          1207 => x"fe",
          1208 => x"e1",
          1209 => x"b9",
          1210 => x"fc",
          1211 => x"aa",
          1212 => x"81",
          1213 => x"05",
          1214 => x"fb",
          1215 => x"53",
          1216 => x"84",
          1217 => x"38",
          1218 => x"05",
          1219 => x"83",
          1220 => x"7b",
          1221 => x"83",
          1222 => x"3f",
          1223 => x"da",
          1224 => x"bc",
          1225 => x"b8",
          1226 => x"05",
          1227 => x"08",
          1228 => x"80",
          1229 => x"5b",
          1230 => x"f2",
          1231 => x"cf",
          1232 => x"ea",
          1233 => x"80",
          1234 => x"49",
          1235 => x"d3",
          1236 => x"83",
          1237 => x"59",
          1238 => x"59",
          1239 => x"94",
          1240 => x"e8",
          1241 => x"83",
          1242 => x"9b",
          1243 => x"92",
          1244 => x"80",
          1245 => x"49",
          1246 => x"5e",
          1247 => x"a0",
          1248 => x"ca",
          1249 => x"83",
          1250 => x"83",
          1251 => x"94",
          1252 => x"ca",
          1253 => x"05",
          1254 => x"08",
          1255 => x"3d",
          1256 => x"87",
          1257 => x"87",
          1258 => x"3f",
          1259 => x"08",
          1260 => x"51",
          1261 => x"08",
          1262 => x"70",
          1263 => x"74",
          1264 => x"08",
          1265 => x"84",
          1266 => x"74",
          1267 => x"8c",
          1268 => x"0c",
          1269 => x"94",
          1270 => x"f1",
          1271 => x"34",
          1272 => x"3d",
          1273 => x"84",
          1274 => x"89",
          1275 => x"51",
          1276 => x"83",
          1277 => x"f2",
          1278 => x"3f",
          1279 => x"53",
          1280 => x"51",
          1281 => x"d2",
          1282 => x"83",
          1283 => x"80",
          1284 => x"e4",
          1285 => x"3d",
          1286 => x"75",
          1287 => x"38",
          1288 => x"52",
          1289 => x"38",
          1290 => x"06",
          1291 => x"38",
          1292 => x"2e",
          1293 => x"2e",
          1294 => x"81",
          1295 => x"2e",
          1296 => x"8b",
          1297 => x"12",
          1298 => x"06",
          1299 => x"06",
          1300 => x"70",
          1301 => x"52",
          1302 => x"72",
          1303 => x"0c",
          1304 => x"87",
          1305 => x"38",
          1306 => x"12",
          1307 => x"06",
          1308 => x"38",
          1309 => x"81",
          1310 => x"81",
          1311 => x"3d",
          1312 => x"80",
          1313 => x"0d",
          1314 => x"51",
          1315 => x"80",
          1316 => x"0c",
          1317 => x"76",
          1318 => x"81",
          1319 => x"83",
          1320 => x"73",
          1321 => x"33",
          1322 => x"fe",
          1323 => x"73",
          1324 => x"33",
          1325 => x"e6",
          1326 => x"74",
          1327 => x"13",
          1328 => x"26",
          1329 => x"98",
          1330 => x"bc",
          1331 => x"b8",
          1332 => x"b4",
          1333 => x"b0",
          1334 => x"ac",
          1335 => x"a8",
          1336 => x"73",
          1337 => x"87",
          1338 => x"84",
          1339 => x"f3",
          1340 => x"9c",
          1341 => x"bc",
          1342 => x"98",
          1343 => x"87",
          1344 => x"1c",
          1345 => x"7b",
          1346 => x"08",
          1347 => x"98",
          1348 => x"87",
          1349 => x"1c",
          1350 => x"79",
          1351 => x"83",
          1352 => x"ff",
          1353 => x"1b",
          1354 => x"1b",
          1355 => x"83",
          1356 => x"51",
          1357 => x"04",
          1358 => x"53",
          1359 => x"80",
          1360 => x"98",
          1361 => x"ff",
          1362 => x"83",
          1363 => x"0c",
          1364 => x"e7",
          1365 => x"2b",
          1366 => x"2e",
          1367 => x"80",
          1368 => x"98",
          1369 => x"ff",
          1370 => x"0d",
          1371 => x"54",
          1372 => x"b9",
          1373 => x"51",
          1374 => x"72",
          1375 => x"25",
          1376 => x"85",
          1377 => x"9b",
          1378 => x"81",
          1379 => x"2e",
          1380 => x"08",
          1381 => x"54",
          1382 => x"91",
          1383 => x"e3",
          1384 => x"72",
          1385 => x"81",
          1386 => x"ff",
          1387 => x"70",
          1388 => x"90",
          1389 => x"c8",
          1390 => x"2a",
          1391 => x"38",
          1392 => x"80",
          1393 => x"06",
          1394 => x"c0",
          1395 => x"81",
          1396 => x"d8",
          1397 => x"33",
          1398 => x"52",
          1399 => x"0d",
          1400 => x"75",
          1401 => x"2e",
          1402 => x"80",
          1403 => x"55",
          1404 => x"c0",
          1405 => x"81",
          1406 => x"8c",
          1407 => x"51",
          1408 => x"81",
          1409 => x"71",
          1410 => x"38",
          1411 => x"94",
          1412 => x"87",
          1413 => x"81",
          1414 => x"9b",
          1415 => x"3d",
          1416 => x"06",
          1417 => x"32",
          1418 => x"38",
          1419 => x"80",
          1420 => x"84",
          1421 => x"53",
          1422 => x"ff",
          1423 => x"70",
          1424 => x"80",
          1425 => x"a4",
          1426 => x"9e",
          1427 => x"c0",
          1428 => x"87",
          1429 => x"0c",
          1430 => x"94",
          1431 => x"f2",
          1432 => x"83",
          1433 => x"08",
          1434 => x"b4",
          1435 => x"9e",
          1436 => x"c0",
          1437 => x"87",
          1438 => x"0c",
          1439 => x"b4",
          1440 => x"71",
          1441 => x"84",
          1442 => x"9e",
          1443 => x"c0",
          1444 => x"81",
          1445 => x"87",
          1446 => x"0a",
          1447 => x"38",
          1448 => x"87",
          1449 => x"0a",
          1450 => x"83",
          1451 => x"34",
          1452 => x"70",
          1453 => x"70",
          1454 => x"83",
          1455 => x"9e",
          1456 => x"51",
          1457 => x"81",
          1458 => x"0b",
          1459 => x"80",
          1460 => x"2e",
          1461 => x"cd",
          1462 => x"08",
          1463 => x"52",
          1464 => x"71",
          1465 => x"c0",
          1466 => x"06",
          1467 => x"38",
          1468 => x"80",
          1469 => x"82",
          1470 => x"80",
          1471 => x"f2",
          1472 => x"90",
          1473 => x"52",
          1474 => x"52",
          1475 => x"87",
          1476 => x"80",
          1477 => x"83",
          1478 => x"34",
          1479 => x"70",
          1480 => x"80",
          1481 => x"f2",
          1482 => x"98",
          1483 => x"71",
          1484 => x"c0",
          1485 => x"51",
          1486 => x"81",
          1487 => x"c0",
          1488 => x"84",
          1489 => x"34",
          1490 => x"70",
          1491 => x"2e",
          1492 => x"d7",
          1493 => x"06",
          1494 => x"3d",
          1495 => x"fb",
          1496 => x"b6",
          1497 => x"73",
          1498 => x"c3",
          1499 => x"74",
          1500 => x"54",
          1501 => x"33",
          1502 => x"cd",
          1503 => x"f2",
          1504 => x"83",
          1505 => x"38",
          1506 => x"85",
          1507 => x"83",
          1508 => x"75",
          1509 => x"54",
          1510 => x"33",
          1511 => x"d1",
          1512 => x"f2",
          1513 => x"83",
          1514 => x"f2",
          1515 => x"ff",
          1516 => x"52",
          1517 => x"3f",
          1518 => x"8c",
          1519 => x"b4",
          1520 => x"22",
          1521 => x"fc",
          1522 => x"84",
          1523 => x"84",
          1524 => x"76",
          1525 => x"08",
          1526 => x"d4",
          1527 => x"b9",
          1528 => x"85",
          1529 => x"c4",
          1530 => x"51",
          1531 => x"bd",
          1532 => x"54",
          1533 => x"90",
          1534 => x"0d",
          1535 => x"84",
          1536 => x"84",
          1537 => x"76",
          1538 => x"08",
          1539 => x"ec",
          1540 => x"80",
          1541 => x"83",
          1542 => x"d9",
          1543 => x"ac",
          1544 => x"b3",
          1545 => x"83",
          1546 => x"83",
          1547 => x"51",
          1548 => x"51",
          1549 => x"52",
          1550 => x"3f",
          1551 => x"c0",
          1552 => x"b9",
          1553 => x"71",
          1554 => x"52",
          1555 => x"3f",
          1556 => x"2e",
          1557 => x"db",
          1558 => x"f2",
          1559 => x"8f",
          1560 => x"51",
          1561 => x"33",
          1562 => x"d6",
          1563 => x"97",
          1564 => x"80",
          1565 => x"dc",
          1566 => x"f2",
          1567 => x"b4",
          1568 => x"52",
          1569 => x"3f",
          1570 => x"2e",
          1571 => x"d8",
          1572 => x"b1",
          1573 => x"74",
          1574 => x"83",
          1575 => x"51",
          1576 => x"33",
          1577 => x"cd",
          1578 => x"98",
          1579 => x"51",
          1580 => x"33",
          1581 => x"c7",
          1582 => x"90",
          1583 => x"51",
          1584 => x"33",
          1585 => x"c1",
          1586 => x"88",
          1587 => x"51",
          1588 => x"33",
          1589 => x"c1",
          1590 => x"a0",
          1591 => x"51",
          1592 => x"33",
          1593 => x"c1",
          1594 => x"a8",
          1595 => x"51",
          1596 => x"33",
          1597 => x"c1",
          1598 => x"94",
          1599 => x"f7",
          1600 => x"80",
          1601 => x"3d",
          1602 => x"85",
          1603 => x"c2",
          1604 => x"de",
          1605 => x"3d",
          1606 => x"af",
          1607 => x"de",
          1608 => x"3d",
          1609 => x"af",
          1610 => x"de",
          1611 => x"3d",
          1612 => x"af",
          1613 => x"88",
          1614 => x"96",
          1615 => x"87",
          1616 => x"0d",
          1617 => x"5a",
          1618 => x"f3",
          1619 => x"84",
          1620 => x"3d",
          1621 => x"54",
          1622 => x"d2",
          1623 => x"2e",
          1624 => x"84",
          1625 => x"80",
          1626 => x"38",
          1627 => x"18",
          1628 => x"70",
          1629 => x"55",
          1630 => x"ff",
          1631 => x"11",
          1632 => x"84",
          1633 => x"2e",
          1634 => x"a9",
          1635 => x"ff",
          1636 => x"81",
          1637 => x"c0",
          1638 => x"3f",
          1639 => x"08",
          1640 => x"51",
          1641 => x"b9",
          1642 => x"3d",
          1643 => x"71",
          1644 => x"57",
          1645 => x"0b",
          1646 => x"10",
          1647 => x"54",
          1648 => x"08",
          1649 => x"89",
          1650 => x"84",
          1651 => x"88",
          1652 => x"16",
          1653 => x"76",
          1654 => x"b9",
          1655 => x"1a",
          1656 => x"ff",
          1657 => x"b9",
          1658 => x"1b",
          1659 => x"3f",
          1660 => x"54",
          1661 => x"70",
          1662 => x"27",
          1663 => x"33",
          1664 => x"e6",
          1665 => x"55",
          1666 => x"fe",
          1667 => x"80",
          1668 => x"39",
          1669 => x"f3",
          1670 => x"3f",
          1671 => x"83",
          1672 => x"77",
          1673 => x"c8",
          1674 => x"ff",
          1675 => x"55",
          1676 => x"9d",
          1677 => x"70",
          1678 => x"53",
          1679 => x"52",
          1680 => x"2e",
          1681 => x"0b",
          1682 => x"04",
          1683 => x"3d",
          1684 => x"80",
          1685 => x"33",
          1686 => x"9e",
          1687 => x"56",
          1688 => x"80",
          1689 => x"06",
          1690 => x"80",
          1691 => x"3d",
          1692 => x"84",
          1693 => x"2c",
          1694 => x"79",
          1695 => x"70",
          1696 => x"80",
          1697 => x"71",
          1698 => x"de",
          1699 => x"52",
          1700 => x"5c",
          1701 => x"cd",
          1702 => x"75",
          1703 => x"05",
          1704 => x"24",
          1705 => x"82",
          1706 => x"d4",
          1707 => x"91",
          1708 => x"70",
          1709 => x"95",
          1710 => x"84",
          1711 => x"2e",
          1712 => x"2b",
          1713 => x"70",
          1714 => x"2c",
          1715 => x"11",
          1716 => x"57",
          1717 => x"76",
          1718 => x"81",
          1719 => x"80",
          1720 => x"98",
          1721 => x"41",
          1722 => x"10",
          1723 => x"0b",
          1724 => x"77",
          1725 => x"15",
          1726 => x"61",
          1727 => x"ff",
          1728 => x"76",
          1729 => x"39",
          1730 => x"76",
          1731 => x"34",
          1732 => x"34",
          1733 => x"26",
          1734 => x"c3",
          1735 => x"de",
          1736 => x"84",
          1737 => x"80",
          1738 => x"56",
          1739 => x"d5",
          1740 => x"8a",
          1741 => x"57",
          1742 => x"39",
          1743 => x"06",
          1744 => x"75",
          1745 => x"ac",
          1746 => x"d1",
          1747 => x"55",
          1748 => x"7c",
          1749 => x"10",
          1750 => x"59",
          1751 => x"88",
          1752 => x"33",
          1753 => x"80",
          1754 => x"52",
          1755 => x"d5",
          1756 => x"8a",
          1757 => x"51",
          1758 => x"33",
          1759 => x"34",
          1760 => x"38",
          1761 => x"84",
          1762 => x"8a",
          1763 => x"8d",
          1764 => x"e0",
          1765 => x"8e",
          1766 => x"2e",
          1767 => x"ec",
          1768 => x"88",
          1769 => x"06",
          1770 => x"ff",
          1771 => x"84",
          1772 => x"2e",
          1773 => x"52",
          1774 => x"d5",
          1775 => x"f2",
          1776 => x"51",
          1777 => x"33",
          1778 => x"34",
          1779 => x"84",
          1780 => x"84",
          1781 => x"79",
          1782 => x"08",
          1783 => x"8c",
          1784 => x"ff",
          1785 => x"70",
          1786 => x"5a",
          1787 => x"38",
          1788 => x"57",
          1789 => x"70",
          1790 => x"84",
          1791 => x"84",
          1792 => x"76",
          1793 => x"84",
          1794 => x"56",
          1795 => x"ff",
          1796 => x"75",
          1797 => x"ff",
          1798 => x"80",
          1799 => x"a0",
          1800 => x"8c",
          1801 => x"84",
          1802 => x"74",
          1803 => x"ac",
          1804 => x"3f",
          1805 => x"0a",
          1806 => x"33",
          1807 => x"e2",
          1808 => x"51",
          1809 => x"0a",
          1810 => x"2c",
          1811 => x"7a",
          1812 => x"39",
          1813 => x"34",
          1814 => x"51",
          1815 => x"0a",
          1816 => x"2c",
          1817 => x"75",
          1818 => x"58",
          1819 => x"ac",
          1820 => x"8a",
          1821 => x"80",
          1822 => x"88",
          1823 => x"ff",
          1824 => x"8c",
          1825 => x"38",
          1826 => x"ff",
          1827 => x"ff",
          1828 => x"76",
          1829 => x"d1",
          1830 => x"34",
          1831 => x"ff",
          1832 => x"7b",
          1833 => x"08",
          1834 => x"38",
          1835 => x"2e",
          1836 => x"70",
          1837 => x"08",
          1838 => x"75",
          1839 => x"e0",
          1840 => x"80",
          1841 => x"7b",
          1842 => x"10",
          1843 => x"41",
          1844 => x"b4",
          1845 => x"83",
          1846 => x"8b",
          1847 => x"34",
          1848 => x"84",
          1849 => x"84",
          1850 => x"b6",
          1851 => x"51",
          1852 => x"08",
          1853 => x"84",
          1854 => x"ae",
          1855 => x"05",
          1856 => x"81",
          1857 => x"d1",
          1858 => x"0b",
          1859 => x"d1",
          1860 => x"34",
          1861 => x"8c",
          1862 => x"84",
          1863 => x"ae",
          1864 => x"a0",
          1865 => x"ac",
          1866 => x"3f",
          1867 => x"7c",
          1868 => x"06",
          1869 => x"51",
          1870 => x"d1",
          1871 => x"34",
          1872 => x"0d",
          1873 => x"ff",
          1874 => x"ca",
          1875 => x"59",
          1876 => x"58",
          1877 => x"ac",
          1878 => x"3f",
          1879 => x"70",
          1880 => x"52",
          1881 => x"38",
          1882 => x"ff",
          1883 => x"70",
          1884 => x"88",
          1885 => x"24",
          1886 => x"52",
          1887 => x"81",
          1888 => x"70",
          1889 => x"51",
          1890 => x"84",
          1891 => x"ac",
          1892 => x"81",
          1893 => x"d1",
          1894 => x"25",
          1895 => x"16",
          1896 => x"d5",
          1897 => x"ac",
          1898 => x"81",
          1899 => x"d1",
          1900 => x"25",
          1901 => x"17",
          1902 => x"52",
          1903 => x"75",
          1904 => x"05",
          1905 => x"43",
          1906 => x"38",
          1907 => x"70",
          1908 => x"2e",
          1909 => x"55",
          1910 => x"2b",
          1911 => x"24",
          1912 => x"81",
          1913 => x"81",
          1914 => x"d1",
          1915 => x"25",
          1916 => x"d1",
          1917 => x"05",
          1918 => x"d1",
          1919 => x"38",
          1920 => x"34",
          1921 => x"81",
          1922 => x"70",
          1923 => x"58",
          1924 => x"38",
          1925 => x"81",
          1926 => x"25",
          1927 => x"52",
          1928 => x"81",
          1929 => x"70",
          1930 => x"57",
          1931 => x"84",
          1932 => x"aa",
          1933 => x"81",
          1934 => x"d1",
          1935 => x"24",
          1936 => x"f2",
          1937 => x"9d",
          1938 => x"84",
          1939 => x"84",
          1940 => x"05",
          1941 => x"be",
          1942 => x"8c",
          1943 => x"c8",
          1944 => x"51",
          1945 => x"08",
          1946 => x"84",
          1947 => x"a9",
          1948 => x"05",
          1949 => x"81",
          1950 => x"80",
          1951 => x"83",
          1952 => x"85",
          1953 => x"77",
          1954 => x"d5",
          1955 => x"52",
          1956 => x"80",
          1957 => x"98",
          1958 => x"57",
          1959 => x"8c",
          1960 => x"79",
          1961 => x"75",
          1962 => x"39",
          1963 => x"fc",
          1964 => x"76",
          1965 => x"84",
          1966 => x"38",
          1967 => x"f3",
          1968 => x"d4",
          1969 => x"83",
          1970 => x"3f",
          1971 => x"3d",
          1972 => x"74",
          1973 => x"0c",
          1974 => x"80",
          1975 => x"75",
          1976 => x"c8",
          1977 => x"c8",
          1978 => x"75",
          1979 => x"93",
          1980 => x"8c",
          1981 => x"f2",
          1982 => x"88",
          1983 => x"ac",
          1984 => x"3f",
          1985 => x"ff",
          1986 => x"ff",
          1987 => x"79",
          1988 => x"7c",
          1989 => x"80",
          1990 => x"b9",
          1991 => x"51",
          1992 => x"08",
          1993 => x"08",
          1994 => x"52",
          1995 => x"1d",
          1996 => x"33",
          1997 => x"56",
          1998 => x"d5",
          1999 => x"f2",
          2000 => x"51",
          2001 => x"08",
          2002 => x"84",
          2003 => x"84",
          2004 => x"55",
          2005 => x"3f",
          2006 => x"34",
          2007 => x"81",
          2008 => x"a9",
          2009 => x"06",
          2010 => x"33",
          2011 => x"f0",
          2012 => x"88",
          2013 => x"ac",
          2014 => x"3f",
          2015 => x"ff",
          2016 => x"ff",
          2017 => x"60",
          2018 => x"51",
          2019 => x"33",
          2020 => x"f2",
          2021 => x"5c",
          2022 => x"c8",
          2023 => x"70",
          2024 => x"08",
          2025 => x"d5",
          2026 => x"ff",
          2027 => x"81",
          2028 => x"93",
          2029 => x"f3",
          2030 => x"fe",
          2031 => x"75",
          2032 => x"b4",
          2033 => x"3f",
          2034 => x"f3",
          2035 => x"80",
          2036 => x"b9",
          2037 => x"53",
          2038 => x"81",
          2039 => x"82",
          2040 => x"3d",
          2041 => x"80",
          2042 => x"3f",
          2043 => x"c8",
          2044 => x"ee",
          2045 => x"a6",
          2046 => x"80",
          2047 => x"e3",
          2048 => x"70",
          2049 => x"81",
          2050 => x"10",
          2051 => x"58",
          2052 => x"76",
          2053 => x"e0",
          2054 => x"80",
          2055 => x"75",
          2056 => x"10",
          2057 => x"40",
          2058 => x"81",
          2059 => x"83",
          2060 => x"81",
          2061 => x"38",
          2062 => x"74",
          2063 => x"b8",
          2064 => x"5b",
          2065 => x"80",
          2066 => x"39",
          2067 => x"f3",
          2068 => x"06",
          2069 => x"54",
          2070 => x"84",
          2071 => x"b8",
          2072 => x"05",
          2073 => x"2e",
          2074 => x"83",
          2075 => x"83",
          2076 => x"e1",
          2077 => x"e7",
          2078 => x"0d",
          2079 => x"05",
          2080 => x"83",
          2081 => x"81",
          2082 => x"38",
          2083 => x"a7",
          2084 => x"70",
          2085 => x"79",
          2086 => x"f8",
          2087 => x"83",
          2088 => x"70",
          2089 => x"88",
          2090 => x"56",
          2091 => x"80",
          2092 => x"73",
          2093 => x"26",
          2094 => x"83",
          2095 => x"79",
          2096 => x"e0",
          2097 => x"05",
          2098 => x"38",
          2099 => x"80",
          2100 => x"10",
          2101 => x"29",
          2102 => x"59",
          2103 => x"bc",
          2104 => x"bb",
          2105 => x"f6",
          2106 => x"75",
          2107 => x"5b",
          2108 => x"74",
          2109 => x"06",
          2110 => x"06",
          2111 => x"ff",
          2112 => x"57",
          2113 => x"38",
          2114 => x"05",
          2115 => x"83",
          2116 => x"38",
          2117 => x"fe",
          2118 => x"55",
          2119 => x"81",
          2120 => x"a0",
          2121 => x"84",
          2122 => x"84",
          2123 => x"83",
          2124 => x"5b",
          2125 => x"78",
          2126 => x"06",
          2127 => x"18",
          2128 => x"bb",
          2129 => x"80",
          2130 => x"f4",
          2131 => x"07",
          2132 => x"7f",
          2133 => x"fd",
          2134 => x"e6",
          2135 => x"ff",
          2136 => x"f9",
          2137 => x"a0",
          2138 => x"5f",
          2139 => x"b7",
          2140 => x"b7",
          2141 => x"f8",
          2142 => x"7c",
          2143 => x"5f",
          2144 => x"26",
          2145 => x"7d",
          2146 => x"06",
          2147 => x"7d",
          2148 => x"06",
          2149 => x"5d",
          2150 => x"75",
          2151 => x"83",
          2152 => x"76",
          2153 => x"fb",
          2154 => x"56",
          2155 => x"ee",
          2156 => x"87",
          2157 => x"34",
          2158 => x"75",
          2159 => x"80",
          2160 => x"34",
          2161 => x"34",
          2162 => x"81",
          2163 => x"a0",
          2164 => x"f8",
          2165 => x"06",
          2166 => x"73",
          2167 => x"07",
          2168 => x"87",
          2169 => x"51",
          2170 => x"73",
          2171 => x"72",
          2172 => x"bc",
          2173 => x"87",
          2174 => x"84",
          2175 => x"02",
          2176 => x"05",
          2177 => x"56",
          2178 => x"38",
          2179 => x"33",
          2180 => x"12",
          2181 => x"f6",
          2182 => x"29",
          2183 => x"f7",
          2184 => x"81",
          2185 => x"22",
          2186 => x"23",
          2187 => x"81",
          2188 => x"5b",
          2189 => x"ff",
          2190 => x"83",
          2191 => x"06",
          2192 => x"79",
          2193 => x"bc",
          2194 => x"54",
          2195 => x"98",
          2196 => x"13",
          2197 => x"81",
          2198 => x"57",
          2199 => x"73",
          2200 => x"a1",
          2201 => x"9a",
          2202 => x"14",
          2203 => x"34",
          2204 => x"eb",
          2205 => x"56",
          2206 => x"78",
          2207 => x"06",
          2208 => x"38",
          2209 => x"bc",
          2210 => x"75",
          2211 => x"a7",
          2212 => x"81",
          2213 => x"5c",
          2214 => x"84",
          2215 => x"33",
          2216 => x"70",
          2217 => x"05",
          2218 => x"34",
          2219 => x"b7",
          2220 => x"5c",
          2221 => x"80",
          2222 => x"3d",
          2223 => x"83",
          2224 => x"06",
          2225 => x"73",
          2226 => x"2e",
          2227 => x"ff",
          2228 => x"72",
          2229 => x"38",
          2230 => x"bc",
          2231 => x"11",
          2232 => x"fe",
          2233 => x"98",
          2234 => x"56",
          2235 => x"75",
          2236 => x"53",
          2237 => x"0b",
          2238 => x"81",
          2239 => x"d8",
          2240 => x"b7",
          2241 => x"83",
          2242 => x"c4",
          2243 => x"33",
          2244 => x"76",
          2245 => x"51",
          2246 => x"10",
          2247 => x"04",
          2248 => x"27",
          2249 => x"80",
          2250 => x"0d",
          2251 => x"83",
          2252 => x"54",
          2253 => x"12",
          2254 => x"0b",
          2255 => x"04",
          2256 => x"70",
          2257 => x"55",
          2258 => x"de",
          2259 => x"84",
          2260 => x"51",
          2261 => x"72",
          2262 => x"b9",
          2263 => x"f8",
          2264 => x"70",
          2265 => x"55",
          2266 => x"84",
          2267 => x"83",
          2268 => x"bc",
          2269 => x"74",
          2270 => x"f8",
          2271 => x"0c",
          2272 => x"f8",
          2273 => x"b7",
          2274 => x"75",
          2275 => x"70",
          2276 => x"ff",
          2277 => x"70",
          2278 => x"83",
          2279 => x"83",
          2280 => x"71",
          2281 => x"84",
          2282 => x"80",
          2283 => x"80",
          2284 => x"0b",
          2285 => x"04",
          2286 => x"90",
          2287 => x"80",
          2288 => x"0d",
          2289 => x"07",
          2290 => x"39",
          2291 => x"86",
          2292 => x"d7",
          2293 => x"34",
          2294 => x"3d",
          2295 => x"fc",
          2296 => x"f4",
          2297 => x"33",
          2298 => x"34",
          2299 => x"81",
          2300 => x"f8",
          2301 => x"f4",
          2302 => x"70",
          2303 => x"83",
          2304 => x"07",
          2305 => x"ef",
          2306 => x"06",
          2307 => x"df",
          2308 => x"06",
          2309 => x"f4",
          2310 => x"33",
          2311 => x"83",
          2312 => x"f8",
          2313 => x"07",
          2314 => x"a7",
          2315 => x"06",
          2316 => x"f4",
          2317 => x"33",
          2318 => x"83",
          2319 => x"f8",
          2320 => x"83",
          2321 => x"f8",
          2322 => x"51",
          2323 => x"39",
          2324 => x"02",
          2325 => x"f8",
          2326 => x"f8",
          2327 => x"41",
          2328 => x"82",
          2329 => x"78",
          2330 => x"b7",
          2331 => x"34",
          2332 => x"f8",
          2333 => x"8f",
          2334 => x"81",
          2335 => x"be",
          2336 => x"82",
          2337 => x"83",
          2338 => x"f6",
          2339 => x"57",
          2340 => x"ba",
          2341 => x"52",
          2342 => x"3f",
          2343 => x"84",
          2344 => x"34",
          2345 => x"f8",
          2346 => x"0b",
          2347 => x"b7",
          2348 => x"34",
          2349 => x"0b",
          2350 => x"33",
          2351 => x"b8",
          2352 => x"7c",
          2353 => x"ff",
          2354 => x"c9",
          2355 => x"38",
          2356 => x"22",
          2357 => x"80",
          2358 => x"06",
          2359 => x"78",
          2360 => x"51",
          2361 => x"be",
          2362 => x"7a",
          2363 => x"f6",
          2364 => x"3d",
          2365 => x"34",
          2366 => x"0b",
          2367 => x"f8",
          2368 => x"23",
          2369 => x"3f",
          2370 => x"f4",
          2371 => x"83",
          2372 => x"78",
          2373 => x"38",
          2374 => x"e3",
          2375 => x"19",
          2376 => x"39",
          2377 => x"a7",
          2378 => x"f8",
          2379 => x"71",
          2380 => x"83",
          2381 => x"71",
          2382 => x"06",
          2383 => x"55",
          2384 => x"38",
          2385 => x"89",
          2386 => x"83",
          2387 => x"38",
          2388 => x"33",
          2389 => x"05",
          2390 => x"33",
          2391 => x"b7",
          2392 => x"f8",
          2393 => x"5a",
          2394 => x"34",
          2395 => x"16",
          2396 => x"a7",
          2397 => x"33",
          2398 => x"22",
          2399 => x"11",
          2400 => x"f4",
          2401 => x"18",
          2402 => x"78",
          2403 => x"33",
          2404 => x"53",
          2405 => x"bf",
          2406 => x"84",
          2407 => x"80",
          2408 => x"0c",
          2409 => x"97",
          2410 => x"75",
          2411 => x"38",
          2412 => x"80",
          2413 => x"39",
          2414 => x"b7",
          2415 => x"2e",
          2416 => x"53",
          2417 => x"81",
          2418 => x"72",
          2419 => x"a0",
          2420 => x"81",
          2421 => x"d8",
          2422 => x"f9",
          2423 => x"51",
          2424 => x"c8",
          2425 => x"ff",
          2426 => x"83",
          2427 => x"55",
          2428 => x"53",
          2429 => x"a0",
          2430 => x"33",
          2431 => x"53",
          2432 => x"83",
          2433 => x"0b",
          2434 => x"51",
          2435 => x"52",
          2436 => x"39",
          2437 => x"33",
          2438 => x"81",
          2439 => x"83",
          2440 => x"38",
          2441 => x"88",
          2442 => x"88",
          2443 => x"f8",
          2444 => x"72",
          2445 => x"c4",
          2446 => x"34",
          2447 => x"33",
          2448 => x"12",
          2449 => x"fa",
          2450 => x"71",
          2451 => x"f4",
          2452 => x"34",
          2453 => x"06",
          2454 => x"33",
          2455 => x"58",
          2456 => x"9a",
          2457 => x"06",
          2458 => x"38",
          2459 => x"f1",
          2460 => x"f9",
          2461 => x"9c",
          2462 => x"8a",
          2463 => x"78",
          2464 => x"db",
          2465 => x"b8",
          2466 => x"f8",
          2467 => x"72",
          2468 => x"c4",
          2469 => x"34",
          2470 => x"33",
          2471 => x"12",
          2472 => x"fa",
          2473 => x"71",
          2474 => x"33",
          2475 => x"b7",
          2476 => x"f8",
          2477 => x"72",
          2478 => x"83",
          2479 => x"05",
          2480 => x"06",
          2481 => x"77",
          2482 => x"b9",
          2483 => x"9b",
          2484 => x"83",
          2485 => x"06",
          2486 => x"f9",
          2487 => x"9c",
          2488 => x"aa",
          2489 => x"84",
          2490 => x"11",
          2491 => x"78",
          2492 => x"ff",
          2493 => x"1a",
          2494 => x"9c",
          2495 => x"e9",
          2496 => x"84",
          2497 => x"83",
          2498 => x"5e",
          2499 => x"86",
          2500 => x"bc",
          2501 => x"f6",
          2502 => x"59",
          2503 => x"83",
          2504 => x"5b",
          2505 => x"b0",
          2506 => x"70",
          2507 => x"83",
          2508 => x"44",
          2509 => x"33",
          2510 => x"1f",
          2511 => x"51",
          2512 => x"f9",
          2513 => x"33",
          2514 => x"06",
          2515 => x"12",
          2516 => x"f6",
          2517 => x"05",
          2518 => x"ce",
          2519 => x"81",
          2520 => x"06",
          2521 => x"38",
          2522 => x"fc",
          2523 => x"34",
          2524 => x"0b",
          2525 => x"b8",
          2526 => x"0c",
          2527 => x"3d",
          2528 => x"b9",
          2529 => x"b9",
          2530 => x"b9",
          2531 => x"0c",
          2532 => x"3d",
          2533 => x"81",
          2534 => x"33",
          2535 => x"06",
          2536 => x"06",
          2537 => x"80",
          2538 => x"72",
          2539 => x"06",
          2540 => x"5c",
          2541 => x"fe",
          2542 => x"58",
          2543 => x"83",
          2544 => x"7a",
          2545 => x"72",
          2546 => x"b7",
          2547 => x"34",
          2548 => x"33",
          2549 => x"12",
          2550 => x"f8",
          2551 => x"60",
          2552 => x"f8",
          2553 => x"34",
          2554 => x"06",
          2555 => x"33",
          2556 => x"5e",
          2557 => x"98",
          2558 => x"ff",
          2559 => x"ea",
          2560 => x"96",
          2561 => x"f8",
          2562 => x"81",
          2563 => x"ac",
          2564 => x"78",
          2565 => x"2e",
          2566 => x"5f",
          2567 => x"56",
          2568 => x"10",
          2569 => x"08",
          2570 => x"80",
          2571 => x"0b",
          2572 => x"04",
          2573 => x"33",
          2574 => x"33",
          2575 => x"11",
          2576 => x"f6",
          2577 => x"70",
          2578 => x"33",
          2579 => x"7f",
          2580 => x"7a",
          2581 => x"7a",
          2582 => x"5c",
          2583 => x"a7",
          2584 => x"33",
          2585 => x"22",
          2586 => x"56",
          2587 => x"83",
          2588 => x"5a",
          2589 => x"b0",
          2590 => x"70",
          2591 => x"83",
          2592 => x"5b",
          2593 => x"33",
          2594 => x"05",
          2595 => x"7a",
          2596 => x"33",
          2597 => x"56",
          2598 => x"70",
          2599 => x"26",
          2600 => x"84",
          2601 => x"72",
          2602 => x"72",
          2603 => x"54",
          2604 => x"e4",
          2605 => x"84",
          2606 => x"83",
          2607 => x"5e",
          2608 => x"fa",
          2609 => x"71",
          2610 => x"33",
          2611 => x"b7",
          2612 => x"f8",
          2613 => x"72",
          2614 => x"83",
          2615 => x"34",
          2616 => x"5b",
          2617 => x"77",
          2618 => x"82",
          2619 => x"84",
          2620 => x"83",
          2621 => x"c4",
          2622 => x"33",
          2623 => x"56",
          2624 => x"ca",
          2625 => x"9c",
          2626 => x"33",
          2627 => x"34",
          2628 => x"33",
          2629 => x"80",
          2630 => x"42",
          2631 => x"51",
          2632 => x"08",
          2633 => x"c9",
          2634 => x"b8",
          2635 => x"41",
          2636 => x"b9",
          2637 => x"f8",
          2638 => x"1c",
          2639 => x"84",
          2640 => x"5b",
          2641 => x"bc",
          2642 => x"f9",
          2643 => x"5b",
          2644 => x"a7",
          2645 => x"33",
          2646 => x"22",
          2647 => x"56",
          2648 => x"f8",
          2649 => x"5e",
          2650 => x"b0",
          2651 => x"70",
          2652 => x"83",
          2653 => x"41",
          2654 => x"33",
          2655 => x"70",
          2656 => x"26",
          2657 => x"58",
          2658 => x"75",
          2659 => x"b8",
          2660 => x"7f",
          2661 => x"c0",
          2662 => x"52",
          2663 => x"84",
          2664 => x"84",
          2665 => x"84",
          2666 => x"84",
          2667 => x"f6",
          2668 => x"33",
          2669 => x"33",
          2670 => x"33",
          2671 => x"84",
          2672 => x"ff",
          2673 => x"7c",
          2674 => x"38",
          2675 => x"83",
          2676 => x"53",
          2677 => x"52",
          2678 => x"fe",
          2679 => x"81",
          2680 => x"76",
          2681 => x"38",
          2682 => x"fd",
          2683 => x"84",
          2684 => x"ff",
          2685 => x"38",
          2686 => x"11",
          2687 => x"a5",
          2688 => x"05",
          2689 => x"33",
          2690 => x"83",
          2691 => x"71",
          2692 => x"72",
          2693 => x"83",
          2694 => x"b8",
          2695 => x"e7",
          2696 => x"70",
          2697 => x"5d",
          2698 => x"38",
          2699 => x"39",
          2700 => x"f8",
          2701 => x"57",
          2702 => x"17",
          2703 => x"9c",
          2704 => x"83",
          2705 => x"ff",
          2706 => x"84",
          2707 => x"f8",
          2708 => x"33",
          2709 => x"83",
          2710 => x"71",
          2711 => x"72",
          2712 => x"83",
          2713 => x"b8",
          2714 => x"c4",
          2715 => x"99",
          2716 => x"84",
          2717 => x"83",
          2718 => x"86",
          2719 => x"22",
          2720 => x"05",
          2721 => x"cc",
          2722 => x"5a",
          2723 => x"92",
          2724 => x"34",
          2725 => x"5a",
          2726 => x"b9",
          2727 => x"81",
          2728 => x"f7",
          2729 => x"c9",
          2730 => x"38",
          2731 => x"33",
          2732 => x"ff",
          2733 => x"83",
          2734 => x"34",
          2735 => x"57",
          2736 => x"b9",
          2737 => x"61",
          2738 => x"59",
          2739 => x"75",
          2740 => x"f4",
          2741 => x"dc",
          2742 => x"57",
          2743 => x"76",
          2744 => x"53",
          2745 => x"bc",
          2746 => x"84",
          2747 => x"39",
          2748 => x"57",
          2749 => x"9c",
          2750 => x"75",
          2751 => x"51",
          2752 => x"b8",
          2753 => x"b7",
          2754 => x"70",
          2755 => x"ff",
          2756 => x"bb",
          2757 => x"40",
          2758 => x"7e",
          2759 => x"f8",
          2760 => x"18",
          2761 => x"77",
          2762 => x"b7",
          2763 => x"60",
          2764 => x"83",
          2765 => x"b8",
          2766 => x"ef",
          2767 => x"bb",
          2768 => x"94",
          2769 => x"bc",
          2770 => x"f9",
          2771 => x"a0",
          2772 => x"40",
          2773 => x"ff",
          2774 => x"59",
          2775 => x"f0",
          2776 => x"7c",
          2777 => x"fe",
          2778 => x"76",
          2779 => x"75",
          2780 => x"06",
          2781 => x"24",
          2782 => x"56",
          2783 => x"16",
          2784 => x"81",
          2785 => x"57",
          2786 => x"75",
          2787 => x"06",
          2788 => x"58",
          2789 => x"b0",
          2790 => x"ff",
          2791 => x"42",
          2792 => x"84",
          2793 => x"33",
          2794 => x"70",
          2795 => x"05",
          2796 => x"34",
          2797 => x"b7",
          2798 => x"40",
          2799 => x"38",
          2800 => x"c4",
          2801 => x"34",
          2802 => x"70",
          2803 => x"b7",
          2804 => x"71",
          2805 => x"78",
          2806 => x"84",
          2807 => x"87",
          2808 => x"33",
          2809 => x"80",
          2810 => x"84",
          2811 => x"79",
          2812 => x"22",
          2813 => x"8b",
          2814 => x"76",
          2815 => x"79",
          2816 => x"ed",
          2817 => x"60",
          2818 => x"06",
          2819 => x"7b",
          2820 => x"76",
          2821 => x"70",
          2822 => x"80",
          2823 => x"b0",
          2824 => x"5d",
          2825 => x"57",
          2826 => x"33",
          2827 => x"71",
          2828 => x"59",
          2829 => x"38",
          2830 => x"7d",
          2831 => x"77",
          2832 => x"84",
          2833 => x"ff",
          2834 => x"f6",
          2835 => x"59",
          2836 => x"76",
          2837 => x"05",
          2838 => x"76",
          2839 => x"f4",
          2840 => x"a0",
          2841 => x"70",
          2842 => x"76",
          2843 => x"e0",
          2844 => x"05",
          2845 => x"27",
          2846 => x"70",
          2847 => x"39",
          2848 => x"06",
          2849 => x"84",
          2850 => x"f0",
          2851 => x"f2",
          2852 => x"70",
          2853 => x"39",
          2854 => x"b7",
          2855 => x"f8",
          2856 => x"f6",
          2857 => x"5f",
          2858 => x"33",
          2859 => x"34",
          2860 => x"56",
          2861 => x"81",
          2862 => x"f8",
          2863 => x"33",
          2864 => x"83",
          2865 => x"f4",
          2866 => x"75",
          2867 => x"f8",
          2868 => x"56",
          2869 => x"39",
          2870 => x"81",
          2871 => x"f4",
          2872 => x"8f",
          2873 => x"ff",
          2874 => x"9f",
          2875 => x"f4",
          2876 => x"33",
          2877 => x"75",
          2878 => x"83",
          2879 => x"c0",
          2880 => x"fe",
          2881 => x"af",
          2882 => x"f4",
          2883 => x"33",
          2884 => x"83",
          2885 => x"f8",
          2886 => x"56",
          2887 => x"39",
          2888 => x"82",
          2889 => x"fe",
          2890 => x"f8",
          2891 => x"fd",
          2892 => x"f0",
          2893 => x"fd",
          2894 => x"f0",
          2895 => x"fd",
          2896 => x"df",
          2897 => x"f8",
          2898 => x"f4",
          2899 => x"75",
          2900 => x"80",
          2901 => x"81",
          2902 => x"84",
          2903 => x"84",
          2904 => x"84",
          2905 => x"f6",
          2906 => x"e8",
          2907 => x"34",
          2908 => x"3d",
          2909 => x"83",
          2910 => x"58",
          2911 => x"b8",
          2912 => x"d8",
          2913 => x"b9",
          2914 => x"08",
          2915 => x"b8",
          2916 => x"0c",
          2917 => x"f9",
          2918 => x"33",
          2919 => x"c9",
          2920 => x"02",
          2921 => x"1e",
          2922 => x"ca",
          2923 => x"80",
          2924 => x"f8",
          2925 => x"ff",
          2926 => x"83",
          2927 => x"d0",
          2928 => x"fe",
          2929 => x"f8",
          2930 => x"9f",
          2931 => x"a6",
          2932 => x"84",
          2933 => x"ee",
          2934 => x"ee",
          2935 => x"05",
          2936 => x"58",
          2937 => x"f8",
          2938 => x"ff",
          2939 => x"f3",
          2940 => x"84",
          2941 => x"58",
          2942 => x"83",
          2943 => x"70",
          2944 => x"71",
          2945 => x"05",
          2946 => x"7e",
          2947 => x"83",
          2948 => x"5f",
          2949 => x"79",
          2950 => x"57",
          2951 => x"b7",
          2952 => x"98",
          2953 => x"f6",
          2954 => x"57",
          2955 => x"84",
          2956 => x"82",
          2957 => x"f8",
          2958 => x"f8",
          2959 => x"76",
          2960 => x"05",
          2961 => x"5c",
          2962 => x"80",
          2963 => x"ff",
          2964 => x"29",
          2965 => x"27",
          2966 => x"57",
          2967 => x"c4",
          2968 => x"34",
          2969 => x"70",
          2970 => x"b7",
          2971 => x"71",
          2972 => x"76",
          2973 => x"33",
          2974 => x"70",
          2975 => x"05",
          2976 => x"34",
          2977 => x"b7",
          2978 => x"41",
          2979 => x"38",
          2980 => x"33",
          2981 => x"34",
          2982 => x"33",
          2983 => x"33",
          2984 => x"76",
          2985 => x"70",
          2986 => x"58",
          2987 => x"79",
          2988 => x"06",
          2989 => x"83",
          2990 => x"34",
          2991 => x"06",
          2992 => x"27",
          2993 => x"f8",
          2994 => x"f9",
          2995 => x"ff",
          2996 => x"ef",
          2997 => x"75",
          2998 => x"38",
          2999 => x"06",
          3000 => x"5d",
          3001 => x"f4",
          3002 => x"56",
          3003 => x"39",
          3004 => x"23",
          3005 => x"75",
          3006 => x"77",
          3007 => x"8d",
          3008 => x"34",
          3009 => x"05",
          3010 => x"38",
          3011 => x"83",
          3012 => x"59",
          3013 => x"d3",
          3014 => x"f8",
          3015 => x"83",
          3016 => x"83",
          3017 => x"0b",
          3018 => x"80",
          3019 => x"39",
          3020 => x"b7",
          3021 => x"83",
          3022 => x"3d",
          3023 => x"be",
          3024 => x"38",
          3025 => x"84",
          3026 => x"76",
          3027 => x"0b",
          3028 => x"04",
          3029 => x"5c",
          3030 => x"81",
          3031 => x"58",
          3032 => x"d6",
          3033 => x"cc",
          3034 => x"0c",
          3035 => x"08",
          3036 => x"38",
          3037 => x"70",
          3038 => x"58",
          3039 => x"80",
          3040 => x"83",
          3041 => x"30",
          3042 => x"5d",
          3043 => x"b7",
          3044 => x"f8",
          3045 => x"a7",
          3046 => x"5b",
          3047 => x"83",
          3048 => x"58",
          3049 => x"8c",
          3050 => x"80",
          3051 => x"88",
          3052 => x"75",
          3053 => x"84",
          3054 => x"34",
          3055 => x"55",
          3056 => x"54",
          3057 => x"ff",
          3058 => x"54",
          3059 => x"72",
          3060 => x"83",
          3061 => x"06",
          3062 => x"38",
          3063 => x"f6",
          3064 => x"34",
          3065 => x"5e",
          3066 => x"f6",
          3067 => x"25",
          3068 => x"34",
          3069 => x"81",
          3070 => x"72",
          3071 => x"83",
          3072 => x"53",
          3073 => x"0b",
          3074 => x"f7",
          3075 => x"f7",
          3076 => x"83",
          3077 => x"5c",
          3078 => x"55",
          3079 => x"f7",
          3080 => x"82",
          3081 => x"53",
          3082 => x"f7",
          3083 => x"38",
          3084 => x"ff",
          3085 => x"33",
          3086 => x"74",
          3087 => x"2e",
          3088 => x"33",
          3089 => x"83",
          3090 => x"c0",
          3091 => x"27",
          3092 => x"98",
          3093 => x"81",
          3094 => x"89",
          3095 => x"f7",
          3096 => x"fe",
          3097 => x"8b",
          3098 => x"05",
          3099 => x"08",
          3100 => x"f4",
          3101 => x"5e",
          3102 => x"0b",
          3103 => x"81",
          3104 => x"f7",
          3105 => x"83",
          3106 => x"58",
          3107 => x"fa",
          3108 => x"33",
          3109 => x"39",
          3110 => x"2e",
          3111 => x"f4",
          3112 => x"54",
          3113 => x"39",
          3114 => x"81",
          3115 => x"81",
          3116 => x"80",
          3117 => x"38",
          3118 => x"27",
          3119 => x"25",
          3120 => x"81",
          3121 => x"81",
          3122 => x"2b",
          3123 => x"24",
          3124 => x"10",
          3125 => x"83",
          3126 => x"54",
          3127 => x"f7",
          3128 => x"59",
          3129 => x"81",
          3130 => x"59",
          3131 => x"9f",
          3132 => x"54",
          3133 => x"7b",
          3134 => x"76",
          3135 => x"7b",
          3136 => x"38",
          3137 => x"53",
          3138 => x"05",
          3139 => x"83",
          3140 => x"06",
          3141 => x"84",
          3142 => x"f9",
          3143 => x"74",
          3144 => x"52",
          3145 => x"b9",
          3146 => x"76",
          3147 => x"72",
          3148 => x"90",
          3149 => x"f7",
          3150 => x"0b",
          3151 => x"83",
          3152 => x"f7",
          3153 => x"81",
          3154 => x"fc",
          3155 => x"55",
          3156 => x"81",
          3157 => x"81",
          3158 => x"08",
          3159 => x"08",
          3160 => x"38",
          3161 => x"9c",
          3162 => x"d7",
          3163 => x"34",
          3164 => x"34",
          3165 => x"9e",
          3166 => x"0b",
          3167 => x"08",
          3168 => x"a4",
          3169 => x"42",
          3170 => x"79",
          3171 => x"38",
          3172 => x"38",
          3173 => x"c0",
          3174 => x"81",
          3175 => x"84",
          3176 => x"38",
          3177 => x"ff",
          3178 => x"b7",
          3179 => x"81",
          3180 => x"59",
          3181 => x"a8",
          3182 => x"0b",
          3183 => x"84",
          3184 => x"ff",
          3185 => x"83",
          3186 => x"23",
          3187 => x"53",
          3188 => x"73",
          3189 => x"33",
          3190 => x"53",
          3191 => x"72",
          3192 => x"b7",
          3193 => x"a5",
          3194 => x"54",
          3195 => x"83",
          3196 => x"81",
          3197 => x"ac",
          3198 => x"0d",
          3199 => x"0d",
          3200 => x"f3",
          3201 => x"33",
          3202 => x"51",
          3203 => x"f3",
          3204 => x"15",
          3205 => x"34",
          3206 => x"d4",
          3207 => x"87",
          3208 => x"98",
          3209 => x"38",
          3210 => x"08",
          3211 => x"71",
          3212 => x"98",
          3213 => x"27",
          3214 => x"2e",
          3215 => x"08",
          3216 => x"98",
          3217 => x"08",
          3218 => x"14",
          3219 => x"52",
          3220 => x"ff",
          3221 => x"08",
          3222 => x"52",
          3223 => x"06",
          3224 => x"74",
          3225 => x"38",
          3226 => x"b9",
          3227 => x"0b",
          3228 => x"04",
          3229 => x"a3",
          3230 => x"f3",
          3231 => x"80",
          3232 => x"51",
          3233 => x"72",
          3234 => x"71",
          3235 => x"72",
          3236 => x"52",
          3237 => x"08",
          3238 => x"83",
          3239 => x"81",
          3240 => x"e8",
          3241 => x"f3",
          3242 => x"53",
          3243 => x"c0",
          3244 => x"f6",
          3245 => x"9c",
          3246 => x"38",
          3247 => x"c0",
          3248 => x"73",
          3249 => x"ff",
          3250 => x"9c",
          3251 => x"c0",
          3252 => x"9c",
          3253 => x"81",
          3254 => x"52",
          3255 => x"81",
          3256 => x"a4",
          3257 => x"ff",
          3258 => x"ff",
          3259 => x"c7",
          3260 => x"fe",
          3261 => x"06",
          3262 => x"7b",
          3263 => x"73",
          3264 => x"53",
          3265 => x"72",
          3266 => x"c8",
          3267 => x"84",
          3268 => x"ff",
          3269 => x"02",
          3270 => x"80",
          3271 => x"2b",
          3272 => x"98",
          3273 => x"83",
          3274 => x"84",
          3275 => x"85",
          3276 => x"83",
          3277 => x"80",
          3278 => x"27",
          3279 => x"33",
          3280 => x"71",
          3281 => x"54",
          3282 => x"08",
          3283 => x"83",
          3284 => x"81",
          3285 => x"e8",
          3286 => x"f3",
          3287 => x"53",
          3288 => x"c0",
          3289 => x"f6",
          3290 => x"9c",
          3291 => x"38",
          3292 => x"c0",
          3293 => x"73",
          3294 => x"ff",
          3295 => x"9c",
          3296 => x"c0",
          3297 => x"9c",
          3298 => x"81",
          3299 => x"52",
          3300 => x"81",
          3301 => x"a4",
          3302 => x"ff",
          3303 => x"ff",
          3304 => x"38",
          3305 => x"d5",
          3306 => x"54",
          3307 => x"76",
          3308 => x"04",
          3309 => x"83",
          3310 => x"34",
          3311 => x"56",
          3312 => x"86",
          3313 => x"9c",
          3314 => x"ce",
          3315 => x"08",
          3316 => x"72",
          3317 => x"87",
          3318 => x"74",
          3319 => x"db",
          3320 => x"ff",
          3321 => x"71",
          3322 => x"87",
          3323 => x"05",
          3324 => x"87",
          3325 => x"2e",
          3326 => x"98",
          3327 => x"87",
          3328 => x"87",
          3329 => x"26",
          3330 => x"16",
          3331 => x"80",
          3332 => x"54",
          3333 => x"3d",
          3334 => x"bf",
          3335 => x"0d",
          3336 => x"83",
          3337 => x"83",
          3338 => x"33",
          3339 => x"77",
          3340 => x"98",
          3341 => x"41",
          3342 => x"57",
          3343 => x"72",
          3344 => x"71",
          3345 => x"05",
          3346 => x"2b",
          3347 => x"52",
          3348 => x"9e",
          3349 => x"71",
          3350 => x"05",
          3351 => x"74",
          3352 => x"54",
          3353 => x"08",
          3354 => x"33",
          3355 => x"5c",
          3356 => x"34",
          3357 => x"08",
          3358 => x"80",
          3359 => x"08",
          3360 => x"14",
          3361 => x"33",
          3362 => x"82",
          3363 => x"58",
          3364 => x"13",
          3365 => x"33",
          3366 => x"83",
          3367 => x"85",
          3368 => x"88",
          3369 => x"58",
          3370 => x"34",
          3371 => x"11",
          3372 => x"71",
          3373 => x"72",
          3374 => x"71",
          3375 => x"55",
          3376 => x"87",
          3377 => x"70",
          3378 => x"07",
          3379 => x"5a",
          3380 => x"81",
          3381 => x"17",
          3382 => x"2b",
          3383 => x"33",
          3384 => x"70",
          3385 => x"05",
          3386 => x"5c",
          3387 => x"34",
          3388 => x"08",
          3389 => x"71",
          3390 => x"05",
          3391 => x"2b",
          3392 => x"2a",
          3393 => x"52",
          3394 => x"84",
          3395 => x"33",
          3396 => x"83",
          3397 => x"12",
          3398 => x"07",
          3399 => x"53",
          3400 => x"33",
          3401 => x"82",
          3402 => x"59",
          3403 => x"34",
          3404 => x"33",
          3405 => x"83",
          3406 => x"83",
          3407 => x"88",
          3408 => x"52",
          3409 => x"15",
          3410 => x"0d",
          3411 => x"76",
          3412 => x"86",
          3413 => x"3d",
          3414 => x"b9",
          3415 => x"b4",
          3416 => x"84",
          3417 => x"84",
          3418 => x"81",
          3419 => x"08",
          3420 => x"85",
          3421 => x"76",
          3422 => x"34",
          3423 => x"22",
          3424 => x"83",
          3425 => x"51",
          3426 => x"89",
          3427 => x"10",
          3428 => x"f8",
          3429 => x"81",
          3430 => x"f7",
          3431 => x"51",
          3432 => x"83",
          3433 => x"06",
          3434 => x"84",
          3435 => x"12",
          3436 => x"59",
          3437 => x"75",
          3438 => x"10",
          3439 => x"71",
          3440 => x"06",
          3441 => x"70",
          3442 => x"52",
          3443 => x"2e",
          3444 => x"12",
          3445 => x"07",
          3446 => x"ff",
          3447 => x"56",
          3448 => x"33",
          3449 => x"70",
          3450 => x"56",
          3451 => x"81",
          3452 => x"8d",
          3453 => x"85",
          3454 => x"74",
          3455 => x"82",
          3456 => x"5c",
          3457 => x"81",
          3458 => x"76",
          3459 => x"34",
          3460 => x"08",
          3461 => x"71",
          3462 => x"ff",
          3463 => x"ff",
          3464 => x"57",
          3465 => x"72",
          3466 => x"34",
          3467 => x"74",
          3468 => x"b8",
          3469 => x"12",
          3470 => x"07",
          3471 => x"75",
          3472 => x"84",
          3473 => x"05",
          3474 => x"88",
          3475 => x"58",
          3476 => x"15",
          3477 => x"84",
          3478 => x"2b",
          3479 => x"5a",
          3480 => x"72",
          3481 => x"70",
          3482 => x"85",
          3483 => x"88",
          3484 => x"15",
          3485 => x"b8",
          3486 => x"b9",
          3487 => x"14",
          3488 => x"71",
          3489 => x"33",
          3490 => x"70",
          3491 => x"52",
          3492 => x"34",
          3493 => x"11",
          3494 => x"71",
          3495 => x"33",
          3496 => x"70",
          3497 => x"5b",
          3498 => x"87",
          3499 => x"70",
          3500 => x"07",
          3501 => x"59",
          3502 => x"81",
          3503 => x"84",
          3504 => x"0d",
          3505 => x"76",
          3506 => x"8a",
          3507 => x"3d",
          3508 => x"84",
          3509 => x"89",
          3510 => x"84",
          3511 => x"b9",
          3512 => x"52",
          3513 => x"3f",
          3514 => x"34",
          3515 => x"b8",
          3516 => x"0b",
          3517 => x"56",
          3518 => x"17",
          3519 => x"b4",
          3520 => x"70",
          3521 => x"58",
          3522 => x"73",
          3523 => x"70",
          3524 => x"05",
          3525 => x"34",
          3526 => x"77",
          3527 => x"39",
          3528 => x"80",
          3529 => x"41",
          3530 => x"80",
          3531 => x"88",
          3532 => x"8f",
          3533 => x"05",
          3534 => x"73",
          3535 => x"83",
          3536 => x"83",
          3537 => x"33",
          3538 => x"70",
          3539 => x"10",
          3540 => x"70",
          3541 => x"07",
          3542 => x"42",
          3543 => x"5c",
          3544 => x"7a",
          3545 => x"83",
          3546 => x"10",
          3547 => x"33",
          3548 => x"53",
          3549 => x"24",
          3550 => x"f6",
          3551 => x"87",
          3552 => x"38",
          3553 => x"be",
          3554 => x"92",
          3555 => x"12",
          3556 => x"07",
          3557 => x"71",
          3558 => x"43",
          3559 => x"60",
          3560 => x"11",
          3561 => x"71",
          3562 => x"33",
          3563 => x"83",
          3564 => x"85",
          3565 => x"88",
          3566 => x"58",
          3567 => x"34",
          3568 => x"08",
          3569 => x"33",
          3570 => x"74",
          3571 => x"71",
          3572 => x"42",
          3573 => x"86",
          3574 => x"b9",
          3575 => x"33",
          3576 => x"06",
          3577 => x"76",
          3578 => x"b9",
          3579 => x"83",
          3580 => x"2b",
          3581 => x"33",
          3582 => x"41",
          3583 => x"79",
          3584 => x"b9",
          3585 => x"12",
          3586 => x"07",
          3587 => x"33",
          3588 => x"41",
          3589 => x"79",
          3590 => x"84",
          3591 => x"33",
          3592 => x"66",
          3593 => x"52",
          3594 => x"fe",
          3595 => x"1e",
          3596 => x"83",
          3597 => x"62",
          3598 => x"84",
          3599 => x"84",
          3600 => x"a0",
          3601 => x"80",
          3602 => x"51",
          3603 => x"08",
          3604 => x"1f",
          3605 => x"84",
          3606 => x"84",
          3607 => x"34",
          3608 => x"b8",
          3609 => x"fe",
          3610 => x"06",
          3611 => x"78",
          3612 => x"84",
          3613 => x"84",
          3614 => x"56",
          3615 => x"15",
          3616 => x"fa",
          3617 => x"38",
          3618 => x"38",
          3619 => x"c8",
          3620 => x"0d",
          3621 => x"71",
          3622 => x"05",
          3623 => x"2b",
          3624 => x"2a",
          3625 => x"34",
          3626 => x"b8",
          3627 => x"75",
          3628 => x"84",
          3629 => x"81",
          3630 => x"83",
          3631 => x"64",
          3632 => x"4a",
          3633 => x"63",
          3634 => x"41",
          3635 => x"b8",
          3636 => x"81",
          3637 => x"05",
          3638 => x"54",
          3639 => x"83",
          3640 => x"39",
          3641 => x"70",
          3642 => x"83",
          3643 => x"10",
          3644 => x"33",
          3645 => x"53",
          3646 => x"73",
          3647 => x"39",
          3648 => x"7a",
          3649 => x"ff",
          3650 => x"38",
          3651 => x"84",
          3652 => x"b9",
          3653 => x"52",
          3654 => x"3f",
          3655 => x"34",
          3656 => x"b8",
          3657 => x"0b",
          3658 => x"58",
          3659 => x"19",
          3660 => x"b4",
          3661 => x"70",
          3662 => x"58",
          3663 => x"34",
          3664 => x"b4",
          3665 => x"b8",
          3666 => x"61",
          3667 => x"34",
          3668 => x"de",
          3669 => x"61",
          3670 => x"39",
          3671 => x"51",
          3672 => x"b9",
          3673 => x"1e",
          3674 => x"8b",
          3675 => x"86",
          3676 => x"2b",
          3677 => x"14",
          3678 => x"07",
          3679 => x"5b",
          3680 => x"64",
          3681 => x"34",
          3682 => x"11",
          3683 => x"71",
          3684 => x"33",
          3685 => x"70",
          3686 => x"59",
          3687 => x"7a",
          3688 => x"08",
          3689 => x"88",
          3690 => x"88",
          3691 => x"34",
          3692 => x"08",
          3693 => x"33",
          3694 => x"74",
          3695 => x"88",
          3696 => x"5e",
          3697 => x"34",
          3698 => x"08",
          3699 => x"71",
          3700 => x"05",
          3701 => x"88",
          3702 => x"40",
          3703 => x"18",
          3704 => x"b8",
          3705 => x"12",
          3706 => x"62",
          3707 => x"5d",
          3708 => x"de",
          3709 => x"05",
          3710 => x"fc",
          3711 => x"b9",
          3712 => x"b4",
          3713 => x"84",
          3714 => x"84",
          3715 => x"81",
          3716 => x"08",
          3717 => x"85",
          3718 => x"7f",
          3719 => x"34",
          3720 => x"22",
          3721 => x"83",
          3722 => x"43",
          3723 => x"89",
          3724 => x"10",
          3725 => x"f8",
          3726 => x"81",
          3727 => x"bd",
          3728 => x"19",
          3729 => x"71",
          3730 => x"33",
          3731 => x"70",
          3732 => x"55",
          3733 => x"85",
          3734 => x"1e",
          3735 => x"8b",
          3736 => x"86",
          3737 => x"2b",
          3738 => x"48",
          3739 => x"05",
          3740 => x"b9",
          3741 => x"33",
          3742 => x"06",
          3743 => x"75",
          3744 => x"b9",
          3745 => x"12",
          3746 => x"07",
          3747 => x"71",
          3748 => x"ff",
          3749 => x"48",
          3750 => x"41",
          3751 => x"34",
          3752 => x"33",
          3753 => x"83",
          3754 => x"12",
          3755 => x"ff",
          3756 => x"5e",
          3757 => x"76",
          3758 => x"ff",
          3759 => x"33",
          3760 => x"83",
          3761 => x"85",
          3762 => x"88",
          3763 => x"78",
          3764 => x"84",
          3765 => x"33",
          3766 => x"83",
          3767 => x"87",
          3768 => x"88",
          3769 => x"55",
          3770 => x"60",
          3771 => x"18",
          3772 => x"2b",
          3773 => x"2a",
          3774 => x"78",
          3775 => x"70",
          3776 => x"8b",
          3777 => x"70",
          3778 => x"07",
          3779 => x"77",
          3780 => x"5f",
          3781 => x"17",
          3782 => x"b8",
          3783 => x"33",
          3784 => x"74",
          3785 => x"88",
          3786 => x"88",
          3787 => x"5d",
          3788 => x"34",
          3789 => x"11",
          3790 => x"71",
          3791 => x"33",
          3792 => x"83",
          3793 => x"85",
          3794 => x"88",
          3795 => x"59",
          3796 => x"1d",
          3797 => x"b8",
          3798 => x"12",
          3799 => x"07",
          3800 => x"33",
          3801 => x"5f",
          3802 => x"77",
          3803 => x"84",
          3804 => x"12",
          3805 => x"ff",
          3806 => x"59",
          3807 => x"84",
          3808 => x"33",
          3809 => x"83",
          3810 => x"15",
          3811 => x"2a",
          3812 => x"55",
          3813 => x"84",
          3814 => x"81",
          3815 => x"2b",
          3816 => x"15",
          3817 => x"2a",
          3818 => x"55",
          3819 => x"34",
          3820 => x"11",
          3821 => x"07",
          3822 => x"42",
          3823 => x"51",
          3824 => x"08",
          3825 => x"70",
          3826 => x"f1",
          3827 => x"33",
          3828 => x"79",
          3829 => x"71",
          3830 => x"48",
          3831 => x"05",
          3832 => x"b9",
          3833 => x"85",
          3834 => x"2b",
          3835 => x"15",
          3836 => x"2a",
          3837 => x"56",
          3838 => x"87",
          3839 => x"70",
          3840 => x"07",
          3841 => x"5c",
          3842 => x"81",
          3843 => x"1f",
          3844 => x"2b",
          3845 => x"33",
          3846 => x"70",
          3847 => x"05",
          3848 => x"58",
          3849 => x"34",
          3850 => x"08",
          3851 => x"71",
          3852 => x"05",
          3853 => x"2b",
          3854 => x"2a",
          3855 => x"5b",
          3856 => x"77",
          3857 => x"39",
          3858 => x"84",
          3859 => x"08",
          3860 => x"52",
          3861 => x"be",
          3862 => x"5b",
          3863 => x"e9",
          3864 => x"84",
          3865 => x"2e",
          3866 => x"73",
          3867 => x"04",
          3868 => x"c8",
          3869 => x"2e",
          3870 => x"b9",
          3871 => x"73",
          3872 => x"04",
          3873 => x"0c",
          3874 => x"82",
          3875 => x"f4",
          3876 => x"b8",
          3877 => x"81",
          3878 => x"76",
          3879 => x"34",
          3880 => x"17",
          3881 => x"b9",
          3882 => x"05",
          3883 => x"ff",
          3884 => x"56",
          3885 => x"34",
          3886 => x"10",
          3887 => x"55",
          3888 => x"83",
          3889 => x"fe",
          3890 => x"0d",
          3891 => x"70",
          3892 => x"11",
          3893 => x"83",
          3894 => x"93",
          3895 => x"26",
          3896 => x"84",
          3897 => x"72",
          3898 => x"34",
          3899 => x"84",
          3900 => x"f7",
          3901 => x"05",
          3902 => x"81",
          3903 => x"b9",
          3904 => x"54",
          3905 => x"85",
          3906 => x"53",
          3907 => x"84",
          3908 => x"74",
          3909 => x"8c",
          3910 => x"26",
          3911 => x"54",
          3912 => x"73",
          3913 => x"3d",
          3914 => x"70",
          3915 => x"78",
          3916 => x"3d",
          3917 => x"af",
          3918 => x"54",
          3919 => x"c4",
          3920 => x"83",
          3921 => x"0b",
          3922 => x"75",
          3923 => x"b9",
          3924 => x"80",
          3925 => x"08",
          3926 => x"d6",
          3927 => x"73",
          3928 => x"55",
          3929 => x"0d",
          3930 => x"81",
          3931 => x"26",
          3932 => x"0d",
          3933 => x"02",
          3934 => x"55",
          3935 => x"84",
          3936 => x"06",
          3937 => x"0b",
          3938 => x"70",
          3939 => x"ad",
          3940 => x"53",
          3941 => x"0d",
          3942 => x"84",
          3943 => x"81",
          3944 => x"c8",
          3945 => x"2b",
          3946 => x"70",
          3947 => x"81",
          3948 => x"38",
          3949 => x"ea",
          3950 => x"70",
          3951 => x"92",
          3952 => x"54",
          3953 => x"08",
          3954 => x"90",
          3955 => x"0b",
          3956 => x"74",
          3957 => x"77",
          3958 => x"38",
          3959 => x"51",
          3960 => x"80",
          3961 => x"b9",
          3962 => x"54",
          3963 => x"53",
          3964 => x"3f",
          3965 => x"2e",
          3966 => x"c8",
          3967 => x"70",
          3968 => x"84",
          3969 => x"74",
          3970 => x"33",
          3971 => x"ff",
          3972 => x"79",
          3973 => x"3f",
          3974 => x"2e",
          3975 => x"18",
          3976 => x"06",
          3977 => x"80",
          3978 => x"05",
          3979 => x"38",
          3980 => x"ff",
          3981 => x"d2",
          3982 => x"34",
          3983 => x"c1",
          3984 => x"84",
          3985 => x"9d",
          3986 => x"19",
          3987 => x"34",
          3988 => x"19",
          3989 => x"a1",
          3990 => x"84",
          3991 => x"7a",
          3992 => x"5b",
          3993 => x"2a",
          3994 => x"90",
          3995 => x"7a",
          3996 => x"34",
          3997 => x"1a",
          3998 => x"52",
          3999 => x"76",
          4000 => x"81",
          4001 => x"b9",
          4002 => x"fd",
          4003 => x"70",
          4004 => x"88",
          4005 => x"38",
          4006 => x"8f",
          4007 => x"58",
          4008 => x"82",
          4009 => x"09",
          4010 => x"16",
          4011 => x"5a",
          4012 => x"2e",
          4013 => x"7b",
          4014 => x"81",
          4015 => x"17",
          4016 => x"c8",
          4017 => x"81",
          4018 => x"9a",
          4019 => x"11",
          4020 => x"1b",
          4021 => x"17",
          4022 => x"83",
          4023 => x"7d",
          4024 => x"81",
          4025 => x"17",
          4026 => x"c8",
          4027 => x"81",
          4028 => x"ca",
          4029 => x"11",
          4030 => x"81",
          4031 => x"59",
          4032 => x"ff",
          4033 => x"0d",
          4034 => x"05",
          4035 => x"38",
          4036 => x"5d",
          4037 => x"81",
          4038 => x"17",
          4039 => x"3f",
          4040 => x"38",
          4041 => x"0c",
          4042 => x"fe",
          4043 => x"33",
          4044 => x"b9",
          4045 => x"04",
          4046 => x"b8",
          4047 => x"05",
          4048 => x"38",
          4049 => x"5e",
          4050 => x"82",
          4051 => x"17",
          4052 => x"3f",
          4053 => x"38",
          4054 => x"0c",
          4055 => x"83",
          4056 => x"11",
          4057 => x"71",
          4058 => x"72",
          4059 => x"ff",
          4060 => x"c8",
          4061 => x"8f",
          4062 => x"08",
          4063 => x"33",
          4064 => x"84",
          4065 => x"06",
          4066 => x"83",
          4067 => x"08",
          4068 => x"7d",
          4069 => x"82",
          4070 => x"81",
          4071 => x"17",
          4072 => x"52",
          4073 => x"7a",
          4074 => x"17",
          4075 => x"18",
          4076 => x"b9",
          4077 => x"82",
          4078 => x"18",
          4079 => x"31",
          4080 => x"38",
          4081 => x"81",
          4082 => x"fb",
          4083 => x"53",
          4084 => x"52",
          4085 => x"b9",
          4086 => x"fd",
          4087 => x"18",
          4088 => x"31",
          4089 => x"a0",
          4090 => x"17",
          4091 => x"06",
          4092 => x"08",
          4093 => x"81",
          4094 => x"5a",
          4095 => x"08",
          4096 => x"33",
          4097 => x"84",
          4098 => x"06",
          4099 => x"83",
          4100 => x"08",
          4101 => x"74",
          4102 => x"82",
          4103 => x"81",
          4104 => x"17",
          4105 => x"52",
          4106 => x"7c",
          4107 => x"17",
          4108 => x"52",
          4109 => x"fa",
          4110 => x"38",
          4111 => x"62",
          4112 => x"76",
          4113 => x"27",
          4114 => x"2e",
          4115 => x"38",
          4116 => x"84",
          4117 => x"75",
          4118 => x"80",
          4119 => x"78",
          4120 => x"7c",
          4121 => x"06",
          4122 => x"b8",
          4123 => x"87",
          4124 => x"85",
          4125 => x"1a",
          4126 => x"75",
          4127 => x"83",
          4128 => x"1f",
          4129 => x"1f",
          4130 => x"84",
          4131 => x"74",
          4132 => x"38",
          4133 => x"58",
          4134 => x"76",
          4135 => x"33",
          4136 => x"81",
          4137 => x"53",
          4138 => x"f1",
          4139 => x"2e",
          4140 => x"b4",
          4141 => x"38",
          4142 => x"05",
          4143 => x"2b",
          4144 => x"07",
          4145 => x"7d",
          4146 => x"7d",
          4147 => x"7d",
          4148 => x"81",
          4149 => x"75",
          4150 => x"1b",
          4151 => x"5a",
          4152 => x"83",
          4153 => x"7d",
          4154 => x"81",
          4155 => x"19",
          4156 => x"c8",
          4157 => x"81",
          4158 => x"7b",
          4159 => x"19",
          4160 => x"5f",
          4161 => x"8f",
          4162 => x"77",
          4163 => x"74",
          4164 => x"7d",
          4165 => x"80",
          4166 => x"76",
          4167 => x"53",
          4168 => x"52",
          4169 => x"b9",
          4170 => x"80",
          4171 => x"1a",
          4172 => x"08",
          4173 => x"08",
          4174 => x"8b",
          4175 => x"2e",
          4176 => x"76",
          4177 => x"3f",
          4178 => x"38",
          4179 => x"0c",
          4180 => x"06",
          4181 => x"56",
          4182 => x"33",
          4183 => x"56",
          4184 => x"1a",
          4185 => x"53",
          4186 => x"52",
          4187 => x"b9",
          4188 => x"fc",
          4189 => x"1a",
          4190 => x"08",
          4191 => x"08",
          4192 => x"fb",
          4193 => x"82",
          4194 => x"81",
          4195 => x"19",
          4196 => x"fb",
          4197 => x"19",
          4198 => x"ee",
          4199 => x"08",
          4200 => x"38",
          4201 => x"b4",
          4202 => x"a0",
          4203 => x"40",
          4204 => x"38",
          4205 => x"09",
          4206 => x"7d",
          4207 => x"51",
          4208 => x"39",
          4209 => x"53",
          4210 => x"3f",
          4211 => x"2e",
          4212 => x"b9",
          4213 => x"08",
          4214 => x"08",
          4215 => x"5e",
          4216 => x"19",
          4217 => x"06",
          4218 => x"53",
          4219 => x"86",
          4220 => x"54",
          4221 => x"33",
          4222 => x"8b",
          4223 => x"7a",
          4224 => x"5f",
          4225 => x"2a",
          4226 => x"39",
          4227 => x"82",
          4228 => x"11",
          4229 => x"0a",
          4230 => x"58",
          4231 => x"88",
          4232 => x"90",
          4233 => x"98",
          4234 => x"cf",
          4235 => x"08",
          4236 => x"90",
          4237 => x"f4",
          4238 => x"ec",
          4239 => x"73",
          4240 => x"2e",
          4241 => x"56",
          4242 => x"82",
          4243 => x"75",
          4244 => x"b9",
          4245 => x"80",
          4246 => x"b1",
          4247 => x"30",
          4248 => x"07",
          4249 => x"38",
          4250 => x"b5",
          4251 => x"0c",
          4252 => x"91",
          4253 => x"39",
          4254 => x"81",
          4255 => x"db",
          4256 => x"b9",
          4257 => x"19",
          4258 => x"38",
          4259 => x"56",
          4260 => x"82",
          4261 => x"3f",
          4262 => x"2e",
          4263 => x"09",
          4264 => x"70",
          4265 => x"51",
          4266 => x"84",
          4267 => x"90",
          4268 => x"a3",
          4269 => x"9b",
          4270 => x"39",
          4271 => x"53",
          4272 => x"84",
          4273 => x"30",
          4274 => x"25",
          4275 => x"74",
          4276 => x"9c",
          4277 => x"56",
          4278 => x"15",
          4279 => x"07",
          4280 => x"74",
          4281 => x"04",
          4282 => x"3d",
          4283 => x"fe",
          4284 => x"38",
          4285 => x"8b",
          4286 => x"a7",
          4287 => x"c8",
          4288 => x"74",
          4289 => x"ff",
          4290 => x"71",
          4291 => x"0a",
          4292 => x"53",
          4293 => x"0c",
          4294 => x"38",
          4295 => x"cc",
          4296 => x"88",
          4297 => x"a9",
          4298 => x"74",
          4299 => x"82",
          4300 => x"89",
          4301 => x"ff",
          4302 => x"80",
          4303 => x"3d",
          4304 => x"0c",
          4305 => x"55",
          4306 => x"17",
          4307 => x"76",
          4308 => x"fe",
          4309 => x"75",
          4310 => x"76",
          4311 => x"53",
          4312 => x"74",
          4313 => x"b9",
          4314 => x"ff",
          4315 => x"c8",
          4316 => x"08",
          4317 => x"ff",
          4318 => x"76",
          4319 => x"0b",
          4320 => x"04",
          4321 => x"12",
          4322 => x"80",
          4323 => x"98",
          4324 => x"56",
          4325 => x"ff",
          4326 => x"94",
          4327 => x"79",
          4328 => x"74",
          4329 => x"18",
          4330 => x"b8",
          4331 => x"84",
          4332 => x"77",
          4333 => x"05",
          4334 => x"38",
          4335 => x"84",
          4336 => x"0b",
          4337 => x"81",
          4338 => x"c6",
          4339 => x"08",
          4340 => x"81",
          4341 => x"51",
          4342 => x"5d",
          4343 => x"2e",
          4344 => x"c8",
          4345 => x"56",
          4346 => x"86",
          4347 => x"33",
          4348 => x"18",
          4349 => x"80",
          4350 => x"19",
          4351 => x"05",
          4352 => x"19",
          4353 => x"76",
          4354 => x"55",
          4355 => x"22",
          4356 => x"81",
          4357 => x"19",
          4358 => x"c8",
          4359 => x"dd",
          4360 => x"84",
          4361 => x"75",
          4362 => x"70",
          4363 => x"86",
          4364 => x"38",
          4365 => x"b4",
          4366 => x"74",
          4367 => x"82",
          4368 => x"81",
          4369 => x"19",
          4370 => x"52",
          4371 => x"fe",
          4372 => x"83",
          4373 => x"09",
          4374 => x"0c",
          4375 => x"5e",
          4376 => x"85",
          4377 => x"b0",
          4378 => x"fc",
          4379 => x"0c",
          4380 => x"64",
          4381 => x"5b",
          4382 => x"5e",
          4383 => x"b8",
          4384 => x"19",
          4385 => x"19",
          4386 => x"09",
          4387 => x"75",
          4388 => x"51",
          4389 => x"80",
          4390 => x"79",
          4391 => x"90",
          4392 => x"58",
          4393 => x"18",
          4394 => x"5b",
          4395 => x"e5",
          4396 => x"30",
          4397 => x"54",
          4398 => x"74",
          4399 => x"2e",
          4400 => x"86",
          4401 => x"51",
          4402 => x"5b",
          4403 => x"98",
          4404 => x"7a",
          4405 => x"04",
          4406 => x"52",
          4407 => x"81",
          4408 => x"09",
          4409 => x"c8",
          4410 => x"a8",
          4411 => x"58",
          4412 => x"b5",
          4413 => x"2e",
          4414 => x"54",
          4415 => x"53",
          4416 => x"de",
          4417 => x"8f",
          4418 => x"76",
          4419 => x"2e",
          4420 => x"bf",
          4421 => x"05",
          4422 => x"ab",
          4423 => x"cc",
          4424 => x"81",
          4425 => x"5b",
          4426 => x"b9",
          4427 => x"5b",
          4428 => x"7d",
          4429 => x"8c",
          4430 => x"33",
          4431 => x"75",
          4432 => x"bf",
          4433 => x"81",
          4434 => x"33",
          4435 => x"71",
          4436 => x"80",
          4437 => x"26",
          4438 => x"76",
          4439 => x"5a",
          4440 => x"38",
          4441 => x"59",
          4442 => x"81",
          4443 => x"61",
          4444 => x"70",
          4445 => x"39",
          4446 => x"81",
          4447 => x"38",
          4448 => x"75",
          4449 => x"05",
          4450 => x"ff",
          4451 => x"e4",
          4452 => x"ff",
          4453 => x"c8",
          4454 => x"0d",
          4455 => x"7b",
          4456 => x"08",
          4457 => x"38",
          4458 => x"ac",
          4459 => x"08",
          4460 => x"2e",
          4461 => x"58",
          4462 => x"81",
          4463 => x"1b",
          4464 => x"3f",
          4465 => x"38",
          4466 => x"0c",
          4467 => x"1c",
          4468 => x"2e",
          4469 => x"06",
          4470 => x"86",
          4471 => x"f2",
          4472 => x"75",
          4473 => x"e2",
          4474 => x"7c",
          4475 => x"57",
          4476 => x"05",
          4477 => x"76",
          4478 => x"59",
          4479 => x"2e",
          4480 => x"06",
          4481 => x"1d",
          4482 => x"33",
          4483 => x"71",
          4484 => x"76",
          4485 => x"2e",
          4486 => x"ac",
          4487 => x"c8",
          4488 => x"b9",
          4489 => x"79",
          4490 => x"04",
          4491 => x"52",
          4492 => x"81",
          4493 => x"09",
          4494 => x"c8",
          4495 => x"a8",
          4496 => x"58",
          4497 => x"ea",
          4498 => x"2e",
          4499 => x"54",
          4500 => x"53",
          4501 => x"b6",
          4502 => x"5a",
          4503 => x"86",
          4504 => x"f2",
          4505 => x"79",
          4506 => x"77",
          4507 => x"7f",
          4508 => x"7d",
          4509 => x"5d",
          4510 => x"84",
          4511 => x"08",
          4512 => x"39",
          4513 => x"ff",
          4514 => x"a2",
          4515 => x"2e",
          4516 => x"08",
          4517 => x"88",
          4518 => x"b3",
          4519 => x"29",
          4520 => x"56",
          4521 => x"81",
          4522 => x"07",
          4523 => x"ed",
          4524 => x"38",
          4525 => x"b9",
          4526 => x"22",
          4527 => x"a0",
          4528 => x"2e",
          4529 => x"56",
          4530 => x"b0",
          4531 => x"06",
          4532 => x"74",
          4533 => x"05",
          4534 => x"38",
          4535 => x"5a",
          4536 => x"c8",
          4537 => x"ff",
          4538 => x"55",
          4539 => x"70",
          4540 => x"06",
          4541 => x"85",
          4542 => x"22",
          4543 => x"38",
          4544 => x"51",
          4545 => x"a0",
          4546 => x"58",
          4547 => x"77",
          4548 => x"55",
          4549 => x"33",
          4550 => x"2e",
          4551 => x"1f",
          4552 => x"8c",
          4553 => x"61",
          4554 => x"59",
          4555 => x"ff",
          4556 => x"27",
          4557 => x"57",
          4558 => x"1a",
          4559 => x"77",
          4560 => x"ff",
          4561 => x"44",
          4562 => x"38",
          4563 => x"18",
          4564 => x"22",
          4565 => x"05",
          4566 => x"07",
          4567 => x"38",
          4568 => x"16",
          4569 => x"56",
          4570 => x"fe",
          4571 => x"78",
          4572 => x"a0",
          4573 => x"78",
          4574 => x"33",
          4575 => x"06",
          4576 => x"77",
          4577 => x"05",
          4578 => x"59",
          4579 => x"87",
          4580 => x"84",
          4581 => x"5b",
          4582 => x"87",
          4583 => x"38",
          4584 => x"c8",
          4585 => x"d6",
          4586 => x"1f",
          4587 => x"db",
          4588 => x"81",
          4589 => x"90",
          4590 => x"8a",
          4591 => x"5b",
          4592 => x"84",
          4593 => x"08",
          4594 => x"b8",
          4595 => x"80",
          4596 => x"f3",
          4597 => x"2e",
          4598 => x"54",
          4599 => x"33",
          4600 => x"08",
          4601 => x"57",
          4602 => x"bc",
          4603 => x"42",
          4604 => x"74",
          4605 => x"5f",
          4606 => x"19",
          4607 => x"81",
          4608 => x"b9",
          4609 => x"80",
          4610 => x"84",
          4611 => x"81",
          4612 => x"f3",
          4613 => x"08",
          4614 => x"78",
          4615 => x"54",
          4616 => x"33",
          4617 => x"08",
          4618 => x"56",
          4619 => x"80",
          4620 => x"57",
          4621 => x"34",
          4622 => x"0b",
          4623 => x"75",
          4624 => x"81",
          4625 => x"ef",
          4626 => x"98",
          4627 => x"81",
          4628 => x"84",
          4629 => x"81",
          4630 => x"57",
          4631 => x"59",
          4632 => x"84",
          4633 => x"08",
          4634 => x"39",
          4635 => x"52",
          4636 => x"84",
          4637 => x"06",
          4638 => x"83",
          4639 => x"08",
          4640 => x"8b",
          4641 => x"2e",
          4642 => x"57",
          4643 => x"1f",
          4644 => x"e9",
          4645 => x"84",
          4646 => x"84",
          4647 => x"74",
          4648 => x"78",
          4649 => x"05",
          4650 => x"56",
          4651 => x"06",
          4652 => x"57",
          4653 => x"b2",
          4654 => x"2e",
          4655 => x"54",
          4656 => x"33",
          4657 => x"08",
          4658 => x"56",
          4659 => x"fe",
          4660 => x"08",
          4661 => x"60",
          4662 => x"34",
          4663 => x"34",
          4664 => x"f3",
          4665 => x"83",
          4666 => x"1f",
          4667 => x"83",
          4668 => x"76",
          4669 => x"88",
          4670 => x"38",
          4671 => x"8c",
          4672 => x"ff",
          4673 => x"70",
          4674 => x"a6",
          4675 => x"1d",
          4676 => x"3f",
          4677 => x"c8",
          4678 => x"40",
          4679 => x"81",
          4680 => x"70",
          4681 => x"96",
          4682 => x"fc",
          4683 => x"1d",
          4684 => x"31",
          4685 => x"a0",
          4686 => x"1c",
          4687 => x"06",
          4688 => x"08",
          4689 => x"81",
          4690 => x"56",
          4691 => x"70",
          4692 => x"2e",
          4693 => x"ff",
          4694 => x"2e",
          4695 => x"80",
          4696 => x"54",
          4697 => x"1c",
          4698 => x"c8",
          4699 => x"38",
          4700 => x"b4",
          4701 => x"74",
          4702 => x"1c",
          4703 => x"84",
          4704 => x"75",
          4705 => x"fa",
          4706 => x"57",
          4707 => x"75",
          4708 => x"39",
          4709 => x"08",
          4710 => x"51",
          4711 => x"54",
          4712 => x"53",
          4713 => x"96",
          4714 => x"7f",
          4715 => x"0b",
          4716 => x"2e",
          4717 => x"2e",
          4718 => x"8c",
          4719 => x"5c",
          4720 => x"54",
          4721 => x"55",
          4722 => x"80",
          4723 => x"5a",
          4724 => x"73",
          4725 => x"58",
          4726 => x"70",
          4727 => x"5c",
          4728 => x"0b",
          4729 => x"59",
          4730 => x"33",
          4731 => x"2e",
          4732 => x"38",
          4733 => x"07",
          4734 => x"26",
          4735 => x"ae",
          4736 => x"18",
          4737 => x"34",
          4738 => x"ba",
          4739 => x"0b",
          4740 => x"72",
          4741 => x"0b",
          4742 => x"94",
          4743 => x"9c",
          4744 => x"73",
          4745 => x"1c",
          4746 => x"34",
          4747 => x"33",
          4748 => x"88",
          4749 => x"07",
          4750 => x"0c",
          4751 => x"71",
          4752 => x"5a",
          4753 => x"99",
          4754 => x"2b",
          4755 => x"8f",
          4756 => x"c0",
          4757 => x"7a",
          4758 => x"7a",
          4759 => x"89",
          4760 => x"ff",
          4761 => x"38",
          4762 => x"88",
          4763 => x"18",
          4764 => x"8c",
          4765 => x"11",
          4766 => x"90",
          4767 => x"30",
          4768 => x"25",
          4769 => x"38",
          4770 => x"80",
          4771 => x"39",
          4772 => x"57",
          4773 => x"96",
          4774 => x"33",
          4775 => x"26",
          4776 => x"33",
          4777 => x"72",
          4778 => x"7d",
          4779 => x"83",
          4780 => x"70",
          4781 => x"16",
          4782 => x"57",
          4783 => x"fd",
          4784 => x"39",
          4785 => x"30",
          4786 => x"a9",
          4787 => x"70",
          4788 => x"57",
          4789 => x"81",
          4790 => x"38",
          4791 => x"16",
          4792 => x"3d",
          4793 => x"27",
          4794 => x"08",
          4795 => x"05",
          4796 => x"38",
          4797 => x"ec",
          4798 => x"38",
          4799 => x"81",
          4800 => x"70",
          4801 => x"71",
          4802 => x"73",
          4803 => x"82",
          4804 => x"38",
          4805 => x"33",
          4806 => x"73",
          4807 => x"2e",
          4808 => x"81",
          4809 => x"38",
          4810 => x"84",
          4811 => x"38",
          4812 => x"81",
          4813 => x"33",
          4814 => x"f0",
          4815 => x"dc",
          4816 => x"07",
          4817 => x"a1",
          4818 => x"74",
          4819 => x"38",
          4820 => x"80",
          4821 => x"e1",
          4822 => x"96",
          4823 => x"9f",
          4824 => x"b5",
          4825 => x"84",
          4826 => x"54",
          4827 => x"84",
          4828 => x"83",
          4829 => x"5c",
          4830 => x"e4",
          4831 => x"80",
          4832 => x"b9",
          4833 => x"3d",
          4834 => x"70",
          4835 => x"55",
          4836 => x"81",
          4837 => x"55",
          4838 => x"80",
          4839 => x"78",
          4840 => x"73",
          4841 => x"5a",
          4842 => x"82",
          4843 => x"76",
          4844 => x"11",
          4845 => x"70",
          4846 => x"5f",
          4847 => x"72",
          4848 => x"38",
          4849 => x"23",
          4850 => x"78",
          4851 => x"58",
          4852 => x"e6",
          4853 => x"72",
          4854 => x"2e",
          4855 => x"22",
          4856 => x"76",
          4857 => x"57",
          4858 => x"70",
          4859 => x"81",
          4860 => x"55",
          4861 => x"34",
          4862 => x"73",
          4863 => x"81",
          4864 => x"2e",
          4865 => x"d0",
          4866 => x"80",
          4867 => x"85",
          4868 => x"59",
          4869 => x"75",
          4870 => x"80",
          4871 => x"54",
          4872 => x"8b",
          4873 => x"8a",
          4874 => x"26",
          4875 => x"7e",
          4876 => x"57",
          4877 => x"18",
          4878 => x"a0",
          4879 => x"83",
          4880 => x"38",
          4881 => x"82",
          4882 => x"83",
          4883 => x"81",
          4884 => x"06",
          4885 => x"90",
          4886 => x"5e",
          4887 => x"07",
          4888 => x"e4",
          4889 => x"1d",
          4890 => x"80",
          4891 => x"08",
          4892 => x"38",
          4893 => x"80",
          4894 => x"81",
          4895 => x"08",
          4896 => x"08",
          4897 => x"16",
          4898 => x"40",
          4899 => x"75",
          4900 => x"07",
          4901 => x"56",
          4902 => x"ac",
          4903 => x"09",
          4904 => x"18",
          4905 => x"1d",
          4906 => x"83",
          4907 => x"05",
          4908 => x"27",
          4909 => x"ab",
          4910 => x"84",
          4911 => x"54",
          4912 => x"74",
          4913 => x"ce",
          4914 => x"81",
          4915 => x"cd",
          4916 => x"60",
          4917 => x"12",
          4918 => x"41",
          4919 => x"d8",
          4920 => x"65",
          4921 => x"55",
          4922 => x"17",
          4923 => x"39",
          4924 => x"fd",
          4925 => x"06",
          4926 => x"2e",
          4927 => x"82",
          4928 => x"a0",
          4929 => x"06",
          4930 => x"0b",
          4931 => x"c8",
          4932 => x"ff",
          4933 => x"80",
          4934 => x"26",
          4935 => x"77",
          4936 => x"79",
          4937 => x"51",
          4938 => x"08",
          4939 => x"81",
          4940 => x"38",
          4941 => x"11",
          4942 => x"ff",
          4943 => x"38",
          4944 => x"33",
          4945 => x"73",
          4946 => x"2e",
          4947 => x"81",
          4948 => x"38",
          4949 => x"d4",
          4950 => x"26",
          4951 => x"ff",
          4952 => x"78",
          4953 => x"70",
          4954 => x"ff",
          4955 => x"1b",
          4956 => x"1b",
          4957 => x"80",
          4958 => x"33",
          4959 => x"80",
          4960 => x"83",
          4961 => x"55",
          4962 => x"39",
          4963 => x"33",
          4964 => x"77",
          4965 => x"95",
          4966 => x"2a",
          4967 => x"7c",
          4968 => x"34",
          4969 => x"83",
          4970 => x"81",
          4971 => x"38",
          4972 => x"06",
          4973 => x"84",
          4974 => x"eb",
          4975 => x"80",
          4976 => x"61",
          4977 => x"42",
          4978 => x"70",
          4979 => x"56",
          4980 => x"74",
          4981 => x"38",
          4982 => x"24",
          4983 => x"d1",
          4984 => x"58",
          4985 => x"61",
          4986 => x"5d",
          4987 => x"17",
          4988 => x"b9",
          4989 => x"06",
          4990 => x"38",
          4991 => x"b9",
          4992 => x"52",
          4993 => x"3f",
          4994 => x"70",
          4995 => x"84",
          4996 => x"75",
          4997 => x"60",
          4998 => x"18",
          4999 => x"7b",
          5000 => x"17",
          5001 => x"ff",
          5002 => x"7b",
          5003 => x"74",
          5004 => x"38",
          5005 => x"33",
          5006 => x"56",
          5007 => x"38",
          5008 => x"bd",
          5009 => x"81",
          5010 => x"8d",
          5011 => x"80",
          5012 => x"71",
          5013 => x"80",
          5014 => x"80",
          5015 => x"71",
          5016 => x"38",
          5017 => x"12",
          5018 => x"07",
          5019 => x"2b",
          5020 => x"43",
          5021 => x"80",
          5022 => x"c8",
          5023 => x"06",
          5024 => x"26",
          5025 => x"76",
          5026 => x"5f",
          5027 => x"77",
          5028 => x"78",
          5029 => x"ca",
          5030 => x"88",
          5031 => x"23",
          5032 => x"58",
          5033 => x"33",
          5034 => x"07",
          5035 => x"17",
          5036 => x"90",
          5037 => x"33",
          5038 => x"71",
          5039 => x"42",
          5040 => x"33",
          5041 => x"58",
          5042 => x"1c",
          5043 => x"26",
          5044 => x"31",
          5045 => x"c8",
          5046 => x"2e",
          5047 => x"80",
          5048 => x"83",
          5049 => x"38",
          5050 => x"eb",
          5051 => x"19",
          5052 => x"70",
          5053 => x"0c",
          5054 => x"38",
          5055 => x"80",
          5056 => x"18",
          5057 => x"8d",
          5058 => x"7a",
          5059 => x"15",
          5060 => x"18",
          5061 => x"18",
          5062 => x"80",
          5063 => x"86",
          5064 => x"a0",
          5065 => x"a0",
          5066 => x"a8",
          5067 => x"18",
          5068 => x"0c",
          5069 => x"b9",
          5070 => x"33",
          5071 => x"57",
          5072 => x"17",
          5073 => x"59",
          5074 => x"7e",
          5075 => x"7c",
          5076 => x"05",
          5077 => x"33",
          5078 => x"99",
          5079 => x"ff",
          5080 => x"77",
          5081 => x"81",
          5082 => x"9f",
          5083 => x"81",
          5084 => x"78",
          5085 => x"9f",
          5086 => x"80",
          5087 => x"1e",
          5088 => x"38",
          5089 => x"2e",
          5090 => x"06",
          5091 => x"80",
          5092 => x"57",
          5093 => x"06",
          5094 => x"32",
          5095 => x"5a",
          5096 => x"81",
          5097 => x"77",
          5098 => x"33",
          5099 => x"38",
          5100 => x"33",
          5101 => x"83",
          5102 => x"2b",
          5103 => x"59",
          5104 => x"84",
          5105 => x"57",
          5106 => x"84",
          5107 => x"9f",
          5108 => x"10",
          5109 => x"44",
          5110 => x"5b",
          5111 => x"38",
          5112 => x"b4",
          5113 => x"ff",
          5114 => x"b8",
          5115 => x"b4",
          5116 => x"2e",
          5117 => x"b4",
          5118 => x"81",
          5119 => x"07",
          5120 => x"d5",
          5121 => x"0b",
          5122 => x"e9",
          5123 => x"32",
          5124 => x"42",
          5125 => x"e8",
          5126 => x"ff",
          5127 => x"1e",
          5128 => x"81",
          5129 => x"27",
          5130 => x"b7",
          5131 => x"83",
          5132 => x"39",
          5133 => x"f8",
          5134 => x"5d",
          5135 => x"71",
          5136 => x"56",
          5137 => x"80",
          5138 => x"18",
          5139 => x"70",
          5140 => x"05",
          5141 => x"5b",
          5142 => x"8e",
          5143 => x"58",
          5144 => x"93",
          5145 => x"3d",
          5146 => x"fe",
          5147 => x"83",
          5148 => x"39",
          5149 => x"3d",
          5150 => x"83",
          5151 => x"81",
          5152 => x"5c",
          5153 => x"57",
          5154 => x"38",
          5155 => x"81",
          5156 => x"58",
          5157 => x"70",
          5158 => x"ff",
          5159 => x"2e",
          5160 => x"38",
          5161 => x"fc",
          5162 => x"80",
          5163 => x"71",
          5164 => x"2e",
          5165 => x"1b",
          5166 => x"2e",
          5167 => x"7a",
          5168 => x"81",
          5169 => x"17",
          5170 => x"b9",
          5171 => x"58",
          5172 => x"f9",
          5173 => x"b7",
          5174 => x"88",
          5175 => x"d5",
          5176 => x"b8",
          5177 => x"71",
          5178 => x"14",
          5179 => x"33",
          5180 => x"5c",
          5181 => x"2e",
          5182 => x"9c",
          5183 => x"71",
          5184 => x"14",
          5185 => x"33",
          5186 => x"5a",
          5187 => x"2e",
          5188 => x"a0",
          5189 => x"71",
          5190 => x"14",
          5191 => x"33",
          5192 => x"a4",
          5193 => x"71",
          5194 => x"14",
          5195 => x"33",
          5196 => x"44",
          5197 => x"56",
          5198 => x"22",
          5199 => x"23",
          5200 => x"0b",
          5201 => x"0c",
          5202 => x"f0",
          5203 => x"95",
          5204 => x"b8",
          5205 => x"59",
          5206 => x"08",
          5207 => x"38",
          5208 => x"b4",
          5209 => x"7f",
          5210 => x"17",
          5211 => x"38",
          5212 => x"39",
          5213 => x"38",
          5214 => x"fc",
          5215 => x"e3",
          5216 => x"88",
          5217 => x"f6",
          5218 => x"f6",
          5219 => x"33",
          5220 => x"88",
          5221 => x"07",
          5222 => x"1e",
          5223 => x"44",
          5224 => x"58",
          5225 => x"58",
          5226 => x"a8",
          5227 => x"59",
          5228 => x"da",
          5229 => x"17",
          5230 => x"52",
          5231 => x"3f",
          5232 => x"80",
          5233 => x"3d",
          5234 => x"75",
          5235 => x"81",
          5236 => x"55",
          5237 => x"ed",
          5238 => x"84",
          5239 => x"80",
          5240 => x"90",
          5241 => x"2e",
          5242 => x"73",
          5243 => x"62",
          5244 => x"80",
          5245 => x"70",
          5246 => x"84",
          5247 => x"c8",
          5248 => x"84",
          5249 => x"75",
          5250 => x"56",
          5251 => x"82",
          5252 => x"5c",
          5253 => x"80",
          5254 => x"5b",
          5255 => x"81",
          5256 => x"5a",
          5257 => x"76",
          5258 => x"81",
          5259 => x"57",
          5260 => x"70",
          5261 => x"70",
          5262 => x"09",
          5263 => x"38",
          5264 => x"07",
          5265 => x"79",
          5266 => x"1d",
          5267 => x"38",
          5268 => x"24",
          5269 => x"fe",
          5270 => x"84",
          5271 => x"89",
          5272 => x"bf",
          5273 => x"53",
          5274 => x"9f",
          5275 => x"b9",
          5276 => x"79",
          5277 => x"0c",
          5278 => x"52",
          5279 => x"3f",
          5280 => x"c8",
          5281 => x"9c",
          5282 => x"38",
          5283 => x"84",
          5284 => x"58",
          5285 => x"81",
          5286 => x"38",
          5287 => x"71",
          5288 => x"58",
          5289 => x"e9",
          5290 => x"0b",
          5291 => x"34",
          5292 => x"56",
          5293 => x"57",
          5294 => x"0b",
          5295 => x"83",
          5296 => x"0b",
          5297 => x"34",
          5298 => x"9f",
          5299 => x"16",
          5300 => x"7e",
          5301 => x"57",
          5302 => x"9c",
          5303 => x"82",
          5304 => x"02",
          5305 => x"5d",
          5306 => x"86",
          5307 => x"b8",
          5308 => x"c2",
          5309 => x"5d",
          5310 => x"2a",
          5311 => x"38",
          5312 => x"38",
          5313 => x"80",
          5314 => x"58",
          5315 => x"67",
          5316 => x"9a",
          5317 => x"33",
          5318 => x"2e",
          5319 => x"9c",
          5320 => x"71",
          5321 => x"14",
          5322 => x"33",
          5323 => x"60",
          5324 => x"5d",
          5325 => x"77",
          5326 => x"34",
          5327 => x"2a",
          5328 => x"ac",
          5329 => x"75",
          5330 => x"89",
          5331 => x"70",
          5332 => x"76",
          5333 => x"06",
          5334 => x"38",
          5335 => x"3f",
          5336 => x"c8",
          5337 => x"84",
          5338 => x"38",
          5339 => x"80",
          5340 => x"95",
          5341 => x"74",
          5342 => x"80",
          5343 => x"80",
          5344 => x"80",
          5345 => x"cd",
          5346 => x"88",
          5347 => x"fc",
          5348 => x"57",
          5349 => x"17",
          5350 => x"07",
          5351 => x"39",
          5352 => x"38",
          5353 => x"3f",
          5354 => x"c8",
          5355 => x"b9",
          5356 => x"84",
          5357 => x"38",
          5358 => x"b2",
          5359 => x"90",
          5360 => x"19",
          5361 => x"ff",
          5362 => x"84",
          5363 => x"18",
          5364 => x"a0",
          5365 => x"17",
          5366 => x"cc",
          5367 => x"71",
          5368 => x"07",
          5369 => x"34",
          5370 => x"90",
          5371 => x"34",
          5372 => x"7e",
          5373 => x"34",
          5374 => x"5d",
          5375 => x"84",
          5376 => x"72",
          5377 => x"7e",
          5378 => x"79",
          5379 => x"81",
          5380 => x"16",
          5381 => x"b9",
          5382 => x"57",
          5383 => x"56",
          5384 => x"7a",
          5385 => x"0c",
          5386 => x"08",
          5387 => x"33",
          5388 => x"b9",
          5389 => x"81",
          5390 => x"17",
          5391 => x"31",
          5392 => x"a0",
          5393 => x"16",
          5394 => x"06",
          5395 => x"08",
          5396 => x"81",
          5397 => x"7c",
          5398 => x"0c",
          5399 => x"1a",
          5400 => x"ff",
          5401 => x"38",
          5402 => x"05",
          5403 => x"df",
          5404 => x"b0",
          5405 => x"2e",
          5406 => x"9c",
          5407 => x"75",
          5408 => x"39",
          5409 => x"39",
          5410 => x"0c",
          5411 => x"fe",
          5412 => x"67",
          5413 => x"0c",
          5414 => x"79",
          5415 => x"75",
          5416 => x"86",
          5417 => x"78",
          5418 => x"74",
          5419 => x"91",
          5420 => x"90",
          5421 => x"76",
          5422 => x"08",
          5423 => x"7b",
          5424 => x"2e",
          5425 => x"ff",
          5426 => x"19",
          5427 => x"5b",
          5428 => x"88",
          5429 => x"85",
          5430 => x"74",
          5431 => x"08",
          5432 => x"41",
          5433 => x"8a",
          5434 => x"08",
          5435 => x"d5",
          5436 => x"57",
          5437 => x"1b",
          5438 => x"7b",
          5439 => x"52",
          5440 => x"3f",
          5441 => x"60",
          5442 => x"2e",
          5443 => x"56",
          5444 => x"76",
          5445 => x"55",
          5446 => x"70",
          5447 => x"74",
          5448 => x"78",
          5449 => x"1e",
          5450 => x"1d",
          5451 => x"80",
          5452 => x"3d",
          5453 => x"92",
          5454 => x"39",
          5455 => x"06",
          5456 => x"78",
          5457 => x"b4",
          5458 => x"0b",
          5459 => x"7f",
          5460 => x"38",
          5461 => x"81",
          5462 => x"84",
          5463 => x"ff",
          5464 => x"7a",
          5465 => x"83",
          5466 => x"b8",
          5467 => x"e6",
          5468 => x"77",
          5469 => x"56",
          5470 => x"70",
          5471 => x"05",
          5472 => x"38",
          5473 => x"08",
          5474 => x"33",
          5475 => x"5b",
          5476 => x"81",
          5477 => x"08",
          5478 => x"1a",
          5479 => x"55",
          5480 => x"38",
          5481 => x"09",
          5482 => x"b4",
          5483 => x"7f",
          5484 => x"fe",
          5485 => x"9c",
          5486 => x"84",
          5487 => x"ff",
          5488 => x"55",
          5489 => x"ff",
          5490 => x"81",
          5491 => x"7a",
          5492 => x"0b",
          5493 => x"c8",
          5494 => x"91",
          5495 => x"0c",
          5496 => x"62",
          5497 => x"80",
          5498 => x"9f",
          5499 => x"97",
          5500 => x"8f",
          5501 => x"59",
          5502 => x"80",
          5503 => x"c4",
          5504 => x"bc",
          5505 => x"81",
          5506 => x"2e",
          5507 => x"11",
          5508 => x"76",
          5509 => x"38",
          5510 => x"a2",
          5511 => x"78",
          5512 => x"38",
          5513 => x"55",
          5514 => x"81",
          5515 => x"86",
          5516 => x"1a",
          5517 => x"60",
          5518 => x"2e",
          5519 => x"05",
          5520 => x"77",
          5521 => x"22",
          5522 => x"56",
          5523 => x"78",
          5524 => x"80",
          5525 => x"76",
          5526 => x"58",
          5527 => x"16",
          5528 => x"b9",
          5529 => x"11",
          5530 => x"27",
          5531 => x"76",
          5532 => x"70",
          5533 => x"05",
          5534 => x"38",
          5535 => x"89",
          5536 => x"1a",
          5537 => x"1b",
          5538 => x"08",
          5539 => x"27",
          5540 => x"0c",
          5541 => x"58",
          5542 => x"1b",
          5543 => x"0c",
          5544 => x"c8",
          5545 => x"33",
          5546 => x"fe",
          5547 => x"56",
          5548 => x"31",
          5549 => x"7a",
          5550 => x"2e",
          5551 => x"71",
          5552 => x"81",
          5553 => x"53",
          5554 => x"ff",
          5555 => x"80",
          5556 => x"76",
          5557 => x"60",
          5558 => x"7a",
          5559 => x"78",
          5560 => x"05",
          5561 => x"34",
          5562 => x"58",
          5563 => x"39",
          5564 => x"16",
          5565 => x"ff",
          5566 => x"c8",
          5567 => x"ab",
          5568 => x"34",
          5569 => x"84",
          5570 => x"17",
          5571 => x"33",
          5572 => x"fe",
          5573 => x"a0",
          5574 => x"16",
          5575 => x"5c",
          5576 => x"8c",
          5577 => x"16",
          5578 => x"7c",
          5579 => x"56",
          5580 => x"f8",
          5581 => x"ff",
          5582 => x"55",
          5583 => x"90",
          5584 => x"52",
          5585 => x"b9",
          5586 => x"fb",
          5587 => x"16",
          5588 => x"17",
          5589 => x"84",
          5590 => x"b9",
          5591 => x"08",
          5592 => x"17",
          5593 => x"33",
          5594 => x"fc",
          5595 => x"a0",
          5596 => x"16",
          5597 => x"56",
          5598 => x"ff",
          5599 => x"81",
          5600 => x"7a",
          5601 => x"54",
          5602 => x"53",
          5603 => x"c6",
          5604 => x"38",
          5605 => x"b4",
          5606 => x"74",
          5607 => x"82",
          5608 => x"81",
          5609 => x"16",
          5610 => x"52",
          5611 => x"3f",
          5612 => x"08",
          5613 => x"91",
          5614 => x"0c",
          5615 => x"1b",
          5616 => x"92",
          5617 => x"58",
          5618 => x"77",
          5619 => x"75",
          5620 => x"86",
          5621 => x"78",
          5622 => x"74",
          5623 => x"90",
          5624 => x"5c",
          5625 => x"7b",
          5626 => x"08",
          5627 => x"5b",
          5628 => x"53",
          5629 => x"ff",
          5630 => x"80",
          5631 => x"78",
          5632 => x"a4",
          5633 => x"5a",
          5634 => x"88",
          5635 => x"5d",
          5636 => x"88",
          5637 => x"17",
          5638 => x"74",
          5639 => x"08",
          5640 => x"5b",
          5641 => x"56",
          5642 => x"59",
          5643 => x"80",
          5644 => x"18",
          5645 => x"80",
          5646 => x"18",
          5647 => x"34",
          5648 => x"b9",
          5649 => x"06",
          5650 => x"84",
          5651 => x"81",
          5652 => x"70",
          5653 => x"93",
          5654 => x"08",
          5655 => x"83",
          5656 => x"08",
          5657 => x"74",
          5658 => x"82",
          5659 => x"81",
          5660 => x"17",
          5661 => x"52",
          5662 => x"3f",
          5663 => x"2a",
          5664 => x"2a",
          5665 => x"08",
          5666 => x"5b",
          5667 => x"56",
          5668 => x"59",
          5669 => x"80",
          5670 => x"18",
          5671 => x"80",
          5672 => x"18",
          5673 => x"34",
          5674 => x"b9",
          5675 => x"06",
          5676 => x"ae",
          5677 => x"a5",
          5678 => x"55",
          5679 => x"56",
          5680 => x"79",
          5681 => x"b9",
          5682 => x"b1",
          5683 => x"38",
          5684 => x"38",
          5685 => x"38",
          5686 => x"52",
          5687 => x"71",
          5688 => x"75",
          5689 => x"3d",
          5690 => x"8f",
          5691 => x"06",
          5692 => x"53",
          5693 => x"7d",
          5694 => x"b2",
          5695 => x"70",
          5696 => x"ac",
          5697 => x"a4",
          5698 => x"71",
          5699 => x"34",
          5700 => x"3d",
          5701 => x"0c",
          5702 => x"11",
          5703 => x"70",
          5704 => x"81",
          5705 => x"76",
          5706 => x"e5",
          5707 => x"57",
          5708 => x"70",
          5709 => x"53",
          5710 => x"e0",
          5711 => x"ff",
          5712 => x"38",
          5713 => x"54",
          5714 => x"71",
          5715 => x"73",
          5716 => x"30",
          5717 => x"59",
          5718 => x"81",
          5719 => x"25",
          5720 => x"39",
          5721 => x"5e",
          5722 => x"80",
          5723 => x"3d",
          5724 => x"08",
          5725 => x"8a",
          5726 => x"3d",
          5727 => x"3d",
          5728 => x"b9",
          5729 => x"80",
          5730 => x"70",
          5731 => x"80",
          5732 => x"84",
          5733 => x"2e",
          5734 => x"9a",
          5735 => x"33",
          5736 => x"2e",
          5737 => x"84",
          5738 => x"84",
          5739 => x"06",
          5740 => x"c8",
          5741 => x"33",
          5742 => x"90",
          5743 => x"5b",
          5744 => x"0c",
          5745 => x"3d",
          5746 => x"e6",
          5747 => x"40",
          5748 => x"3d",
          5749 => x"51",
          5750 => x"59",
          5751 => x"60",
          5752 => x"11",
          5753 => x"db",
          5754 => x"82",
          5755 => x"40",
          5756 => x"aa",
          5757 => x"b9",
          5758 => x"df",
          5759 => x"77",
          5760 => x"83",
          5761 => x"38",
          5762 => x"81",
          5763 => x"84",
          5764 => x"ff",
          5765 => x"78",
          5766 => x"9b",
          5767 => x"2b",
          5768 => x"56",
          5769 => x"76",
          5770 => x"51",
          5771 => x"08",
          5772 => x"38",
          5773 => x"3f",
          5774 => x"c8",
          5775 => x"9b",
          5776 => x"2b",
          5777 => x"5e",
          5778 => x"76",
          5779 => x"08",
          5780 => x"84",
          5781 => x"08",
          5782 => x"2e",
          5783 => x"80",
          5784 => x"51",
          5785 => x"05",
          5786 => x"38",
          5787 => x"70",
          5788 => x"81",
          5789 => x"38",
          5790 => x"82",
          5791 => x"08",
          5792 => x"56",
          5793 => x"38",
          5794 => x"5f",
          5795 => x"08",
          5796 => x"2e",
          5797 => x"a4",
          5798 => x"05",
          5799 => x"5e",
          5800 => x"1a",
          5801 => x"74",
          5802 => x"26",
          5803 => x"94",
          5804 => x"70",
          5805 => x"79",
          5806 => x"81",
          5807 => x"81",
          5808 => x"7c",
          5809 => x"e4",
          5810 => x"17",
          5811 => x"07",
          5812 => x"39",
          5813 => x"98",
          5814 => x"80",
          5815 => x"7a",
          5816 => x"c8",
          5817 => x"2e",
          5818 => x"54",
          5819 => x"53",
          5820 => x"fe",
          5821 => x"fc",
          5822 => x"17",
          5823 => x"31",
          5824 => x"a0",
          5825 => x"16",
          5826 => x"06",
          5827 => x"08",
          5828 => x"81",
          5829 => x"7c",
          5830 => x"e6",
          5831 => x"34",
          5832 => x"10",
          5833 => x"70",
          5834 => x"7a",
          5835 => x"fd",
          5836 => x"81",
          5837 => x"81",
          5838 => x"8e",
          5839 => x"19",
          5840 => x"05",
          5841 => x"fd",
          5842 => x"78",
          5843 => x"0d",
          5844 => x"55",
          5845 => x"74",
          5846 => x"73",
          5847 => x"86",
          5848 => x"78",
          5849 => x"72",
          5850 => x"91",
          5851 => x"8c",
          5852 => x"b9",
          5853 => x"76",
          5854 => x"11",
          5855 => x"73",
          5856 => x"ff",
          5857 => x"b9",
          5858 => x"53",
          5859 => x"b9",
          5860 => x"75",
          5861 => x"77",
          5862 => x"59",
          5863 => x"77",
          5864 => x"94",
          5865 => x"16",
          5866 => x"5a",
          5867 => x"73",
          5868 => x"84",
          5869 => x"08",
          5870 => x"2e",
          5871 => x"38",
          5872 => x"82",
          5873 => x"ae",
          5874 => x"53",
          5875 => x"0d",
          5876 => x"81",
          5877 => x"75",
          5878 => x"76",
          5879 => x"38",
          5880 => x"54",
          5881 => x"16",
          5882 => x"57",
          5883 => x"06",
          5884 => x"15",
          5885 => x"16",
          5886 => x"8b",
          5887 => x"0c",
          5888 => x"80",
          5889 => x"80",
          5890 => x"84",
          5891 => x"17",
          5892 => x"56",
          5893 => x"15",
          5894 => x"56",
          5895 => x"16",
          5896 => x"05",
          5897 => x"78",
          5898 => x"08",
          5899 => x"51",
          5900 => x"08",
          5901 => x"51",
          5902 => x"08",
          5903 => x"72",
          5904 => x"73",
          5905 => x"84",
          5906 => x"08",
          5907 => x"08",
          5908 => x"c8",
          5909 => x"0c",
          5910 => x"34",
          5911 => x"3d",
          5912 => x"89",
          5913 => x"53",
          5914 => x"84",
          5915 => x"c8",
          5916 => x"2e",
          5917 => x"73",
          5918 => x"04",
          5919 => x"ff",
          5920 => x"55",
          5921 => x"ab",
          5922 => x"80",
          5923 => x"70",
          5924 => x"80",
          5925 => x"9b",
          5926 => x"2b",
          5927 => x"55",
          5928 => x"88",
          5929 => x"84",
          5930 => x"99",
          5931 => x"74",
          5932 => x"ff",
          5933 => x"39",
          5934 => x"39",
          5935 => x"98",
          5936 => x"88",
          5937 => x"fa",
          5938 => x"80",
          5939 => x"80",
          5940 => x"80",
          5941 => x"16",
          5942 => x"38",
          5943 => x"73",
          5944 => x"88",
          5945 => x"fe",
          5946 => x"81",
          5947 => x"08",
          5948 => x"7a",
          5949 => x"2e",
          5950 => x"2e",
          5951 => x"2e",
          5952 => x"22",
          5953 => x"38",
          5954 => x"80",
          5955 => x"38",
          5956 => x"3f",
          5957 => x"c8",
          5958 => x"c8",
          5959 => x"ff",
          5960 => x"ff",
          5961 => x"84",
          5962 => x"2c",
          5963 => x"54",
          5964 => x"0d",
          5965 => x"ff",
          5966 => x"ff",
          5967 => x"84",
          5968 => x"2c",
          5969 => x"54",
          5970 => x"96",
          5971 => x"b9",
          5972 => x"14",
          5973 => x"b9",
          5974 => x"d8",
          5975 => x"d2",
          5976 => x"53",
          5977 => x"56",
          5978 => x"55",
          5979 => x"38",
          5980 => x"0d",
          5981 => x"a9",
          5982 => x"b9",
          5983 => x"05",
          5984 => x"74",
          5985 => x"38",
          5986 => x"3f",
          5987 => x"0d",
          5988 => x"95",
          5989 => x"68",
          5990 => x"05",
          5991 => x"84",
          5992 => x"08",
          5993 => x"9c",
          5994 => x"59",
          5995 => x"38",
          5996 => x"0c",
          5997 => x"08",
          5998 => x"82",
          5999 => x"b9",
          6000 => x"c1",
          6001 => x"56",
          6002 => x"38",
          6003 => x"81",
          6004 => x"17",
          6005 => x"b7",
          6006 => x"85",
          6007 => x"18",
          6008 => x"cc",
          6009 => x"82",
          6010 => x"11",
          6011 => x"71",
          6012 => x"72",
          6013 => x"ff",
          6014 => x"70",
          6015 => x"83",
          6016 => x"43",
          6017 => x"56",
          6018 => x"7a",
          6019 => x"07",
          6020 => x"b9",
          6021 => x"54",
          6022 => x"53",
          6023 => x"a6",
          6024 => x"fe",
          6025 => x"18",
          6026 => x"31",
          6027 => x"a0",
          6028 => x"17",
          6029 => x"06",
          6030 => x"08",
          6031 => x"81",
          6032 => x"77",
          6033 => x"92",
          6034 => x"ff",
          6035 => x"ff",
          6036 => x"08",
          6037 => x"c8",
          6038 => x"07",
          6039 => x"5a",
          6040 => x"26",
          6041 => x"18",
          6042 => x"77",
          6043 => x"17",
          6044 => x"71",
          6045 => x"25",
          6046 => x"1f",
          6047 => x"78",
          6048 => x"5a",
          6049 => x"7a",
          6050 => x"17",
          6051 => x"34",
          6052 => x"e7",
          6053 => x"56",
          6054 => x"55",
          6055 => x"54",
          6056 => x"22",
          6057 => x"2e",
          6058 => x"75",
          6059 => x"75",
          6060 => x"81",
          6061 => x"73",
          6062 => x"08",
          6063 => x"38",
          6064 => x"77",
          6065 => x"38",
          6066 => x"82",
          6067 => x"17",
          6068 => x"07",
          6069 => x"2e",
          6070 => x"55",
          6071 => x"0d",
          6072 => x"ff",
          6073 => x"ca",
          6074 => x"b9",
          6075 => x"84",
          6076 => x"38",
          6077 => x"e5",
          6078 => x"ff",
          6079 => x"82",
          6080 => x"94",
          6081 => x"27",
          6082 => x"0c",
          6083 => x"84",
          6084 => x"ff",
          6085 => x"51",
          6086 => x"08",
          6087 => x"73",
          6088 => x"80",
          6089 => x"56",
          6090 => x"39",
          6091 => x"fd",
          6092 => x"2e",
          6093 => x"81",
          6094 => x"38",
          6095 => x"19",
          6096 => x"c8",
          6097 => x"56",
          6098 => x"27",
          6099 => x"9c",
          6100 => x"80",
          6101 => x"75",
          6102 => x"c8",
          6103 => x"e3",
          6104 => x"d2",
          6105 => x"b9",
          6106 => x"84",
          6107 => x"38",
          6108 => x"fe",
          6109 => x"ff",
          6110 => x"80",
          6111 => x"94",
          6112 => x"27",
          6113 => x"84",
          6114 => x"17",
          6115 => x"a1",
          6116 => x"33",
          6117 => x"bb",
          6118 => x"56",
          6119 => x"82",
          6120 => x"86",
          6121 => x"33",
          6122 => x"90",
          6123 => x"84",
          6124 => x"56",
          6125 => x"53",
          6126 => x"3d",
          6127 => x"c8",
          6128 => x"2e",
          6129 => x"a7",
          6130 => x"08",
          6131 => x"ab",
          6132 => x"84",
          6133 => x"93",
          6134 => x"59",
          6135 => x"98",
          6136 => x"02",
          6137 => x"5d",
          6138 => x"7d",
          6139 => x"12",
          6140 => x"41",
          6141 => x"80",
          6142 => x"57",
          6143 => x"56",
          6144 => x"38",
          6145 => x"08",
          6146 => x"8b",
          6147 => x"84",
          6148 => x"b9",
          6149 => x"b4",
          6150 => x"b9",
          6151 => x"b9",
          6152 => x"16",
          6153 => x"71",
          6154 => x"5d",
          6155 => x"84",
          6156 => x"fe",
          6157 => x"08",
          6158 => x"d3",
          6159 => x"92",
          6160 => x"b9",
          6161 => x"30",
          6162 => x"7a",
          6163 => x"95",
          6164 => x"7b",
          6165 => x"26",
          6166 => x"d2",
          6167 => x"84",
          6168 => x"a7",
          6169 => x"19",
          6170 => x"76",
          6171 => x"7a",
          6172 => x"06",
          6173 => x"b8",
          6174 => x"f1",
          6175 => x"2e",
          6176 => x"b4",
          6177 => x"9c",
          6178 => x"0b",
          6179 => x"27",
          6180 => x"ff",
          6181 => x"56",
          6182 => x"96",
          6183 => x"fe",
          6184 => x"81",
          6185 => x"81",
          6186 => x"81",
          6187 => x"09",
          6188 => x"c8",
          6189 => x"a8",
          6190 => x"59",
          6191 => x"eb",
          6192 => x"2e",
          6193 => x"54",
          6194 => x"53",
          6195 => x"f1",
          6196 => x"79",
          6197 => x"74",
          6198 => x"84",
          6199 => x"08",
          6200 => x"c8",
          6201 => x"b9",
          6202 => x"80",
          6203 => x"9b",
          6204 => x"9c",
          6205 => x"58",
          6206 => x"38",
          6207 => x"33",
          6208 => x"79",
          6209 => x"80",
          6210 => x"f7",
          6211 => x"95",
          6212 => x"3d",
          6213 => x"05",
          6214 => x"3f",
          6215 => x"c8",
          6216 => x"b9",
          6217 => x"43",
          6218 => x"ff",
          6219 => x"56",
          6220 => x"0b",
          6221 => x"04",
          6222 => x"81",
          6223 => x"33",
          6224 => x"86",
          6225 => x"74",
          6226 => x"83",
          6227 => x"57",
          6228 => x"87",
          6229 => x"80",
          6230 => x"2e",
          6231 => x"7d",
          6232 => x"5d",
          6233 => x"19",
          6234 => x"80",
          6235 => x"17",
          6236 => x"05",
          6237 => x"17",
          6238 => x"76",
          6239 => x"55",
          6240 => x"22",
          6241 => x"81",
          6242 => x"17",
          6243 => x"b9",
          6244 => x"58",
          6245 => x"81",
          6246 => x"70",
          6247 => x"ee",
          6248 => x"08",
          6249 => x"18",
          6250 => x"31",
          6251 => x"ee",
          6252 => x"2e",
          6253 => x"54",
          6254 => x"53",
          6255 => x"ed",
          6256 => x"7b",
          6257 => x"fd",
          6258 => x"fd",
          6259 => x"f2",
          6260 => x"84",
          6261 => x"38",
          6262 => x"8d",
          6263 => x"fd",
          6264 => x"51",
          6265 => x"08",
          6266 => x"11",
          6267 => x"7b",
          6268 => x"0c",
          6269 => x"84",
          6270 => x"ff",
          6271 => x"9f",
          6272 => x"74",
          6273 => x"76",
          6274 => x"38",
          6275 => x"75",
          6276 => x"56",
          6277 => x"b8",
          6278 => x"c3",
          6279 => x"1a",
          6280 => x"0b",
          6281 => x"80",
          6282 => x"ff",
          6283 => x"34",
          6284 => x"17",
          6285 => x"81",
          6286 => x"d8",
          6287 => x"70",
          6288 => x"05",
          6289 => x"38",
          6290 => x"34",
          6291 => x"5b",
          6292 => x"78",
          6293 => x"34",
          6294 => x"f0",
          6295 => x"34",
          6296 => x"b9",
          6297 => x"fd",
          6298 => x"08",
          6299 => x"97",
          6300 => x"80",
          6301 => x"58",
          6302 => x"2a",
          6303 => x"5a",
          6304 => x"55",
          6305 => x"81",
          6306 => x"ed",
          6307 => x"75",
          6308 => x"04",
          6309 => x"17",
          6310 => x"ed",
          6311 => x"2a",
          6312 => x"88",
          6313 => x"7d",
          6314 => x"1b",
          6315 => x"90",
          6316 => x"88",
          6317 => x"55",
          6318 => x"81",
          6319 => x"ec",
          6320 => x"ff",
          6321 => x"b4",
          6322 => x"80",
          6323 => x"5b",
          6324 => x"ba",
          6325 => x"75",
          6326 => x"b1",
          6327 => x"51",
          6328 => x"08",
          6329 => x"8a",
          6330 => x"3d",
          6331 => x"3d",
          6332 => x"ff",
          6333 => x"56",
          6334 => x"81",
          6335 => x"86",
          6336 => x"3d",
          6337 => x"70",
          6338 => x"05",
          6339 => x"38",
          6340 => x"58",
          6341 => x"77",
          6342 => x"55",
          6343 => x"77",
          6344 => x"c8",
          6345 => x"d8",
          6346 => x"cb",
          6347 => x"b1",
          6348 => x"70",
          6349 => x"89",
          6350 => x"ff",
          6351 => x"2e",
          6352 => x"e5",
          6353 => x"5f",
          6354 => x"79",
          6355 => x"12",
          6356 => x"38",
          6357 => x"55",
          6358 => x"89",
          6359 => x"58",
          6360 => x"55",
          6361 => x"38",
          6362 => x"70",
          6363 => x"07",
          6364 => x"38",
          6365 => x"83",
          6366 => x"5a",
          6367 => x"fd",
          6368 => x"b1",
          6369 => x"51",
          6370 => x"08",
          6371 => x"38",
          6372 => x"2e",
          6373 => x"51",
          6374 => x"08",
          6375 => x"38",
          6376 => x"88",
          6377 => x"75",
          6378 => x"81",
          6379 => x"ef",
          6380 => x"19",
          6381 => x"81",
          6382 => x"a0",
          6383 => x"5d",
          6384 => x"33",
          6385 => x"75",
          6386 => x"08",
          6387 => x"19",
          6388 => x"07",
          6389 => x"83",
          6390 => x"18",
          6391 => x"27",
          6392 => x"71",
          6393 => x"75",
          6394 => x"5d",
          6395 => x"38",
          6396 => x"38",
          6397 => x"81",
          6398 => x"84",
          6399 => x"ff",
          6400 => x"7f",
          6401 => x"7b",
          6402 => x"79",
          6403 => x"6a",
          6404 => x"7b",
          6405 => x"58",
          6406 => x"5b",
          6407 => x"38",
          6408 => x"18",
          6409 => x"ed",
          6410 => x"18",
          6411 => x"3d",
          6412 => x"95",
          6413 => x"a2",
          6414 => x"b9",
          6415 => x"5c",
          6416 => x"16",
          6417 => x"33",
          6418 => x"81",
          6419 => x"53",
          6420 => x"fe",
          6421 => x"80",
          6422 => x"76",
          6423 => x"38",
          6424 => x"81",
          6425 => x"7b",
          6426 => x"fe",
          6427 => x"55",
          6428 => x"98",
          6429 => x"e1",
          6430 => x"7f",
          6431 => x"c8",
          6432 => x"0d",
          6433 => x"b1",
          6434 => x"19",
          6435 => x"07",
          6436 => x"39",
          6437 => x"fe",
          6438 => x"fe",
          6439 => x"b1",
          6440 => x"08",
          6441 => x"fe",
          6442 => x"c8",
          6443 => x"db",
          6444 => x"34",
          6445 => x"84",
          6446 => x"17",
          6447 => x"33",
          6448 => x"fe",
          6449 => x"a0",
          6450 => x"16",
          6451 => x"58",
          6452 => x"08",
          6453 => x"33",
          6454 => x"5c",
          6455 => x"84",
          6456 => x"17",
          6457 => x"c8",
          6458 => x"27",
          6459 => x"7c",
          6460 => x"38",
          6461 => x"08",
          6462 => x"51",
          6463 => x"e8",
          6464 => x"05",
          6465 => x"33",
          6466 => x"05",
          6467 => x"3f",
          6468 => x"c8",
          6469 => x"b9",
          6470 => x"5a",
          6471 => x"ff",
          6472 => x"56",
          6473 => x"80",
          6474 => x"86",
          6475 => x"61",
          6476 => x"7a",
          6477 => x"73",
          6478 => x"83",
          6479 => x"3f",
          6480 => x"0c",
          6481 => x"67",
          6482 => x"52",
          6483 => x"84",
          6484 => x"08",
          6485 => x"c8",
          6486 => x"66",
          6487 => x"95",
          6488 => x"84",
          6489 => x"cf",
          6490 => x"55",
          6491 => x"86",
          6492 => x"59",
          6493 => x"2a",
          6494 => x"2a",
          6495 => x"2a",
          6496 => x"81",
          6497 => x"e1",
          6498 => x"b9",
          6499 => x"3d",
          6500 => x"9a",
          6501 => x"ff",
          6502 => x"84",
          6503 => x"c8",
          6504 => x"7a",
          6505 => x"06",
          6506 => x"30",
          6507 => x"7b",
          6508 => x"76",
          6509 => x"80",
          6510 => x"80",
          6511 => x"f6",
          6512 => x"74",
          6513 => x"38",
          6514 => x"81",
          6515 => x"84",
          6516 => x"ff",
          6517 => x"78",
          6518 => x"56",
          6519 => x"8b",
          6520 => x"83",
          6521 => x"83",
          6522 => x"2b",
          6523 => x"70",
          6524 => x"07",
          6525 => x"56",
          6526 => x"0d",
          6527 => x"8e",
          6528 => x"3f",
          6529 => x"c8",
          6530 => x"84",
          6531 => x"80",
          6532 => x"77",
          6533 => x"70",
          6534 => x"dc",
          6535 => x"08",
          6536 => x"38",
          6537 => x"b4",
          6538 => x"b9",
          6539 => x"08",
          6540 => x"55",
          6541 => x"a0",
          6542 => x"17",
          6543 => x"33",
          6544 => x"81",
          6545 => x"16",
          6546 => x"b9",
          6547 => x"fe",
          6548 => x"f8",
          6549 => x"84",
          6550 => x"b9",
          6551 => x"5c",
          6552 => x"1b",
          6553 => x"81",
          6554 => x"8b",
          6555 => x"77",
          6556 => x"7b",
          6557 => x"a0",
          6558 => x"57",
          6559 => x"53",
          6560 => x"3d",
          6561 => x"c8",
          6562 => x"a6",
          6563 => x"55",
          6564 => x"ff",
          6565 => x"3d",
          6566 => x"5b",
          6567 => x"b7",
          6568 => x"75",
          6569 => x"74",
          6570 => x"83",
          6571 => x"51",
          6572 => x"b9",
          6573 => x"b9",
          6574 => x"76",
          6575 => x"d8",
          6576 => x"ff",
          6577 => x"81",
          6578 => x"99",
          6579 => x"ff",
          6580 => x"89",
          6581 => x"e9",
          6582 => x"81",
          6583 => x"f8",
          6584 => x"81",
          6585 => x"2a",
          6586 => x"34",
          6587 => x"05",
          6588 => x"70",
          6589 => x"58",
          6590 => x"8f",
          6591 => x"e5",
          6592 => x"38",
          6593 => x"33",
          6594 => x"06",
          6595 => x"38",
          6596 => x"3d",
          6597 => x"84",
          6598 => x"08",
          6599 => x"84",
          6600 => x"83",
          6601 => x"84",
          6602 => x"55",
          6603 => x"84",
          6604 => x"83",
          6605 => x"81",
          6606 => x"84",
          6607 => x"08",
          6608 => x"c4",
          6609 => x"76",
          6610 => x"81",
          6611 => x"ef",
          6612 => x"34",
          6613 => x"b9",
          6614 => x"39",
          6615 => x"56",
          6616 => x"84",
          6617 => x"80",
          6618 => x"75",
          6619 => x"ee",
          6620 => x"84",
          6621 => x"06",
          6622 => x"b8",
          6623 => x"80",
          6624 => x"38",
          6625 => x"09",
          6626 => x"76",
          6627 => x"51",
          6628 => x"08",
          6629 => x"59",
          6630 => x"be",
          6631 => x"57",
          6632 => x"9e",
          6633 => x"07",
          6634 => x"38",
          6635 => x"38",
          6636 => x"3f",
          6637 => x"c8",
          6638 => x"55",
          6639 => x"55",
          6640 => x"55",
          6641 => x"ff",
          6642 => x"88",
          6643 => x"59",
          6644 => x"33",
          6645 => x"15",
          6646 => x"76",
          6647 => x"81",
          6648 => x"da",
          6649 => x"7a",
          6650 => x"34",
          6651 => x"b9",
          6652 => x"57",
          6653 => x"08",
          6654 => x"fe",
          6655 => x"79",
          6656 => x"84",
          6657 => x"18",
          6658 => x"a0",
          6659 => x"33",
          6660 => x"b9",
          6661 => x"5a",
          6662 => x"3f",
          6663 => x"c8",
          6664 => x"ae",
          6665 => x"2e",
          6666 => x"54",
          6667 => x"53",
          6668 => x"d3",
          6669 => x"0d",
          6670 => x"05",
          6671 => x"80",
          6672 => x"80",
          6673 => x"80",
          6674 => x"18",
          6675 => x"c2",
          6676 => x"a5",
          6677 => x"9d",
          6678 => x"8c",
          6679 => x"33",
          6680 => x"74",
          6681 => x"11",
          6682 => x"54",
          6683 => x"ff",
          6684 => x"07",
          6685 => x"90",
          6686 => x"58",
          6687 => x"08",
          6688 => x"78",
          6689 => x"51",
          6690 => x"55",
          6691 => x"38",
          6692 => x"2e",
          6693 => x"ff",
          6694 => x"08",
          6695 => x"7d",
          6696 => x"81",
          6697 => x"73",
          6698 => x"04",
          6699 => x"3d",
          6700 => x"d0",
          6701 => x"06",
          6702 => x"08",
          6703 => x"2e",
          6704 => x"7c",
          6705 => x"74",
          6706 => x"77",
          6707 => x"84",
          6708 => x"08",
          6709 => x"17",
          6710 => x"7e",
          6711 => x"ff",
          6712 => x"8c",
          6713 => x"07",
          6714 => x"08",
          6715 => x"76",
          6716 => x"31",
          6717 => x"07",
          6718 => x"fe",
          6719 => x"74",
          6720 => x"54",
          6721 => x"39",
          6722 => x"b9",
          6723 => x"08",
          6724 => x"87",
          6725 => x"a2",
          6726 => x"80",
          6727 => x"05",
          6728 => x"75",
          6729 => x"38",
          6730 => x"d1",
          6731 => x"e5",
          6732 => x"05",
          6733 => x"84",
          6734 => x"b9",
          6735 => x"33",
          6736 => x"fe",
          6737 => x"81",
          6738 => x"83",
          6739 => x"2a",
          6740 => x"9f",
          6741 => x"52",
          6742 => x"b9",
          6743 => x"74",
          6744 => x"80",
          6745 => x"75",
          6746 => x"80",
          6747 => x"83",
          6748 => x"83",
          6749 => x"74",
          6750 => x"3d",
          6751 => x"59",
          6752 => x"ab",
          6753 => x"07",
          6754 => x"38",
          6755 => x"54",
          6756 => x"cd",
          6757 => x"08",
          6758 => x"33",
          6759 => x"2b",
          6760 => x"d4",
          6761 => x"38",
          6762 => x"11",
          6763 => x"e7",
          6764 => x"82",
          6765 => x"2b",
          6766 => x"88",
          6767 => x"1f",
          6768 => x"90",
          6769 => x"33",
          6770 => x"71",
          6771 => x"3d",
          6772 => x"45",
          6773 => x"8e",
          6774 => x"38",
          6775 => x"87",
          6776 => x"45",
          6777 => x"61",
          6778 => x"38",
          6779 => x"38",
          6780 => x"7a",
          6781 => x"7a",
          6782 => x"0b",
          6783 => x"80",
          6784 => x"38",
          6785 => x"17",
          6786 => x"2e",
          6787 => x"77",
          6788 => x"84",
          6789 => x"84",
          6790 => x"38",
          6791 => x"84",
          6792 => x"2a",
          6793 => x"15",
          6794 => x"7b",
          6795 => x"ff",
          6796 => x"4e",
          6797 => x"38",
          6798 => x"70",
          6799 => x"82",
          6800 => x"78",
          6801 => x"80",
          6802 => x"62",
          6803 => x"2e",
          6804 => x"ff",
          6805 => x"82",
          6806 => x"18",
          6807 => x"38",
          6808 => x"76",
          6809 => x"84",
          6810 => x"fe",
          6811 => x"9f",
          6812 => x"7c",
          6813 => x"57",
          6814 => x"82",
          6815 => x"5d",
          6816 => x"80",
          6817 => x"08",
          6818 => x"5c",
          6819 => x"ff",
          6820 => x"26",
          6821 => x"06",
          6822 => x"99",
          6823 => x"ff",
          6824 => x"2a",
          6825 => x"06",
          6826 => x"7a",
          6827 => x"2a",
          6828 => x"2e",
          6829 => x"5f",
          6830 => x"7f",
          6831 => x"05",
          6832 => x"dd",
          6833 => x"fe",
          6834 => x"84",
          6835 => x"38",
          6836 => x"75",
          6837 => x"59",
          6838 => x"39",
          6839 => x"7a",
          6840 => x"61",
          6841 => x"2e",
          6842 => x"4a",
          6843 => x"c8",
          6844 => x"8b",
          6845 => x"27",
          6846 => x"b9",
          6847 => x"d4",
          6848 => x"86",
          6849 => x"38",
          6850 => x"fd",
          6851 => x"80",
          6852 => x"15",
          6853 => x"e5",
          6854 => x"05",
          6855 => x"34",
          6856 => x"8b",
          6857 => x"8c",
          6858 => x"7b",
          6859 => x"8e",
          6860 => x"61",
          6861 => x"34",
          6862 => x"80",
          6863 => x"82",
          6864 => x"6c",
          6865 => x"ad",
          6866 => x"74",
          6867 => x"4c",
          6868 => x"95",
          6869 => x"80",
          6870 => x"05",
          6871 => x"61",
          6872 => x"67",
          6873 => x"4c",
          6874 => x"2a",
          6875 => x"08",
          6876 => x"85",
          6877 => x"80",
          6878 => x"05",
          6879 => x"7c",
          6880 => x"96",
          6881 => x"61",
          6882 => x"05",
          6883 => x"61",
          6884 => x"55",
          6885 => x"70",
          6886 => x"74",
          6887 => x"80",
          6888 => x"4b",
          6889 => x"53",
          6890 => x"3f",
          6891 => x"e7",
          6892 => x"87",
          6893 => x"76",
          6894 => x"55",
          6895 => x"62",
          6896 => x"ff",
          6897 => x"f8",
          6898 => x"7c",
          6899 => x"46",
          6900 => x"70",
          6901 => x"56",
          6902 => x"76",
          6903 => x"54",
          6904 => x"c5",
          6905 => x"e6",
          6906 => x"76",
          6907 => x"55",
          6908 => x"31",
          6909 => x"05",
          6910 => x"77",
          6911 => x"56",
          6912 => x"75",
          6913 => x"79",
          6914 => x"c8",
          6915 => x"76",
          6916 => x"58",
          6917 => x"6c",
          6918 => x"58",
          6919 => x"7d",
          6920 => x"06",
          6921 => x"61",
          6922 => x"57",
          6923 => x"80",
          6924 => x"60",
          6925 => x"81",
          6926 => x"05",
          6927 => x"67",
          6928 => x"c1",
          6929 => x"3f",
          6930 => x"c8",
          6931 => x"67",
          6932 => x"67",
          6933 => x"05",
          6934 => x"6b",
          6935 => x"d4",
          6936 => x"61",
          6937 => x"45",
          6938 => x"90",
          6939 => x"34",
          6940 => x"cd",
          6941 => x"52",
          6942 => x"57",
          6943 => x"80",
          6944 => x"dd",
          6945 => x"f7",
          6946 => x"b9",
          6947 => x"d4",
          6948 => x"74",
          6949 => x"39",
          6950 => x"81",
          6951 => x"74",
          6952 => x"98",
          6953 => x"82",
          6954 => x"80",
          6955 => x"38",
          6956 => x"3f",
          6957 => x"87",
          6958 => x"5c",
          6959 => x"80",
          6960 => x"0a",
          6961 => x"f8",
          6962 => x"ff",
          6963 => x"d3",
          6964 => x"bf",
          6965 => x"81",
          6966 => x"38",
          6967 => x"a0",
          6968 => x"61",
          6969 => x"7a",
          6970 => x"57",
          6971 => x"39",
          6972 => x"61",
          6973 => x"c5",
          6974 => x"05",
          6975 => x"88",
          6976 => x"7c",
          6977 => x"34",
          6978 => x"05",
          6979 => x"61",
          6980 => x"34",
          6981 => x"b0",
          6982 => x"86",
          6983 => x"05",
          6984 => x"34",
          6985 => x"61",
          6986 => x"57",
          6987 => x"76",
          6988 => x"55",
          6989 => x"70",
          6990 => x"05",
          6991 => x"38",
          6992 => x"60",
          6993 => x"81",
          6994 => x"38",
          6995 => x"62",
          6996 => x"b9",
          6997 => x"fe",
          6998 => x"0b",
          6999 => x"84",
          7000 => x"7b",
          7001 => x"34",
          7002 => x"ff",
          7003 => x"ff",
          7004 => x"05",
          7005 => x"61",
          7006 => x"34",
          7007 => x"34",
          7008 => x"86",
          7009 => x"be",
          7010 => x"80",
          7011 => x"17",
          7012 => x"d2",
          7013 => x"55",
          7014 => x"34",
          7015 => x"34",
          7016 => x"83",
          7017 => x"e5",
          7018 => x"05",
          7019 => x"34",
          7020 => x"e8",
          7021 => x"61",
          7022 => x"56",
          7023 => x"98",
          7024 => x"34",
          7025 => x"61",
          7026 => x"ee",
          7027 => x"34",
          7028 => x"34",
          7029 => x"79",
          7030 => x"81",
          7031 => x"bd",
          7032 => x"a6",
          7033 => x"5b",
          7034 => x"57",
          7035 => x"59",
          7036 => x"78",
          7037 => x"7b",
          7038 => x"8d",
          7039 => x"38",
          7040 => x"81",
          7041 => x"77",
          7042 => x"7a",
          7043 => x"84",
          7044 => x"f7",
          7045 => x"05",
          7046 => x"d5",
          7047 => x"24",
          7048 => x"8c",
          7049 => x"16",
          7050 => x"84",
          7051 => x"8b",
          7052 => x"54",
          7053 => x"51",
          7054 => x"70",
          7055 => x"30",
          7056 => x"0c",
          7057 => x"76",
          7058 => x"e3",
          7059 => x"8d",
          7060 => x"55",
          7061 => x"ff",
          7062 => x"08",
          7063 => x"38",
          7064 => x"38",
          7065 => x"77",
          7066 => x"24",
          7067 => x"19",
          7068 => x"24",
          7069 => x"55",
          7070 => x"51",
          7071 => x"08",
          7072 => x"ff",
          7073 => x"0d",
          7074 => x"75",
          7075 => x"ff",
          7076 => x"30",
          7077 => x"52",
          7078 => x"52",
          7079 => x"39",
          7080 => x"0d",
          7081 => x"05",
          7082 => x"72",
          7083 => x"ff",
          7084 => x"0c",
          7085 => x"73",
          7086 => x"81",
          7087 => x"38",
          7088 => x"2e",
          7089 => x"ff",
          7090 => x"8d",
          7091 => x"70",
          7092 => x"12",
          7093 => x"0c",
          7094 => x"0d",
          7095 => x"96",
          7096 => x"80",
          7097 => x"84",
          7098 => x"71",
          7099 => x"38",
          7100 => x"10",
          7101 => x"b9",
          7102 => x"fb",
          7103 => x"ff",
          7104 => x"ff",
          7105 => x"9f",
          7106 => x"82",
          7107 => x"80",
          7108 => x"53",
          7109 => x"05",
          7110 => x"56",
          7111 => x"70",
          7112 => x"73",
          7113 => x"22",
          7114 => x"79",
          7115 => x"2e",
          7116 => x"c8",
          7117 => x"80",
          7118 => x"ea",
          7119 => x"05",
          7120 => x"70",
          7121 => x"51",
          7122 => x"ff",
          7123 => x"16",
          7124 => x"e6",
          7125 => x"06",
          7126 => x"83",
          7127 => x"e0",
          7128 => x"51",
          7129 => x"ff",
          7130 => x"73",
          7131 => x"83",
          7132 => x"a6",
          7133 => x"70",
          7134 => x"00",
          7135 => x"ff",
          7136 => x"00",
          7137 => x"80",
          7138 => x"6a",
          7139 => x"54",
          7140 => x"3e",
          7141 => x"28",
          7142 => x"12",
          7143 => x"fc",
          7144 => x"e6",
          7145 => x"d0",
          7146 => x"ba",
          7147 => x"59",
          7148 => x"59",
          7149 => x"59",
          7150 => x"59",
          7151 => x"59",
          7152 => x"59",
          7153 => x"59",
          7154 => x"59",
          7155 => x"59",
          7156 => x"59",
          7157 => x"59",
          7158 => x"59",
          7159 => x"59",
          7160 => x"59",
          7161 => x"59",
          7162 => x"59",
          7163 => x"59",
          7164 => x"59",
          7165 => x"59",
          7166 => x"59",
          7167 => x"59",
          7168 => x"71",
          7169 => x"59",
          7170 => x"59",
          7171 => x"59",
          7172 => x"59",
          7173 => x"59",
          7174 => x"59",
          7175 => x"59",
          7176 => x"59",
          7177 => x"06",
          7178 => x"8a",
          7179 => x"67",
          7180 => x"ce",
          7181 => x"59",
          7182 => x"59",
          7183 => x"59",
          7184 => x"59",
          7185 => x"59",
          7186 => x"59",
          7187 => x"59",
          7188 => x"59",
          7189 => x"59",
          7190 => x"59",
          7191 => x"59",
          7192 => x"59",
          7193 => x"59",
          7194 => x"59",
          7195 => x"59",
          7196 => x"59",
          7197 => x"59",
          7198 => x"59",
          7199 => x"59",
          7200 => x"59",
          7201 => x"59",
          7202 => x"59",
          7203 => x"59",
          7204 => x"59",
          7205 => x"59",
          7206 => x"59",
          7207 => x"70",
          7208 => x"59",
          7209 => x"59",
          7210 => x"59",
          7211 => x"59",
          7212 => x"58",
          7213 => x"41",
          7214 => x"51",
          7215 => x"3a",
          7216 => x"3a",
          7217 => x"52",
          7218 => x"2e",
          7219 => x"85",
          7220 => x"4f",
          7221 => x"de",
          7222 => x"74",
          7223 => x"a3",
          7224 => x"2a",
          7225 => x"01",
          7226 => x"9b",
          7227 => x"de",
          7228 => x"a3",
          7229 => x"4f",
          7230 => x"95",
          7231 => x"db",
          7232 => x"00",
          7233 => x"a5",
          7234 => x"62",
          7235 => x"62",
          7236 => x"62",
          7237 => x"62",
          7238 => x"62",
          7239 => x"62",
          7240 => x"62",
          7241 => x"62",
          7242 => x"62",
          7243 => x"62",
          7244 => x"62",
          7245 => x"62",
          7246 => x"62",
          7247 => x"62",
          7248 => x"7a",
          7249 => x"55",
          7250 => x"6c",
          7251 => x"1d",
          7252 => x"62",
          7253 => x"0d",
          7254 => x"b6",
          7255 => x"fb",
          7256 => x"d7",
          7257 => x"62",
          7258 => x"08",
          7259 => x"49",
          7260 => x"7d",
          7261 => x"32",
          7262 => x"89",
          7263 => x"cb",
          7264 => x"89",
          7265 => x"89",
          7266 => x"89",
          7267 => x"b3",
          7268 => x"89",
          7269 => x"89",
          7270 => x"89",
          7271 => x"89",
          7272 => x"89",
          7273 => x"89",
          7274 => x"89",
          7275 => x"89",
          7276 => x"89",
          7277 => x"89",
          7278 => x"89",
          7279 => x"89",
          7280 => x"d9",
          7281 => x"89",
          7282 => x"89",
          7283 => x"60",
          7284 => x"43",
          7285 => x"21",
          7286 => x"21",
          7287 => x"21",
          7288 => x"fc",
          7289 => x"21",
          7290 => x"21",
          7291 => x"21",
          7292 => x"21",
          7293 => x"21",
          7294 => x"21",
          7295 => x"21",
          7296 => x"21",
          7297 => x"21",
          7298 => x"21",
          7299 => x"21",
          7300 => x"06",
          7301 => x"e0",
          7302 => x"91",
          7303 => x"6e",
          7304 => x"5e",
          7305 => x"3c",
          7306 => x"18",
          7307 => x"78",
          7308 => x"50",
          7309 => x"9a",
          7310 => x"d7",
          7311 => x"d7",
          7312 => x"d7",
          7313 => x"d7",
          7314 => x"d7",
          7315 => x"d7",
          7316 => x"d7",
          7317 => x"d7",
          7318 => x"d7",
          7319 => x"d7",
          7320 => x"c5",
          7321 => x"d7",
          7322 => x"d7",
          7323 => x"d8",
          7324 => x"e5",
          7325 => x"c6",
          7326 => x"b0",
          7327 => x"9a",
          7328 => x"80",
          7329 => x"fd",
          7330 => x"49",
          7331 => x"fd",
          7332 => x"fd",
          7333 => x"fd",
          7334 => x"fd",
          7335 => x"7f",
          7336 => x"fd",
          7337 => x"fd",
          7338 => x"fd",
          7339 => x"fd",
          7340 => x"fd",
          7341 => x"fd",
          7342 => x"fd",
          7343 => x"fd",
          7344 => x"fd",
          7345 => x"fd",
          7346 => x"fd",
          7347 => x"fd",
          7348 => x"fd",
          7349 => x"fd",
          7350 => x"fd",
          7351 => x"fd",
          7352 => x"fd",
          7353 => x"fd",
          7354 => x"1d",
          7355 => x"fd",
          7356 => x"fd",
          7357 => x"fd",
          7358 => x"fd",
          7359 => x"fd",
          7360 => x"fd",
          7361 => x"fd",
          7362 => x"2b",
          7363 => x"b8",
          7364 => x"b8",
          7365 => x"e1",
          7366 => x"fd",
          7367 => x"fd",
          7368 => x"16",
          7369 => x"fd",
          7370 => x"58",
          7371 => x"18",
          7372 => x"fd",
          7373 => x"69",
          7374 => x"63",
          7375 => x"69",
          7376 => x"61",
          7377 => x"65",
          7378 => x"65",
          7379 => x"70",
          7380 => x"66",
          7381 => x"6d",
          7382 => x"00",
          7383 => x"00",
          7384 => x"00",
          7385 => x"00",
          7386 => x"00",
          7387 => x"74",
          7388 => x"65",
          7389 => x"6f",
          7390 => x"74",
          7391 => x"00",
          7392 => x"73",
          7393 => x"73",
          7394 => x"6f",
          7395 => x"00",
          7396 => x"20",
          7397 => x"00",
          7398 => x"65",
          7399 => x"72",
          7400 => x"00",
          7401 => x"79",
          7402 => x"69",
          7403 => x"00",
          7404 => x"63",
          7405 => x"6d",
          7406 => x"00",
          7407 => x"20",
          7408 => x"00",
          7409 => x"2c",
          7410 => x"69",
          7411 => x"65",
          7412 => x"00",
          7413 => x"61",
          7414 => x"00",
          7415 => x"61",
          7416 => x"69",
          7417 => x"6d",
          7418 => x"6f",
          7419 => x"00",
          7420 => x"74",
          7421 => x"64",
          7422 => x"76",
          7423 => x"72",
          7424 => x"61",
          7425 => x"00",
          7426 => x"72",
          7427 => x"74",
          7428 => x"00",
          7429 => x"6e",
          7430 => x"61",
          7431 => x"00",
          7432 => x"72",
          7433 => x"69",
          7434 => x"00",
          7435 => x"64",
          7436 => x"00",
          7437 => x"20",
          7438 => x"65",
          7439 => x"70",
          7440 => x"6e",
          7441 => x"66",
          7442 => x"6e",
          7443 => x"6b",
          7444 => x"61",
          7445 => x"65",
          7446 => x"72",
          7447 => x"6b",
          7448 => x"00",
          7449 => x"2e",
          7450 => x"75",
          7451 => x"25",
          7452 => x"75",
          7453 => x"73",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"58",
          7458 => x"00",
          7459 => x"00",
          7460 => x"00",
          7461 => x"20",
          7462 => x"00",
          7463 => x"00",
          7464 => x"30",
          7465 => x"32",
          7466 => x"55",
          7467 => x"30",
          7468 => x"25",
          7469 => x"00",
          7470 => x"20",
          7471 => x"64",
          7472 => x"20",
          7473 => x"20",
          7474 => x"78",
          7475 => x"20",
          7476 => x"72",
          7477 => x"20",
          7478 => x"20",
          7479 => x"78",
          7480 => x"20",
          7481 => x"70",
          7482 => x"65",
          7483 => x"54",
          7484 => x"74",
          7485 => x"00",
          7486 => x"58",
          7487 => x"75",
          7488 => x"54",
          7489 => x"74",
          7490 => x"00",
          7491 => x"58",
          7492 => x"75",
          7493 => x"54",
          7494 => x"74",
          7495 => x"00",
          7496 => x"44",
          7497 => x"75",
          7498 => x"20",
          7499 => x"70",
          7500 => x"65",
          7501 => x"72",
          7502 => x"74",
          7503 => x"74",
          7504 => x"00",
          7505 => x"67",
          7506 => x"2e",
          7507 => x"6f",
          7508 => x"74",
          7509 => x"5f",
          7510 => x"00",
          7511 => x"74",
          7512 => x"61",
          7513 => x"20",
          7514 => x"20",
          7515 => x"69",
          7516 => x"75",
          7517 => x"00",
          7518 => x"5c",
          7519 => x"00",
          7520 => x"6d",
          7521 => x"00",
          7522 => x"00",
          7523 => x"25",
          7524 => x"00",
          7525 => x"62",
          7526 => x"2e",
          7527 => x"74",
          7528 => x"61",
          7529 => x"69",
          7530 => x"00",
          7531 => x"20",
          7532 => x"25",
          7533 => x"2e",
          7534 => x"6c",
          7535 => x"65",
          7536 => x"28",
          7537 => x"00",
          7538 => x"6e",
          7539 => x"40",
          7540 => x"2e",
          7541 => x"6c",
          7542 => x"2d",
          7543 => x"6c",
          7544 => x"00",
          7545 => x"6e",
          7546 => x"00",
          7547 => x"30",
          7548 => x"38",
          7549 => x"29",
          7550 => x"79",
          7551 => x"00",
          7552 => x"30",
          7553 => x"61",
          7554 => x"2e",
          7555 => x"70",
          7556 => x"00",
          7557 => x"74",
          7558 => x"5c",
          7559 => x"00",
          7560 => x"65",
          7561 => x"64",
          7562 => x"74",
          7563 => x"73",
          7564 => x"64",
          7565 => x"00",
          7566 => x"64",
          7567 => x"25",
          7568 => x"00",
          7569 => x"66",
          7570 => x"6f",
          7571 => x"65",
          7572 => x"6d",
          7573 => x"65",
          7574 => x"72",
          7575 => x"00",
          7576 => x"20",
          7577 => x"65",
          7578 => x"64",
          7579 => x"25",
          7580 => x"00",
          7581 => x"20",
          7582 => x"53",
          7583 => x"64",
          7584 => x"25",
          7585 => x"00",
          7586 => x"63",
          7587 => x"20",
          7588 => x"20",
          7589 => x"25",
          7590 => x"00",
          7591 => x"00",
          7592 => x"20",
          7593 => x"20",
          7594 => x"20",
          7595 => x"25",
          7596 => x"00",
          7597 => x"74",
          7598 => x"6b",
          7599 => x"20",
          7600 => x"25",
          7601 => x"48",
          7602 => x"20",
          7603 => x"65",
          7604 => x"43",
          7605 => x"65",
          7606 => x"30",
          7607 => x"00",
          7608 => x"41",
          7609 => x"20",
          7610 => x"20",
          7611 => x"25",
          7612 => x"48",
          7613 => x"20",
          7614 => x"20",
          7615 => x"20",
          7616 => x"00",
          7617 => x"49",
          7618 => x"20",
          7619 => x"45",
          7620 => x"00",
          7621 => x"52",
          7622 => x"43",
          7623 => x"3d",
          7624 => x"00",
          7625 => x"45",
          7626 => x"54",
          7627 => x"3d",
          7628 => x"00",
          7629 => x"43",
          7630 => x"44",
          7631 => x"3d",
          7632 => x"00",
          7633 => x"20",
          7634 => x"25",
          7635 => x"58",
          7636 => x"20",
          7637 => x"20",
          7638 => x"3a",
          7639 => x"00",
          7640 => x"4e",
          7641 => x"25",
          7642 => x"58",
          7643 => x"20",
          7644 => x"20",
          7645 => x"3a",
          7646 => x"00",
          7647 => x"53",
          7648 => x"25",
          7649 => x"58",
          7650 => x"72",
          7651 => x"63",
          7652 => x"00",
          7653 => x"00",
          7654 => x"00",
          7655 => x"00",
          7656 => x"00",
          7657 => x"00",
          7658 => x"ac",
          7659 => x"02",
          7660 => x"00",
          7661 => x"a4",
          7662 => x"04",
          7663 => x"00",
          7664 => x"9c",
          7665 => x"06",
          7666 => x"00",
          7667 => x"94",
          7668 => x"01",
          7669 => x"00",
          7670 => x"8c",
          7671 => x"0b",
          7672 => x"00",
          7673 => x"84",
          7674 => x"0a",
          7675 => x"00",
          7676 => x"7c",
          7677 => x"0c",
          7678 => x"00",
          7679 => x"74",
          7680 => x"0f",
          7681 => x"00",
          7682 => x"6c",
          7683 => x"10",
          7684 => x"00",
          7685 => x"64",
          7686 => x"12",
          7687 => x"00",
          7688 => x"5c",
          7689 => x"14",
          7690 => x"00",
          7691 => x"00",
          7692 => x"00",
          7693 => x"7e",
          7694 => x"7e",
          7695 => x"7e",
          7696 => x"7e",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"6e",
          7703 => x"2f",
          7704 => x"68",
          7705 => x"66",
          7706 => x"73",
          7707 => x"00",
          7708 => x"00",
          7709 => x"00",
          7710 => x"6c",
          7711 => x"00",
          7712 => x"74",
          7713 => x"20",
          7714 => x"74",
          7715 => x"65",
          7716 => x"2e",
          7717 => x"0a",
          7718 => x"7e",
          7719 => x"00",
          7720 => x"00",
          7721 => x"30",
          7722 => x"31",
          7723 => x"32",
          7724 => x"33",
          7725 => x"34",
          7726 => x"35",
          7727 => x"37",
          7728 => x"38",
          7729 => x"39",
          7730 => x"30",
          7731 => x"7e",
          7732 => x"7e",
          7733 => x"00",
          7734 => x"00",
          7735 => x"00",
          7736 => x"2c",
          7737 => x"64",
          7738 => x"78",
          7739 => x"64",
          7740 => x"25",
          7741 => x"2c",
          7742 => x"00",
          7743 => x"00",
          7744 => x"00",
          7745 => x"64",
          7746 => x"6f",
          7747 => x"6f",
          7748 => x"25",
          7749 => x"78",
          7750 => x"25",
          7751 => x"78",
          7752 => x"25",
          7753 => x"00",
          7754 => x"20",
          7755 => x"2e",
          7756 => x"00",
          7757 => x"7f",
          7758 => x"3d",
          7759 => x"00",
          7760 => x"00",
          7761 => x"53",
          7762 => x"4e",
          7763 => x"46",
          7764 => x"00",
          7765 => x"20",
          7766 => x"32",
          7767 => x"60",
          7768 => x"00",
          7769 => x"07",
          7770 => x"1c",
          7771 => x"41",
          7772 => x"49",
          7773 => x"4f",
          7774 => x"9b",
          7775 => x"55",
          7776 => x"ab",
          7777 => x"b3",
          7778 => x"bb",
          7779 => x"c3",
          7780 => x"cb",
          7781 => x"d3",
          7782 => x"db",
          7783 => x"e3",
          7784 => x"eb",
          7785 => x"f3",
          7786 => x"fb",
          7787 => x"3b",
          7788 => x"3a",
          7789 => x"00",
          7790 => x"40",
          7791 => x"00",
          7792 => x"08",
          7793 => x"00",
          7794 => x"e2",
          7795 => x"e7",
          7796 => x"ef",
          7797 => x"c5",
          7798 => x"f4",
          7799 => x"f9",
          7800 => x"a2",
          7801 => x"92",
          7802 => x"fa",
          7803 => x"ba",
          7804 => x"bd",
          7805 => x"bb",
          7806 => x"02",
          7807 => x"56",
          7808 => x"57",
          7809 => x"10",
          7810 => x"1c",
          7811 => x"5f",
          7812 => x"66",
          7813 => x"67",
          7814 => x"59",
          7815 => x"6b",
          7816 => x"88",
          7817 => x"80",
          7818 => x"c0",
          7819 => x"c4",
          7820 => x"b4",
          7821 => x"29",
          7822 => x"64",
          7823 => x"48",
          7824 => x"1a",
          7825 => x"a0",
          7826 => x"17",
          7827 => x"01",
          7828 => x"32",
          7829 => x"4a",
          7830 => x"80",
          7831 => x"82",
          7832 => x"86",
          7833 => x"8a",
          7834 => x"8e",
          7835 => x"91",
          7836 => x"96",
          7837 => x"3d",
          7838 => x"20",
          7839 => x"a2",
          7840 => x"a6",
          7841 => x"aa",
          7842 => x"ae",
          7843 => x"b2",
          7844 => x"b5",
          7845 => x"ba",
          7846 => x"be",
          7847 => x"c2",
          7848 => x"c4",
          7849 => x"ca",
          7850 => x"10",
          7851 => x"de",
          7852 => x"f1",
          7853 => x"28",
          7854 => x"09",
          7855 => x"3d",
          7856 => x"41",
          7857 => x"53",
          7858 => x"55",
          7859 => x"8f",
          7860 => x"5d",
          7861 => x"61",
          7862 => x"65",
          7863 => x"96",
          7864 => x"6d",
          7865 => x"71",
          7866 => x"9f",
          7867 => x"79",
          7868 => x"64",
          7869 => x"81",
          7870 => x"85",
          7871 => x"44",
          7872 => x"8d",
          7873 => x"91",
          7874 => x"fd",
          7875 => x"04",
          7876 => x"8a",
          7877 => x"02",
          7878 => x"08",
          7879 => x"8e",
          7880 => x"f2",
          7881 => x"f4",
          7882 => x"f7",
          7883 => x"30",
          7884 => x"60",
          7885 => x"c1",
          7886 => x"c0",
          7887 => x"26",
          7888 => x"01",
          7889 => x"a0",
          7890 => x"10",
          7891 => x"30",
          7892 => x"51",
          7893 => x"5b",
          7894 => x"5f",
          7895 => x"0e",
          7896 => x"c9",
          7897 => x"db",
          7898 => x"eb",
          7899 => x"08",
          7900 => x"08",
          7901 => x"b9",
          7902 => x"01",
          7903 => x"e0",
          7904 => x"ec",
          7905 => x"4e",
          7906 => x"10",
          7907 => x"d0",
          7908 => x"60",
          7909 => x"75",
          7910 => x"00",
          7911 => x"00",
          7912 => x"68",
          7913 => x"00",
          7914 => x"70",
          7915 => x"00",
          7916 => x"78",
          7917 => x"00",
          7918 => x"80",
          7919 => x"00",
          7920 => x"88",
          7921 => x"00",
          7922 => x"90",
          7923 => x"00",
          7924 => x"98",
          7925 => x"00",
          7926 => x"a0",
          7927 => x"00",
          7928 => x"a8",
          7929 => x"00",
          7930 => x"b0",
          7931 => x"00",
          7932 => x"b4",
          7933 => x"00",
          7934 => x"b8",
          7935 => x"00",
          7936 => x"bc",
          7937 => x"00",
          7938 => x"c0",
          7939 => x"00",
          7940 => x"c4",
          7941 => x"00",
          7942 => x"c8",
          7943 => x"00",
          7944 => x"cc",
          7945 => x"00",
          7946 => x"d4",
          7947 => x"00",
          7948 => x"d8",
          7949 => x"00",
          7950 => x"e0",
          7951 => x"00",
          7952 => x"e8",
          7953 => x"00",
          7954 => x"f0",
          7955 => x"00",
          7956 => x"f8",
          7957 => x"00",
          7958 => x"fc",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"08",
          7963 => x"00",
          7964 => x"10",
          7965 => x"00",
          7966 => x"18",
          7967 => x"00",
          7968 => x"00",
          7969 => x"ff",
          7970 => x"ff",
          7971 => x"ff",
          7972 => x"00",
          7973 => x"ff",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"01",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"00",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"fd",
          7996 => x"5b",
          7997 => x"74",
          7998 => x"6c",
          7999 => x"64",
          8000 => x"34",
          8001 => x"20",
          8002 => x"f4",
          8003 => x"f0",
          8004 => x"83",
          8005 => x"fd",
          8006 => x"5b",
          8007 => x"54",
          8008 => x"4c",
          8009 => x"44",
          8010 => x"34",
          8011 => x"20",
          8012 => x"f4",
          8013 => x"f0",
          8014 => x"83",
          8015 => x"fd",
          8016 => x"7b",
          8017 => x"54",
          8018 => x"4c",
          8019 => x"44",
          8020 => x"24",
          8021 => x"20",
          8022 => x"e1",
          8023 => x"f0",
          8024 => x"88",
          8025 => x"fa",
          8026 => x"1b",
          8027 => x"14",
          8028 => x"0c",
          8029 => x"04",
          8030 => x"f0",
          8031 => x"f0",
          8032 => x"f0",
          8033 => x"f0",
          8034 => x"83",
          8035 => x"c9",
          8036 => x"b3",
          8037 => x"31",
          8038 => x"56",
          8039 => x"48",
          8040 => x"3b",
          8041 => x"00",
          8042 => x"c1",
          8043 => x"f0",
          8044 => x"83",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"30",
          8060 => x"38",
          8061 => x"3c",
          8062 => x"40",
          8063 => x"44",
          8064 => x"48",
          8065 => x"50",
          8066 => x"58",
          8067 => x"60",
          8068 => x"68",
          8069 => x"70",
          8070 => x"78",
          8071 => x"80",
          8072 => x"88",
          8073 => x"90",
          8074 => x"98",
          8075 => x"a0",
          8076 => x"a8",
          8077 => x"ac",
          8078 => x"b4",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"19",
          9080 => x"00",
          9081 => x"f7",
          9082 => x"ff",
          9083 => x"e2",
          9084 => x"f4",
          9085 => x"67",
          9086 => x"2d",
          9087 => x"27",
          9088 => x"49",
          9089 => x"07",
          9090 => x"0f",
          9091 => x"17",
          9092 => x"3c",
          9093 => x"87",
          9094 => x"8f",
          9095 => x"97",
          9096 => x"c0",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"01",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"e9",
             2 => x"00",
             3 => x"00",
             4 => x"8c",
             5 => x"90",
             6 => x"00",
             7 => x"00",
             8 => x"06",
             9 => x"82",
            10 => x"06",
            11 => x"00",
            12 => x"06",
            13 => x"09",
            14 => x"09",
            15 => x"0b",
            16 => x"81",
            17 => x"09",
            18 => x"81",
            19 => x"00",
            20 => x"24",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"05",
            26 => x"0a",
            27 => x"53",
            28 => x"26",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"9f",
            45 => x"93",
            46 => x"00",
            47 => x"00",
            48 => x"2a",
            49 => x"09",
            50 => x"53",
            51 => x"00",
            52 => x"53",
            53 => x"81",
            54 => x"07",
            55 => x"00",
            56 => x"81",
            57 => x"09",
            58 => x"00",
            59 => x"00",
            60 => x"81",
            61 => x"09",
            62 => x"04",
            63 => x"00",
            64 => x"81",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"09",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"72",
            73 => x"51",
            74 => x"00",
            75 => x"00",
            76 => x"06",
            77 => x"83",
            78 => x"06",
            79 => x"00",
            80 => x"06",
            81 => x"83",
            82 => x"0b",
            83 => x"00",
            84 => x"8c",
            85 => x"0b",
            86 => x"56",
            87 => x"04",
            88 => x"8c",
            89 => x"0b",
            90 => x"56",
            91 => x"04",
            92 => x"70",
            93 => x"ff",
            94 => x"72",
            95 => x"51",
            96 => x"70",
            97 => x"06",
            98 => x"09",
            99 => x"51",
           100 => x"05",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"05",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"05",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"05",
           125 => x"04",
           126 => x"ff",
           127 => x"ff",
           128 => x"06",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"85",
           134 => x"0b",
           135 => x"0b",
           136 => x"c6",
           137 => x"0b",
           138 => x"0b",
           139 => x"86",
           140 => x"0b",
           141 => x"0b",
           142 => x"c6",
           143 => x"0b",
           144 => x"0b",
           145 => x"8a",
           146 => x"0b",
           147 => x"0b",
           148 => x"ce",
           149 => x"0b",
           150 => x"0b",
           151 => x"92",
           152 => x"0b",
           153 => x"0b",
           154 => x"d6",
           155 => x"0b",
           156 => x"0b",
           157 => x"9a",
           158 => x"0b",
           159 => x"0b",
           160 => x"de",
           161 => x"0b",
           162 => x"0b",
           163 => x"a2",
           164 => x"0b",
           165 => x"0b",
           166 => x"e6",
           167 => x"0b",
           168 => x"0b",
           169 => x"aa",
           170 => x"0b",
           171 => x"0b",
           172 => x"ed",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"8c",
           193 => x"d6",
           194 => x"c0",
           195 => x"a2",
           196 => x"c0",
           197 => x"a0",
           198 => x"c0",
           199 => x"a0",
           200 => x"c0",
           201 => x"94",
           202 => x"c0",
           203 => x"a1",
           204 => x"c0",
           205 => x"af",
           206 => x"c0",
           207 => x"ad",
           208 => x"c0",
           209 => x"94",
           210 => x"c0",
           211 => x"95",
           212 => x"c0",
           213 => x"95",
           214 => x"c0",
           215 => x"b1",
           216 => x"c0",
           217 => x"80",
           218 => x"80",
           219 => x"0c",
           220 => x"08",
           221 => x"d4",
           222 => x"d4",
           223 => x"b9",
           224 => x"b9",
           225 => x"84",
           226 => x"84",
           227 => x"04",
           228 => x"2d",
           229 => x"90",
           230 => x"9e",
           231 => x"80",
           232 => x"d7",
           233 => x"c0",
           234 => x"82",
           235 => x"80",
           236 => x"0c",
           237 => x"08",
           238 => x"d4",
           239 => x"d4",
           240 => x"b9",
           241 => x"b9",
           242 => x"84",
           243 => x"84",
           244 => x"04",
           245 => x"2d",
           246 => x"90",
           247 => x"a2",
           248 => x"80",
           249 => x"fe",
           250 => x"c0",
           251 => x"83",
           252 => x"80",
           253 => x"0c",
           254 => x"08",
           255 => x"d4",
           256 => x"d4",
           257 => x"b9",
           258 => x"b9",
           259 => x"84",
           260 => x"84",
           261 => x"04",
           262 => x"2d",
           263 => x"90",
           264 => x"8e",
           265 => x"80",
           266 => x"f6",
           267 => x"c0",
           268 => x"83",
           269 => x"80",
           270 => x"0c",
           271 => x"08",
           272 => x"d4",
           273 => x"d4",
           274 => x"b9",
           275 => x"b9",
           276 => x"84",
           277 => x"84",
           278 => x"04",
           279 => x"2d",
           280 => x"90",
           281 => x"c5",
           282 => x"80",
           283 => x"f3",
           284 => x"c0",
           285 => x"81",
           286 => x"80",
           287 => x"0c",
           288 => x"08",
           289 => x"d4",
           290 => x"d4",
           291 => x"b9",
           292 => x"b9",
           293 => x"84",
           294 => x"84",
           295 => x"04",
           296 => x"84",
           297 => x"04",
           298 => x"2d",
           299 => x"90",
           300 => x"bc",
           301 => x"80",
           302 => x"f1",
           303 => x"c0",
           304 => x"81",
           305 => x"80",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"04",
           311 => x"83",
           312 => x"10",
           313 => x"51",
           314 => x"06",
           315 => x"10",
           316 => x"ed",
           317 => x"b9",
           318 => x"38",
           319 => x"0b",
           320 => x"51",
           321 => x"0d",
           322 => x"08",
           323 => x"08",
           324 => x"04",
           325 => x"11",
           326 => x"25",
           327 => x"72",
           328 => x"38",
           329 => x"30",
           330 => x"55",
           331 => x"71",
           332 => x"fa",
           333 => x"b9",
           334 => x"b9",
           335 => x"34",
           336 => x"70",
           337 => x"54",
           338 => x"34",
           339 => x"88",
           340 => x"c8",
           341 => x"0d",
           342 => x"05",
           343 => x"3d",
           344 => x"e4",
           345 => x"80",
           346 => x"3d",
           347 => x"52",
           348 => x"04",
           349 => x"5d",
           350 => x"1e",
           351 => x"06",
           352 => x"2e",
           353 => x"33",
           354 => x"81",
           355 => x"80",
           356 => x"7e",
           357 => x"32",
           358 => x"55",
           359 => x"38",
           360 => x"06",
           361 => x"7a",
           362 => x"76",
           363 => x"73",
           364 => x"04",
           365 => x"10",
           366 => x"98",
           367 => x"8b",
           368 => x"5b",
           369 => x"38",
           370 => x"38",
           371 => x"f7",
           372 => x"09",
           373 => x"5a",
           374 => x"76",
           375 => x"52",
           376 => x"57",
           377 => x"7a",
           378 => x"78",
           379 => x"54",
           380 => x"80",
           381 => x"83",
           382 => x"73",
           383 => x"27",
           384 => x"eb",
           385 => x"fe",
           386 => x"59",
           387 => x"84",
           388 => x"06",
           389 => x"5e",
           390 => x"84",
           391 => x"b9",
           392 => x"72",
           393 => x"08",
           394 => x"05",
           395 => x"ca",
           396 => x"b9",
           397 => x"d8",
           398 => x"56",
           399 => x"80",
           400 => x"90",
           401 => x"81",
           402 => x"38",
           403 => x"80",
           404 => x"77",
           405 => x"05",
           406 => x"2a",
           407 => x"2e",
           408 => x"ff",
           409 => x"cc",
           410 => x"83",
           411 => x"74",
           412 => x"f0",
           413 => x"90",
           414 => x"53",
           415 => x"81",
           416 => x"38",
           417 => x"86",
           418 => x"54",
           419 => x"54",
           420 => x"81",
           421 => x"77",
           422 => x"80",
           423 => x"80",
           424 => x"51",
           425 => x"80",
           426 => x"2c",
           427 => x"38",
           428 => x"b2",
           429 => x"81",
           430 => x"55",
           431 => x"52",
           432 => x"81",
           433 => x"70",
           434 => x"24",
           435 => x"06",
           436 => x"38",
           437 => x"76",
           438 => x"80",
           439 => x"b9",
           440 => x"1e",
           441 => x"7d",
           442 => x"ec",
           443 => x"2e",
           444 => x"80",
           445 => x"2c",
           446 => x"91",
           447 => x"3f",
           448 => x"a0",
           449 => x"87",
           450 => x"07",
           451 => x"84",
           452 => x"06",
           453 => x"39",
           454 => x"0a",
           455 => x"72",
           456 => x"80",
           457 => x"5a",
           458 => x"70",
           459 => x"38",
           460 => x"80",
           461 => x"5f",
           462 => x"52",
           463 => x"ff",
           464 => x"57",
           465 => x"38",
           466 => x"33",
           467 => x"1a",
           468 => x"79",
           469 => x"7c",
           470 => x"51",
           471 => x"0a",
           472 => x"80",
           473 => x"90",
           474 => x"87",
           475 => x"7a",
           476 => x"60",
           477 => x"41",
           478 => x"7a",
           479 => x"d8",
           480 => x"7c",
           481 => x"f8",
           482 => x"7c",
           483 => x"f8",
           484 => x"08",
           485 => x"72",
           486 => x"3f",
           487 => x"06",
           488 => x"72",
           489 => x"80",
           490 => x"f7",
           491 => x"84",
           492 => x"58",
           493 => x"51",
           494 => x"83",
           495 => x"2b",
           496 => x"07",
           497 => x"38",
           498 => x"80",
           499 => x"2c",
           500 => x"d6",
           501 => x"3f",
           502 => x"bb",
           503 => x"fa",
           504 => x"ab",
           505 => x"7e",
           506 => x"39",
           507 => x"2b",
           508 => x"57",
           509 => x"ff",
           510 => x"fb",
           511 => x"2e",
           512 => x"52",
           513 => x"74",
           514 => x"f1",
           515 => x"98",
           516 => x"b7",
           517 => x"3f",
           518 => x"bb",
           519 => x"51",
           520 => x"83",
           521 => x"2b",
           522 => x"07",
           523 => x"52",
           524 => x"0d",
           525 => x"74",
           526 => x"04",
           527 => x"84",
           528 => x"81",
           529 => x"56",
           530 => x"2e",
           531 => x"70",
           532 => x"2e",
           533 => x"72",
           534 => x"84",
           535 => x"ff",
           536 => x"53",
           537 => x"ac",
           538 => x"08",
           539 => x"51",
           540 => x"b9",
           541 => x"57",
           542 => x"88",
           543 => x"7a",
           544 => x"70",
           545 => x"51",
           546 => x"2e",
           547 => x"81",
           548 => x"09",
           549 => x"84",
           550 => x"73",
           551 => x"80",
           552 => x"90",
           553 => x"c8",
           554 => x"70",
           555 => x"e3",
           556 => x"d5",
           557 => x"83",
           558 => x"7a",
           559 => x"32",
           560 => x"56",
           561 => x"06",
           562 => x"15",
           563 => x"91",
           564 => x"74",
           565 => x"08",
           566 => x"56",
           567 => x"0d",
           568 => x"51",
           569 => x"56",
           570 => x"15",
           571 => x"56",
           572 => x"11",
           573 => x"32",
           574 => x"54",
           575 => x"06",
           576 => x"81",
           577 => x"38",
           578 => x"80",
           579 => x"0c",
           580 => x"0c",
           581 => x"b9",
           582 => x"ff",
           583 => x"8c",
           584 => x"84",
           585 => x"3d",
           586 => x"55",
           587 => x"84",
           588 => x"38",
           589 => x"52",
           590 => x"38",
           591 => x"34",
           592 => x"87",
           593 => x"72",
           594 => x"fd",
           595 => x"54",
           596 => x"70",
           597 => x"81",
           598 => x"81",
           599 => x"84",
           600 => x"fc",
           601 => x"55",
           602 => x"73",
           603 => x"93",
           604 => x"73",
           605 => x"51",
           606 => x"0c",
           607 => x"73",
           608 => x"53",
           609 => x"71",
           610 => x"80",
           611 => x"53",
           612 => x"51",
           613 => x"0d",
           614 => x"05",
           615 => x"12",
           616 => x"51",
           617 => x"75",
           618 => x"81",
           619 => x"81",
           620 => x"84",
           621 => x"fd",
           622 => x"55",
           623 => x"71",
           624 => x"81",
           625 => x"ef",
           626 => x"3d",
           627 => x"7a",
           628 => x"38",
           629 => x"33",
           630 => x"06",
           631 => x"2e",
           632 => x"38",
           633 => x"86",
           634 => x"38",
           635 => x"2e",
           636 => x"51",
           637 => x"31",
           638 => x"04",
           639 => x"0d",
           640 => x"70",
           641 => x"c8",
           642 => x"52",
           643 => x"c8",
           644 => x"2e",
           645 => x"54",
           646 => x"84",
           647 => x"84",
           648 => x"c8",
           649 => x"0d",
           650 => x"54",
           651 => x"81",
           652 => x"8c",
           653 => x"09",
           654 => x"75",
           655 => x"0c",
           656 => x"75",
           657 => x"70",
           658 => x"81",
           659 => x"f4",
           660 => x"3d",
           661 => x"58",
           662 => x"38",
           663 => x"c8",
           664 => x"2e",
           665 => x"71",
           666 => x"52",
           667 => x"52",
           668 => x"13",
           669 => x"71",
           670 => x"74",
           671 => x"9f",
           672 => x"72",
           673 => x"06",
           674 => x"1c",
           675 => x"53",
           676 => x"52",
           677 => x"0d",
           678 => x"80",
           679 => x"80",
           680 => x"75",
           681 => x"70",
           682 => x"71",
           683 => x"06",
           684 => x"84",
           685 => x"75",
           686 => x"70",
           687 => x"71",
           688 => x"81",
           689 => x"75",
           690 => x"52",
           691 => x"55",
           692 => x"51",
           693 => x"04",
           694 => x"71",
           695 => x"b9",
           696 => x"84",
           697 => x"04",
           698 => x"a0",
           699 => x"51",
           700 => x"53",
           701 => x"38",
           702 => x"b9",
           703 => x"9f",
           704 => x"9f",
           705 => x"2a",
           706 => x"54",
           707 => x"a8",
           708 => x"74",
           709 => x"11",
           710 => x"06",
           711 => x"52",
           712 => x"38",
           713 => x"0d",
           714 => x"7a",
           715 => x"7c",
           716 => x"71",
           717 => x"59",
           718 => x"84",
           719 => x"84",
           720 => x"f7",
           721 => x"70",
           722 => x"56",
           723 => x"8f",
           724 => x"33",
           725 => x"73",
           726 => x"2e",
           727 => x"56",
           728 => x"58",
           729 => x"38",
           730 => x"14",
           731 => x"14",
           732 => x"73",
           733 => x"ff",
           734 => x"89",
           735 => x"77",
           736 => x"0c",
           737 => x"26",
           738 => x"38",
           739 => x"56",
           740 => x"0d",
           741 => x"70",
           742 => x"09",
           743 => x"70",
           744 => x"80",
           745 => x"80",
           746 => x"74",
           747 => x"56",
           748 => x"38",
           749 => x"0d",
           750 => x"0c",
           751 => x"ca",
           752 => x"8b",
           753 => x"7d",
           754 => x"08",
           755 => x"2e",
           756 => x"70",
           757 => x"a0",
           758 => x"f5",
           759 => x"d0",
           760 => x"80",
           761 => x"74",
           762 => x"27",
           763 => x"06",
           764 => x"06",
           765 => x"f9",
           766 => x"89",
           767 => x"27",
           768 => x"81",
           769 => x"56",
           770 => x"78",
           771 => x"75",
           772 => x"c8",
           773 => x"16",
           774 => x"59",
           775 => x"ff",
           776 => x"33",
           777 => x"38",
           778 => x"38",
           779 => x"d0",
           780 => x"73",
           781 => x"c8",
           782 => x"81",
           783 => x"55",
           784 => x"84",
           785 => x"80",
           786 => x"81",
           787 => x"ff",
           788 => x"8c",
           789 => x"05",
           790 => x"51",
           791 => x"83",
           792 => x"3d",
           793 => x"a8",
           794 => x"dc",
           795 => x"04",
           796 => x"83",
           797 => x"ef",
           798 => x"cf",
           799 => x"0d",
           800 => x"3f",
           801 => x"51",
           802 => x"83",
           803 => x"3d",
           804 => x"d0",
           805 => x"a4",
           806 => x"04",
           807 => x"83",
           808 => x"ee",
           809 => x"d0",
           810 => x"0d",
           811 => x"3f",
           812 => x"51",
           813 => x"83",
           814 => x"3d",
           815 => x"f8",
           816 => x"b8",
           817 => x"04",
           818 => x"83",
           819 => x"02",
           820 => x"58",
           821 => x"73",
           822 => x"75",
           823 => x"74",
           824 => x"55",
           825 => x"53",
           826 => x"82",
           827 => x"57",
           828 => x"d0",
           829 => x"76",
           830 => x"30",
           831 => x"57",
           832 => x"c0",
           833 => x"26",
           834 => x"e8",
           835 => x"c8",
           836 => x"52",
           837 => x"76",
           838 => x"04",
           839 => x"88",
           840 => x"3d",
           841 => x"52",
           842 => x"b9",
           843 => x"ff",
           844 => x"ff",
           845 => x"59",
           846 => x"f4",
           847 => x"78",
           848 => x"08",
           849 => x"83",
           850 => x"97",
           851 => x"05",
           852 => x"80",
           853 => x"3f",
           854 => x"80",
           855 => x"38",
           856 => x"0d",
           857 => x"61",
           858 => x"7f",
           859 => x"c8",
           860 => x"0d",
           861 => x"02",
           862 => x"73",
           863 => x"5d",
           864 => x"7a",
           865 => x"3f",
           866 => x"80",
           867 => x"90",
           868 => x"82",
           869 => x"27",
           870 => x"d2",
           871 => x"84",
           872 => x"ec",
           873 => x"83",
           874 => x"56",
           875 => x"18",
           876 => x"7a",
           877 => x"9f",
           878 => x"73",
           879 => x"74",
           880 => x"27",
           881 => x"52",
           882 => x"56",
           883 => x"94",
           884 => x"1c",
           885 => x"84",
           886 => x"2c",
           887 => x"38",
           888 => x"1e",
           889 => x"ff",
           890 => x"0d",
           891 => x"3f",
           892 => x"54",
           893 => x"26",
           894 => x"d2",
           895 => x"84",
           896 => x"ea",
           897 => x"38",
           898 => x"38",
           899 => x"db",
           900 => x"08",
           901 => x"78",
           902 => x"83",
           903 => x"14",
           904 => x"51",
           905 => x"ff",
           906 => x"df",
           907 => x"51",
           908 => x"ac",
           909 => x"3f",
           910 => x"39",
           911 => x"e9",
           912 => x"39",
           913 => x"08",
           914 => x"a8",
           915 => x"80",
           916 => x"38",
           917 => x"9b",
           918 => x"2b",
           919 => x"30",
           920 => x"07",
           921 => x"59",
           922 => x"e8",
           923 => x"b9",
           924 => x"70",
           925 => x"70",
           926 => x"06",
           927 => x"80",
           928 => x"39",
           929 => x"3d",
           930 => x"96",
           931 => x"51",
           932 => x"9d",
           933 => x"72",
           934 => x"71",
           935 => x"81",
           936 => x"72",
           937 => x"71",
           938 => x"81",
           939 => x"72",
           940 => x"71",
           941 => x"81",
           942 => x"72",
           943 => x"71",
           944 => x"53",
           945 => x"3d",
           946 => x"83",
           947 => x"51",
           948 => x"3d",
           949 => x"83",
           950 => x"51",
           951 => x"06",
           952 => x"39",
           953 => x"80",
           954 => x"d2",
           955 => x"51",
           956 => x"c2",
           957 => x"d4",
           958 => x"9b",
           959 => x"06",
           960 => x"38",
           961 => x"3f",
           962 => x"80",
           963 => x"70",
           964 => x"fe",
           965 => x"9a",
           966 => x"8a",
           967 => x"84",
           968 => x"80",
           969 => x"81",
           970 => x"51",
           971 => x"3f",
           972 => x"52",
           973 => x"bd",
           974 => x"d4",
           975 => x"9a",
           976 => x"06",
           977 => x"38",
           978 => x"70",
           979 => x"0c",
           980 => x"8c",
           981 => x"06",
           982 => x"84",
           983 => x"b8",
           984 => x"51",
           985 => x"53",
           986 => x"0b",
           987 => x"ff",
           988 => x"f1",
           989 => x"78",
           990 => x"83",
           991 => x"80",
           992 => x"7b",
           993 => x"81",
           994 => x"2e",
           995 => x"be",
           996 => x"05",
           997 => x"84",
           998 => x"54",
           999 => x"da",
          1000 => x"84",
          1001 => x"80",
          1002 => x"5d",
          1003 => x"3d",
          1004 => x"38",
          1005 => x"3f",
          1006 => x"c8",
          1007 => x"b9",
          1008 => x"05",
          1009 => x"08",
          1010 => x"2e",
          1011 => x"51",
          1012 => x"8f",
          1013 => x"3d",
          1014 => x"38",
          1015 => x"81",
          1016 => x"53",
          1017 => x"dd",
          1018 => x"f8",
          1019 => x"90",
          1020 => x"7c",
          1021 => x"08",
          1022 => x"70",
          1023 => x"42",
          1024 => x"81",
          1025 => x"2e",
          1026 => x"06",
          1027 => x"81",
          1028 => x"81",
          1029 => x"38",
          1030 => x"d5",
          1031 => x"80",
          1032 => x"bc",
          1033 => x"70",
          1034 => x"91",
          1035 => x"84",
          1036 => x"84",
          1037 => x"0b",
          1038 => x"d0",
          1039 => x"82",
          1040 => x"80",
          1041 => x"51",
          1042 => x"bc",
          1043 => x"7d",
          1044 => x"38",
          1045 => x"a1",
          1046 => x"ee",
          1047 => x"f8",
          1048 => x"70",
          1049 => x"39",
          1050 => x"59",
          1051 => x"78",
          1052 => x"79",
          1053 => x"52",
          1054 => x"7e",
          1055 => x"84",
          1056 => x"09",
          1057 => x"9a",
          1058 => x"83",
          1059 => x"51",
          1060 => x"83",
          1061 => x"90",
          1062 => x"7c",
          1063 => x"81",
          1064 => x"f8",
          1065 => x"51",
          1066 => x"8d",
          1067 => x"a4",
          1068 => x"04",
          1069 => x"d0",
          1070 => x"ff",
          1071 => x"ec",
          1072 => x"2e",
          1073 => x"d4",
          1074 => x"2d",
          1075 => x"a4",
          1076 => x"d6",
          1077 => x"39",
          1078 => x"80",
          1079 => x"c8",
          1080 => x"52",
          1081 => x"68",
          1082 => x"11",
          1083 => x"3f",
          1084 => x"dc",
          1085 => x"ff",
          1086 => x"b9",
          1087 => x"78",
          1088 => x"51",
          1089 => x"53",
          1090 => x"3f",
          1091 => x"2e",
          1092 => x"d3",
          1093 => x"cf",
          1094 => x"ff",
          1095 => x"b9",
          1096 => x"b8",
          1097 => x"05",
          1098 => x"08",
          1099 => x"53",
          1100 => x"a5",
          1101 => x"f8",
          1102 => x"48",
          1103 => x"c4",
          1104 => x"64",
          1105 => x"b8",
          1106 => x"05",
          1107 => x"08",
          1108 => x"fe",
          1109 => x"e9",
          1110 => x"2e",
          1111 => x"11",
          1112 => x"3f",
          1113 => x"f4",
          1114 => x"3f",
          1115 => x"83",
          1116 => x"5f",
          1117 => x"7a",
          1118 => x"52",
          1119 => x"66",
          1120 => x"47",
          1121 => x"11",
          1122 => x"3f",
          1123 => x"a4",
          1124 => x"ff",
          1125 => x"b9",
          1126 => x"b8",
          1127 => x"05",
          1128 => x"08",
          1129 => x"f0",
          1130 => x"67",
          1131 => x"70",
          1132 => x"81",
          1133 => x"84",
          1134 => x"93",
          1135 => x"f6",
          1136 => x"53",
          1137 => x"84",
          1138 => x"33",
          1139 => x"ed",
          1140 => x"f8",
          1141 => x"48",
          1142 => x"8c",
          1143 => x"68",
          1144 => x"02",
          1145 => x"81",
          1146 => x"53",
          1147 => x"84",
          1148 => x"38",
          1149 => x"79",
          1150 => x"fe",
          1151 => x"e7",
          1152 => x"bd",
          1153 => x"84",
          1154 => x"f3",
          1155 => x"f5",
          1156 => x"53",
          1157 => x"84",
          1158 => x"38",
          1159 => x"80",
          1160 => x"c8",
          1161 => x"46",
          1162 => x"68",
          1163 => x"38",
          1164 => x"5b",
          1165 => x"51",
          1166 => x"3d",
          1167 => x"84",
          1168 => x"05",
          1169 => x"84",
          1170 => x"83",
          1171 => x"f4",
          1172 => x"e7",
          1173 => x"ff",
          1174 => x"e5",
          1175 => x"38",
          1176 => x"2e",
          1177 => x"49",
          1178 => x"80",
          1179 => x"c8",
          1180 => x"5a",
          1181 => x"f2",
          1182 => x"11",
          1183 => x"3f",
          1184 => x"38",
          1185 => x"83",
          1186 => x"30",
          1187 => x"5c",
          1188 => x"7a",
          1189 => x"d8",
          1190 => x"68",
          1191 => x"eb",
          1192 => x"b0",
          1193 => x"0c",
          1194 => x"fe",
          1195 => x"e2",
          1196 => x"2e",
          1197 => x"59",
          1198 => x"f0",
          1199 => x"87",
          1200 => x"f2",
          1201 => x"05",
          1202 => x"7d",
          1203 => x"ff",
          1204 => x"b9",
          1205 => x"64",
          1206 => x"70",
          1207 => x"3d",
          1208 => x"51",
          1209 => x"ff",
          1210 => x"fe",
          1211 => x"e3",
          1212 => x"2e",
          1213 => x"db",
          1214 => x"49",
          1215 => x"11",
          1216 => x"3f",
          1217 => x"98",
          1218 => x"84",
          1219 => x"7a",
          1220 => x"38",
          1221 => x"53",
          1222 => x"f5",
          1223 => x"51",
          1224 => x"d8",
          1225 => x"39",
          1226 => x"80",
          1227 => x"c8",
          1228 => x"02",
          1229 => x"05",
          1230 => x"83",
          1231 => x"80",
          1232 => x"fc",
          1233 => x"7b",
          1234 => x"08",
          1235 => x"51",
          1236 => x"39",
          1237 => x"64",
          1238 => x"33",
          1239 => x"f2",
          1240 => x"d8",
          1241 => x"39",
          1242 => x"2e",
          1243 => x"fc",
          1244 => x"7d",
          1245 => x"08",
          1246 => x"33",
          1247 => x"f2",
          1248 => x"f2",
          1249 => x"38",
          1250 => x"39",
          1251 => x"2e",
          1252 => x"fb",
          1253 => x"80",
          1254 => x"b4",
          1255 => x"f3",
          1256 => x"34",
          1257 => x"57",
          1258 => x"d2",
          1259 => x"77",
          1260 => x"75",
          1261 => x"c8",
          1262 => x"9c",
          1263 => x"52",
          1264 => x"c8",
          1265 => x"87",
          1266 => x"3f",
          1267 => x"0c",
          1268 => x"84",
          1269 => x"94",
          1270 => x"c7",
          1271 => x"05",
          1272 => x"89",
          1273 => x"0c",
          1274 => x"3f",
          1275 => x"8d",
          1276 => x"52",
          1277 => x"83",
          1278 => x"97",
          1279 => x"c8",
          1280 => x"d0",
          1281 => x"83",
          1282 => x"52",
          1283 => x"90",
          1284 => x"c3",
          1285 => x"fb",
          1286 => x"80",
          1287 => x"83",
          1288 => x"52",
          1289 => x"91",
          1290 => x"ff",
          1291 => x"f1",
          1292 => x"a2",
          1293 => x"81",
          1294 => x"70",
          1295 => x"a0",
          1296 => x"2e",
          1297 => x"81",
          1298 => x"ff",
          1299 => x"81",
          1300 => x"32",
          1301 => x"52",
          1302 => x"80",
          1303 => x"76",
          1304 => x"0c",
          1305 => x"c4",
          1306 => x"81",
          1307 => x"ff",
          1308 => x"e4",
          1309 => x"55",
          1310 => x"09",
          1311 => x"fc",
          1312 => x"38",
          1313 => x"3d",
          1314 => x"72",
          1315 => x"08",
          1316 => x"c8",
          1317 => x"0d",
          1318 => x"53",
          1319 => x"38",
          1320 => x"52",
          1321 => x"13",
          1322 => x"80",
          1323 => x"52",
          1324 => x"13",
          1325 => x"80",
          1326 => x"52",
          1327 => x"8a",
          1328 => x"e7",
          1329 => x"c0",
          1330 => x"98",
          1331 => x"98",
          1332 => x"98",
          1333 => x"98",
          1334 => x"98",
          1335 => x"98",
          1336 => x"0c",
          1337 => x"0b",
          1338 => x"71",
          1339 => x"04",
          1340 => x"98",
          1341 => x"98",
          1342 => x"c0",
          1343 => x"34",
          1344 => x"83",
          1345 => x"5c",
          1346 => x"ac",
          1347 => x"c0",
          1348 => x"34",
          1349 => x"88",
          1350 => x"5a",
          1351 => x"79",
          1352 => x"ff",
          1353 => x"85",
          1354 => x"83",
          1355 => x"7d",
          1356 => x"ec",
          1357 => x"0d",
          1358 => x"33",
          1359 => x"51",
          1360 => x"08",
          1361 => x"71",
          1362 => x"72",
          1363 => x"c8",
          1364 => x"80",
          1365 => x"98",
          1366 => x"ff",
          1367 => x"51",
          1368 => x"08",
          1369 => x"71",
          1370 => x"3d",
          1371 => x"2b",
          1372 => x"84",
          1373 => x"2c",
          1374 => x"73",
          1375 => x"73",
          1376 => x"0c",
          1377 => x"02",
          1378 => x"70",
          1379 => x"80",
          1380 => x"94",
          1381 => x"53",
          1382 => x"71",
          1383 => x"70",
          1384 => x"53",
          1385 => x"2a",
          1386 => x"81",
          1387 => x"52",
          1388 => x"94",
          1389 => x"b9",
          1390 => x"91",
          1391 => x"97",
          1392 => x"72",
          1393 => x"81",
          1394 => x"87",
          1395 => x"70",
          1396 => x"38",
          1397 => x"05",
          1398 => x"52",
          1399 => x"3d",
          1400 => x"80",
          1401 => x"77",
          1402 => x"f2",
          1403 => x"57",
          1404 => x"87",
          1405 => x"70",
          1406 => x"2e",
          1407 => x"06",
          1408 => x"32",
          1409 => x"38",
          1410 => x"cf",
          1411 => x"c0",
          1412 => x"38",
          1413 => x"0c",
          1414 => x"ff",
          1415 => x"88",
          1416 => x"81",
          1417 => x"81",
          1418 => x"c1",
          1419 => x"71",
          1420 => x"94",
          1421 => x"06",
          1422 => x"39",
          1423 => x"08",
          1424 => x"70",
          1425 => x"9e",
          1426 => x"c0",
          1427 => x"87",
          1428 => x"0c",
          1429 => x"90",
          1430 => x"f2",
          1431 => x"83",
          1432 => x"08",
          1433 => x"b0",
          1434 => x"9e",
          1435 => x"c0",
          1436 => x"87",
          1437 => x"0c",
          1438 => x"b0",
          1439 => x"f2",
          1440 => x"52",
          1441 => x"9e",
          1442 => x"c0",
          1443 => x"87",
          1444 => x"0c",
          1445 => x"0b",
          1446 => x"80",
          1447 => x"fb",
          1448 => x"0b",
          1449 => x"80",
          1450 => x"2e",
          1451 => x"ca",
          1452 => x"08",
          1453 => x"52",
          1454 => x"71",
          1455 => x"c0",
          1456 => x"06",
          1457 => x"38",
          1458 => x"80",
          1459 => x"a0",
          1460 => x"80",
          1461 => x"f2",
          1462 => x"90",
          1463 => x"52",
          1464 => x"52",
          1465 => x"87",
          1466 => x"80",
          1467 => x"83",
          1468 => x"34",
          1469 => x"70",
          1470 => x"70",
          1471 => x"83",
          1472 => x"9e",
          1473 => x"51",
          1474 => x"81",
          1475 => x"0b",
          1476 => x"c0",
          1477 => x"2e",
          1478 => x"d2",
          1479 => x"08",
          1480 => x"70",
          1481 => x"83",
          1482 => x"08",
          1483 => x"51",
          1484 => x"87",
          1485 => x"06",
          1486 => x"38",
          1487 => x"87",
          1488 => x"70",
          1489 => x"d6",
          1490 => x"08",
          1491 => x"80",
          1492 => x"f2",
          1493 => x"87",
          1494 => x"83",
          1495 => x"39",
          1496 => x"ff",
          1497 => x"54",
          1498 => x"51",
          1499 => x"55",
          1500 => x"33",
          1501 => x"cc",
          1502 => x"f2",
          1503 => x"83",
          1504 => x"38",
          1505 => x"a8",
          1506 => x"84",
          1507 => x"74",
          1508 => x"56",
          1509 => x"33",
          1510 => x"d0",
          1511 => x"f2",
          1512 => x"83",
          1513 => x"38",
          1514 => x"83",
          1515 => x"51",
          1516 => x"08",
          1517 => x"9d",
          1518 => x"da",
          1519 => x"da",
          1520 => x"b8",
          1521 => x"b4",
          1522 => x"bd",
          1523 => x"3f",
          1524 => x"29",
          1525 => x"c8",
          1526 => x"b4",
          1527 => x"74",
          1528 => x"74",
          1529 => x"f2",
          1530 => x"75",
          1531 => x"08",
          1532 => x"54",
          1533 => x"db",
          1534 => x"3d",
          1535 => x"bd",
          1536 => x"3f",
          1537 => x"29",
          1538 => x"c8",
          1539 => x"b3",
          1540 => x"74",
          1541 => x"39",
          1542 => x"83",
          1543 => x"f2",
          1544 => x"ff",
          1545 => x"52",
          1546 => x"3f",
          1547 => x"8c",
          1548 => x"b4",
          1549 => x"22",
          1550 => x"95",
          1551 => x"84",
          1552 => x"84",
          1553 => x"76",
          1554 => x"08",
          1555 => x"ed",
          1556 => x"80",
          1557 => x"83",
          1558 => x"83",
          1559 => x"fd",
          1560 => x"f8",
          1561 => x"d1",
          1562 => x"38",
          1563 => x"bf",
          1564 => x"74",
          1565 => x"83",
          1566 => x"83",
          1567 => x"fc",
          1568 => x"33",
          1569 => x"fd",
          1570 => x"80",
          1571 => x"f2",
          1572 => x"ff",
          1573 => x"55",
          1574 => x"39",
          1575 => x"e4",
          1576 => x"d7",
          1577 => x"38",
          1578 => x"f2",
          1579 => x"84",
          1580 => x"d3",
          1581 => x"38",
          1582 => x"f2",
          1583 => x"a0",
          1584 => x"ce",
          1585 => x"38",
          1586 => x"f2",
          1587 => x"bc",
          1588 => x"cd",
          1589 => x"38",
          1590 => x"f2",
          1591 => x"d8",
          1592 => x"cc",
          1593 => x"38",
          1594 => x"f2",
          1595 => x"f4",
          1596 => x"cf",
          1597 => x"38",
          1598 => x"b0",
          1599 => x"bc",
          1600 => x"74",
          1601 => x"ff",
          1602 => x"71",
          1603 => x"83",
          1604 => x"83",
          1605 => x"83",
          1606 => x"ff",
          1607 => x"83",
          1608 => x"83",
          1609 => x"ff",
          1610 => x"83",
          1611 => x"83",
          1612 => x"ff",
          1613 => x"71",
          1614 => x"c0",
          1615 => x"08",
          1616 => x"3d",
          1617 => x"5a",
          1618 => x"83",
          1619 => x"3f",
          1620 => x"8b",
          1621 => x"08",
          1622 => x"82",
          1623 => x"80",
          1624 => x"3f",
          1625 => x"55",
          1626 => x"8e",
          1627 => x"70",
          1628 => x"09",
          1629 => x"51",
          1630 => x"73",
          1631 => x"8c",
          1632 => x"3f",
          1633 => x"76",
          1634 => x"0c",
          1635 => x"51",
          1636 => x"09",
          1637 => x"51",
          1638 => x"f5",
          1639 => x"c8",
          1640 => x"a8",
          1641 => x"84",
          1642 => x"d8",
          1643 => x"08",
          1644 => x"5a",
          1645 => x"80",
          1646 => x"10",
          1647 => x"52",
          1648 => x"c8",
          1649 => x"c0",
          1650 => x"38",
          1651 => x"81",
          1652 => x"81",
          1653 => x"82",
          1654 => x"84",
          1655 => x"81",
          1656 => x"53",
          1657 => x"84",
          1658 => x"ff",
          1659 => x"a6",
          1660 => x"06",
          1661 => x"16",
          1662 => x"76",
          1663 => x"78",
          1664 => x"fe",
          1665 => x"33",
          1666 => x"06",
          1667 => x"38",
          1668 => x"cd",
          1669 => x"83",
          1670 => x"ea",
          1671 => x"38",
          1672 => x"52",
          1673 => x"b9",
          1674 => x"51",
          1675 => x"08",
          1676 => x"25",
          1677 => x"05",
          1678 => x"77",
          1679 => x"f0",
          1680 => x"ff",
          1681 => x"81",
          1682 => x"0d",
          1683 => x"b7",
          1684 => x"5c",
          1685 => x"b8",
          1686 => x"74",
          1687 => x"56",
          1688 => x"77",
          1689 => x"77",
          1690 => x"77",
          1691 => x"b4",
          1692 => x"3f",
          1693 => x"98",
          1694 => x"38",
          1695 => x"33",
          1696 => x"d1",
          1697 => x"2c",
          1698 => x"83",
          1699 => x"33",
          1700 => x"58",
          1701 => x"80",
          1702 => x"38",
          1703 => x"0a",
          1704 => x"76",
          1705 => x"70",
          1706 => x"de",
          1707 => x"25",
          1708 => x"18",
          1709 => x"81",
          1710 => x"75",
          1711 => x"80",
          1712 => x"98",
          1713 => x"33",
          1714 => x"98",
          1715 => x"d4",
          1716 => x"5d",
          1717 => x"38",
          1718 => x"39",
          1719 => x"81",
          1720 => x"70",
          1721 => x"57",
          1722 => x"75",
          1723 => x"80",
          1724 => x"57",
          1725 => x"d0",
          1726 => x"78",
          1727 => x"2e",
          1728 => x"57",
          1729 => x"e7",
          1730 => x"57",
          1731 => x"84",
          1732 => x"7e",
          1733 => x"95",
          1734 => x"83",
          1735 => x"83",
          1736 => x"0b",
          1737 => x"d1",
          1738 => x"33",
          1739 => x"84",
          1740 => x"b6",
          1741 => x"05",
          1742 => x"eb",
          1743 => x"ff",
          1744 => x"55",
          1745 => x"d5",
          1746 => x"84",
          1747 => x"52",
          1748 => x"39",
          1749 => x"10",
          1750 => x"57",
          1751 => x"d1",
          1752 => x"88",
          1753 => x"74",
          1754 => x"08",
          1755 => x"84",
          1756 => x"b5",
          1757 => x"88",
          1758 => x"8c",
          1759 => x"8c",
          1760 => x"cc",
          1761 => x"75",
          1762 => x"7c",
          1763 => x"75",
          1764 => x"f2",
          1765 => x"75",
          1766 => x"80",
          1767 => x"b7",
          1768 => x"d1",
          1769 => x"ff",
          1770 => x"51",
          1771 => x"33",
          1772 => x"80",
          1773 => x"08",
          1774 => x"84",
          1775 => x"b3",
          1776 => x"88",
          1777 => x"8c",
          1778 => x"8c",
          1779 => x"39",
          1780 => x"06",
          1781 => x"75",
          1782 => x"ac",
          1783 => x"d1",
          1784 => x"55",
          1785 => x"33",
          1786 => x"33",
          1787 => x"83",
          1788 => x"15",
          1789 => x"16",
          1790 => x"3f",
          1791 => x"06",
          1792 => x"77",
          1793 => x"39",
          1794 => x"33",
          1795 => x"38",
          1796 => x"34",
          1797 => x"81",
          1798 => x"24",
          1799 => x"52",
          1800 => x"d1",
          1801 => x"2c",
          1802 => x"41",
          1803 => x"d5",
          1804 => x"8b",
          1805 => x"80",
          1806 => x"88",
          1807 => x"f8",
          1808 => x"88",
          1809 => x"80",
          1810 => x"98",
          1811 => x"5a",
          1812 => x"bb",
          1813 => x"78",
          1814 => x"33",
          1815 => x"80",
          1816 => x"98",
          1817 => x"55",
          1818 => x"16",
          1819 => x"d5",
          1820 => x"b1",
          1821 => x"81",
          1822 => x"d1",
          1823 => x"24",
          1824 => x"d1",
          1825 => x"d3",
          1826 => x"51",
          1827 => x"33",
          1828 => x"34",
          1829 => x"84",
          1830 => x"7f",
          1831 => x"51",
          1832 => x"52",
          1833 => x"c8",
          1834 => x"cf",
          1835 => x"80",
          1836 => x"33",
          1837 => x"70",
          1838 => x"38",
          1839 => x"f2",
          1840 => x"5b",
          1841 => x"08",
          1842 => x"10",
          1843 => x"57",
          1844 => x"f3",
          1845 => x"38",
          1846 => x"2e",
          1847 => x"8c",
          1848 => x"7b",
          1849 => x"04",
          1850 => x"2e",
          1851 => x"88",
          1852 => x"ac",
          1853 => x"3f",
          1854 => x"ff",
          1855 => x"ff",
          1856 => x"75",
          1857 => x"83",
          1858 => x"80",
          1859 => x"84",
          1860 => x"7c",
          1861 => x"d1",
          1862 => x"38",
          1863 => x"ff",
          1864 => x"52",
          1865 => x"d5",
          1866 => x"9b",
          1867 => x"5d",
          1868 => x"ff",
          1869 => x"f0",
          1870 => x"84",
          1871 => x"88",
          1872 => x"3d",
          1873 => x"81",
          1874 => x"f4",
          1875 => x"05",
          1876 => x"16",
          1877 => x"d5",
          1878 => x"bb",
          1879 => x"2b",
          1880 => x"5a",
          1881 => x"ef",
          1882 => x"51",
          1883 => x"33",
          1884 => x"d1",
          1885 => x"7a",
          1886 => x"08",
          1887 => x"74",
          1888 => x"05",
          1889 => x"5b",
          1890 => x"38",
          1891 => x"ff",
          1892 => x"29",
          1893 => x"84",
          1894 => x"75",
          1895 => x"7b",
          1896 => x"84",
          1897 => x"ff",
          1898 => x"29",
          1899 => x"84",
          1900 => x"61",
          1901 => x"81",
          1902 => x"08",
          1903 => x"3f",
          1904 => x"0a",
          1905 => x"33",
          1906 => x"a7",
          1907 => x"33",
          1908 => x"60",
          1909 => x"33",
          1910 => x"98",
          1911 => x"76",
          1912 => x"33",
          1913 => x"29",
          1914 => x"84",
          1915 => x"78",
          1916 => x"84",
          1917 => x"7c",
          1918 => x"84",
          1919 => x"8b",
          1920 => x"88",
          1921 => x"70",
          1922 => x"05",
          1923 => x"44",
          1924 => x"ef",
          1925 => x"78",
          1926 => x"7a",
          1927 => x"08",
          1928 => x"75",
          1929 => x"05",
          1930 => x"57",
          1931 => x"38",
          1932 => x"ff",
          1933 => x"29",
          1934 => x"84",
          1935 => x"76",
          1936 => x"83",
          1937 => x"f4",
          1938 => x"3f",
          1939 => x"34",
          1940 => x"81",
          1941 => x"ad",
          1942 => x"d1",
          1943 => x"f4",
          1944 => x"88",
          1945 => x"ac",
          1946 => x"3f",
          1947 => x"ff",
          1948 => x"ff",
          1949 => x"7a",
          1950 => x"51",
          1951 => x"08",
          1952 => x"08",
          1953 => x"34",
          1954 => x"84",
          1955 => x"33",
          1956 => x"81",
          1957 => x"70",
          1958 => x"57",
          1959 => x"d1",
          1960 => x"2c",
          1961 => x"58",
          1962 => x"e4",
          1963 => x"ee",
          1964 => x"56",
          1965 => x"16",
          1966 => x"f0",
          1967 => x"83",
          1968 => x"ee",
          1969 => x"3f",
          1970 => x"fe",
          1971 => x"93",
          1972 => x"39",
          1973 => x"77",
          1974 => x"75",
          1975 => x"39",
          1976 => x"b9",
          1977 => x"b9",
          1978 => x"53",
          1979 => x"3f",
          1980 => x"d1",
          1981 => x"2e",
          1982 => x"52",
          1983 => x"d5",
          1984 => x"eb",
          1985 => x"51",
          1986 => x"33",
          1987 => x"34",
          1988 => x"80",
          1989 => x"34",
          1990 => x"84",
          1991 => x"75",
          1992 => x"c8",
          1993 => x"c8",
          1994 => x"75",
          1995 => x"81",
          1996 => x"88",
          1997 => x"5e",
          1998 => x"84",
          1999 => x"a5",
          2000 => x"a0",
          2001 => x"ac",
          2002 => x"3f",
          2003 => x"76",
          2004 => x"06",
          2005 => x"fd",
          2006 => x"88",
          2007 => x"06",
          2008 => x"ff",
          2009 => x"ff",
          2010 => x"8c",
          2011 => x"2e",
          2012 => x"52",
          2013 => x"d5",
          2014 => x"fb",
          2015 => x"51",
          2016 => x"33",
          2017 => x"34",
          2018 => x"74",
          2019 => x"b8",
          2020 => x"83",
          2021 => x"52",
          2022 => x"b9",
          2023 => x"33",
          2024 => x"70",
          2025 => x"f4",
          2026 => x"51",
          2027 => x"33",
          2028 => x"56",
          2029 => x"83",
          2030 => x"3d",
          2031 => x"52",
          2032 => x"f3",
          2033 => x"88",
          2034 => x"df",
          2035 => x"34",
          2036 => x"84",
          2037 => x"93",
          2038 => x"51",
          2039 => x"08",
          2040 => x"96",
          2041 => x"53",
          2042 => x"f2",
          2043 => x"b9",
          2044 => x"e9",
          2045 => x"ff",
          2046 => x"56",
          2047 => x"80",
          2048 => x"05",
          2049 => x"75",
          2050 => x"70",
          2051 => x"08",
          2052 => x"38",
          2053 => x"f2",
          2054 => x"55",
          2055 => x"08",
          2056 => x"10",
          2057 => x"57",
          2058 => x"70",
          2059 => x"27",
          2060 => x"09",
          2061 => x"ed",
          2062 => x"52",
          2063 => x"f3",
          2064 => x"06",
          2065 => x"38",
          2066 => x"bd",
          2067 => x"83",
          2068 => x"fc",
          2069 => x"70",
          2070 => x"3f",
          2071 => x"f3",
          2072 => x"e0",
          2073 => x"80",
          2074 => x"76",
          2075 => x"75",
          2076 => x"83",
          2077 => x"77",
          2078 => x"3d",
          2079 => x"84",
          2080 => x"72",
          2081 => x"2e",
          2082 => x"9e",
          2083 => x"86",
          2084 => x"80",
          2085 => x"58",
          2086 => x"f8",
          2087 => x"75",
          2088 => x"33",
          2089 => x"71",
          2090 => x"56",
          2091 => x"38",
          2092 => x"74",
          2093 => x"74",
          2094 => x"38",
          2095 => x"17",
          2096 => x"0b",
          2097 => x"81",
          2098 => x"ee",
          2099 => x"a0",
          2100 => x"10",
          2101 => x"90",
          2102 => x"40",
          2103 => x"b7",
          2104 => x"b7",
          2105 => x"f8",
          2106 => x"70",
          2107 => x"57",
          2108 => x"72",
          2109 => x"ff",
          2110 => x"ff",
          2111 => x"81",
          2112 => x"42",
          2113 => x"8f",
          2114 => x"31",
          2115 => x"76",
          2116 => x"9c",
          2117 => x"26",
          2118 => x"05",
          2119 => x"70",
          2120 => x"a7",
          2121 => x"70",
          2122 => x"06",
          2123 => x"06",
          2124 => x"5d",
          2125 => x"74",
          2126 => x"ff",
          2127 => x"29",
          2128 => x"fd",
          2129 => x"34",
          2130 => x"f8",
          2131 => x"2b",
          2132 => x"7a",
          2133 => x"26",
          2134 => x"fc",
          2135 => x"81",
          2136 => x"f8",
          2137 => x"a7",
          2138 => x"56",
          2139 => x"84",
          2140 => x"84",
          2141 => x"83",
          2142 => x"06",
          2143 => x"41",
          2144 => x"73",
          2145 => x"70",
          2146 => x"ff",
          2147 => x"29",
          2148 => x"ff",
          2149 => x"5c",
          2150 => x"77",
          2151 => x"79",
          2152 => x"38",
          2153 => x"38",
          2154 => x"29",
          2155 => x"86",
          2156 => x"34",
          2157 => x"73",
          2158 => x"f4",
          2159 => x"ee",
          2160 => x"76",
          2161 => x"74",
          2162 => x"34",
          2163 => x"86",
          2164 => x"81",
          2165 => x"77",
          2166 => x"34",
          2167 => x"c0",
          2168 => x"a0",
          2169 => x"07",
          2170 => x"34",
          2171 => x"53",
          2172 => x"b7",
          2173 => x"0c",
          2174 => x"33",
          2175 => x"0d",
          2176 => x"b3",
          2177 => x"59",
          2178 => x"da",
          2179 => x"f9",
          2180 => x"29",
          2181 => x"f8",
          2182 => x"7c",
          2183 => x"83",
          2184 => x"72",
          2185 => x"f6",
          2186 => x"f6",
          2187 => x"70",
          2188 => x"55",
          2189 => x"38",
          2190 => x"34",
          2191 => x"ff",
          2192 => x"57",
          2193 => x"b7",
          2194 => x"80",
          2195 => x"84",
          2196 => x"e0",
          2197 => x"70",
          2198 => x"05",
          2199 => x"b9",
          2200 => x"26",
          2201 => x"98",
          2202 => x"e0",
          2203 => x"55",
          2204 => x"27",
          2205 => x"05",
          2206 => x"57",
          2207 => x"ff",
          2208 => x"fd",
          2209 => x"b7",
          2210 => x"57",
          2211 => x"86",
          2212 => x"75",
          2213 => x"5c",
          2214 => x"38",
          2215 => x"14",
          2216 => x"78",
          2217 => x"81",
          2218 => x"59",
          2219 => x"84",
          2220 => x"56",
          2221 => x"38",
          2222 => x"8b",
          2223 => x"34",
          2224 => x"ff",
          2225 => x"57",
          2226 => x"80",
          2227 => x"06",
          2228 => x"53",
          2229 => x"c8",
          2230 => x"b7",
          2231 => x"29",
          2232 => x"27",
          2233 => x"84",
          2234 => x"56",
          2235 => x"75",
          2236 => x"13",
          2237 => x"a0",
          2238 => x"70",
          2239 => x"72",
          2240 => x"84",
          2241 => x"39",
          2242 => x"b7",
          2243 => x"bb",
          2244 => x"0d",
          2245 => x"53",
          2246 => x"10",
          2247 => x"08",
          2248 => x"71",
          2249 => x"34",
          2250 => x"3d",
          2251 => x"34",
          2252 => x"06",
          2253 => x"ff",
          2254 => x"80",
          2255 => x"0d",
          2256 => x"31",
          2257 => x"54",
          2258 => x"34",
          2259 => x"05",
          2260 => x"56",
          2261 => x"53",
          2262 => x"84",
          2263 => x"83",
          2264 => x"09",
          2265 => x"53",
          2266 => x"0b",
          2267 => x"04",
          2268 => x"b7",
          2269 => x"70",
          2270 => x"83",
          2271 => x"c8",
          2272 => x"83",
          2273 => x"84",
          2274 => x"71",
          2275 => x"51",
          2276 => x"39",
          2277 => x"51",
          2278 => x"10",
          2279 => x"04",
          2280 => x"06",
          2281 => x"72",
          2282 => x"71",
          2283 => x"38",
          2284 => x"80",
          2285 => x"0d",
          2286 => x"06",
          2287 => x"34",
          2288 => x"3d",
          2289 => x"f0",
          2290 => x"e8",
          2291 => x"06",
          2292 => x"34",
          2293 => x"f4",
          2294 => x"83",
          2295 => x"81",
          2296 => x"f8",
          2297 => x"f4",
          2298 => x"f4",
          2299 => x"33",
          2300 => x"83",
          2301 => x"f8",
          2302 => x"51",
          2303 => x"39",
          2304 => x"81",
          2305 => x"fe",
          2306 => x"f8",
          2307 => x"fe",
          2308 => x"df",
          2309 => x"f8",
          2310 => x"f4",
          2311 => x"70",
          2312 => x"83",
          2313 => x"e0",
          2314 => x"fe",
          2315 => x"cf",
          2316 => x"f8",
          2317 => x"f4",
          2318 => x"70",
          2319 => x"83",
          2320 => x"70",
          2321 => x"83",
          2322 => x"07",
          2323 => x"e0",
          2324 => x"33",
          2325 => x"83",
          2326 => x"83",
          2327 => x"43",
          2328 => x"2e",
          2329 => x"38",
          2330 => x"84",
          2331 => x"c0",
          2332 => x"83",
          2333 => x"34",
          2334 => x"09",
          2335 => x"b7",
          2336 => x"34",
          2337 => x"0b",
          2338 => x"f8",
          2339 => x"33",
          2340 => x"b7",
          2341 => x"7a",
          2342 => x"d5",
          2343 => x"0b",
          2344 => x"f8",
          2345 => x"83",
          2346 => x"80",
          2347 => x"84",
          2348 => x"f8",
          2349 => x"80",
          2350 => x"cb",
          2351 => x"84",
          2352 => x"54",
          2353 => x"51",
          2354 => x"b8",
          2355 => x"a5",
          2356 => x"70",
          2357 => x"ff",
          2358 => x"ff",
          2359 => x"59",
          2360 => x"a4",
          2361 => x"b7",
          2362 => x"34",
          2363 => x"f8",
          2364 => x"8f",
          2365 => x"be",
          2366 => x"81",
          2367 => x"83",
          2368 => x"f6",
          2369 => x"9d",
          2370 => x"e3",
          2371 => x"59",
          2372 => x"3f",
          2373 => x"a6",
          2374 => x"83",
          2375 => x"81",
          2376 => x"d8",
          2377 => x"05",
          2378 => x"83",
          2379 => x"72",
          2380 => x"11",
          2381 => x"5c",
          2382 => x"ff",
          2383 => x"51",
          2384 => x"e9",
          2385 => x"75",
          2386 => x"2e",
          2387 => x"d5",
          2388 => x"f8",
          2389 => x"29",
          2390 => x"16",
          2391 => x"84",
          2392 => x"83",
          2393 => x"5a",
          2394 => x"18",
          2395 => x"29",
          2396 => x"86",
          2397 => x"bc",
          2398 => x"f6",
          2399 => x"29",
          2400 => x"f8",
          2401 => x"81",
          2402 => x"73",
          2403 => x"bd",
          2404 => x"17",
          2405 => x"b7",
          2406 => x"38",
          2407 => x"2e",
          2408 => x"c8",
          2409 => x"2e",
          2410 => x"38",
          2411 => x"c1",
          2412 => x"3f",
          2413 => x"be",
          2414 => x"84",
          2415 => x"89",
          2416 => x"80",
          2417 => x"3f",
          2418 => x"54",
          2419 => x"52",
          2420 => x"70",
          2421 => x"27",
          2422 => x"f8",
          2423 => x"83",
          2424 => x"b9",
          2425 => x"80",
          2426 => x"38",
          2427 => x"06",
          2428 => x"73",
          2429 => x"52",
          2430 => x"f9",
          2431 => x"05",
          2432 => x"72",
          2433 => x"80",
          2434 => x"81",
          2435 => x"80",
          2436 => x"86",
          2437 => x"05",
          2438 => x"75",
          2439 => x"2e",
          2440 => x"b5",
          2441 => x"78",
          2442 => x"2e",
          2443 => x"83",
          2444 => x"72",
          2445 => x"b7",
          2446 => x"17",
          2447 => x"f9",
          2448 => x"29",
          2449 => x"f8",
          2450 => x"60",
          2451 => x"f8",
          2452 => x"05",
          2453 => x"ff",
          2454 => x"f9",
          2455 => x"5d",
          2456 => x"98",
          2457 => x"ff",
          2458 => x"b8",
          2459 => x"86",
          2460 => x"f8",
          2461 => x"0c",
          2462 => x"84",
          2463 => x"38",
          2464 => x"80",
          2465 => x"84",
          2466 => x"83",
          2467 => x"72",
          2468 => x"b7",
          2469 => x"1d",
          2470 => x"f9",
          2471 => x"29",
          2472 => x"f8",
          2473 => x"76",
          2474 => x"f4",
          2475 => x"84",
          2476 => x"83",
          2477 => x"72",
          2478 => x"59",
          2479 => x"9a",
          2480 => x"ff",
          2481 => x"38",
          2482 => x"84",
          2483 => x"78",
          2484 => x"24",
          2485 => x"81",
          2486 => x"f8",
          2487 => x"0c",
          2488 => x"82",
          2489 => x"26",
          2490 => x"81",
          2491 => x"34",
          2492 => x"81",
          2493 => x"cc",
          2494 => x"0c",
          2495 => x"fd",
          2496 => x"0c",
          2497 => x"33",
          2498 => x"05",
          2499 => x"33",
          2500 => x"b7",
          2501 => x"f8",
          2502 => x"5f",
          2503 => x"34",
          2504 => x"19",
          2505 => x"a7",
          2506 => x"33",
          2507 => x"22",
          2508 => x"11",
          2509 => x"f4",
          2510 => x"81",
          2511 => x"81",
          2512 => x"f8",
          2513 => x"bc",
          2514 => x"ff",
          2515 => x"29",
          2516 => x"f8",
          2517 => x"29",
          2518 => x"f7",
          2519 => x"75",
          2520 => x"ff",
          2521 => x"95",
          2522 => x"34",
          2523 => x"c8",
          2524 => x"80",
          2525 => x"84",
          2526 => x"c4",
          2527 => x"9c",
          2528 => x"84",
          2529 => x"84",
          2530 => x"84",
          2531 => x"c4",
          2532 => x"9c",
          2533 => x"09",
          2534 => x"f8",
          2535 => x"ff",
          2536 => x"ff",
          2537 => x"a0",
          2538 => x"40",
          2539 => x"ff",
          2540 => x"43",
          2541 => x"85",
          2542 => x"1a",
          2543 => x"76",
          2544 => x"06",
          2545 => x"06",
          2546 => x"84",
          2547 => x"1e",
          2548 => x"f9",
          2549 => x"29",
          2550 => x"83",
          2551 => x"33",
          2552 => x"83",
          2553 => x"1a",
          2554 => x"ff",
          2555 => x"f9",
          2556 => x"5a",
          2557 => x"84",
          2558 => x"81",
          2559 => x"95",
          2560 => x"79",
          2561 => x"83",
          2562 => x"70",
          2563 => x"fd",
          2564 => x"38",
          2565 => x"bf",
          2566 => x"33",
          2567 => x"19",
          2568 => x"75",
          2569 => x"77",
          2570 => x"34",
          2571 => x"80",
          2572 => x"0d",
          2573 => x"bc",
          2574 => x"f9",
          2575 => x"29",
          2576 => x"f8",
          2577 => x"05",
          2578 => x"ce",
          2579 => x"5b",
          2580 => x"5c",
          2581 => x"06",
          2582 => x"05",
          2583 => x"86",
          2584 => x"bc",
          2585 => x"f6",
          2586 => x"5e",
          2587 => x"34",
          2588 => x"1e",
          2589 => x"a7",
          2590 => x"33",
          2591 => x"22",
          2592 => x"11",
          2593 => x"f4",
          2594 => x"81",
          2595 => x"7e",
          2596 => x"bd",
          2597 => x"19",
          2598 => x"1c",
          2599 => x"83",
          2600 => x"33",
          2601 => x"33",
          2602 => x"06",
          2603 => x"05",
          2604 => x"b7",
          2605 => x"34",
          2606 => x"33",
          2607 => x"12",
          2608 => x"f8",
          2609 => x"76",
          2610 => x"f4",
          2611 => x"84",
          2612 => x"83",
          2613 => x"72",
          2614 => x"59",
          2615 => x"18",
          2616 => x"06",
          2617 => x"38",
          2618 => x"39",
          2619 => x"0b",
          2620 => x"04",
          2621 => x"b7",
          2622 => x"f9",
          2623 => x"05",
          2624 => x"b8",
          2625 => x"0c",
          2626 => x"17",
          2627 => x"7c",
          2628 => x"bc",
          2629 => x"5b",
          2630 => x"cc",
          2631 => x"05",
          2632 => x"c8",
          2633 => x"b8",
          2634 => x"84",
          2635 => x"06",
          2636 => x"84",
          2637 => x"83",
          2638 => x"c4",
          2639 => x"33",
          2640 => x"33",
          2641 => x"b7",
          2642 => x"f8",
          2643 => x"5d",
          2644 => x"86",
          2645 => x"bc",
          2646 => x"f6",
          2647 => x"5b",
          2648 => x"83",
          2649 => x"41",
          2650 => x"a7",
          2651 => x"33",
          2652 => x"22",
          2653 => x"11",
          2654 => x"f4",
          2655 => x"1c",
          2656 => x"7b",
          2657 => x"33",
          2658 => x"56",
          2659 => x"84",
          2660 => x"40",
          2661 => x"b7",
          2662 => x"78",
          2663 => x"0b",
          2664 => x"04",
          2665 => x"34",
          2666 => x"34",
          2667 => x"f8",
          2668 => x"f8",
          2669 => x"f9",
          2670 => x"f7",
          2671 => x"39",
          2672 => x"2e",
          2673 => x"5d",
          2674 => x"85",
          2675 => x"55",
          2676 => x"9b",
          2677 => x"70",
          2678 => x"51",
          2679 => x"08",
          2680 => x"57",
          2681 => x"cd",
          2682 => x"fe",
          2683 => x"0b",
          2684 => x"81",
          2685 => x"ad",
          2686 => x"81",
          2687 => x"8a",
          2688 => x"a4",
          2689 => x"c9",
          2690 => x"38",
          2691 => x"33",
          2692 => x"2c",
          2693 => x"75",
          2694 => x"84",
          2695 => x"8e",
          2696 => x"05",
          2697 => x"33",
          2698 => x"c5",
          2699 => x"bd",
          2700 => x"83",
          2701 => x"5d",
          2702 => x"ff",
          2703 => x"fd",
          2704 => x"34",
          2705 => x"33",
          2706 => x"fd",
          2707 => x"f8",
          2708 => x"c9",
          2709 => x"38",
          2710 => x"33",
          2711 => x"2c",
          2712 => x"75",
          2713 => x"84",
          2714 => x"fc",
          2715 => x"60",
          2716 => x"38",
          2717 => x"33",
          2718 => x"12",
          2719 => x"f6",
          2720 => x"29",
          2721 => x"f7",
          2722 => x"42",
          2723 => x"2e",
          2724 => x"cd",
          2725 => x"33",
          2726 => x"84",
          2727 => x"09",
          2728 => x"83",
          2729 => x"b8",
          2730 => x"be",
          2731 => x"f9",
          2732 => x"33",
          2733 => x"25",
          2734 => x"f9",
          2735 => x"33",
          2736 => x"84",
          2737 => x"42",
          2738 => x"11",
          2739 => x"38",
          2740 => x"fa",
          2741 => x"e8",
          2742 => x"33",
          2743 => x"38",
          2744 => x"22",
          2745 => x"e8",
          2746 => x"06",
          2747 => x"da",
          2748 => x"5f",
          2749 => x"b9",
          2750 => x"38",
          2751 => x"06",
          2752 => x"84",
          2753 => x"8e",
          2754 => x"05",
          2755 => x"33",
          2756 => x"b7",
          2757 => x"11",
          2758 => x"77",
          2759 => x"83",
          2760 => x"ff",
          2761 => x"38",
          2762 => x"84",
          2763 => x"7a",
          2764 => x"75",
          2765 => x"84",
          2766 => x"8a",
          2767 => x"b7",
          2768 => x"f9",
          2769 => x"b7",
          2770 => x"f8",
          2771 => x"a7",
          2772 => x"5f",
          2773 => x"ff",
          2774 => x"52",
          2775 => x"84",
          2776 => x"70",
          2777 => x"8e",
          2778 => x"76",
          2779 => x"56",
          2780 => x"ff",
          2781 => x"60",
          2782 => x"33",
          2783 => x"ff",
          2784 => x"7e",
          2785 => x"57",
          2786 => x"38",
          2787 => x"ff",
          2788 => x"79",
          2789 => x"a7",
          2790 => x"81",
          2791 => x"58",
          2792 => x"38",
          2793 => x"17",
          2794 => x"7b",
          2795 => x"81",
          2796 => x"5e",
          2797 => x"84",
          2798 => x"43",
          2799 => x"9d",
          2800 => x"b7",
          2801 => x"5d",
          2802 => x"7c",
          2803 => x"84",
          2804 => x"71",
          2805 => x"7f",
          2806 => x"39",
          2807 => x"2e",
          2808 => x"9d",
          2809 => x"39",
          2810 => x"11",
          2811 => x"58",
          2812 => x"9c",
          2813 => x"06",
          2814 => x"58",
          2815 => x"33",
          2816 => x"81",
          2817 => x"7a",
          2818 => x"ff",
          2819 => x"38",
          2820 => x"57",
          2821 => x"1b",
          2822 => x"a0",
          2823 => x"a7",
          2824 => x"51",
          2825 => x"06",
          2826 => x"f4",
          2827 => x"07",
          2828 => x"7f",
          2829 => x"9e",
          2830 => x"0c",
          2831 => x"79",
          2832 => x"33",
          2833 => x"81",
          2834 => x"f8",
          2835 => x"59",
          2836 => x"38",
          2837 => x"62",
          2838 => x"57",
          2839 => x"f8",
          2840 => x"5a",
          2841 => x"78",
          2842 => x"57",
          2843 => x"0b",
          2844 => x"81",
          2845 => x"77",
          2846 => x"1f",
          2847 => x"8a",
          2848 => x"f0",
          2849 => x"71",
          2850 => x"80",
          2851 => x"80",
          2852 => x"18",
          2853 => x"b6",
          2854 => x"84",
          2855 => x"f8",
          2856 => x"f8",
          2857 => x"5c",
          2858 => x"f4",
          2859 => x"f4",
          2860 => x"59",
          2861 => x"33",
          2862 => x"83",
          2863 => x"f4",
          2864 => x"75",
          2865 => x"f8",
          2866 => x"56",
          2867 => x"83",
          2868 => x"07",
          2869 => x"b1",
          2870 => x"34",
          2871 => x"56",
          2872 => x"81",
          2873 => x"34",
          2874 => x"81",
          2875 => x"f8",
          2876 => x"f4",
          2877 => x"56",
          2878 => x"39",
          2879 => x"80",
          2880 => x"34",
          2881 => x"81",
          2882 => x"f8",
          2883 => x"f4",
          2884 => x"75",
          2885 => x"83",
          2886 => x"07",
          2887 => x"a1",
          2888 => x"06",
          2889 => x"34",
          2890 => x"81",
          2891 => x"34",
          2892 => x"80",
          2893 => x"34",
          2894 => x"80",
          2895 => x"34",
          2896 => x"81",
          2897 => x"83",
          2898 => x"f8",
          2899 => x"56",
          2900 => x"39",
          2901 => x"52",
          2902 => x"39",
          2903 => x"34",
          2904 => x"34",
          2905 => x"f8",
          2906 => x"0c",
          2907 => x"cb",
          2908 => x"9c",
          2909 => x"34",
          2910 => x"06",
          2911 => x"84",
          2912 => x"53",
          2913 => x"84",
          2914 => x"c8",
          2915 => x"84",
          2916 => x"c8",
          2917 => x"f8",
          2918 => x"c9",
          2919 => x"b8",
          2920 => x"5d",
          2921 => x"9c",
          2922 => x"34",
          2923 => x"34",
          2924 => x"83",
          2925 => x"58",
          2926 => x"0b",
          2927 => x"51",
          2928 => x"51",
          2929 => x"83",
          2930 => x"70",
          2931 => x"f2",
          2932 => x"39",
          2933 => x"27",
          2934 => x"34",
          2935 => x"ff",
          2936 => x"06",
          2937 => x"f8",
          2938 => x"33",
          2939 => x"25",
          2940 => x"39",
          2941 => x"06",
          2942 => x"38",
          2943 => x"33",
          2944 => x"33",
          2945 => x"80",
          2946 => x"71",
          2947 => x"06",
          2948 => x"42",
          2949 => x"38",
          2950 => x"5c",
          2951 => x"84",
          2952 => x"83",
          2953 => x"f8",
          2954 => x"11",
          2955 => x"38",
          2956 => x"27",
          2957 => x"83",
          2958 => x"83",
          2959 => x"76",
          2960 => x"81",
          2961 => x"29",
          2962 => x"a0",
          2963 => x"81",
          2964 => x"71",
          2965 => x"7e",
          2966 => x"1a",
          2967 => x"b7",
          2968 => x"5d",
          2969 => x"7d",
          2970 => x"84",
          2971 => x"71",
          2972 => x"77",
          2973 => x"17",
          2974 => x"7b",
          2975 => x"81",
          2976 => x"5f",
          2977 => x"84",
          2978 => x"59",
          2979 => x"99",
          2980 => x"17",
          2981 => x"7b",
          2982 => x"bc",
          2983 => x"bb",
          2984 => x"39",
          2985 => x"33",
          2986 => x"42",
          2987 => x"5a",
          2988 => x"ff",
          2989 => x"27",
          2990 => x"f8",
          2991 => x"ff",
          2992 => x"78",
          2993 => x"83",
          2994 => x"f8",
          2995 => x"33",
          2996 => x"25",
          2997 => x"39",
          2998 => x"c0",
          2999 => x"ff",
          3000 => x"5d",
          3001 => x"06",
          3002 => x"1d",
          3003 => x"93",
          3004 => x"f6",
          3005 => x"56",
          3006 => x"39",
          3007 => x"f5",
          3008 => x"58",
          3009 => x"81",
          3010 => x"ec",
          3011 => x"34",
          3012 => x"05",
          3013 => x"f4",
          3014 => x"83",
          3015 => x"0b",
          3016 => x"7e",
          3017 => x"80",
          3018 => x"39",
          3019 => x"a7",
          3020 => x"84",
          3021 => x"0b",
          3022 => x"fd",
          3023 => x"b7",
          3024 => x"90",
          3025 => x"0b",
          3026 => x"04",
          3027 => x"80",
          3028 => x"0d",
          3029 => x"33",
          3030 => x"70",
          3031 => x"33",
          3032 => x"80",
          3033 => x"f7",
          3034 => x"c8",
          3035 => x"a8",
          3036 => x"91",
          3037 => x"07",
          3038 => x"5e",
          3039 => x"59",
          3040 => x"06",
          3041 => x"70",
          3042 => x"5c",
          3043 => x"84",
          3044 => x"83",
          3045 => x"86",
          3046 => x"22",
          3047 => x"70",
          3048 => x"33",
          3049 => x"83",
          3050 => x"ee",
          3051 => x"98",
          3052 => x"56",
          3053 => x"80",
          3054 => x"15",
          3055 => x"55",
          3056 => x"80",
          3057 => x"81",
          3058 => x"58",
          3059 => x"38",
          3060 => x"74",
          3061 => x"ff",
          3062 => x"cd",
          3063 => x"83",
          3064 => x"15",
          3065 => x"55",
          3066 => x"83",
          3067 => x"80",
          3068 => x"a0",
          3069 => x"2a",
          3070 => x"58",
          3071 => x"0b",
          3072 => x"06",
          3073 => x"81",
          3074 => x"83",
          3075 => x"83",
          3076 => x"33",
          3077 => x"5e",
          3078 => x"33",
          3079 => x"83",
          3080 => x"2e",
          3081 => x"33",
          3082 => x"83",
          3083 => x"ec",
          3084 => x"81",
          3085 => x"16",
          3086 => x"38",
          3087 => x"ff",
          3088 => x"16",
          3089 => x"38",
          3090 => x"87",
          3091 => x"73",
          3092 => x"c0",
          3093 => x"58",
          3094 => x"54",
          3095 => x"83",
          3096 => x"34",
          3097 => x"82",
          3098 => x"ec",
          3099 => x"d0",
          3100 => x"83",
          3101 => x"5e",
          3102 => x"80",
          3103 => x"72",
          3104 => x"83",
          3105 => x"08",
          3106 => x"06",
          3107 => x"f8",
          3108 => x"14",
          3109 => x"a5",
          3110 => x"80",
          3111 => x"83",
          3112 => x"f0",
          3113 => x"e0",
          3114 => x"7c",
          3115 => x"09",
          3116 => x"2e",
          3117 => x"d7",
          3118 => x"77",
          3119 => x"80",
          3120 => x"38",
          3121 => x"10",
          3122 => x"98",
          3123 => x"73",
          3124 => x"79",
          3125 => x"05",
          3126 => x"56",
          3127 => x"83",
          3128 => x"80",
          3129 => x"79",
          3130 => x"82",
          3131 => x"fa",
          3132 => x"33",
          3133 => x"38",
          3134 => x"25",
          3135 => x"38",
          3136 => x"cc",
          3137 => x"80",
          3138 => x"d4",
          3139 => x"2e",
          3140 => x"ff",
          3141 => x"38",
          3142 => x"2e",
          3143 => x"55",
          3144 => x"06",
          3145 => x"84",
          3146 => x"be",
          3147 => x"39",
          3148 => x"f7",
          3149 => x"83",
          3150 => x"80",
          3151 => x"0b",
          3152 => x"83",
          3153 => x"74",
          3154 => x"2e",
          3155 => x"33",
          3156 => x"77",
          3157 => x"09",
          3158 => x"9c",
          3159 => x"9c",
          3160 => x"e8",
          3161 => x"f7",
          3162 => x"fb",
          3163 => x"15",
          3164 => x"a1",
          3165 => x"fa",
          3166 => x"80",
          3167 => x"a8",
          3168 => x"f7",
          3169 => x"5d",
          3170 => x"39",
          3171 => x"cb",
          3172 => x"ce",
          3173 => x"fc",
          3174 => x"34",
          3175 => x"0b",
          3176 => x"83",
          3177 => x"34",
          3178 => x"84",
          3179 => x"38",
          3180 => x"ff",
          3181 => x"f7",
          3182 => x"84",
          3183 => x"39",
          3184 => x"06",
          3185 => x"27",
          3186 => x"f6",
          3187 => x"55",
          3188 => x"54",
          3189 => x"bc",
          3190 => x"05",
          3191 => x"53",
          3192 => x"f6",
          3193 => x"ba",
          3194 => x"72",
          3195 => x"52",
          3196 => x"3f",
          3197 => x"f7",
          3198 => x"3d",
          3199 => x"3d",
          3200 => x"83",
          3201 => x"05",
          3202 => x"08",
          3203 => x"83",
          3204 => x"81",
          3205 => x"e8",
          3206 => x"f3",
          3207 => x"53",
          3208 => x"c0",
          3209 => x"f6",
          3210 => x"9c",
          3211 => x"38",
          3212 => x"c0",
          3213 => x"73",
          3214 => x"ff",
          3215 => x"9c",
          3216 => x"c0",
          3217 => x"9c",
          3218 => x"81",
          3219 => x"52",
          3220 => x"81",
          3221 => x"a4",
          3222 => x"ff",
          3223 => x"ff",
          3224 => x"38",
          3225 => x"d5",
          3226 => x"84",
          3227 => x"81",
          3228 => x"0d",
          3229 => x"05",
          3230 => x"83",
          3231 => x"fc",
          3232 => x"07",
          3233 => x"34",
          3234 => x"34",
          3235 => x"34",
          3236 => x"08",
          3237 => x"d4",
          3238 => x"0b",
          3239 => x"0b",
          3240 => x"80",
          3241 => x"83",
          3242 => x"05",
          3243 => x"87",
          3244 => x"2e",
          3245 => x"98",
          3246 => x"87",
          3247 => x"87",
          3248 => x"70",
          3249 => x"71",
          3250 => x"98",
          3251 => x"87",
          3252 => x"98",
          3253 => x"38",
          3254 => x"08",
          3255 => x"71",
          3256 => x"98",
          3257 => x"38",
          3258 => x"81",
          3259 => x"80",
          3260 => x"71",
          3261 => x"ff",
          3262 => x"14",
          3263 => x"70",
          3264 => x"05",
          3265 => x"34",
          3266 => x"b9",
          3267 => x"0b",
          3268 => x"04",
          3269 => x"79",
          3270 => x"56",
          3271 => x"88",
          3272 => x"79",
          3273 => x"75",
          3274 => x"70",
          3275 => x"71",
          3276 => x"7a",
          3277 => x"84",
          3278 => x"73",
          3279 => x"52",
          3280 => x"72",
          3281 => x"08",
          3282 => x"d4",
          3283 => x"0b",
          3284 => x"0b",
          3285 => x"80",
          3286 => x"83",
          3287 => x"05",
          3288 => x"87",
          3289 => x"2e",
          3290 => x"98",
          3291 => x"87",
          3292 => x"87",
          3293 => x"70",
          3294 => x"71",
          3295 => x"98",
          3296 => x"87",
          3297 => x"98",
          3298 => x"38",
          3299 => x"08",
          3300 => x"71",
          3301 => x"98",
          3302 => x"38",
          3303 => x"81",
          3304 => x"a1",
          3305 => x"fe",
          3306 => x"06",
          3307 => x"57",
          3308 => x"0d",
          3309 => x"0d",
          3310 => x"71",
          3311 => x"56",
          3312 => x"0b",
          3313 => x"98",
          3314 => x"80",
          3315 => x"9c",
          3316 => x"53",
          3317 => x"33",
          3318 => x"70",
          3319 => x"2e",
          3320 => x"51",
          3321 => x"38",
          3322 => x"38",
          3323 => x"90",
          3324 => x"52",
          3325 => x"72",
          3326 => x"c0",
          3327 => x"27",
          3328 => x"38",
          3329 => x"71",
          3330 => x"ff",
          3331 => x"75",
          3332 => x"06",
          3333 => x"80",
          3334 => x"d0",
          3335 => x"3d",
          3336 => x"31",
          3337 => x"70",
          3338 => x"12",
          3339 => x"07",
          3340 => x"71",
          3341 => x"54",
          3342 => x"56",
          3343 => x"38",
          3344 => x"33",
          3345 => x"76",
          3346 => x"98",
          3347 => x"5c",
          3348 => x"83",
          3349 => x"33",
          3350 => x"75",
          3351 => x"57",
          3352 => x"06",
          3353 => x"b8",
          3354 => x"13",
          3355 => x"2a",
          3356 => x"14",
          3357 => x"b8",
          3358 => x"34",
          3359 => x"b8",
          3360 => x"85",
          3361 => x"70",
          3362 => x"07",
          3363 => x"58",
          3364 => x"81",
          3365 => x"12",
          3366 => x"71",
          3367 => x"33",
          3368 => x"70",
          3369 => x"58",
          3370 => x"12",
          3371 => x"84",
          3372 => x"2b",
          3373 => x"52",
          3374 => x"33",
          3375 => x"52",
          3376 => x"72",
          3377 => x"15",
          3378 => x"2b",
          3379 => x"2a",
          3380 => x"77",
          3381 => x"70",
          3382 => x"8b",
          3383 => x"70",
          3384 => x"07",
          3385 => x"77",
          3386 => x"54",
          3387 => x"14",
          3388 => x"b8",
          3389 => x"33",
          3390 => x"74",
          3391 => x"88",
          3392 => x"88",
          3393 => x"54",
          3394 => x"34",
          3395 => x"11",
          3396 => x"71",
          3397 => x"81",
          3398 => x"2b",
          3399 => x"53",
          3400 => x"71",
          3401 => x"07",
          3402 => x"59",
          3403 => x"16",
          3404 => x"70",
          3405 => x"71",
          3406 => x"33",
          3407 => x"70",
          3408 => x"56",
          3409 => x"83",
          3410 => x"3d",
          3411 => x"58",
          3412 => x"2e",
          3413 => x"89",
          3414 => x"84",
          3415 => x"b9",
          3416 => x"52",
          3417 => x"3f",
          3418 => x"34",
          3419 => x"b8",
          3420 => x"0b",
          3421 => x"56",
          3422 => x"17",
          3423 => x"b4",
          3424 => x"70",
          3425 => x"58",
          3426 => x"73",
          3427 => x"70",
          3428 => x"05",
          3429 => x"34",
          3430 => x"39",
          3431 => x"81",
          3432 => x"12",
          3433 => x"ff",
          3434 => x"06",
          3435 => x"85",
          3436 => x"52",
          3437 => x"54",
          3438 => x"10",
          3439 => x"33",
          3440 => x"ff",
          3441 => x"06",
          3442 => x"54",
          3443 => x"80",
          3444 => x"84",
          3445 => x"2b",
          3446 => x"81",
          3447 => x"54",
          3448 => x"70",
          3449 => x"07",
          3450 => x"5d",
          3451 => x"38",
          3452 => x"82",
          3453 => x"82",
          3454 => x"38",
          3455 => x"74",
          3456 => x"5b",
          3457 => x"78",
          3458 => x"15",
          3459 => x"14",
          3460 => x"b8",
          3461 => x"33",
          3462 => x"8f",
          3463 => x"ff",
          3464 => x"53",
          3465 => x"34",
          3466 => x"12",
          3467 => x"75",
          3468 => x"b9",
          3469 => x"87",
          3470 => x"2b",
          3471 => x"57",
          3472 => x"34",
          3473 => x"78",
          3474 => x"71",
          3475 => x"54",
          3476 => x"87",
          3477 => x"19",
          3478 => x"8b",
          3479 => x"58",
          3480 => x"34",
          3481 => x"08",
          3482 => x"33",
          3483 => x"70",
          3484 => x"84",
          3485 => x"b9",
          3486 => x"84",
          3487 => x"86",
          3488 => x"2b",
          3489 => x"17",
          3490 => x"07",
          3491 => x"54",
          3492 => x"12",
          3493 => x"84",
          3494 => x"2b",
          3495 => x"14",
          3496 => x"07",
          3497 => x"56",
          3498 => x"76",
          3499 => x"18",
          3500 => x"2b",
          3501 => x"2a",
          3502 => x"74",
          3503 => x"18",
          3504 => x"3d",
          3505 => x"58",
          3506 => x"77",
          3507 => x"89",
          3508 => x"3f",
          3509 => x"0c",
          3510 => x"0b",
          3511 => x"84",
          3512 => x"76",
          3513 => x"b4",
          3514 => x"75",
          3515 => x"b9",
          3516 => x"81",
          3517 => x"08",
          3518 => x"87",
          3519 => x"b9",
          3520 => x"07",
          3521 => x"2a",
          3522 => x"34",
          3523 => x"22",
          3524 => x"08",
          3525 => x"15",
          3526 => x"54",
          3527 => x"e3",
          3528 => x"5f",
          3529 => x"45",
          3530 => x"7e",
          3531 => x"2e",
          3532 => x"27",
          3533 => x"82",
          3534 => x"58",
          3535 => x"31",
          3536 => x"70",
          3537 => x"12",
          3538 => x"31",
          3539 => x"10",
          3540 => x"11",
          3541 => x"2b",
          3542 => x"53",
          3543 => x"44",
          3544 => x"80",
          3545 => x"33",
          3546 => x"70",
          3547 => x"12",
          3548 => x"07",
          3549 => x"74",
          3550 => x"82",
          3551 => x"2e",
          3552 => x"f9",
          3553 => x"87",
          3554 => x"24",
          3555 => x"81",
          3556 => x"2b",
          3557 => x"33",
          3558 => x"47",
          3559 => x"80",
          3560 => x"82",
          3561 => x"2b",
          3562 => x"11",
          3563 => x"71",
          3564 => x"33",
          3565 => x"70",
          3566 => x"41",
          3567 => x"1d",
          3568 => x"b8",
          3569 => x"12",
          3570 => x"07",
          3571 => x"33",
          3572 => x"5f",
          3573 => x"77",
          3574 => x"84",
          3575 => x"12",
          3576 => x"ff",
          3577 => x"59",
          3578 => x"84",
          3579 => x"33",
          3580 => x"83",
          3581 => x"15",
          3582 => x"2a",
          3583 => x"55",
          3584 => x"84",
          3585 => x"81",
          3586 => x"2b",
          3587 => x"15",
          3588 => x"2a",
          3589 => x"55",
          3590 => x"34",
          3591 => x"11",
          3592 => x"07",
          3593 => x"42",
          3594 => x"51",
          3595 => x"08",
          3596 => x"70",
          3597 => x"7a",
          3598 => x"73",
          3599 => x"04",
          3600 => x"0c",
          3601 => x"82",
          3602 => x"f4",
          3603 => x"b8",
          3604 => x"81",
          3605 => x"60",
          3606 => x"34",
          3607 => x"1d",
          3608 => x"b9",
          3609 => x"05",
          3610 => x"ff",
          3611 => x"57",
          3612 => x"34",
          3613 => x"10",
          3614 => x"55",
          3615 => x"83",
          3616 => x"7e",
          3617 => x"8c",
          3618 => x"df",
          3619 => x"b9",
          3620 => x"3d",
          3621 => x"08",
          3622 => x"7f",
          3623 => x"88",
          3624 => x"88",
          3625 => x"7b",
          3626 => x"b9",
          3627 => x"58",
          3628 => x"34",
          3629 => x"33",
          3630 => x"70",
          3631 => x"05",
          3632 => x"2a",
          3633 => x"63",
          3634 => x"06",
          3635 => x"b9",
          3636 => x"60",
          3637 => x"08",
          3638 => x"7e",
          3639 => x"70",
          3640 => x"ac",
          3641 => x"31",
          3642 => x"33",
          3643 => x"70",
          3644 => x"12",
          3645 => x"07",
          3646 => x"54",
          3647 => x"bc",
          3648 => x"80",
          3649 => x"ff",
          3650 => x"dd",
          3651 => x"0b",
          3652 => x"84",
          3653 => x"7e",
          3654 => x"cc",
          3655 => x"7a",
          3656 => x"b9",
          3657 => x"81",
          3658 => x"08",
          3659 => x"87",
          3660 => x"b9",
          3661 => x"07",
          3662 => x"2a",
          3663 => x"05",
          3664 => x"b9",
          3665 => x"b9",
          3666 => x"7e",
          3667 => x"05",
          3668 => x"83",
          3669 => x"5b",
          3670 => x"f2",
          3671 => x"7e",
          3672 => x"84",
          3673 => x"76",
          3674 => x"71",
          3675 => x"11",
          3676 => x"8b",
          3677 => x"84",
          3678 => x"2b",
          3679 => x"56",
          3680 => x"78",
          3681 => x"05",
          3682 => x"84",
          3683 => x"2b",
          3684 => x"14",
          3685 => x"07",
          3686 => x"5d",
          3687 => x"34",
          3688 => x"b8",
          3689 => x"71",
          3690 => x"70",
          3691 => x"7d",
          3692 => x"b8",
          3693 => x"12",
          3694 => x"07",
          3695 => x"71",
          3696 => x"5c",
          3697 => x"7c",
          3698 => x"b8",
          3699 => x"33",
          3700 => x"74",
          3701 => x"71",
          3702 => x"47",
          3703 => x"82",
          3704 => x"b9",
          3705 => x"83",
          3706 => x"57",
          3707 => x"58",
          3708 => x"bd",
          3709 => x"84",
          3710 => x"5f",
          3711 => x"84",
          3712 => x"b9",
          3713 => x"52",
          3714 => x"3f",
          3715 => x"34",
          3716 => x"b8",
          3717 => x"0b",
          3718 => x"54",
          3719 => x"15",
          3720 => x"b4",
          3721 => x"70",
          3722 => x"45",
          3723 => x"60",
          3724 => x"70",
          3725 => x"05",
          3726 => x"34",
          3727 => x"e7",
          3728 => x"86",
          3729 => x"2b",
          3730 => x"1c",
          3731 => x"07",
          3732 => x"59",
          3733 => x"61",
          3734 => x"70",
          3735 => x"71",
          3736 => x"05",
          3737 => x"88",
          3738 => x"48",
          3739 => x"86",
          3740 => x"84",
          3741 => x"12",
          3742 => x"ff",
          3743 => x"58",
          3744 => x"84",
          3745 => x"81",
          3746 => x"2b",
          3747 => x"33",
          3748 => x"8f",
          3749 => x"2a",
          3750 => x"44",
          3751 => x"17",
          3752 => x"70",
          3753 => x"71",
          3754 => x"81",
          3755 => x"ff",
          3756 => x"5e",
          3757 => x"34",
          3758 => x"ff",
          3759 => x"15",
          3760 => x"71",
          3761 => x"33",
          3762 => x"70",
          3763 => x"5d",
          3764 => x"34",
          3765 => x"11",
          3766 => x"71",
          3767 => x"33",
          3768 => x"70",
          3769 => x"42",
          3770 => x"75",
          3771 => x"08",
          3772 => x"88",
          3773 => x"88",
          3774 => x"34",
          3775 => x"08",
          3776 => x"71",
          3777 => x"05",
          3778 => x"2b",
          3779 => x"06",
          3780 => x"5f",
          3781 => x"82",
          3782 => x"b9",
          3783 => x"12",
          3784 => x"07",
          3785 => x"71",
          3786 => x"70",
          3787 => x"59",
          3788 => x"1d",
          3789 => x"82",
          3790 => x"2b",
          3791 => x"11",
          3792 => x"71",
          3793 => x"33",
          3794 => x"70",
          3795 => x"42",
          3796 => x"84",
          3797 => x"b9",
          3798 => x"85",
          3799 => x"2b",
          3800 => x"15",
          3801 => x"2a",
          3802 => x"57",
          3803 => x"34",
          3804 => x"81",
          3805 => x"ff",
          3806 => x"5e",
          3807 => x"34",
          3808 => x"11",
          3809 => x"71",
          3810 => x"81",
          3811 => x"88",
          3812 => x"55",
          3813 => x"34",
          3814 => x"33",
          3815 => x"83",
          3816 => x"83",
          3817 => x"88",
          3818 => x"55",
          3819 => x"1a",
          3820 => x"82",
          3821 => x"2b",
          3822 => x"2b",
          3823 => x"05",
          3824 => x"b8",
          3825 => x"1c",
          3826 => x"5f",
          3827 => x"1a",
          3828 => x"07",
          3829 => x"33",
          3830 => x"40",
          3831 => x"84",
          3832 => x"84",
          3833 => x"33",
          3834 => x"83",
          3835 => x"87",
          3836 => x"88",
          3837 => x"41",
          3838 => x"64",
          3839 => x"1d",
          3840 => x"2b",
          3841 => x"2a",
          3842 => x"7c",
          3843 => x"70",
          3844 => x"8b",
          3845 => x"70",
          3846 => x"07",
          3847 => x"77",
          3848 => x"49",
          3849 => x"1e",
          3850 => x"b8",
          3851 => x"33",
          3852 => x"74",
          3853 => x"88",
          3854 => x"88",
          3855 => x"5e",
          3856 => x"34",
          3857 => x"83",
          3858 => x"3f",
          3859 => x"c8",
          3860 => x"73",
          3861 => x"b5",
          3862 => x"61",
          3863 => x"f0",
          3864 => x"29",
          3865 => x"80",
          3866 => x"38",
          3867 => x"0d",
          3868 => x"b9",
          3869 => x"80",
          3870 => x"84",
          3871 => x"3f",
          3872 => x"0d",
          3873 => x"b8",
          3874 => x"23",
          3875 => x"ff",
          3876 => x"b9",
          3877 => x"0b",
          3878 => x"54",
          3879 => x"15",
          3880 => x"86",
          3881 => x"84",
          3882 => x"ff",
          3883 => x"ff",
          3884 => x"55",
          3885 => x"17",
          3886 => x"10",
          3887 => x"05",
          3888 => x"0b",
          3889 => x"2e",
          3890 => x"3d",
          3891 => x"52",
          3892 => x"c4",
          3893 => x"0c",
          3894 => x"02",
          3895 => x"81",
          3896 => x"3f",
          3897 => x"53",
          3898 => x"13",
          3899 => x"72",
          3900 => x"04",
          3901 => x"8c",
          3902 => x"59",
          3903 => x"84",
          3904 => x"06",
          3905 => x"58",
          3906 => x"78",
          3907 => x"3f",
          3908 => x"55",
          3909 => x"98",
          3910 => x"78",
          3911 => x"06",
          3912 => x"54",
          3913 => x"8b",
          3914 => x"19",
          3915 => x"79",
          3916 => x"f7",
          3917 => x"05",
          3918 => x"81",
          3919 => x"b9",
          3920 => x"54",
          3921 => x"85",
          3922 => x"53",
          3923 => x"84",
          3924 => x"74",
          3925 => x"8c",
          3926 => x"26",
          3927 => x"54",
          3928 => x"73",
          3929 => x"3d",
          3930 => x"70",
          3931 => x"78",
          3932 => x"3d",
          3933 => x"33",
          3934 => x"53",
          3935 => x"38",
          3936 => x"81",
          3937 => x"85",
          3938 => x"53",
          3939 => x"25",
          3940 => x"84",
          3941 => x"3d",
          3942 => x"73",
          3943 => x"04",
          3944 => x"b9",
          3945 => x"84",
          3946 => x"54",
          3947 => x"2a",
          3948 => x"8a",
          3949 => x"74",
          3950 => x"51",
          3951 => x"c0",
          3952 => x"06",
          3953 => x"71",
          3954 => x"ff",
          3955 => x"80",
          3956 => x"57",
          3957 => x"38",
          3958 => x"87",
          3959 => x"33",
          3960 => x"08",
          3961 => x"84",
          3962 => x"81",
          3963 => x"70",
          3964 => x"ff",
          3965 => x"77",
          3966 => x"b9",
          3967 => x"08",
          3968 => x"08",
          3969 => x"5b",
          3970 => x"18",
          3971 => x"06",
          3972 => x"53",
          3973 => x"b7",
          3974 => x"83",
          3975 => x"84",
          3976 => x"81",
          3977 => x"84",
          3978 => x"81",
          3979 => x"f4",
          3980 => x"34",
          3981 => x"80",
          3982 => x"19",
          3983 => x"80",
          3984 => x"0b",
          3985 => x"84",
          3986 => x"9e",
          3987 => x"19",
          3988 => x"a0",
          3989 => x"84",
          3990 => x"75",
          3991 => x"5b",
          3992 => x"08",
          3993 => x"88",
          3994 => x"7a",
          3995 => x"34",
          3996 => x"19",
          3997 => x"b4",
          3998 => x"79",
          3999 => x"3f",
          4000 => x"52",
          4001 => x"84",
          4002 => x"38",
          4003 => x"60",
          4004 => x"27",
          4005 => x"8c",
          4006 => x"0c",
          4007 => x"56",
          4008 => x"74",
          4009 => x"2e",
          4010 => x"2a",
          4011 => x"05",
          4012 => x"79",
          4013 => x"7b",
          4014 => x"38",
          4015 => x"81",
          4016 => x"b9",
          4017 => x"59",
          4018 => x"ff",
          4019 => x"b8",
          4020 => x"a8",
          4021 => x"b4",
          4022 => x"0b",
          4023 => x"74",
          4024 => x"38",
          4025 => x"81",
          4026 => x"b9",
          4027 => x"59",
          4028 => x"fe",
          4029 => x"b8",
          4030 => x"78",
          4031 => x"59",
          4032 => x"9f",
          4033 => x"3d",
          4034 => x"08",
          4035 => x"b5",
          4036 => x"5c",
          4037 => x"06",
          4038 => x"b8",
          4039 => x"a8",
          4040 => x"85",
          4041 => x"18",
          4042 => x"83",
          4043 => x"11",
          4044 => x"84",
          4045 => x"0d",
          4046 => x"fd",
          4047 => x"08",
          4048 => x"b5",
          4049 => x"5c",
          4050 => x"06",
          4051 => x"b8",
          4052 => x"c0",
          4053 => x"85",
          4054 => x"18",
          4055 => x"2b",
          4056 => x"83",
          4057 => x"2b",
          4058 => x"70",
          4059 => x"80",
          4060 => x"b9",
          4061 => x"56",
          4062 => x"17",
          4063 => x"18",
          4064 => x"5a",
          4065 => x"81",
          4066 => x"08",
          4067 => x"18",
          4068 => x"5e",
          4069 => x"38",
          4070 => x"09",
          4071 => x"b4",
          4072 => x"7b",
          4073 => x"3f",
          4074 => x"b4",
          4075 => x"81",
          4076 => x"84",
          4077 => x"06",
          4078 => x"83",
          4079 => x"08",
          4080 => x"8b",
          4081 => x"2e",
          4082 => x"5b",
          4083 => x"08",
          4084 => x"33",
          4085 => x"84",
          4086 => x"06",
          4087 => x"83",
          4088 => x"08",
          4089 => x"7d",
          4090 => x"82",
          4091 => x"81",
          4092 => x"17",
          4093 => x"52",
          4094 => x"7a",
          4095 => x"17",
          4096 => x"18",
          4097 => x"5a",
          4098 => x"81",
          4099 => x"08",
          4100 => x"18",
          4101 => x"55",
          4102 => x"38",
          4103 => x"09",
          4104 => x"b4",
          4105 => x"7d",
          4106 => x"3f",
          4107 => x"b4",
          4108 => x"7b",
          4109 => x"3f",
          4110 => x"bb",
          4111 => x"60",
          4112 => x"81",
          4113 => x"08",
          4114 => x"78",
          4115 => x"80",
          4116 => x"77",
          4117 => x"04",
          4118 => x"58",
          4119 => x"76",
          4120 => x"33",
          4121 => x"81",
          4122 => x"53",
          4123 => x"f2",
          4124 => x"2e",
          4125 => x"b4",
          4126 => x"38",
          4127 => x"7b",
          4128 => x"b8",
          4129 => x"b9",
          4130 => x"77",
          4131 => x"04",
          4132 => x"ff",
          4133 => x"05",
          4134 => x"5c",
          4135 => x"19",
          4136 => x"09",
          4137 => x"77",
          4138 => x"51",
          4139 => x"80",
          4140 => x"77",
          4141 => x"b7",
          4142 => x"79",
          4143 => x"98",
          4144 => x"06",
          4145 => x"34",
          4146 => x"34",
          4147 => x"34",
          4148 => x"34",
          4149 => x"39",
          4150 => x"a8",
          4151 => x"59",
          4152 => x"0b",
          4153 => x"74",
          4154 => x"38",
          4155 => x"81",
          4156 => x"b9",
          4157 => x"58",
          4158 => x"58",
          4159 => x"06",
          4160 => x"06",
          4161 => x"2e",
          4162 => x"06",
          4163 => x"5a",
          4164 => x"34",
          4165 => x"56",
          4166 => x"74",
          4167 => x"74",
          4168 => x"33",
          4169 => x"84",
          4170 => x"06",
          4171 => x"83",
          4172 => x"1b",
          4173 => x"c8",
          4174 => x"27",
          4175 => x"82",
          4176 => x"53",
          4177 => x"d8",
          4178 => x"85",
          4179 => x"1a",
          4180 => x"ff",
          4181 => x"56",
          4182 => x"76",
          4183 => x"07",
          4184 => x"83",
          4185 => x"76",
          4186 => x"33",
          4187 => x"84",
          4188 => x"06",
          4189 => x"83",
          4190 => x"1b",
          4191 => x"c8",
          4192 => x"27",
          4193 => x"74",
          4194 => x"38",
          4195 => x"81",
          4196 => x"5a",
          4197 => x"b8",
          4198 => x"57",
          4199 => x"c8",
          4200 => x"ae",
          4201 => x"34",
          4202 => x"31",
          4203 => x"5f",
          4204 => x"f0",
          4205 => x"2e",
          4206 => x"54",
          4207 => x"33",
          4208 => x"d0",
          4209 => x"70",
          4210 => x"cf",
          4211 => x"7c",
          4212 => x"84",
          4213 => x"19",
          4214 => x"1b",
          4215 => x"40",
          4216 => x"82",
          4217 => x"81",
          4218 => x"1e",
          4219 => x"ed",
          4220 => x"81",
          4221 => x"19",
          4222 => x"fd",
          4223 => x"06",
          4224 => x"59",
          4225 => x"88",
          4226 => x"fa",
          4227 => x"76",
          4228 => x"b8",
          4229 => x"8f",
          4230 => x"42",
          4231 => x"7d",
          4232 => x"7d",
          4233 => x"7d",
          4234 => x"fa",
          4235 => x"71",
          4236 => x"38",
          4237 => x"80",
          4238 => x"80",
          4239 => x"54",
          4240 => x"7b",
          4241 => x"16",
          4242 => x"38",
          4243 => x"38",
          4244 => x"84",
          4245 => x"38",
          4246 => x"2e",
          4247 => x"70",
          4248 => x"7b",
          4249 => x"aa",
          4250 => x"ff",
          4251 => x"c8",
          4252 => x"ff",
          4253 => x"ca",
          4254 => x"3f",
          4255 => x"27",
          4256 => x"84",
          4257 => x"9c",
          4258 => x"c4",
          4259 => x"1b",
          4260 => x"38",
          4261 => x"eb",
          4262 => x"81",
          4263 => x"08",
          4264 => x"25",
          4265 => x"54",
          4266 => x"38",
          4267 => x"38",
          4268 => x"fe",
          4269 => x"fe",
          4270 => x"96",
          4271 => x"ff",
          4272 => x"3f",
          4273 => x"08",
          4274 => x"80",
          4275 => x"38",
          4276 => x"0c",
          4277 => x"08",
          4278 => x"ff",
          4279 => x"81",
          4280 => x"55",
          4281 => x"0d",
          4282 => x"8c",
          4283 => x"58",
          4284 => x"b8",
          4285 => x"f5",
          4286 => x"ff",
          4287 => x"b9",
          4288 => x"56",
          4289 => x"55",
          4290 => x"7c",
          4291 => x"80",
          4292 => x"06",
          4293 => x"19",
          4294 => x"df",
          4295 => x"80",
          4296 => x"0b",
          4297 => x"27",
          4298 => x"0c",
          4299 => x"53",
          4300 => x"73",
          4301 => x"83",
          4302 => x"0c",
          4303 => x"8a",
          4304 => x"c8",
          4305 => x"08",
          4306 => x"8a",
          4307 => x"73",
          4308 => x"53",
          4309 => x"59",
          4310 => x"22",
          4311 => x"5a",
          4312 => x"39",
          4313 => x"84",
          4314 => x"08",
          4315 => x"b9",
          4316 => x"17",
          4317 => x"27",
          4318 => x"73",
          4319 => x"81",
          4320 => x"0d",
          4321 => x"90",
          4322 => x"f0",
          4323 => x"0b",
          4324 => x"84",
          4325 => x"83",
          4326 => x"15",
          4327 => x"38",
          4328 => x"55",
          4329 => x"98",
          4330 => x"1b",
          4331 => x"75",
          4332 => x"04",
          4333 => x"ff",
          4334 => x"da",
          4335 => x"3f",
          4336 => x"81",
          4337 => x"38",
          4338 => x"2e",
          4339 => x"c8",
          4340 => x"2e",
          4341 => x"76",
          4342 => x"08",
          4343 => x"80",
          4344 => x"b9",
          4345 => x"81",
          4346 => x"ff",
          4347 => x"1a",
          4348 => x"fe",
          4349 => x"56",
          4350 => x"8a",
          4351 => x"08",
          4352 => x"b8",
          4353 => x"80",
          4354 => x"15",
          4355 => x"19",
          4356 => x"38",
          4357 => x"81",
          4358 => x"b9",
          4359 => x"56",
          4360 => x"0b",
          4361 => x"04",
          4362 => x"19",
          4363 => x"e4",
          4364 => x"f3",
          4365 => x"34",
          4366 => x"55",
          4367 => x"38",
          4368 => x"09",
          4369 => x"b4",
          4370 => x"75",
          4371 => x"3f",
          4372 => x"74",
          4373 => x"2e",
          4374 => x"18",
          4375 => x"05",
          4376 => x"fd",
          4377 => x"29",
          4378 => x"5c",
          4379 => x"c8",
          4380 => x"0d",
          4381 => x"5a",
          4382 => x"58",
          4383 => x"38",
          4384 => x"b4",
          4385 => x"83",
          4386 => x"2e",
          4387 => x"54",
          4388 => x"33",
          4389 => x"08",
          4390 => x"57",
          4391 => x"82",
          4392 => x"58",
          4393 => x"8b",
          4394 => x"06",
          4395 => x"81",
          4396 => x"70",
          4397 => x"07",
          4398 => x"38",
          4399 => x"88",
          4400 => x"81",
          4401 => x"7b",
          4402 => x"08",
          4403 => x"38",
          4404 => x"38",
          4405 => x"0d",
          4406 => x"7e",
          4407 => x"3f",
          4408 => x"2e",
          4409 => x"b9",
          4410 => x"08",
          4411 => x"08",
          4412 => x"fe",
          4413 => x"82",
          4414 => x"81",
          4415 => x"05",
          4416 => x"e0",
          4417 => x"79",
          4418 => x"38",
          4419 => x"80",
          4420 => x"81",
          4421 => x"ac",
          4422 => x"2e",
          4423 => x"fe",
          4424 => x"09",
          4425 => x"84",
          4426 => x"84",
          4427 => x"77",
          4428 => x"57",
          4429 => x"38",
          4430 => x"1a",
          4431 => x"41",
          4432 => x"81",
          4433 => x"5a",
          4434 => x"17",
          4435 => x"33",
          4436 => x"7a",
          4437 => x"fe",
          4438 => x"05",
          4439 => x"1a",
          4440 => x"cc",
          4441 => x"06",
          4442 => x"79",
          4443 => x"10",
          4444 => x"1d",
          4445 => x"9d",
          4446 => x"38",
          4447 => x"a8",
          4448 => x"2a",
          4449 => x"81",
          4450 => x"81",
          4451 => x"76",
          4452 => x"38",
          4453 => x"b9",
          4454 => x"3d",
          4455 => x"52",
          4456 => x"c8",
          4457 => x"80",
          4458 => x"0b",
          4459 => x"1c",
          4460 => x"76",
          4461 => x"78",
          4462 => x"06",
          4463 => x"b8",
          4464 => x"e0",
          4465 => x"85",
          4466 => x"1c",
          4467 => x"9c",
          4468 => x"80",
          4469 => x"bf",
          4470 => x"77",
          4471 => x"80",
          4472 => x"55",
          4473 => x"80",
          4474 => x"38",
          4475 => x"8b",
          4476 => x"29",
          4477 => x"57",
          4478 => x"19",
          4479 => x"7f",
          4480 => x"81",
          4481 => x"a0",
          4482 => x"5a",
          4483 => x"71",
          4484 => x"40",
          4485 => x"80",
          4486 => x"0b",
          4487 => x"f5",
          4488 => x"84",
          4489 => x"38",
          4490 => x"0d",
          4491 => x"7d",
          4492 => x"3f",
          4493 => x"2e",
          4494 => x"b9",
          4495 => x"08",
          4496 => x"08",
          4497 => x"fd",
          4498 => x"82",
          4499 => x"81",
          4500 => x"05",
          4501 => x"db",
          4502 => x"77",
          4503 => x"70",
          4504 => x"fe",
          4505 => x"5a",
          4506 => x"33",
          4507 => x"08",
          4508 => x"76",
          4509 => x"74",
          4510 => x"3f",
          4511 => x"c8",
          4512 => x"c8",
          4513 => x"81",
          4514 => x"fe",
          4515 => x"77",
          4516 => x"1b",
          4517 => x"71",
          4518 => x"ff",
          4519 => x"8d",
          4520 => x"59",
          4521 => x"05",
          4522 => x"2b",
          4523 => x"80",
          4524 => x"84",
          4525 => x"84",
          4526 => x"70",
          4527 => x"81",
          4528 => x"08",
          4529 => x"76",
          4530 => x"ff",
          4531 => x"81",
          4532 => x"38",
          4533 => x"60",
          4534 => x"b4",
          4535 => x"5e",
          4536 => x"b9",
          4537 => x"83",
          4538 => x"ff",
          4539 => x"68",
          4540 => x"a0",
          4541 => x"74",
          4542 => x"70",
          4543 => x"8e",
          4544 => x"22",
          4545 => x"3d",
          4546 => x"58",
          4547 => x"33",
          4548 => x"15",
          4549 => x"05",
          4550 => x"80",
          4551 => x"ab",
          4552 => x"5b",
          4553 => x"7a",
          4554 => x"05",
          4555 => x"34",
          4556 => x"7b",
          4557 => x"56",
          4558 => x"82",
          4559 => x"06",
          4560 => x"83",
          4561 => x"06",
          4562 => x"87",
          4563 => x"ff",
          4564 => x"78",
          4565 => x"84",
          4566 => x"b0",
          4567 => x"84",
          4568 => x"ff",
          4569 => x"59",
          4570 => x"80",
          4571 => x"80",
          4572 => x"74",
          4573 => x"75",
          4574 => x"70",
          4575 => x"81",
          4576 => x"55",
          4577 => x"78",
          4578 => x"57",
          4579 => x"27",
          4580 => x"3f",
          4581 => x"1b",
          4582 => x"38",
          4583 => x"e7",
          4584 => x"b9",
          4585 => x"82",
          4586 => x"ab",
          4587 => x"80",
          4588 => x"2a",
          4589 => x"2e",
          4590 => x"fe",
          4591 => x"1b",
          4592 => x"3f",
          4593 => x"c8",
          4594 => x"08",
          4595 => x"56",
          4596 => x"85",
          4597 => x"77",
          4598 => x"81",
          4599 => x"18",
          4600 => x"c8",
          4601 => x"81",
          4602 => x"76",
          4603 => x"56",
          4604 => x"38",
          4605 => x"56",
          4606 => x"81",
          4607 => x"38",
          4608 => x"84",
          4609 => x"08",
          4610 => x"75",
          4611 => x"75",
          4612 => x"81",
          4613 => x"1c",
          4614 => x"33",
          4615 => x"81",
          4616 => x"1c",
          4617 => x"c8",
          4618 => x"81",
          4619 => x"75",
          4620 => x"08",
          4621 => x"58",
          4622 => x"8b",
          4623 => x"55",
          4624 => x"70",
          4625 => x"74",
          4626 => x"33",
          4627 => x"34",
          4628 => x"75",
          4629 => x"04",
          4630 => x"07",
          4631 => x"74",
          4632 => x"3f",
          4633 => x"c8",
          4634 => x"bd",
          4635 => x"7c",
          4636 => x"3f",
          4637 => x"81",
          4638 => x"08",
          4639 => x"19",
          4640 => x"27",
          4641 => x"82",
          4642 => x"08",
          4643 => x"90",
          4644 => x"51",
          4645 => x"58",
          4646 => x"79",
          4647 => x"57",
          4648 => x"05",
          4649 => x"76",
          4650 => x"59",
          4651 => x"ff",
          4652 => x"08",
          4653 => x"2e",
          4654 => x"76",
          4655 => x"81",
          4656 => x"1c",
          4657 => x"c8",
          4658 => x"81",
          4659 => x"75",
          4660 => x"1f",
          4661 => x"5f",
          4662 => x"1c",
          4663 => x"1c",
          4664 => x"29",
          4665 => x"76",
          4666 => x"10",
          4667 => x"56",
          4668 => x"55",
          4669 => x"76",
          4670 => x"85",
          4671 => x"58",
          4672 => x"ff",
          4673 => x"1f",
          4674 => x"81",
          4675 => x"83",
          4676 => x"e1",
          4677 => x"b9",
          4678 => x"05",
          4679 => x"39",
          4680 => x"1c",
          4681 => x"d0",
          4682 => x"08",
          4683 => x"83",
          4684 => x"08",
          4685 => x"60",
          4686 => x"82",
          4687 => x"81",
          4688 => x"1c",
          4689 => x"52",
          4690 => x"77",
          4691 => x"08",
          4692 => x"e5",
          4693 => x"fb",
          4694 => x"80",
          4695 => x"7c",
          4696 => x"81",
          4697 => x"81",
          4698 => x"b9",
          4699 => x"bc",
          4700 => x"34",
          4701 => x"55",
          4702 => x"82",
          4703 => x"38",
          4704 => x"39",
          4705 => x"2e",
          4706 => x"1a",
          4707 => x"56",
          4708 => x"fd",
          4709 => x"1d",
          4710 => x"33",
          4711 => x"81",
          4712 => x"05",
          4713 => x"ce",
          4714 => x"0d",
          4715 => x"80",
          4716 => x"80",
          4717 => x"ff",
          4718 => x"60",
          4719 => x"5b",
          4720 => x"77",
          4721 => x"5b",
          4722 => x"d0",
          4723 => x"58",
          4724 => x"38",
          4725 => x"5d",
          4726 => x"30",
          4727 => x"5a",
          4728 => x"80",
          4729 => x"1f",
          4730 => x"70",
          4731 => x"a0",
          4732 => x"bc",
          4733 => x"72",
          4734 => x"8b",
          4735 => x"38",
          4736 => x"81",
          4737 => x"59",
          4738 => x"ff",
          4739 => x"80",
          4740 => x"53",
          4741 => x"bf",
          4742 => x"17",
          4743 => x"34",
          4744 => x"53",
          4745 => x"9c",
          4746 => x"1e",
          4747 => x"11",
          4748 => x"71",
          4749 => x"72",
          4750 => x"64",
          4751 => x"33",
          4752 => x"40",
          4753 => x"23",
          4754 => x"88",
          4755 => x"23",
          4756 => x"fe",
          4757 => x"ff",
          4758 => x"52",
          4759 => x"91",
          4760 => x"ff",
          4761 => x"ad",
          4762 => x"74",
          4763 => x"97",
          4764 => x"0b",
          4765 => x"75",
          4766 => x"fd",
          4767 => x"76",
          4768 => x"80",
          4769 => x"f9",
          4770 => x"58",
          4771 => x"cd",
          4772 => x"57",
          4773 => x"7c",
          4774 => x"14",
          4775 => x"99",
          4776 => x"11",
          4777 => x"38",
          4778 => x"5e",
          4779 => x"70",
          4780 => x"78",
          4781 => x"81",
          4782 => x"5e",
          4783 => x"38",
          4784 => x"cc",
          4785 => x"70",
          4786 => x"fc",
          4787 => x"08",
          4788 => x"33",
          4789 => x"38",
          4790 => x"df",
          4791 => x"98",
          4792 => x"96",
          4793 => x"75",
          4794 => x"16",
          4795 => x"81",
          4796 => x"df",
          4797 => x"81",
          4798 => x"8b",
          4799 => x"23",
          4800 => x"06",
          4801 => x"27",
          4802 => x"55",
          4803 => x"2e",
          4804 => x"b2",
          4805 => x"e4",
          4806 => x"56",
          4807 => x"75",
          4808 => x"70",
          4809 => x"ee",
          4810 => x"81",
          4811 => x"fd",
          4812 => x"23",
          4813 => x"52",
          4814 => x"fe",
          4815 => x"80",
          4816 => x"73",
          4817 => x"2e",
          4818 => x"80",
          4819 => x"dd",
          4820 => x"70",
          4821 => x"72",
          4822 => x"33",
          4823 => x"74",
          4824 => x"83",
          4825 => x"3f",
          4826 => x"06",
          4827 => x"73",
          4828 => x"04",
          4829 => x"06",
          4830 => x"38",
          4831 => x"34",
          4832 => x"84",
          4833 => x"93",
          4834 => x"32",
          4835 => x"41",
          4836 => x"38",
          4837 => x"55",
          4838 => x"72",
          4839 => x"25",
          4840 => x"38",
          4841 => x"2b",
          4842 => x"76",
          4843 => x"59",
          4844 => x"78",
          4845 => x"32",
          4846 => x"56",
          4847 => x"38",
          4848 => x"dd",
          4849 => x"76",
          4850 => x"80",
          4851 => x"72",
          4852 => x"82",
          4853 => x"53",
          4854 => x"80",
          4855 => x"70",
          4856 => x"38",
          4857 => x"17",
          4858 => x"14",
          4859 => x"09",
          4860 => x"1d",
          4861 => x"56",
          4862 => x"72",
          4863 => x"22",
          4864 => x"80",
          4865 => x"83",
          4866 => x"70",
          4867 => x"2e",
          4868 => x"72",
          4869 => x"59",
          4870 => x"07",
          4871 => x"54",
          4872 => x"7c",
          4873 => x"2e",
          4874 => x"77",
          4875 => x"8b",
          4876 => x"18",
          4877 => x"81",
          4878 => x"38",
          4879 => x"2e",
          4880 => x"e3",
          4881 => x"2e",
          4882 => x"74",
          4883 => x"2a",
          4884 => x"81",
          4885 => x"79",
          4886 => x"06",
          4887 => x"88",
          4888 => x"51",
          4889 => x"ab",
          4890 => x"08",
          4891 => x"c8",
          4892 => x"f7",
          4893 => x"79",
          4894 => x"2a",
          4895 => x"7b",
          4896 => x"16",
          4897 => x"81",
          4898 => x"40",
          4899 => x"38",
          4900 => x"83",
          4901 => x"22",
          4902 => x"fc",
          4903 => x"2e",
          4904 => x"10",
          4905 => x"a0",
          4906 => x"26",
          4907 => x"81",
          4908 => x"73",
          4909 => x"77",
          4910 => x"3f",
          4911 => x"56",
          4912 => x"38",
          4913 => x"fa",
          4914 => x"2a",
          4915 => x"83",
          4916 => x"06",
          4917 => x"d2",
          4918 => x"33",
          4919 => x"82",
          4920 => x"08",
          4921 => x"22",
          4922 => x"76",
          4923 => x"ab",
          4924 => x"5a",
          4925 => x"fc",
          4926 => x"8c",
          4927 => x"79",
          4928 => x"0b",
          4929 => x"81",
          4930 => x"80",
          4931 => x"b9",
          4932 => x"80",
          4933 => x"27",
          4934 => x"7b",
          4935 => x"7d",
          4936 => x"39",
          4937 => x"74",
          4938 => x"c8",
          4939 => x"2a",
          4940 => x"c4",
          4941 => x"d8",
          4942 => x"26",
          4943 => x"85",
          4944 => x"f0",
          4945 => x"59",
          4946 => x"75",
          4947 => x"70",
          4948 => x"ee",
          4949 => x"80",
          4950 => x"99",
          4951 => x"81",
          4952 => x"59",
          4953 => x"07",
          4954 => x"83",
          4955 => x"7b",
          4956 => x"81",
          4957 => x"39",
          4958 => x"f0",
          4959 => x"78",
          4960 => x"7a",
          4961 => x"5b",
          4962 => x"d2",
          4963 => x"15",
          4964 => x"07",
          4965 => x"fd",
          4966 => x"88",
          4967 => x"1b",
          4968 => x"79",
          4969 => x"79",
          4970 => x"76",
          4971 => x"a3",
          4972 => x"81",
          4973 => x"0b",
          4974 => x"04",
          4975 => x"05",
          4976 => x"80",
          4977 => x"5b",
          4978 => x"79",
          4979 => x"26",
          4980 => x"38",
          4981 => x"c7",
          4982 => x"76",
          4983 => x"84",
          4984 => x"8c",
          4985 => x"76",
          4986 => x"33",
          4987 => x"81",
          4988 => x"84",
          4989 => x"81",
          4990 => x"96",
          4991 => x"84",
          4992 => x"81",
          4993 => x"a4",
          4994 => x"06",
          4995 => x"7f",
          4996 => x"38",
          4997 => x"58",
          4998 => x"83",
          4999 => x"7a",
          5000 => x"b8",
          5001 => x"58",
          5002 => x"08",
          5003 => x"59",
          5004 => x"99",
          5005 => x"18",
          5006 => x"83",
          5007 => x"a5",
          5008 => x"b9",
          5009 => x"38",
          5010 => x"38",
          5011 => x"38",
          5012 => x"33",
          5013 => x"84",
          5014 => x"38",
          5015 => x"33",
          5016 => x"a4",
          5017 => x"82",
          5018 => x"2b",
          5019 => x"88",
          5020 => x"45",
          5021 => x"0c",
          5022 => x"80",
          5023 => x"ff",
          5024 => x"81",
          5025 => x"06",
          5026 => x"5a",
          5027 => x"59",
          5028 => x"18",
          5029 => x"80",
          5030 => x"71",
          5031 => x"18",
          5032 => x"8d",
          5033 => x"17",
          5034 => x"2b",
          5035 => x"d8",
          5036 => x"71",
          5037 => x"14",
          5038 => x"33",
          5039 => x"42",
          5040 => x"18",
          5041 => x"8d",
          5042 => x"7d",
          5043 => x"75",
          5044 => x"7a",
          5045 => x"b9",
          5046 => x"80",
          5047 => x"08",
          5048 => x"38",
          5049 => x"83",
          5050 => x"85",
          5051 => x"9c",
          5052 => x"1d",
          5053 => x"1a",
          5054 => x"87",
          5055 => x"7b",
          5056 => x"ac",
          5057 => x"2e",
          5058 => x"2a",
          5059 => x"ff",
          5060 => x"a0",
          5061 => x"94",
          5062 => x"ff",
          5063 => x"2e",
          5064 => x"d1",
          5065 => x"d1",
          5066 => x"d1",
          5067 => x"98",
          5068 => x"c8",
          5069 => x"84",
          5070 => x"76",
          5071 => x"57",
          5072 => x"82",
          5073 => x"5d",
          5074 => x"80",
          5075 => x"5c",
          5076 => x"81",
          5077 => x"5b",
          5078 => x"77",
          5079 => x"81",
          5080 => x"58",
          5081 => x"70",
          5082 => x"70",
          5083 => x"09",
          5084 => x"38",
          5085 => x"07",
          5086 => x"7a",
          5087 => x"84",
          5088 => x"98",
          5089 => x"80",
          5090 => x"81",
          5091 => x"38",
          5092 => x"33",
          5093 => x"81",
          5094 => x"eb",
          5095 => x"07",
          5096 => x"75",
          5097 => x"3d",
          5098 => x"16",
          5099 => x"a5",
          5100 => x"17",
          5101 => x"07",
          5102 => x"88",
          5103 => x"52",
          5104 => x"70",
          5105 => x"17",
          5106 => x"38",
          5107 => x"70",
          5108 => x"71",
          5109 => x"1c",
          5110 => x"08",
          5111 => x"fb",
          5112 => x"0b",
          5113 => x"7a",
          5114 => x"53",
          5115 => x"ff",
          5116 => x"76",
          5117 => x"74",
          5118 => x"38",
          5119 => x"2b",
          5120 => x"d4",
          5121 => x"80",
          5122 => x"81",
          5123 => x"eb",
          5124 => x"07",
          5125 => x"81",
          5126 => x"81",
          5127 => x"bd",
          5128 => x"09",
          5129 => x"76",
          5130 => x"f8",
          5131 => x"5a",
          5132 => x"a8",
          5133 => x"e4",
          5134 => x"05",
          5135 => x"33",
          5136 => x"56",
          5137 => x"75",
          5138 => x"8a",
          5139 => x"7b",
          5140 => x"81",
          5141 => x"1b",
          5142 => x"85",
          5143 => x"82",
          5144 => x"fa",
          5145 => x"97",
          5146 => x"2e",
          5147 => x"18",
          5148 => x"b7",
          5149 => x"97",
          5150 => x"18",
          5151 => x"70",
          5152 => x"05",
          5153 => x"5b",
          5154 => x"d1",
          5155 => x"0b",
          5156 => x"5a",
          5157 => x"7a",
          5158 => x"31",
          5159 => x"80",
          5160 => x"e1",
          5161 => x"59",
          5162 => x"39",
          5163 => x"33",
          5164 => x"81",
          5165 => x"81",
          5166 => x"78",
          5167 => x"7a",
          5168 => x"38",
          5169 => x"81",
          5170 => x"84",
          5171 => x"ff",
          5172 => x"79",
          5173 => x"84",
          5174 => x"71",
          5175 => x"d4",
          5176 => x"38",
          5177 => x"33",
          5178 => x"81",
          5179 => x"75",
          5180 => x"42",
          5181 => x"d2",
          5182 => x"84",
          5183 => x"33",
          5184 => x"81",
          5185 => x"75",
          5186 => x"5c",
          5187 => x"f2",
          5188 => x"84",
          5189 => x"33",
          5190 => x"81",
          5191 => x"75",
          5192 => x"84",
          5193 => x"33",
          5194 => x"81",
          5195 => x"75",
          5196 => x"59",
          5197 => x"5b",
          5198 => x"a0",
          5199 => x"a0",
          5200 => x"a8",
          5201 => x"18",
          5202 => x"f8",
          5203 => x"f2",
          5204 => x"53",
          5205 => x"52",
          5206 => x"c8",
          5207 => x"a4",
          5208 => x"34",
          5209 => x"40",
          5210 => x"82",
          5211 => x"8d",
          5212 => x"a0",
          5213 => x"91",
          5214 => x"e4",
          5215 => x"80",
          5216 => x"71",
          5217 => x"7d",
          5218 => x"61",
          5219 => x"11",
          5220 => x"71",
          5221 => x"72",
          5222 => x"ac",
          5223 => x"43",
          5224 => x"75",
          5225 => x"82",
          5226 => x"f2",
          5227 => x"83",
          5228 => x"f5",
          5229 => x"b4",
          5230 => x"78",
          5231 => x"e7",
          5232 => x"02",
          5233 => x"93",
          5234 => x"40",
          5235 => x"70",
          5236 => x"55",
          5237 => x"73",
          5238 => x"38",
          5239 => x"24",
          5240 => x"d1",
          5241 => x"80",
          5242 => x"54",
          5243 => x"34",
          5244 => x"7c",
          5245 => x"3d",
          5246 => x"3f",
          5247 => x"b9",
          5248 => x"0b",
          5249 => x"04",
          5250 => x"06",
          5251 => x"38",
          5252 => x"05",
          5253 => x"38",
          5254 => x"5f",
          5255 => x"70",
          5256 => x"05",
          5257 => x"55",
          5258 => x"70",
          5259 => x"16",
          5260 => x"16",
          5261 => x"30",
          5262 => x"2e",
          5263 => x"be",
          5264 => x"72",
          5265 => x"54",
          5266 => x"84",
          5267 => x"99",
          5268 => x"83",
          5269 => x"54",
          5270 => x"02",
          5271 => x"59",
          5272 => x"74",
          5273 => x"05",
          5274 => x"ed",
          5275 => x"84",
          5276 => x"80",
          5277 => x"c8",
          5278 => x"6d",
          5279 => x"9a",
          5280 => x"b9",
          5281 => x"77",
          5282 => x"ca",
          5283 => x"76",
          5284 => x"07",
          5285 => x"2a",
          5286 => x"d1",
          5287 => x"33",
          5288 => x"42",
          5289 => x"84",
          5290 => x"80",
          5291 => x"17",
          5292 => x"66",
          5293 => x"67",
          5294 => x"80",
          5295 => x"7c",
          5296 => x"80",
          5297 => x"1c",
          5298 => x"0b",
          5299 => x"83",
          5300 => x"38",
          5301 => x"53",
          5302 => x"38",
          5303 => x"38",
          5304 => x"39",
          5305 => x"2b",
          5306 => x"38",
          5307 => x"fe",
          5308 => x"80",
          5309 => x"06",
          5310 => x"81",
          5311 => x"89",
          5312 => x"f6",
          5313 => x"75",
          5314 => x"07",
          5315 => x"0c",
          5316 => x"33",
          5317 => x"73",
          5318 => x"83",
          5319 => x"0c",
          5320 => x"33",
          5321 => x"81",
          5322 => x"75",
          5323 => x"0c",
          5324 => x"57",
          5325 => x"23",
          5326 => x"1a",
          5327 => x"85",
          5328 => x"84",
          5329 => x"38",
          5330 => x"70",
          5331 => x"30",
          5332 => x"79",
          5333 => x"76",
          5334 => x"86",
          5335 => x"db",
          5336 => x"b9",
          5337 => x"57",
          5338 => x"cb",
          5339 => x"02",
          5340 => x"7d",
          5341 => x"55",
          5342 => x"57",
          5343 => x"57",
          5344 => x"57",
          5345 => x"51",
          5346 => x"78",
          5347 => x"38",
          5348 => x"57",
          5349 => x"94",
          5350 => x"2b",
          5351 => x"fc",
          5352 => x"bd",
          5353 => x"cb",
          5354 => x"b9",
          5355 => x"84",
          5356 => x"38",
          5357 => x"99",
          5358 => x"ff",
          5359 => x"83",
          5360 => x"94",
          5361 => x"27",
          5362 => x"0c",
          5363 => x"84",
          5364 => x"ff",
          5365 => x"94",
          5366 => x"fb",
          5367 => x"33",
          5368 => x"7e",
          5369 => x"17",
          5370 => x"0b",
          5371 => x"17",
          5372 => x"34",
          5373 => x"17",
          5374 => x"33",
          5375 => x"fb",
          5376 => x"7f",
          5377 => x"08",
          5378 => x"5a",
          5379 => x"38",
          5380 => x"81",
          5381 => x"84",
          5382 => x"ff",
          5383 => x"7e",
          5384 => x"57",
          5385 => x"79",
          5386 => x"16",
          5387 => x"17",
          5388 => x"84",
          5389 => x"06",
          5390 => x"83",
          5391 => x"08",
          5392 => x"74",
          5393 => x"82",
          5394 => x"81",
          5395 => x"16",
          5396 => x"52",
          5397 => x"3f",
          5398 => x"1a",
          5399 => x"98",
          5400 => x"83",
          5401 => x"9a",
          5402 => x"fe",
          5403 => x"f9",
          5404 => x"29",
          5405 => x"80",
          5406 => x"15",
          5407 => x"39",
          5408 => x"e4",
          5409 => x"da",
          5410 => x"79",
          5411 => x"5b",
          5412 => x"65",
          5413 => x"7e",
          5414 => x"38",
          5415 => x"38",
          5416 => x"38",
          5417 => x"59",
          5418 => x"55",
          5419 => x"38",
          5420 => x"38",
          5421 => x"56",
          5422 => x"1a",
          5423 => x"56",
          5424 => x"80",
          5425 => x"83",
          5426 => x"8a",
          5427 => x"06",
          5428 => x"38",
          5429 => x"84",
          5430 => x"38",
          5431 => x"1a",
          5432 => x"05",
          5433 => x"38",
          5434 => x"1b",
          5435 => x"83",
          5436 => x"59",
          5437 => x"77",
          5438 => x"75",
          5439 => x"7c",
          5440 => x"e0",
          5441 => x"38",
          5442 => x"80",
          5443 => x"31",
          5444 => x"80",
          5445 => x"58",
          5446 => x"77",
          5447 => x"55",
          5448 => x"7b",
          5449 => x"78",
          5450 => x"94",
          5451 => x"38",
          5452 => x"92",
          5453 => x"0c",
          5454 => x"8e",
          5455 => x"ff",
          5456 => x"7b",
          5457 => x"56",
          5458 => x"80",
          5459 => x"5f",
          5460 => x"e4",
          5461 => x"52",
          5462 => x"3f",
          5463 => x"38",
          5464 => x"0c",
          5465 => x"08",
          5466 => x"58",
          5467 => x"fe",
          5468 => x"33",
          5469 => x"16",
          5470 => x"74",
          5471 => x"81",
          5472 => x"da",
          5473 => x"19",
          5474 => x"1a",
          5475 => x"81",
          5476 => x"09",
          5477 => x"c8",
          5478 => x"a8",
          5479 => x"5c",
          5480 => x"e1",
          5481 => x"2e",
          5482 => x"54",
          5483 => x"53",
          5484 => x"9d",
          5485 => x"76",
          5486 => x"fe",
          5487 => x"51",
          5488 => x"08",
          5489 => x"51",
          5490 => x"08",
          5491 => x"74",
          5492 => x"81",
          5493 => x"b9",
          5494 => x"0b",
          5495 => x"c8",
          5496 => x"0d",
          5497 => x"5a",
          5498 => x"2e",
          5499 => x"2e",
          5500 => x"2e",
          5501 => x"22",
          5502 => x"38",
          5503 => x"82",
          5504 => x"82",
          5505 => x"2a",
          5506 => x"80",
          5507 => x"7b",
          5508 => x"38",
          5509 => x"81",
          5510 => x"82",
          5511 => x"05",
          5512 => x"aa",
          5513 => x"08",
          5514 => x"74",
          5515 => x"2e",
          5516 => x"88",
          5517 => x"0c",
          5518 => x"08",
          5519 => x"fe",
          5520 => x"58",
          5521 => x"16",
          5522 => x"05",
          5523 => x"38",
          5524 => x"77",
          5525 => x"5f",
          5526 => x"31",
          5527 => x"81",
          5528 => x"84",
          5529 => x"b4",
          5530 => x"78",
          5531 => x"18",
          5532 => x"74",
          5533 => x"81",
          5534 => x"ef",
          5535 => x"77",
          5536 => x"08",
          5537 => x"08",
          5538 => x"1e",
          5539 => x"75",
          5540 => x"1b",
          5541 => x"33",
          5542 => x"90",
          5543 => x"c8",
          5544 => x"b9",
          5545 => x"16",
          5546 => x"56",
          5547 => x"59",
          5548 => x"71",
          5549 => x"38",
          5550 => x"78",
          5551 => x"33",
          5552 => x"09",
          5553 => x"77",
          5554 => x"51",
          5555 => x"08",
          5556 => x"5c",
          5557 => x"38",
          5558 => x"11",
          5559 => x"58",
          5560 => x"81",
          5561 => x"57",
          5562 => x"60",
          5563 => x"a3",
          5564 => x"b8",
          5565 => x"40",
          5566 => x"b9",
          5567 => x"ff",
          5568 => x"17",
          5569 => x"31",
          5570 => x"a0",
          5571 => x"16",
          5572 => x"06",
          5573 => x"08",
          5574 => x"81",
          5575 => x"7e",
          5576 => x"57",
          5577 => x"83",
          5578 => x"60",
          5579 => x"58",
          5580 => x"fd",
          5581 => x"51",
          5582 => x"08",
          5583 => x"38",
          5584 => x"76",
          5585 => x"84",
          5586 => x"08",
          5587 => x"b4",
          5588 => x"81",
          5589 => x"3f",
          5590 => x"84",
          5591 => x"16",
          5592 => x"a0",
          5593 => x"16",
          5594 => x"06",
          5595 => x"08",
          5596 => x"81",
          5597 => x"60",
          5598 => x"51",
          5599 => x"08",
          5600 => x"74",
          5601 => x"81",
          5602 => x"70",
          5603 => x"96",
          5604 => x"c6",
          5605 => x"34",
          5606 => x"55",
          5607 => x"38",
          5608 => x"09",
          5609 => x"b4",
          5610 => x"76",
          5611 => x"87",
          5612 => x"1b",
          5613 => x"0b",
          5614 => x"c8",
          5615 => x"91",
          5616 => x"0c",
          5617 => x"7d",
          5618 => x"38",
          5619 => x"38",
          5620 => x"38",
          5621 => x"59",
          5622 => x"55",
          5623 => x"38",
          5624 => x"06",
          5625 => x"38",
          5626 => x"17",
          5627 => x"33",
          5628 => x"78",
          5629 => x"51",
          5630 => x"08",
          5631 => x"56",
          5632 => x"38",
          5633 => x"07",
          5634 => x"08",
          5635 => x"06",
          5636 => x"7a",
          5637 => x"9c",
          5638 => x"5b",
          5639 => x"18",
          5640 => x"2a",
          5641 => x"2a",
          5642 => x"2a",
          5643 => x"34",
          5644 => x"98",
          5645 => x"34",
          5646 => x"93",
          5647 => x"1c",
          5648 => x"84",
          5649 => x"bf",
          5650 => x"75",
          5651 => x"04",
          5652 => x"17",
          5653 => x"ff",
          5654 => x"c8",
          5655 => x"08",
          5656 => x"18",
          5657 => x"55",
          5658 => x"38",
          5659 => x"09",
          5660 => x"b4",
          5661 => x"7a",
          5662 => x"ef",
          5663 => x"90",
          5664 => x"88",
          5665 => x"18",
          5666 => x"2a",
          5667 => x"2a",
          5668 => x"2a",
          5669 => x"34",
          5670 => x"98",
          5671 => x"34",
          5672 => x"93",
          5673 => x"1c",
          5674 => x"84",
          5675 => x"bf",
          5676 => x"fe",
          5677 => x"90",
          5678 => x"06",
          5679 => x"08",
          5680 => x"0d",
          5681 => x"84",
          5682 => x"08",
          5683 => x"9e",
          5684 => x"96",
          5685 => x"8e",
          5686 => x"58",
          5687 => x"52",
          5688 => x"75",
          5689 => x"89",
          5690 => x"ff",
          5691 => x"81",
          5692 => x"08",
          5693 => x"ff",
          5694 => x"2e",
          5695 => x"33",
          5696 => x"2e",
          5697 => x"2e",
          5698 => x"80",
          5699 => x"a4",
          5700 => x"8c",
          5701 => x"c8",
          5702 => x"d0",
          5703 => x"53",
          5704 => x"73",
          5705 => x"73",
          5706 => x"83",
          5707 => x"56",
          5708 => x"75",
          5709 => x"12",
          5710 => x"38",
          5711 => x"54",
          5712 => x"89",
          5713 => x"54",
          5714 => x"51",
          5715 => x"38",
          5716 => x"70",
          5717 => x"07",
          5718 => x"38",
          5719 => x"78",
          5720 => x"cf",
          5721 => x"76",
          5722 => x"0d",
          5723 => x"99",
          5724 => x"c8",
          5725 => x"2e",
          5726 => x"98",
          5727 => x"98",
          5728 => x"84",
          5729 => x"08",
          5730 => x"33",
          5731 => x"24",
          5732 => x"70",
          5733 => x"80",
          5734 => x"33",
          5735 => x"73",
          5736 => x"83",
          5737 => x"74",
          5738 => x"04",
          5739 => x"81",
          5740 => x"b9",
          5741 => x"16",
          5742 => x"71",
          5743 => x"0c",
          5744 => x"12",
          5745 => x"98",
          5746 => x"80",
          5747 => x"5d",
          5748 => x"e4",
          5749 => x"3d",
          5750 => x"08",
          5751 => x"38",
          5752 => x"98",
          5753 => x"80",
          5754 => x"2e",
          5755 => x"3d",
          5756 => x"a4",
          5757 => x"84",
          5758 => x"80",
          5759 => x"08",
          5760 => x"08",
          5761 => x"c7",
          5762 => x"52",
          5763 => x"3f",
          5764 => x"38",
          5765 => x"0c",
          5766 => x"08",
          5767 => x"88",
          5768 => x"59",
          5769 => x"38",
          5770 => x"7a",
          5771 => x"c8",
          5772 => x"9f",
          5773 => x"f5",
          5774 => x"b9",
          5775 => x"08",
          5776 => x"88",
          5777 => x"59",
          5778 => x"38",
          5779 => x"c8",
          5780 => x"3f",
          5781 => x"c8",
          5782 => x"84",
          5783 => x"38",
          5784 => x"7a",
          5785 => x"82",
          5786 => x"90",
          5787 => x"17",
          5788 => x"38",
          5789 => x"95",
          5790 => x"17",
          5791 => x"3d",
          5792 => x"59",
          5793 => x"eb",
          5794 => x"11",
          5795 => x"3d",
          5796 => x"60",
          5797 => x"d1",
          5798 => x"b8",
          5799 => x"59",
          5800 => x"81",
          5801 => x"5a",
          5802 => x"78",
          5803 => x"27",
          5804 => x"7c",
          5805 => x"57",
          5806 => x"70",
          5807 => x"09",
          5808 => x"80",
          5809 => x"80",
          5810 => x"94",
          5811 => x"2b",
          5812 => x"f0",
          5813 => x"71",
          5814 => x"07",
          5815 => x"52",
          5816 => x"b9",
          5817 => x"80",
          5818 => x"81",
          5819 => x"70",
          5820 => x"88",
          5821 => x"08",
          5822 => x"83",
          5823 => x"08",
          5824 => x"74",
          5825 => x"82",
          5826 => x"81",
          5827 => x"16",
          5828 => x"52",
          5829 => x"3f",
          5830 => x"80",
          5831 => x"7b",
          5832 => x"70",
          5833 => x"08",
          5834 => x"7e",
          5835 => x"38",
          5836 => x"18",
          5837 => x"70",
          5838 => x"fe",
          5839 => x"81",
          5840 => x"81",
          5841 => x"38",
          5842 => x"34",
          5843 => x"3d",
          5844 => x"58",
          5845 => x"38",
          5846 => x"38",
          5847 => x"38",
          5848 => x"59",
          5849 => x"53",
          5850 => x"38",
          5851 => x"38",
          5852 => x"81",
          5853 => x"58",
          5854 => x"8a",
          5855 => x"56",
          5856 => x"52",
          5857 => x"84",
          5858 => x"70",
          5859 => x"84",
          5860 => x"38",
          5861 => x"0c",
          5862 => x"58",
          5863 => x"75",
          5864 => x"31",
          5865 => x"90",
          5866 => x"51",
          5867 => x"38",
          5868 => x"3f",
          5869 => x"c8",
          5870 => x"ff",
          5871 => x"b4",
          5872 => x"27",
          5873 => x"ff",
          5874 => x"81",
          5875 => x"3d",
          5876 => x"2a",
          5877 => x"38",
          5878 => x"58",
          5879 => x"b6",
          5880 => x"08",
          5881 => x"8c",
          5882 => x"07",
          5883 => x"ff",
          5884 => x"9c",
          5885 => x"9c",
          5886 => x"0c",
          5887 => x"16",
          5888 => x"2e",
          5889 => x"73",
          5890 => x"39",
          5891 => x"08",
          5892 => x"06",
          5893 => x"fe",
          5894 => x"55",
          5895 => x"8a",
          5896 => x"08",
          5897 => x"53",
          5898 => x"15",
          5899 => x"74",
          5900 => x"c8",
          5901 => x"33",
          5902 => x"c8",
          5903 => x"38",
          5904 => x"39",
          5905 => x"3f",
          5906 => x"c8",
          5907 => x"c8",
          5908 => x"b9",
          5909 => x"16",
          5910 => x"16",
          5911 => x"8b",
          5912 => x"56",
          5913 => x"80",
          5914 => x"3d",
          5915 => x"b9",
          5916 => x"80",
          5917 => x"54",
          5918 => x"0d",
          5919 => x"51",
          5920 => x"08",
          5921 => x"38",
          5922 => x"59",
          5923 => x"33",
          5924 => x"79",
          5925 => x"08",
          5926 => x"88",
          5927 => x"5a",
          5928 => x"77",
          5929 => x"22",
          5930 => x"ff",
          5931 => x"55",
          5932 => x"2e",
          5933 => x"fe",
          5934 => x"f6",
          5935 => x"71",
          5936 => x"07",
          5937 => x"39",
          5938 => x"74",
          5939 => x"72",
          5940 => x"71",
          5941 => x"84",
          5942 => x"94",
          5943 => x"38",
          5944 => x"0c",
          5945 => x"51",
          5946 => x"08",
          5947 => x"75",
          5948 => x"0d",
          5949 => x"80",
          5950 => x"80",
          5951 => x"80",
          5952 => x"16",
          5953 => x"97",
          5954 => x"75",
          5955 => x"f3",
          5956 => x"bd",
          5957 => x"b9",
          5958 => x"b9",
          5959 => x"51",
          5960 => x"51",
          5961 => x"08",
          5962 => x"9f",
          5963 => x"57",
          5964 => x"3d",
          5965 => x"53",
          5966 => x"51",
          5967 => x"08",
          5968 => x"9f",
          5969 => x"57",
          5970 => x"ff",
          5971 => x"84",
          5972 => x"81",
          5973 => x"84",
          5974 => x"fe",
          5975 => x"fe",
          5976 => x"80",
          5977 => x"52",
          5978 => x"08",
          5979 => x"8a",
          5980 => x"3d",
          5981 => x"b5",
          5982 => x"84",
          5983 => x"cb",
          5984 => x"80",
          5985 => x"d1",
          5986 => x"bd",
          5987 => x"3d",
          5988 => x"0c",
          5989 => x"66",
          5990 => x"ec",
          5991 => x"3f",
          5992 => x"c8",
          5993 => x"08",
          5994 => x"08",
          5995 => x"8d",
          5996 => x"c8",
          5997 => x"c8",
          5998 => x"2e",
          5999 => x"84",
          6000 => x"80",
          6001 => x"5d",
          6002 => x"ef",
          6003 => x"7c",
          6004 => x"b8",
          6005 => x"fc",
          6006 => x"2e",
          6007 => x"b4",
          6008 => x"80",
          6009 => x"2e",
          6010 => x"83",
          6011 => x"2b",
          6012 => x"70",
          6013 => x"80",
          6014 => x"30",
          6015 => x"05",
          6016 => x"41",
          6017 => x"5e",
          6018 => x"0c",
          6019 => x"81",
          6020 => x"84",
          6021 => x"81",
          6022 => x"70",
          6023 => x"fc",
          6024 => x"08",
          6025 => x"83",
          6026 => x"08",
          6027 => x"74",
          6028 => x"82",
          6029 => x"81",
          6030 => x"17",
          6031 => x"52",
          6032 => x"3f",
          6033 => x"42",
          6034 => x"51",
          6035 => x"08",
          6036 => x"c8",
          6037 => x"b9",
          6038 => x"08",
          6039 => x"62",
          6040 => x"76",
          6041 => x"94",
          6042 => x"58",
          6043 => x"77",
          6044 => x"33",
          6045 => x"80",
          6046 => x"ff",
          6047 => x"55",
          6048 => x"77",
          6049 => x"5a",
          6050 => x"84",
          6051 => x"18",
          6052 => x"5a",
          6053 => x"89",
          6054 => x"08",
          6055 => x"33",
          6056 => x"15",
          6057 => x"78",
          6058 => x"5a",
          6059 => x"56",
          6060 => x"70",
          6061 => x"55",
          6062 => x"17",
          6063 => x"b7",
          6064 => x"08",
          6065 => x"88",
          6066 => x"38",
          6067 => x"94",
          6068 => x"c0",
          6069 => x"80",
          6070 => x"75",
          6071 => x"3d",
          6072 => x"80",
          6073 => x"fe",
          6074 => x"84",
          6075 => x"38",
          6076 => x"d8",
          6077 => x"82",
          6078 => x"51",
          6079 => x"08",
          6080 => x"11",
          6081 => x"74",
          6082 => x"17",
          6083 => x"73",
          6084 => x"26",
          6085 => x"33",
          6086 => x"c8",
          6087 => x"38",
          6088 => x"39",
          6089 => x"73",
          6090 => x"c7",
          6091 => x"fe",
          6092 => x"ff",
          6093 => x"08",
          6094 => x"ae",
          6095 => x"9c",
          6096 => x"b9",
          6097 => x"58",
          6098 => x"08",
          6099 => x"08",
          6100 => x"74",
          6101 => x"52",
          6102 => x"b9",
          6103 => x"80",
          6104 => x"fc",
          6105 => x"84",
          6106 => x"38",
          6107 => x"dc",
          6108 => x"80",
          6109 => x"51",
          6110 => x"08",
          6111 => x"11",
          6112 => x"74",
          6113 => x"0c",
          6114 => x"84",
          6115 => x"ff",
          6116 => x"17",
          6117 => x"fe",
          6118 => x"59",
          6119 => x"39",
          6120 => x"fe",
          6121 => x"18",
          6122 => x"0b",
          6123 => x"39",
          6124 => x"81",
          6125 => x"82",
          6126 => x"a8",
          6127 => x"b9",
          6128 => x"80",
          6129 => x"0c",
          6130 => x"3d",
          6131 => x"ff",
          6132 => x"56",
          6133 => x"81",
          6134 => x"06",
          6135 => x"76",
          6136 => x"38",
          6137 => x"06",
          6138 => x"38",
          6139 => x"9a",
          6140 => x"33",
          6141 => x"2e",
          6142 => x"06",
          6143 => x"87",
          6144 => x"83",
          6145 => x"c8",
          6146 => x"ff",
          6147 => x"56",
          6148 => x"84",
          6149 => x"91",
          6150 => x"84",
          6151 => x"84",
          6152 => x"95",
          6153 => x"2b",
          6154 => x"5d",
          6155 => x"08",
          6156 => x"08",
          6157 => x"3d",
          6158 => x"80",
          6159 => x"8b",
          6160 => x"84",
          6161 => x"75",
          6162 => x"5a",
          6163 => x"2e",
          6164 => x"81",
          6165 => x"7b",
          6166 => x"fd",
          6167 => x"3f",
          6168 => x"0c",
          6169 => x"98",
          6170 => x"08",
          6171 => x"33",
          6172 => x"81",
          6173 => x"53",
          6174 => x"fe",
          6175 => x"80",
          6176 => x"75",
          6177 => x"38",
          6178 => x"81",
          6179 => x"7c",
          6180 => x"51",
          6181 => x"08",
          6182 => x"ff",
          6183 => x"06",
          6184 => x"39",
          6185 => x"52",
          6186 => x"3f",
          6187 => x"2e",
          6188 => x"b9",
          6189 => x"08",
          6190 => x"08",
          6191 => x"fe",
          6192 => x"82",
          6193 => x"81",
          6194 => x"05",
          6195 => x"fe",
          6196 => x"39",
          6197 => x"38",
          6198 => x"3f",
          6199 => x"c8",
          6200 => x"b9",
          6201 => x"84",
          6202 => x"38",
          6203 => x"fd",
          6204 => x"38",
          6205 => x"08",
          6206 => x"b0",
          6207 => x"17",
          6208 => x"34",
          6209 => x"38",
          6210 => x"fd",
          6211 => x"fd",
          6212 => x"e3",
          6213 => x"bc",
          6214 => x"c0",
          6215 => x"b9",
          6216 => x"84",
          6217 => x"7d",
          6218 => x"5a",
          6219 => x"08",
          6220 => x"88",
          6221 => x"0d",
          6222 => x"09",
          6223 => x"05",
          6224 => x"58",
          6225 => x"5f",
          6226 => x"ff",
          6227 => x"75",
          6228 => x"38",
          6229 => x"2e",
          6230 => x"ff",
          6231 => x"38",
          6232 => x"33",
          6233 => x"fe",
          6234 => x"56",
          6235 => x"8a",
          6236 => x"08",
          6237 => x"b8",
          6238 => x"80",
          6239 => x"15",
          6240 => x"17",
          6241 => x"38",
          6242 => x"81",
          6243 => x"84",
          6244 => x"18",
          6245 => x"39",
          6246 => x"17",
          6247 => x"fe",
          6248 => x"c8",
          6249 => x"83",
          6250 => x"08",
          6251 => x"fe",
          6252 => x"82",
          6253 => x"75",
          6254 => x"05",
          6255 => x"fe",
          6256 => x"56",
          6257 => x"27",
          6258 => x"27",
          6259 => x"fe",
          6260 => x"5a",
          6261 => x"96",
          6262 => x"fd",
          6263 => x"2e",
          6264 => x"76",
          6265 => x"c8",
          6266 => x"fe",
          6267 => x"77",
          6268 => x"18",
          6269 => x"7b",
          6270 => x"26",
          6271 => x"0c",
          6272 => x"55",
          6273 => x"56",
          6274 => x"f0",
          6275 => x"a0",
          6276 => x"16",
          6277 => x"0b",
          6278 => x"80",
          6279 => x"ce",
          6280 => x"a1",
          6281 => x"0b",
          6282 => x"ff",
          6283 => x"17",
          6284 => x"d3",
          6285 => x"2e",
          6286 => x"80",
          6287 => x"74",
          6288 => x"81",
          6289 => x"ef",
          6290 => x"17",
          6291 => x"06",
          6292 => x"34",
          6293 => x"17",
          6294 => x"80",
          6295 => x"1c",
          6296 => x"84",
          6297 => x"08",
          6298 => x"c8",
          6299 => x"08",
          6300 => x"34",
          6301 => x"6a",
          6302 => x"88",
          6303 => x"33",
          6304 => x"69",
          6305 => x"57",
          6306 => x"fe",
          6307 => x"56",
          6308 => x"0d",
          6309 => x"ec",
          6310 => x"80",
          6311 => x"90",
          6312 => x"7a",
          6313 => x"34",
          6314 => x"b8",
          6315 => x"7b",
          6316 => x"77",
          6317 => x"69",
          6318 => x"57",
          6319 => x"fe",
          6320 => x"56",
          6321 => x"3d",
          6322 => x"79",
          6323 => x"05",
          6324 => x"75",
          6325 => x"38",
          6326 => x"53",
          6327 => x"3d",
          6328 => x"c8",
          6329 => x"2e",
          6330 => x"b1",
          6331 => x"b2",
          6332 => x"59",
          6333 => x"08",
          6334 => x"02",
          6335 => x"5d",
          6336 => x"92",
          6337 => x"75",
          6338 => x"81",
          6339 => x"ef",
          6340 => x"58",
          6341 => x"33",
          6342 => x"15",
          6343 => x"52",
          6344 => x"b9",
          6345 => x"85",
          6346 => x"81",
          6347 => x"0c",
          6348 => x"11",
          6349 => x"74",
          6350 => x"81",
          6351 => x"7a",
          6352 => x"83",
          6353 => x"5f",
          6354 => x"33",
          6355 => x"9f",
          6356 => x"89",
          6357 => x"57",
          6358 => x"26",
          6359 => x"06",
          6360 => x"59",
          6361 => x"85",
          6362 => x"32",
          6363 => x"7a",
          6364 => x"95",
          6365 => x"7b",
          6366 => x"7e",
          6367 => x"24",
          6368 => x"53",
          6369 => x"3d",
          6370 => x"c8",
          6371 => x"b2",
          6372 => x"08",
          6373 => x"77",
          6374 => x"c8",
          6375 => x"92",
          6376 => x"02",
          6377 => x"5a",
          6378 => x"70",
          6379 => x"79",
          6380 => x"8b",
          6381 => x"2a",
          6382 => x"75",
          6383 => x"7f",
          6384 => x"18",
          6385 => x"5c",
          6386 => x"3d",
          6387 => x"9b",
          6388 => x"2b",
          6389 => x"7d",
          6390 => x"9c",
          6391 => x"7d",
          6392 => x"76",
          6393 => x"5e",
          6394 => x"7a",
          6395 => x"aa",
          6396 => x"bc",
          6397 => x"52",
          6398 => x"3f",
          6399 => x"38",
          6400 => x"0c",
          6401 => x"56",
          6402 => x"5a",
          6403 => x"38",
          6404 => x"56",
          6405 => x"2a",
          6406 => x"33",
          6407 => x"93",
          6408 => x"ec",
          6409 => x"80",
          6410 => x"83",
          6411 => x"b2",
          6412 => x"2e",
          6413 => x"fb",
          6414 => x"84",
          6415 => x"16",
          6416 => x"b4",
          6417 => x"16",
          6418 => x"09",
          6419 => x"76",
          6420 => x"51",
          6421 => x"08",
          6422 => x"58",
          6423 => x"aa",
          6424 => x"34",
          6425 => x"08",
          6426 => x"51",
          6427 => x"08",
          6428 => x"ff",
          6429 => x"f9",
          6430 => x"38",
          6431 => x"b9",
          6432 => x"3d",
          6433 => x"0c",
          6434 => x"94",
          6435 => x"2b",
          6436 => x"8d",
          6437 => x"fb",
          6438 => x"2e",
          6439 => x"0c",
          6440 => x"16",
          6441 => x"51",
          6442 => x"b9",
          6443 => x"fe",
          6444 => x"17",
          6445 => x"31",
          6446 => x"a0",
          6447 => x"16",
          6448 => x"06",
          6449 => x"08",
          6450 => x"81",
          6451 => x"79",
          6452 => x"17",
          6453 => x"18",
          6454 => x"81",
          6455 => x"38",
          6456 => x"b4",
          6457 => x"b9",
          6458 => x"08",
          6459 => x"5d",
          6460 => x"81",
          6461 => x"18",
          6462 => x"33",
          6463 => x"fb",
          6464 => x"df",
          6465 => x"05",
          6466 => x"cc",
          6467 => x"d8",
          6468 => x"b9",
          6469 => x"84",
          6470 => x"78",
          6471 => x"51",
          6472 => x"08",
          6473 => x"02",
          6474 => x"54",
          6475 => x"06",
          6476 => x"06",
          6477 => x"55",
          6478 => x"0b",
          6479 => x"9a",
          6480 => x"c8",
          6481 => x"0d",
          6482 => x"05",
          6483 => x"3f",
          6484 => x"c8",
          6485 => x"b9",
          6486 => x"5a",
          6487 => x"ff",
          6488 => x"55",
          6489 => x"80",
          6490 => x"86",
          6491 => x"22",
          6492 => x"59",
          6493 => x"88",
          6494 => x"90",
          6495 => x"98",
          6496 => x"57",
          6497 => x"fe",
          6498 => x"84",
          6499 => x"e8",
          6500 => x"53",
          6501 => x"51",
          6502 => x"08",
          6503 => x"b9",
          6504 => x"57",
          6505 => x"76",
          6506 => x"76",
          6507 => x"5b",
          6508 => x"70",
          6509 => x"81",
          6510 => x"56",
          6511 => x"82",
          6512 => x"55",
          6513 => x"98",
          6514 => x"52",
          6515 => x"3f",
          6516 => x"38",
          6517 => x"0c",
          6518 => x"33",
          6519 => x"2e",
          6520 => x"2e",
          6521 => x"05",
          6522 => x"90",
          6523 => x"33",
          6524 => x"71",
          6525 => x"59",
          6526 => x"3d",
          6527 => x"52",
          6528 => x"8b",
          6529 => x"b9",
          6530 => x"76",
          6531 => x"38",
          6532 => x"39",
          6533 => x"16",
          6534 => x"fe",
          6535 => x"c8",
          6536 => x"e8",
          6537 => x"34",
          6538 => x"84",
          6539 => x"17",
          6540 => x"33",
          6541 => x"fe",
          6542 => x"a0",
          6543 => x"16",
          6544 => x"59",
          6545 => x"81",
          6546 => x"84",
          6547 => x"38",
          6548 => x"fe",
          6549 => x"57",
          6550 => x"84",
          6551 => x"66",
          6552 => x"7c",
          6553 => x"34",
          6554 => x"38",
          6555 => x"34",
          6556 => x"18",
          6557 => x"79",
          6558 => x"79",
          6559 => x"82",
          6560 => x"a2",
          6561 => x"b9",
          6562 => x"82",
          6563 => x"57",
          6564 => x"34",
          6565 => x"a3",
          6566 => x"06",
          6567 => x"81",
          6568 => x"5c",
          6569 => x"55",
          6570 => x"74",
          6571 => x"74",
          6572 => x"84",
          6573 => x"84",
          6574 => x"57",
          6575 => x"e6",
          6576 => x"81",
          6577 => x"2e",
          6578 => x"2e",
          6579 => x"81",
          6580 => x"2e",
          6581 => x"06",
          6582 => x"78",
          6583 => x"81",
          6584 => x"38",
          6585 => x"88",
          6586 => x"5d",
          6587 => x"81",
          6588 => x"08",
          6589 => x"58",
          6590 => x"38",
          6591 => x"81",
          6592 => x"99",
          6593 => x"70",
          6594 => x"81",
          6595 => x"ed",
          6596 => x"95",
          6597 => x"3f",
          6598 => x"c8",
          6599 => x"75",
          6600 => x"04",
          6601 => x"3f",
          6602 => x"06",
          6603 => x"75",
          6604 => x"04",
          6605 => x"39",
          6606 => x"3f",
          6607 => x"c8",
          6608 => x"82",
          6609 => x"55",
          6610 => x"70",
          6611 => x"74",
          6612 => x"1e",
          6613 => x"84",
          6614 => x"87",
          6615 => x"86",
          6616 => x"08",
          6617 => x"38",
          6618 => x"38",
          6619 => x"fe",
          6620 => x"57",
          6621 => x"81",
          6622 => x"08",
          6623 => x"57",
          6624 => x"b2",
          6625 => x"2e",
          6626 => x"54",
          6627 => x"33",
          6628 => x"c8",
          6629 => x"81",
          6630 => x"78",
          6631 => x"33",
          6632 => x"81",
          6633 => x"78",
          6634 => x"d7",
          6635 => x"a5",
          6636 => x"a1",
          6637 => x"b9",
          6638 => x"87",
          6639 => x"76",
          6640 => x"57",
          6641 => x"34",
          6642 => x"56",
          6643 => x"7e",
          6644 => x"58",
          6645 => x"ff",
          6646 => x"38",
          6647 => x"70",
          6648 => x"74",
          6649 => x"e5",
          6650 => x"1e",
          6651 => x"84",
          6652 => x"81",
          6653 => x"18",
          6654 => x"51",
          6655 => x"08",
          6656 => x"38",
          6657 => x"b4",
          6658 => x"7b",
          6659 => x"18",
          6660 => x"84",
          6661 => x"74",
          6662 => x"d1",
          6663 => x"b9",
          6664 => x"fe",
          6665 => x"80",
          6666 => x"81",
          6667 => x"05",
          6668 => x"fe",
          6669 => x"3d",
          6670 => x"cb",
          6671 => x"76",
          6672 => x"74",
          6673 => x"73",
          6674 => x"84",
          6675 => x"81",
          6676 => x"81",
          6677 => x"81",
          6678 => x"38",
          6679 => x"17",
          6680 => x"5d",
          6681 => x"8a",
          6682 => x"7c",
          6683 => x"3f",
          6684 => x"72",
          6685 => x"05",
          6686 => x"55",
          6687 => x"19",
          6688 => x"77",
          6689 => x"76",
          6690 => x"7f",
          6691 => x"83",
          6692 => x"81",
          6693 => x"08",
          6694 => x"c8",
          6695 => x"78",
          6696 => x"09",
          6697 => x"54",
          6698 => x"0d",
          6699 => x"90",
          6700 => x"fe",
          6701 => x"81",
          6702 => x"77",
          6703 => x"80",
          6704 => x"58",
          6705 => x"54",
          6706 => x"53",
          6707 => x"3f",
          6708 => x"c8",
          6709 => x"ff",
          6710 => x"7e",
          6711 => x"2e",
          6712 => x"79",
          6713 => x"c0",
          6714 => x"15",
          6715 => x"5a",
          6716 => x"7d",
          6717 => x"81",
          6718 => x"54",
          6719 => x"39",
          6720 => x"82",
          6721 => x"c0",
          6722 => x"84",
          6723 => x"3d",
          6724 => x"81",
          6725 => x"0b",
          6726 => x"79",
          6727 => x"81",
          6728 => x"56",
          6729 => x"ed",
          6730 => x"84",
          6731 => x"84",
          6732 => x"90",
          6733 => x"2e",
          6734 => x"84",
          6735 => x"12",
          6736 => x"51",
          6737 => x"08",
          6738 => x"56",
          6739 => x"82",
          6740 => x"84",
          6741 => x"83",
          6742 => x"84",
          6743 => x"55",
          6744 => x"82",
          6745 => x"15",
          6746 => x"7e",
          6747 => x"26",
          6748 => x"26",
          6749 => x"55",
          6750 => x"a6",
          6751 => x"77",
          6752 => x"85",
          6753 => x"77",
          6754 => x"b0",
          6755 => x"81",
          6756 => x"fe",
          6757 => x"c8",
          6758 => x"05",
          6759 => x"88",
          6760 => x"82",
          6761 => x"f8",
          6762 => x"b2",
          6763 => x"82",
          6764 => x"33",
          6765 => x"88",
          6766 => x"07",
          6767 => x"ba",
          6768 => x"71",
          6769 => x"14",
          6770 => x"33",
          6771 => x"a3",
          6772 => x"54",
          6773 => x"4d",
          6774 => x"90",
          6775 => x"82",
          6776 => x"06",
          6777 => x"38",
          6778 => x"89",
          6779 => x"f4",
          6780 => x"43",
          6781 => x"38",
          6782 => x"81",
          6783 => x"74",
          6784 => x"98",
          6785 => x"82",
          6786 => x"80",
          6787 => x"38",
          6788 => x"3f",
          6789 => x"55",
          6790 => x"96",
          6791 => x"10",
          6792 => x"72",
          6793 => x"ff",
          6794 => x"47",
          6795 => x"11",
          6796 => x"58",
          6797 => x"b8",
          6798 => x"16",
          6799 => x"26",
          6800 => x"31",
          6801 => x"fd",
          6802 => x"40",
          6803 => x"82",
          6804 => x"83",
          6805 => x"27",
          6806 => x"77",
          6807 => x"ef",
          6808 => x"57",
          6809 => x"0d",
          6810 => x"fb",
          6811 => x"0c",
          6812 => x"04",
          6813 => x"06",
          6814 => x"38",
          6815 => x"05",
          6816 => x"38",
          6817 => x"7d",
          6818 => x"05",
          6819 => x"33",
          6820 => x"99",
          6821 => x"ff",
          6822 => x"64",
          6823 => x"81",
          6824 => x"9f",
          6825 => x"81",
          6826 => x"75",
          6827 => x"9f",
          6828 => x"80",
          6829 => x"1f",
          6830 => x"38",
          6831 => x"f8",
          6832 => x"ca",
          6833 => x"08",
          6834 => x"06",
          6835 => x"83",
          6836 => x"7e",
          6837 => x"31",
          6838 => x"d2",
          6839 => x"7b",
          6840 => x"39",
          6841 => x"80",
          6842 => x"30",
          6843 => x"b9",
          6844 => x"7a",
          6845 => x"7b",
          6846 => x"84",
          6847 => x"b9",
          6848 => x"2e",
          6849 => x"8b",
          6850 => x"7a",
          6851 => x"55",
          6852 => x"ff",
          6853 => x"83",
          6854 => x"81",
          6855 => x"58",
          6856 => x"60",
          6857 => x"61",
          6858 => x"34",
          6859 => x"61",
          6860 => x"7b",
          6861 => x"05",
          6862 => x"48",
          6863 => x"2a",
          6864 => x"34",
          6865 => x"86",
          6866 => x"55",
          6867 => x"2a",
          6868 => x"61",
          6869 => x"34",
          6870 => x"9a",
          6871 => x"7e",
          6872 => x"48",
          6873 => x"2a",
          6874 => x"98",
          6875 => x"d4",
          6876 => x"2e",
          6877 => x"34",
          6878 => x"a9",
          6879 => x"34",
          6880 => x"61",
          6881 => x"6a",
          6882 => x"a4",
          6883 => x"93",
          6884 => x"57",
          6885 => x"76",
          6886 => x"55",
          6887 => x"49",
          6888 => x"05",
          6889 => x"7e",
          6890 => x"8f",
          6891 => x"fa",
          6892 => x"2e",
          6893 => x"80",
          6894 => x"15",
          6895 => x"5b",
          6896 => x"ff",
          6897 => x"38",
          6898 => x"2a",
          6899 => x"05",
          6900 => x"64",
          6901 => x"2a",
          6902 => x"59",
          6903 => x"78",
          6904 => x"fe",
          6905 => x"85",
          6906 => x"80",
          6907 => x"15",
          6908 => x"7a",
          6909 => x"81",
          6910 => x"38",
          6911 => x"66",
          6912 => x"38",
          6913 => x"52",
          6914 => x"b9",
          6915 => x"76",
          6916 => x"8c",
          6917 => x"58",
          6918 => x"84",
          6919 => x"58",
          6920 => x"81",
          6921 => x"80",
          6922 => x"05",
          6923 => x"38",
          6924 => x"34",
          6925 => x"34",
          6926 => x"82",
          6927 => x"77",
          6928 => x"fd",
          6929 => x"9a",
          6930 => x"b9",
          6931 => x"76",
          6932 => x"08",
          6933 => x"c6",
          6934 => x"34",
          6935 => x"b9",
          6936 => x"62",
          6937 => x"2a",
          6938 => x"62",
          6939 => x"05",
          6940 => x"83",
          6941 => x"60",
          6942 => x"81",
          6943 => x"38",
          6944 => x"c3",
          6945 => x"08",
          6946 => x"84",
          6947 => x"b9",
          6948 => x"39",
          6949 => x"c4",
          6950 => x"57",
          6951 => x"58",
          6952 => x"26",
          6953 => x"10",
          6954 => x"74",
          6955 => x"ee",
          6956 => x"c2",
          6957 => x"84",
          6958 => x"a0",
          6959 => x"fc",
          6960 => x"f0",
          6961 => x"57",
          6962 => x"83",
          6963 => x"f8",
          6964 => x"f4",
          6965 => x"68",
          6966 => x"af",
          6967 => x"61",
          6968 => x"68",
          6969 => x"5b",
          6970 => x"2a",
          6971 => x"c6",
          6972 => x"80",
          6973 => x"80",
          6974 => x"c6",
          6975 => x"7c",
          6976 => x"34",
          6977 => x"05",
          6978 => x"a7",
          6979 => x"80",
          6980 => x"05",
          6981 => x"61",
          6982 => x"34",
          6983 => x"b3",
          6984 => x"05",
          6985 => x"93",
          6986 => x"59",
          6987 => x"33",
          6988 => x"15",
          6989 => x"76",
          6990 => x"81",
          6991 => x"da",
          6992 => x"53",
          6993 => x"3f",
          6994 => x"b0",
          6995 => x"77",
          6996 => x"84",
          6997 => x"51",
          6998 => x"81",
          6999 => x"0d",
          7000 => x"34",
          7001 => x"4c",
          7002 => x"34",
          7003 => x"34",
          7004 => x"86",
          7005 => x"ff",
          7006 => x"05",
          7007 => x"65",
          7008 => x"54",
          7009 => x"fe",
          7010 => x"57",
          7011 => x"ff",
          7012 => x"80",
          7013 => x"7b",
          7014 => x"57",
          7015 => x"57",
          7016 => x"61",
          7017 => x"83",
          7018 => x"e6",
          7019 => x"05",
          7020 => x"83",
          7021 => x"78",
          7022 => x"2a",
          7023 => x"7a",
          7024 => x"05",
          7025 => x"76",
          7026 => x"83",
          7027 => x"05",
          7028 => x"6b",
          7029 => x"52",
          7030 => x"54",
          7031 => x"fe",
          7032 => x"f7",
          7033 => x"5b",
          7034 => x"57",
          7035 => x"3d",
          7036 => x"53",
          7037 => x"3f",
          7038 => x"38",
          7039 => x"90",
          7040 => x"34",
          7041 => x"38",
          7042 => x"34",
          7043 => x"74",
          7044 => x"04",
          7045 => x"b3",
          7046 => x"80",
          7047 => x"76",
          7048 => x"17",
          7049 => x"81",
          7050 => x"74",
          7051 => x"0c",
          7052 => x"05",
          7053 => x"08",
          7054 => x"32",
          7055 => x"70",
          7056 => x"1b",
          7057 => x"52",
          7058 => x"39",
          7059 => x"33",
          7060 => x"57",
          7061 => x"34",
          7062 => x"3d",
          7063 => x"f7",
          7064 => x"c0",
          7065 => x"59",
          7066 => x"bb",
          7067 => x"81",
          7068 => x"75",
          7069 => x"11",
          7070 => x"08",
          7071 => x"c8",
          7072 => x"38",
          7073 => x"3d",
          7074 => x"55",
          7075 => x"51",
          7076 => x"70",
          7077 => x"30",
          7078 => x"8d",
          7079 => x"81",
          7080 => x"3d",
          7081 => x"84",
          7082 => x"52",
          7083 => x"83",
          7084 => x"c8",
          7085 => x"ff",
          7086 => x"09",
          7087 => x"e4",
          7088 => x"71",
          7089 => x"ff",
          7090 => x"26",
          7091 => x"05",
          7092 => x"80",
          7093 => x"c8",
          7094 => x"3d",
          7095 => x"05",
          7096 => x"70",
          7097 => x"72",
          7098 => x"04",
          7099 => x"ef",
          7100 => x"70",
          7101 => x"84",
          7102 => x"04",
          7103 => x"ff",
          7104 => x"ff",
          7105 => x"75",
          7106 => x"70",
          7107 => x"70",
          7108 => x"56",
          7109 => x"82",
          7110 => x"54",
          7111 => x"54",
          7112 => x"38",
          7113 => x"52",
          7114 => x"75",
          7115 => x"80",
          7116 => x"b9",
          7117 => x"ed",
          7118 => x"26",
          7119 => x"e0",
          7120 => x"16",
          7121 => x"75",
          7122 => x"83",
          7123 => x"88",
          7124 => x"51",
          7125 => x"ff",
          7126 => x"70",
          7127 => x"39",
          7128 => x"57",
          7129 => x"ff",
          7130 => x"75",
          7131 => x"70",
          7132 => x"ff",
          7133 => x"05",
          7134 => x"00",
          7135 => x"ff",
          7136 => x"ff",
          7137 => x"19",
          7138 => x"19",
          7139 => x"19",
          7140 => x"19",
          7141 => x"19",
          7142 => x"19",
          7143 => x"18",
          7144 => x"18",
          7145 => x"18",
          7146 => x"18",
          7147 => x"1f",
          7148 => x"1f",
          7149 => x"1f",
          7150 => x"1f",
          7151 => x"1f",
          7152 => x"1f",
          7153 => x"1f",
          7154 => x"1f",
          7155 => x"1f",
          7156 => x"1f",
          7157 => x"1f",
          7158 => x"1f",
          7159 => x"1f",
          7160 => x"1f",
          7161 => x"1f",
          7162 => x"1f",
          7163 => x"1f",
          7164 => x"1f",
          7165 => x"1f",
          7166 => x"1f",
          7167 => x"1f",
          7168 => x"24",
          7169 => x"1f",
          7170 => x"1f",
          7171 => x"1f",
          7172 => x"1f",
          7173 => x"1f",
          7174 => x"1f",
          7175 => x"1f",
          7176 => x"1f",
          7177 => x"23",
          7178 => x"22",
          7179 => x"23",
          7180 => x"21",
          7181 => x"1f",
          7182 => x"1f",
          7183 => x"1f",
          7184 => x"1f",
          7185 => x"1f",
          7186 => x"1f",
          7187 => x"1f",
          7188 => x"1f",
          7189 => x"1f",
          7190 => x"1f",
          7191 => x"1f",
          7192 => x"1f",
          7193 => x"1f",
          7194 => x"1f",
          7195 => x"1f",
          7196 => x"1f",
          7197 => x"1f",
          7198 => x"1f",
          7199 => x"1f",
          7200 => x"1f",
          7201 => x"1f",
          7202 => x"1f",
          7203 => x"1f",
          7204 => x"1f",
          7205 => x"1f",
          7206 => x"1f",
          7207 => x"21",
          7208 => x"1f",
          7209 => x"1f",
          7210 => x"1f",
          7211 => x"1f",
          7212 => x"21",
          7213 => x"21",
          7214 => x"21",
          7215 => x"21",
          7216 => x"32",
          7217 => x"32",
          7218 => x"32",
          7219 => x"3a",
          7220 => x"36",
          7221 => x"34",
          7222 => x"36",
          7223 => x"36",
          7224 => x"39",
          7225 => x"39",
          7226 => x"37",
          7227 => x"34",
          7228 => x"36",
          7229 => x"36",
          7230 => x"46",
          7231 => x"46",
          7232 => x"47",
          7233 => x"47",
          7234 => x"47",
          7235 => x"47",
          7236 => x"47",
          7237 => x"47",
          7238 => x"47",
          7239 => x"47",
          7240 => x"47",
          7241 => x"47",
          7242 => x"47",
          7243 => x"47",
          7244 => x"47",
          7245 => x"47",
          7246 => x"47",
          7247 => x"47",
          7248 => x"48",
          7249 => x"48",
          7250 => x"47",
          7251 => x"48",
          7252 => x"47",
          7253 => x"48",
          7254 => x"47",
          7255 => x"47",
          7256 => x"47",
          7257 => x"47",
          7258 => x"54",
          7259 => x"55",
          7260 => x"54",
          7261 => x"54",
          7262 => x"52",
          7263 => x"57",
          7264 => x"52",
          7265 => x"52",
          7266 => x"52",
          7267 => x"57",
          7268 => x"52",
          7269 => x"52",
          7270 => x"52",
          7271 => x"52",
          7272 => x"52",
          7273 => x"52",
          7274 => x"52",
          7275 => x"52",
          7276 => x"52",
          7277 => x"52",
          7278 => x"52",
          7279 => x"52",
          7280 => x"53",
          7281 => x"52",
          7282 => x"52",
          7283 => x"53",
          7284 => x"53",
          7285 => x"59",
          7286 => x"59",
          7287 => x"59",
          7288 => x"58",
          7289 => x"59",
          7290 => x"59",
          7291 => x"59",
          7292 => x"59",
          7293 => x"59",
          7294 => x"59",
          7295 => x"59",
          7296 => x"59",
          7297 => x"59",
          7298 => x"59",
          7299 => x"59",
          7300 => x"5a",
          7301 => x"59",
          7302 => x"5a",
          7303 => x"5a",
          7304 => x"5a",
          7305 => x"5a",
          7306 => x"5a",
          7307 => x"59",
          7308 => x"59",
          7309 => x"59",
          7310 => x"61",
          7311 => x"61",
          7312 => x"61",
          7313 => x"61",
          7314 => x"61",
          7315 => x"61",
          7316 => x"61",
          7317 => x"61",
          7318 => x"61",
          7319 => x"61",
          7320 => x"63",
          7321 => x"61",
          7322 => x"61",
          7323 => x"5e",
          7324 => x"de",
          7325 => x"de",
          7326 => x"de",
          7327 => x"de",
          7328 => x"de",
          7329 => x"0b",
          7330 => x"0f",
          7331 => x"0b",
          7332 => x"0b",
          7333 => x"0b",
          7334 => x"0d",
          7335 => x"0f",
          7336 => x"0b",
          7337 => x"0b",
          7338 => x"0b",
          7339 => x"0b",
          7340 => x"0b",
          7341 => x"0b",
          7342 => x"0b",
          7343 => x"0b",
          7344 => x"0b",
          7345 => x"0b",
          7346 => x"0b",
          7347 => x"0b",
          7348 => x"0b",
          7349 => x"0b",
          7350 => x"0b",
          7351 => x"0b",
          7352 => x"0b",
          7353 => x"0b",
          7354 => x"0f",
          7355 => x"0b",
          7356 => x"0b",
          7357 => x"0b",
          7358 => x"0b",
          7359 => x"0b",
          7360 => x"0b",
          7361 => x"0b",
          7362 => x"0e",
          7363 => x"0e",
          7364 => x"0e",
          7365 => x"0e",
          7366 => x"0b",
          7367 => x"0b",
          7368 => x"0c",
          7369 => x"0b",
          7370 => x"0f",
          7371 => x"0c",
          7372 => x"0b",
          7373 => x"6e",
          7374 => x"6f",
          7375 => x"6e",
          7376 => x"6f",
          7377 => x"78",
          7378 => x"6c",
          7379 => x"6f",
          7380 => x"69",
          7381 => x"75",
          7382 => x"62",
          7383 => x"77",
          7384 => x"65",
          7385 => x"65",
          7386 => x"00",
          7387 => x"73",
          7388 => x"73",
          7389 => x"66",
          7390 => x"73",
          7391 => x"73",
          7392 => x"61",
          7393 => x"61",
          7394 => x"6c",
          7395 => x"00",
          7396 => x"6e",
          7397 => x"00",
          7398 => x"74",
          7399 => x"6f",
          7400 => x"00",
          7401 => x"6e",
          7402 => x"66",
          7403 => x"00",
          7404 => x"69",
          7405 => x"65",
          7406 => x"00",
          7407 => x"73",
          7408 => x"2e",
          7409 => x"74",
          7410 => x"74",
          7411 => x"63",
          7412 => x"00",
          7413 => x"20",
          7414 => x"2e",
          7415 => x"70",
          7416 => x"66",
          7417 => x"65",
          7418 => x"20",
          7419 => x"2e",
          7420 => x"6f",
          7421 => x"65",
          7422 => x"69",
          7423 => x"65",
          7424 => x"76",
          7425 => x"00",
          7426 => x"77",
          7427 => x"6f",
          7428 => x"00",
          7429 => x"61",
          7430 => x"76",
          7431 => x"00",
          7432 => x"6c",
          7433 => x"78",
          7434 => x"00",
          7435 => x"20",
          7436 => x"00",
          7437 => x"64",
          7438 => x"6d",
          7439 => x"20",
          7440 => x"75",
          7441 => x"20",
          7442 => x"75",
          7443 => x"73",
          7444 => x"65",
          7445 => x"74",
          7446 => x"72",
          7447 => x"73",
          7448 => x"00",
          7449 => x"73",
          7450 => x"6c",
          7451 => x"20",
          7452 => x"6c",
          7453 => x"2f",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"32",
          7458 => x"00",
          7459 => x"00",
          7460 => x"00",
          7461 => x"20",
          7462 => x"53",
          7463 => x"28",
          7464 => x"32",
          7465 => x"2e",
          7466 => x"50",
          7467 => x"25",
          7468 => x"20",
          7469 => x"00",
          7470 => x"20",
          7471 => x"64",
          7472 => x"20",
          7473 => x"20",
          7474 => x"6c",
          7475 => x"20",
          7476 => x"64",
          7477 => x"20",
          7478 => x"20",
          7479 => x"6c",
          7480 => x"55",
          7481 => x"75",
          7482 => x"6c",
          7483 => x"52",
          7484 => x"6e",
          7485 => x"00",
          7486 => x"52",
          7487 => x"72",
          7488 => x"52",
          7489 => x"6e",
          7490 => x"00",
          7491 => x"52",
          7492 => x"72",
          7493 => x"43",
          7494 => x"6e",
          7495 => x"00",
          7496 => x"52",
          7497 => x"72",
          7498 => x"32",
          7499 => x"75",
          7500 => x"6d",
          7501 => x"72",
          7502 => x"74",
          7503 => x"20",
          7504 => x"2e",
          7505 => x"6e",
          7506 => x"2e",
          7507 => x"74",
          7508 => x"61",
          7509 => x"53",
          7510 => x"74",
          7511 => x"20",
          7512 => x"69",
          7513 => x"64",
          7514 => x"2c",
          7515 => x"20",
          7516 => x"6e",
          7517 => x"00",
          7518 => x"3a",
          7519 => x"00",
          7520 => x"6d",
          7521 => x"00",
          7522 => x"6e",
          7523 => x"5c",
          7524 => x"00",
          7525 => x"65",
          7526 => x"2e",
          7527 => x"73",
          7528 => x"20",
          7529 => x"74",
          7530 => x"00",
          7531 => x"67",
          7532 => x"20",
          7533 => x"2e",
          7534 => x"6c",
          7535 => x"6e",
          7536 => x"20",
          7537 => x"00",
          7538 => x"69",
          7539 => x"20",
          7540 => x"20",
          7541 => x"38",
          7542 => x"58",
          7543 => x"38",
          7544 => x"2d",
          7545 => x"69",
          7546 => x"00",
          7547 => x"25",
          7548 => x"30",
          7549 => x"78",
          7550 => x"70",
          7551 => x"00",
          7552 => x"25",
          7553 => x"65",
          7554 => x"2e",
          7555 => x"6d",
          7556 => x"79",
          7557 => x"65",
          7558 => x"3a",
          7559 => x"00",
          7560 => x"20",
          7561 => x"65",
          7562 => x"6f",
          7563 => x"73",
          7564 => x"6e",
          7565 => x"3f",
          7566 => x"25",
          7567 => x"3a",
          7568 => x"0a",
          7569 => x"6e",
          7570 => x"69",
          7571 => x"44",
          7572 => x"69",
          7573 => x"74",
          7574 => x"64",
          7575 => x"00",
          7576 => x"55",
          7577 => x"56",
          7578 => x"64",
          7579 => x"20",
          7580 => x"00",
          7581 => x"55",
          7582 => x"20",
          7583 => x"64",
          7584 => x"20",
          7585 => x"00",
          7586 => x"61",
          7587 => x"74",
          7588 => x"73",
          7589 => x"20",
          7590 => x"00",
          7591 => x"00",
          7592 => x"55",
          7593 => x"20",
          7594 => x"20",
          7595 => x"20",
          7596 => x"00",
          7597 => x"73",
          7598 => x"63",
          7599 => x"20",
          7600 => x"20",
          7601 => x"4d",
          7602 => x"20",
          7603 => x"6e",
          7604 => x"20",
          7605 => x"72",
          7606 => x"25",
          7607 => x"00",
          7608 => x"52",
          7609 => x"6b",
          7610 => x"20",
          7611 => x"20",
          7612 => x"4d",
          7613 => x"20",
          7614 => x"20",
          7615 => x"20",
          7616 => x"00",
          7617 => x"20",
          7618 => x"20",
          7619 => x"4e",
          7620 => x"00",
          7621 => x"54",
          7622 => x"28",
          7623 => x"73",
          7624 => x"0a",
          7625 => x"4d",
          7626 => x"28",
          7627 => x"20",
          7628 => x"0a",
          7629 => x"20",
          7630 => x"28",
          7631 => x"20",
          7632 => x"0a",
          7633 => x"4d",
          7634 => x"28",
          7635 => x"38",
          7636 => x"20",
          7637 => x"20",
          7638 => x"58",
          7639 => x"0a",
          7640 => x"53",
          7641 => x"28",
          7642 => x"38",
          7643 => x"20",
          7644 => x"20",
          7645 => x"58",
          7646 => x"0a",
          7647 => x"20",
          7648 => x"28",
          7649 => x"38",
          7650 => x"66",
          7651 => x"20",
          7652 => x"00",
          7653 => x"6e",
          7654 => x"00",
          7655 => x"00",
          7656 => x"00",
          7657 => x"00",
          7658 => x"f0",
          7659 => x"00",
          7660 => x"00",
          7661 => x"f0",
          7662 => x"00",
          7663 => x"00",
          7664 => x"f0",
          7665 => x"00",
          7666 => x"00",
          7667 => x"f0",
          7668 => x"00",
          7669 => x"00",
          7670 => x"f0",
          7671 => x"00",
          7672 => x"00",
          7673 => x"f0",
          7674 => x"00",
          7675 => x"00",
          7676 => x"f0",
          7677 => x"00",
          7678 => x"00",
          7679 => x"f0",
          7680 => x"00",
          7681 => x"00",
          7682 => x"f0",
          7683 => x"00",
          7684 => x"00",
          7685 => x"f0",
          7686 => x"00",
          7687 => x"00",
          7688 => x"f0",
          7689 => x"00",
          7690 => x"00",
          7691 => x"44",
          7692 => x"42",
          7693 => x"36",
          7694 => x"34",
          7695 => x"33",
          7696 => x"31",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"6e",
          7703 => x"6e",
          7704 => x"20",
          7705 => x"20",
          7706 => x"69",
          7707 => x"2e",
          7708 => x"79",
          7709 => x"00",
          7710 => x"36",
          7711 => x"00",
          7712 => x"20",
          7713 => x"74",
          7714 => x"73",
          7715 => x"6c",
          7716 => x"46",
          7717 => x"73",
          7718 => x"31",
          7719 => x"41",
          7720 => x"43",
          7721 => x"31",
          7722 => x"31",
          7723 => x"31",
          7724 => x"31",
          7725 => x"31",
          7726 => x"31",
          7727 => x"31",
          7728 => x"31",
          7729 => x"31",
          7730 => x"32",
          7731 => x"32",
          7732 => x"33",
          7733 => x"46",
          7734 => x"00",
          7735 => x"00",
          7736 => x"64",
          7737 => x"25",
          7738 => x"32",
          7739 => x"25",
          7740 => x"3a",
          7741 => x"64",
          7742 => x"2c",
          7743 => x"00",
          7744 => x"00",
          7745 => x"25",
          7746 => x"70",
          7747 => x"73",
          7748 => x"3a",
          7749 => x"32",
          7750 => x"3a",
          7751 => x"32",
          7752 => x"3a",
          7753 => x"00",
          7754 => x"74",
          7755 => x"64",
          7756 => x"00",
          7757 => x"7c",
          7758 => x"3b",
          7759 => x"54",
          7760 => x"00",
          7761 => x"4f",
          7762 => x"20",
          7763 => x"20",
          7764 => x"20",
          7765 => x"45",
          7766 => x"33",
          7767 => x"f2",
          7768 => x"00",
          7769 => x"05",
          7770 => x"18",
          7771 => x"45",
          7772 => x"45",
          7773 => x"92",
          7774 => x"9a",
          7775 => x"4f",
          7776 => x"aa",
          7777 => x"b2",
          7778 => x"ba",
          7779 => x"c2",
          7780 => x"ca",
          7781 => x"d2",
          7782 => x"da",
          7783 => x"e2",
          7784 => x"ea",
          7785 => x"f2",
          7786 => x"fa",
          7787 => x"2c",
          7788 => x"2a",
          7789 => x"00",
          7790 => x"00",
          7791 => x"00",
          7792 => x"00",
          7793 => x"00",
          7794 => x"00",
          7795 => x"00",
          7796 => x"00",
          7797 => x"00",
          7798 => x"00",
          7799 => x"00",
          7800 => x"00",
          7801 => x"01",
          7802 => x"00",
          7803 => x"00",
          7804 => x"00",
          7805 => x"00",
          7806 => x"25",
          7807 => x"25",
          7808 => x"25",
          7809 => x"25",
          7810 => x"25",
          7811 => x"25",
          7812 => x"25",
          7813 => x"25",
          7814 => x"25",
          7815 => x"25",
          7816 => x"25",
          7817 => x"25",
          7818 => x"03",
          7819 => x"03",
          7820 => x"03",
          7821 => x"22",
          7822 => x"22",
          7823 => x"22",
          7824 => x"22",
          7825 => x"00",
          7826 => x"03",
          7827 => x"00",
          7828 => x"01",
          7829 => x"01",
          7830 => x"01",
          7831 => x"01",
          7832 => x"01",
          7833 => x"01",
          7834 => x"01",
          7835 => x"01",
          7836 => x"01",
          7837 => x"02",
          7838 => x"02",
          7839 => x"01",
          7840 => x"01",
          7841 => x"01",
          7842 => x"01",
          7843 => x"01",
          7844 => x"01",
          7845 => x"01",
          7846 => x"01",
          7847 => x"01",
          7848 => x"01",
          7849 => x"01",
          7850 => x"01",
          7851 => x"01",
          7852 => x"01",
          7853 => x"01",
          7854 => x"00",
          7855 => x"02",
          7856 => x"02",
          7857 => x"02",
          7858 => x"02",
          7859 => x"01",
          7860 => x"02",
          7861 => x"02",
          7862 => x"02",
          7863 => x"01",
          7864 => x"02",
          7865 => x"02",
          7866 => x"01",
          7867 => x"02",
          7868 => x"2c",
          7869 => x"02",
          7870 => x"02",
          7871 => x"02",
          7872 => x"02",
          7873 => x"02",
          7874 => x"03",
          7875 => x"00",
          7876 => x"03",
          7877 => x"00",
          7878 => x"03",
          7879 => x"03",
          7880 => x"03",
          7881 => x"03",
          7882 => x"03",
          7883 => x"04",
          7884 => x"04",
          7885 => x"04",
          7886 => x"04",
          7887 => x"04",
          7888 => x"00",
          7889 => x"1e",
          7890 => x"1f",
          7891 => x"1f",
          7892 => x"1f",
          7893 => x"1f",
          7894 => x"1f",
          7895 => x"00",
          7896 => x"1f",
          7897 => x"1f",
          7898 => x"1f",
          7899 => x"06",
          7900 => x"06",
          7901 => x"1f",
          7902 => x"00",
          7903 => x"1f",
          7904 => x"1f",
          7905 => x"21",
          7906 => x"02",
          7907 => x"24",
          7908 => x"2c",
          7909 => x"2c",
          7910 => x"2d",
          7911 => x"00",
          7912 => x"e6",
          7913 => x"00",
          7914 => x"e6",
          7915 => x"00",
          7916 => x"e6",
          7917 => x"00",
          7918 => x"e6",
          7919 => x"00",
          7920 => x"e6",
          7921 => x"00",
          7922 => x"e6",
          7923 => x"00",
          7924 => x"e6",
          7925 => x"00",
          7926 => x"e6",
          7927 => x"00",
          7928 => x"e6",
          7929 => x"00",
          7930 => x"e6",
          7931 => x"00",
          7932 => x"e6",
          7933 => x"00",
          7934 => x"e6",
          7935 => x"00",
          7936 => x"e6",
          7937 => x"00",
          7938 => x"e6",
          7939 => x"00",
          7940 => x"e6",
          7941 => x"00",
          7942 => x"e6",
          7943 => x"00",
          7944 => x"e6",
          7945 => x"00",
          7946 => x"e6",
          7947 => x"00",
          7948 => x"e6",
          7949 => x"00",
          7950 => x"e6",
          7951 => x"00",
          7952 => x"e6",
          7953 => x"00",
          7954 => x"e6",
          7955 => x"00",
          7956 => x"e6",
          7957 => x"00",
          7958 => x"e6",
          7959 => x"00",
          7960 => x"e7",
          7961 => x"00",
          7962 => x"e7",
          7963 => x"00",
          7964 => x"e7",
          7965 => x"00",
          7966 => x"e7",
          7967 => x"00",
          7968 => x"00",
          7969 => x"7f",
          7970 => x"7f",
          7971 => x"7f",
          7972 => x"00",
          7973 => x"ff",
          7974 => x"00",
          7975 => x"00",
          7976 => x"e1",
          7977 => x"00",
          7978 => x"01",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"00",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"5f",
          7996 => x"40",
          7997 => x"73",
          7998 => x"6b",
          7999 => x"63",
          8000 => x"33",
          8001 => x"2d",
          8002 => x"f3",
          8003 => x"f0",
          8004 => x"82",
          8005 => x"58",
          8006 => x"40",
          8007 => x"53",
          8008 => x"4b",
          8009 => x"43",
          8010 => x"33",
          8011 => x"2d",
          8012 => x"f3",
          8013 => x"f0",
          8014 => x"82",
          8015 => x"58",
          8016 => x"60",
          8017 => x"53",
          8018 => x"4b",
          8019 => x"43",
          8020 => x"23",
          8021 => x"3d",
          8022 => x"e0",
          8023 => x"f0",
          8024 => x"87",
          8025 => x"1e",
          8026 => x"00",
          8027 => x"13",
          8028 => x"0b",
          8029 => x"03",
          8030 => x"f0",
          8031 => x"f0",
          8032 => x"f0",
          8033 => x"f0",
          8034 => x"82",
          8035 => x"cf",
          8036 => x"d7",
          8037 => x"41",
          8038 => x"6c",
          8039 => x"d9",
          8040 => x"7e",
          8041 => x"d1",
          8042 => x"c2",
          8043 => x"f0",
          8044 => x"82",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"f1",
          8060 => x"f1",
          8061 => x"f1",
          8062 => x"f1",
          8063 => x"f1",
          8064 => x"f1",
          8065 => x"f1",
          8066 => x"f1",
          8067 => x"f1",
          8068 => x"f1",
          8069 => x"f1",
          8070 => x"f1",
          8071 => x"f1",
          8072 => x"f1",
          8073 => x"f1",
          8074 => x"f1",
          8075 => x"f1",
          8076 => x"f1",
          8077 => x"f1",
          8078 => x"f1",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"32",
          9080 => x"00",
          9081 => x"f6",
          9082 => x"fe",
          9083 => x"c6",
          9084 => x"ef",
          9085 => x"66",
          9086 => x"2e",
          9087 => x"26",
          9088 => x"57",
          9089 => x"06",
          9090 => x"0e",
          9091 => x"16",
          9092 => x"be",
          9093 => x"86",
          9094 => x"8e",
          9095 => x"96",
          9096 => x"a5",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"01",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"93",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"2d",
             6 => x"00",
             7 => x"00",
             8 => x"fd",
             9 => x"05",
            10 => x"ff",
            11 => x"00",
            12 => x"fd",
            13 => x"06",
            14 => x"2b",
            15 => x"0b",
            16 => x"09",
            17 => x"06",
            18 => x"0a",
            19 => x"00",
            20 => x"72",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"73",
            25 => x"81",
            26 => x"10",
            27 => x"51",
            28 => x"72",
            29 => x"04",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"0a",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"72",
            45 => x"0b",
            46 => x"00",
            47 => x"00",
            48 => x"72",
            49 => x"74",
            50 => x"07",
            51 => x"00",
            52 => x"71",
            53 => x"09",
            54 => x"2b",
            55 => x"04",
            56 => x"09",
            57 => x"05",
            58 => x"04",
            59 => x"00",
            60 => x"09",
            61 => x"05",
            62 => x"51",
            63 => x"00",
            64 => x"09",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"72",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"09",
            73 => x"53",
            74 => x"00",
            75 => x"00",
            76 => x"fc",
            77 => x"05",
            78 => x"ff",
            79 => x"00",
            80 => x"fc",
            81 => x"73",
            82 => x"0b",
            83 => x"00",
            84 => x"08",
            85 => x"0b",
            86 => x"08",
            87 => x"51",
            88 => x"08",
            89 => x"0b",
            90 => x"08",
            91 => x"51",
            92 => x"09",
            93 => x"06",
            94 => x"09",
            95 => x"51",
            96 => x"09",
            97 => x"81",
            98 => x"73",
            99 => x"07",
           100 => x"ff",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"81",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"84",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"0d",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"8c",
           134 => x"04",
           135 => x"0b",
           136 => x"8c",
           137 => x"04",
           138 => x"0b",
           139 => x"8d",
           140 => x"04",
           141 => x"0b",
           142 => x"8d",
           143 => x"04",
           144 => x"0b",
           145 => x"8e",
           146 => x"04",
           147 => x"0b",
           148 => x"8e",
           149 => x"04",
           150 => x"0b",
           151 => x"8f",
           152 => x"04",
           153 => x"0b",
           154 => x"8f",
           155 => x"04",
           156 => x"0b",
           157 => x"90",
           158 => x"04",
           159 => x"0b",
           160 => x"90",
           161 => x"04",
           162 => x"0b",
           163 => x"91",
           164 => x"04",
           165 => x"0b",
           166 => x"91",
           167 => x"04",
           168 => x"0b",
           169 => x"92",
           170 => x"04",
           171 => x"0b",
           172 => x"92",
           173 => x"04",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"00",
           193 => x"80",
           194 => x"80",
           195 => x"0c",
           196 => x"80",
           197 => x"0c",
           198 => x"80",
           199 => x"0c",
           200 => x"80",
           201 => x"0c",
           202 => x"80",
           203 => x"0c",
           204 => x"80",
           205 => x"0c",
           206 => x"80",
           207 => x"0c",
           208 => x"80",
           209 => x"0c",
           210 => x"80",
           211 => x"0c",
           212 => x"80",
           213 => x"0c",
           214 => x"80",
           215 => x"0c",
           216 => x"80",
           217 => x"0c",
           218 => x"08",
           219 => x"d4",
           220 => x"d4",
           221 => x"b9",
           222 => x"b9",
           223 => x"84",
           224 => x"84",
           225 => x"04",
           226 => x"2d",
           227 => x"90",
           228 => x"80",
           229 => x"80",
           230 => x"d2",
           231 => x"c0",
           232 => x"82",
           233 => x"80",
           234 => x"0c",
           235 => x"08",
           236 => x"d4",
           237 => x"d4",
           238 => x"b9",
           239 => x"b9",
           240 => x"84",
           241 => x"84",
           242 => x"04",
           243 => x"2d",
           244 => x"90",
           245 => x"e0",
           246 => x"80",
           247 => x"84",
           248 => x"c0",
           249 => x"82",
           250 => x"80",
           251 => x"0c",
           252 => x"08",
           253 => x"d4",
           254 => x"d4",
           255 => x"b9",
           256 => x"b9",
           257 => x"84",
           258 => x"84",
           259 => x"04",
           260 => x"2d",
           261 => x"90",
           262 => x"e7",
           263 => x"80",
           264 => x"e7",
           265 => x"c0",
           266 => x"82",
           267 => x"80",
           268 => x"0c",
           269 => x"08",
           270 => x"d4",
           271 => x"d4",
           272 => x"b9",
           273 => x"b9",
           274 => x"84",
           275 => x"84",
           276 => x"04",
           277 => x"2d",
           278 => x"90",
           279 => x"93",
           280 => x"80",
           281 => x"b7",
           282 => x"c0",
           283 => x"81",
           284 => x"80",
           285 => x"0c",
           286 => x"08",
           287 => x"d4",
           288 => x"d4",
           289 => x"b9",
           290 => x"b9",
           291 => x"84",
           292 => x"84",
           293 => x"04",
           294 => x"2d",
           295 => x"90",
           296 => x"2d",
           297 => x"90",
           298 => x"81",
           299 => x"80",
           300 => x"dc",
           301 => x"c0",
           302 => x"81",
           303 => x"80",
           304 => x"0c",
           305 => x"08",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"51",
           311 => x"73",
           312 => x"10",
           313 => x"0c",
           314 => x"81",
           315 => x"71",
           316 => x"72",
           317 => x"84",
           318 => x"8e",
           319 => x"0c",
           320 => x"81",
           321 => x"3d",
           322 => x"52",
           323 => x"ac",
           324 => x"0d",
           325 => x"85",
           326 => x"73",
           327 => x"52",
           328 => x"d3",
           329 => x"70",
           330 => x"55",
           331 => x"38",
           332 => x"8e",
           333 => x"84",
           334 => x"84",
           335 => x"57",
           336 => x"30",
           337 => x"54",
           338 => x"75",
           339 => x"0c",
           340 => x"b9",
           341 => x"3d",
           342 => x"99",
           343 => x"8e",
           344 => x"3d",
           345 => x"54",
           346 => x"fd",
           347 => x"76",
           348 => x"0d",
           349 => x"42",
           350 => x"85",
           351 => x"81",
           352 => x"7b",
           353 => x"7b",
           354 => x"38",
           355 => x"72",
           356 => x"5f",
           357 => x"b0",
           358 => x"54",
           359 => x"a9",
           360 => x"81",
           361 => x"38",
           362 => x"57",
           363 => x"54",
           364 => x"0d",
           365 => x"10",
           366 => x"70",
           367 => x"29",
           368 => x"5a",
           369 => x"86",
           370 => x"bd",
           371 => x"fe",
           372 => x"2e",
           373 => x"74",
           374 => x"5a",
           375 => x"7c",
           376 => x"33",
           377 => x"39",
           378 => x"55",
           379 => x"40",
           380 => x"72",
           381 => x"10",
           382 => x"04",
           383 => x"73",
           384 => x"8a",
           385 => x"76",
           386 => x"ff",
           387 => x"60",
           388 => x"cf",
           389 => x"d8",
           390 => x"3f",
           391 => x"84",
           392 => x"53",
           393 => x"c8",
           394 => x"81",
           395 => x"90",
           396 => x"84",
           397 => x"b9",
           398 => x"40",
           399 => x"84",
           400 => x"70",
           401 => x"70",
           402 => x"9e",
           403 => x"80",
           404 => x"38",
           405 => x"80",
           406 => x"83",
           407 => x"80",
           408 => x"81",
           409 => x"86",
           410 => x"70",
           411 => x"5b",
           412 => x"85",
           413 => x"70",
           414 => x"59",
           415 => x"7a",
           416 => x"eb",
           417 => x"73",
           418 => x"06",
           419 => x"06",
           420 => x"2a",
           421 => x"38",
           422 => x"80",
           423 => x"54",
           424 => x"b0",
           425 => x"80",
           426 => x"90",
           427 => x"e5",
           428 => x"2e",
           429 => x"29",
           430 => x"5b",
           431 => x"7c",
           432 => x"79",
           433 => x"05",
           434 => x"80",
           435 => x"81",
           436 => x"b9",
           437 => x"38",
           438 => x"76",
           439 => x"84",
           440 => x"ff",
           441 => x"3f",
           442 => x"06",
           443 => x"80",
           444 => x"80",
           445 => x"90",
           446 => x"fc",
           447 => x"f4",
           448 => x"7a",
           449 => x"fa",
           450 => x"c0",
           451 => x"61",
           452 => x"cf",
           453 => x"fd",
           454 => x"80",
           455 => x"2b",
           456 => x"fc",
           457 => x"52",
           458 => x"2a",
           459 => x"c9",
           460 => x"fc",
           461 => x"54",
           462 => x"7c",
           463 => x"39",
           464 => x"5b",
           465 => x"ca",
           466 => x"57",
           467 => x"ff",
           468 => x"54",
           469 => x"38",
           470 => x"33",
           471 => x"fc",
           472 => x"84",
           473 => x"70",
           474 => x"7b",
           475 => x"57",
           476 => x"7f",
           477 => x"40",
           478 => x"38",
           479 => x"b9",
           480 => x"07",
           481 => x"38",
           482 => x"80",
           483 => x"38",
           484 => x"71",
           485 => x"5f",
           486 => x"f6",
           487 => x"ff",
           488 => x"5a",
           489 => x"7a",
           490 => x"76",
           491 => x"60",
           492 => x"5d",
           493 => x"75",
           494 => x"08",
           495 => x"90",
           496 => x"80",
           497 => x"88",
           498 => x"80",
           499 => x"90",
           500 => x"fa",
           501 => x"c4",
           502 => x"83",
           503 => x"06",
           504 => x"83",
           505 => x"5f",
           506 => x"d8",
           507 => x"90",
           508 => x"06",
           509 => x"38",
           510 => x"82",
           511 => x"80",
           512 => x"7c",
           513 => x"3f",
           514 => x"f7",
           515 => x"31",
           516 => x"f9",
           517 => x"c4",
           518 => x"82",
           519 => x"75",
           520 => x"08",
           521 => x"90",
           522 => x"82",
           523 => x"06",
           524 => x"3d",
           525 => x"52",
           526 => x"0d",
           527 => x"0b",
           528 => x"70",
           529 => x"51",
           530 => x"77",
           531 => x"74",
           532 => x"77",
           533 => x"52",
           534 => x"2d",
           535 => x"38",
           536 => x"33",
           537 => x"d5",
           538 => x"ac",
           539 => x"8a",
           540 => x"84",
           541 => x"ff",
           542 => x"0c",
           543 => x"78",
           544 => x"33",
           545 => x"06",
           546 => x"77",
           547 => x"70",
           548 => x"2e",
           549 => x"75",
           550 => x"04",
           551 => x"72",
           552 => x"51",
           553 => x"b9",
           554 => x"74",
           555 => x"72",
           556 => x"84",
           557 => x"3f",
           558 => x"78",
           559 => x"81",
           560 => x"ff",
           561 => x"81",
           562 => x"8c",
           563 => x"25",
           564 => x"34",
           565 => x"15",
           566 => x"76",
           567 => x"3d",
           568 => x"06",
           569 => x"ff",
           570 => x"8c",
           571 => x"76",
           572 => x"85",
           573 => x"81",
           574 => x"ff",
           575 => x"81",
           576 => x"2a",
           577 => x"c3",
           578 => x"71",
           579 => x"76",
           580 => x"17",
           581 => x"84",
           582 => x"74",
           583 => x"34",
           584 => x"0c",
           585 => x"87",
           586 => x"08",
           587 => x"52",
           588 => x"b9",
           589 => x"54",
           590 => x"85",
           591 => x"17",
           592 => x"0c",
           593 => x"53",
           594 => x"39",
           595 => x"54",
           596 => x"51",
           597 => x"70",
           598 => x"70",
           599 => x"73",
           600 => x"04",
           601 => x"55",
           602 => x"38",
           603 => x"2e",
           604 => x"33",
           605 => x"11",
           606 => x"c8",
           607 => x"55",
           608 => x"75",
           609 => x"53",
           610 => x"70",
           611 => x"13",
           612 => x"11",
           613 => x"3d",
           614 => x"81",
           615 => x"ff",
           616 => x"0c",
           617 => x"0d",
           618 => x"70",
           619 => x"70",
           620 => x"73",
           621 => x"04",
           622 => x"55",
           623 => x"38",
           624 => x"70",
           625 => x"70",
           626 => x"85",
           627 => x"78",
           628 => x"a1",
           629 => x"57",
           630 => x"81",
           631 => x"80",
           632 => x"e1",
           633 => x"0c",
           634 => x"f1",
           635 => x"80",
           636 => x"81",
           637 => x"72",
           638 => x"0d",
           639 => x"3d",
           640 => x"53",
           641 => x"b9",
           642 => x"05",
           643 => x"b9",
           644 => x"80",
           645 => x"15",
           646 => x"52",
           647 => x"3f",
           648 => x"b9",
           649 => x"3d",
           650 => x"53",
           651 => x"70",
           652 => x"2e",
           653 => x"2e",
           654 => x"70",
           655 => x"c8",
           656 => x"0d",
           657 => x"54",
           658 => x"70",
           659 => x"70",
           660 => x"85",
           661 => x"7a",
           662 => x"8b",
           663 => x"b9",
           664 => x"80",
           665 => x"3f",
           666 => x"80",
           667 => x"73",
           668 => x"81",
           669 => x"76",
           670 => x"56",
           671 => x"74",
           672 => x"78",
           673 => x"81",
           674 => x"ff",
           675 => x"55",
           676 => x"07",
           677 => x"3d",
           678 => x"fc",
           679 => x"07",
           680 => x"31",
           681 => x"06",
           682 => x"88",
           683 => x"f0",
           684 => x"2b",
           685 => x"53",
           686 => x"30",
           687 => x"77",
           688 => x"70",
           689 => x"06",
           690 => x"51",
           691 => x"53",
           692 => x"56",
           693 => x"0d",
           694 => x"54",
           695 => x"84",
           696 => x"31",
           697 => x"0d",
           698 => x"54",
           699 => x"76",
           700 => x"08",
           701 => x"8d",
           702 => x"84",
           703 => x"71",
           704 => x"71",
           705 => x"71",
           706 => x"57",
           707 => x"2e",
           708 => x"07",
           709 => x"ff",
           710 => x"72",
           711 => x"56",
           712 => x"da",
           713 => x"3d",
           714 => x"2c",
           715 => x"32",
           716 => x"32",
           717 => x"56",
           718 => x"3f",
           719 => x"31",
           720 => x"04",
           721 => x"80",
           722 => x"56",
           723 => x"06",
           724 => x"70",
           725 => x"38",
           726 => x"b0",
           727 => x"80",
           728 => x"8a",
           729 => x"c4",
           730 => x"e0",
           731 => x"d0",
           732 => x"90",
           733 => x"81",
           734 => x"81",
           735 => x"38",
           736 => x"79",
           737 => x"a0",
           738 => x"84",
           739 => x"81",
           740 => x"3d",
           741 => x"0c",
           742 => x"2e",
           743 => x"15",
           744 => x"73",
           745 => x"73",
           746 => x"a0",
           747 => x"80",
           748 => x"e1",
           749 => x"3d",
           750 => x"78",
           751 => x"fe",
           752 => x"0c",
           753 => x"7b",
           754 => x"77",
           755 => x"a0",
           756 => x"15",
           757 => x"73",
           758 => x"80",
           759 => x"38",
           760 => x"26",
           761 => x"a0",
           762 => x"74",
           763 => x"ff",
           764 => x"ff",
           765 => x"38",
           766 => x"54",
           767 => x"78",
           768 => x"13",
           769 => x"56",
           770 => x"38",
           771 => x"56",
           772 => x"b9",
           773 => x"70",
           774 => x"56",
           775 => x"fe",
           776 => x"70",
           777 => x"a6",
           778 => x"a0",
           779 => x"38",
           780 => x"89",
           781 => x"b9",
           782 => x"58",
           783 => x"55",
           784 => x"0b",
           785 => x"04",
           786 => x"08",
           787 => x"04",
           788 => x"26",
           789 => x"84",
           790 => x"9c",
           791 => x"04",
           792 => x"83",
           793 => x"ef",
           794 => x"ce",
           795 => x"0d",
           796 => x"3f",
           797 => x"51",
           798 => x"83",
           799 => x"3d",
           800 => x"f1",
           801 => x"dc",
           802 => x"04",
           803 => x"83",
           804 => x"ee",
           805 => x"d0",
           806 => x"0d",
           807 => x"3f",
           808 => x"51",
           809 => x"83",
           810 => x"3d",
           811 => x"99",
           812 => x"88",
           813 => x"04",
           814 => x"83",
           815 => x"ed",
           816 => x"d1",
           817 => x"0d",
           818 => x"3f",
           819 => x"66",
           820 => x"5b",
           821 => x"07",
           822 => x"57",
           823 => x"57",
           824 => x"51",
           825 => x"81",
           826 => x"58",
           827 => x"08",
           828 => x"80",
           829 => x"3f",
           830 => x"7b",
           831 => x"57",
           832 => x"87",
           833 => x"e7",
           834 => x"87",
           835 => x"b9",
           836 => x"78",
           837 => x"3f",
           838 => x"0d",
           839 => x"98",
           840 => x"96",
           841 => x"75",
           842 => x"84",
           843 => x"08",
           844 => x"2e",
           845 => x"57",
           846 => x"51",
           847 => x"52",
           848 => x"c8",
           849 => x"52",
           850 => x"ff",
           851 => x"84",
           852 => x"58",
           853 => x"ec",
           854 => x"76",
           855 => x"8a",
           856 => x"3d",
           857 => x"56",
           858 => x"53",
           859 => x"b9",
           860 => x"3d",
           861 => x"63",
           862 => x"73",
           863 => x"5f",
           864 => x"38",
           865 => x"fe",
           866 => x"3f",
           867 => x"7c",
           868 => x"2e",
           869 => x"7a",
           870 => x"83",
           871 => x"14",
           872 => x"51",
           873 => x"38",
           874 => x"80",
           875 => x"75",
           876 => x"72",
           877 => x"53",
           878 => x"74",
           879 => x"57",
           880 => x"74",
           881 => x"08",
           882 => x"16",
           883 => x"d2",
           884 => x"79",
           885 => x"3f",
           886 => x"98",
           887 => x"ee",
           888 => x"7b",
           889 => x"38",
           890 => x"3d",
           891 => x"ae",
           892 => x"53",
           893 => x"74",
           894 => x"83",
           895 => x"14",
           896 => x"51",
           897 => x"c0",
           898 => x"df",
           899 => x"51",
           900 => x"ac",
           901 => x"3f",
           902 => x"39",
           903 => x"84",
           904 => x"a0",
           905 => x"fd",
           906 => x"27",
           907 => x"fc",
           908 => x"d5",
           909 => x"84",
           910 => x"d8",
           911 => x"51",
           912 => x"91",
           913 => x"c8",
           914 => x"72",
           915 => x"72",
           916 => x"e0",
           917 => x"51",
           918 => x"98",
           919 => x"70",
           920 => x"72",
           921 => x"58",
           922 => x"fd",
           923 => x"84",
           924 => x"2c",
           925 => x"32",
           926 => x"07",
           927 => x"53",
           928 => x"b9",
           929 => x"8f",
           930 => x"c0",
           931 => x"81",
           932 => x"51",
           933 => x"3f",
           934 => x"52",
           935 => x"70",
           936 => x"38",
           937 => x"52",
           938 => x"70",
           939 => x"38",
           940 => x"52",
           941 => x"70",
           942 => x"38",
           943 => x"52",
           944 => x"06",
           945 => x"84",
           946 => x"3f",
           947 => x"80",
           948 => x"84",
           949 => x"3f",
           950 => x"80",
           951 => x"81",
           952 => x"cb",
           953 => x"d4",
           954 => x"9b",
           955 => x"06",
           956 => x"38",
           957 => x"83",
           958 => x"51",
           959 => x"81",
           960 => x"f0",
           961 => x"9b",
           962 => x"3f",
           963 => x"2a",
           964 => x"2e",
           965 => x"51",
           966 => x"9b",
           967 => x"72",
           968 => x"71",
           969 => x"39",
           970 => x"d0",
           971 => x"cb",
           972 => x"51",
           973 => x"ff",
           974 => x"83",
           975 => x"51",
           976 => x"81",
           977 => x"b8",
           978 => x"80",
           979 => x"d4",
           980 => x"b6",
           981 => x"ff",
           982 => x"2e",
           983 => x"e3",
           984 => x"ec",
           985 => x"f8",
           986 => x"3f",
           987 => x"81",
           988 => x"82",
           989 => x"38",
           990 => x"2e",
           991 => x"79",
           992 => x"5c",
           993 => x"38",
           994 => x"a0",
           995 => x"26",
           996 => x"c0",
           997 => x"3f",
           998 => x"08",
           999 => x"e8",
          1000 => x"38",
          1001 => x"83",
          1002 => x"06",
          1003 => x"9a",
          1004 => x"dd",
          1005 => x"92",
          1006 => x"b9",
          1007 => x"84",
          1008 => x"80",
          1009 => x"c8",
          1010 => x"80",
          1011 => x"08",
          1012 => x"08",
          1013 => x"a5",
          1014 => x"85",
          1015 => x"7a",
          1016 => x"80",
          1017 => x"d5",
          1018 => x"b9",
          1019 => x"54",
          1020 => x"52",
          1021 => x"c8",
          1022 => x"30",
          1023 => x"5b",
          1024 => x"38",
          1025 => x"80",
          1026 => x"ff",
          1027 => x"7f",
          1028 => x"7c",
          1029 => x"e8",
          1030 => x"83",
          1031 => x"48",
          1032 => x"e8",
          1033 => x"33",
          1034 => x"fd",
          1035 => x"52",
          1036 => x"3f",
          1037 => x"81",
          1038 => x"84",
          1039 => x"51",
          1040 => x"08",
          1041 => x"08",
          1042 => x"ee",
          1043 => x"59",
          1044 => x"d3",
          1045 => x"82",
          1046 => x"83",
          1047 => x"80",
          1048 => x"67",
          1049 => x"90",
          1050 => x"33",
          1051 => x"38",
          1052 => x"5a",
          1053 => x"f8",
          1054 => x"53",
          1055 => x"85",
          1056 => x"2e",
          1057 => x"70",
          1058 => x"39",
          1059 => x"7d",
          1060 => x"39",
          1061 => x"d6",
          1062 => x"52",
          1063 => x"39",
          1064 => x"9a",
          1065 => x"83",
          1066 => x"81",
          1067 => x"d6",
          1068 => x"78",
          1069 => x"3f",
          1070 => x"3d",
          1071 => x"51",
          1072 => x"80",
          1073 => x"d6",
          1074 => x"79",
          1075 => x"fa",
          1076 => x"83",
          1077 => x"95",
          1078 => x"ff",
          1079 => x"b9",
          1080 => x"68",
          1081 => x"3f",
          1082 => x"f4",
          1083 => x"a8",
          1084 => x"f9",
          1085 => x"53",
          1086 => x"84",
          1087 => x"59",
          1088 => x"a8",
          1089 => x"08",
          1090 => x"91",
          1091 => x"ae",
          1092 => x"87",
          1093 => x"59",
          1094 => x"53",
          1095 => x"84",
          1096 => x"38",
          1097 => x"80",
          1098 => x"c8",
          1099 => x"22",
          1100 => x"cf",
          1101 => x"80",
          1102 => x"7e",
          1103 => x"f8",
          1104 => x"38",
          1105 => x"39",
          1106 => x"80",
          1107 => x"c8",
          1108 => x"3d",
          1109 => x"51",
          1110 => x"80",
          1111 => x"f8",
          1112 => x"c4",
          1113 => x"f7",
          1114 => x"b6",
          1115 => x"27",
          1116 => x"33",
          1117 => x"38",
          1118 => x"78",
          1119 => x"3f",
          1120 => x"1b",
          1121 => x"84",
          1122 => x"f4",
          1123 => x"f7",
          1124 => x"53",
          1125 => x"84",
          1126 => x"38",
          1127 => x"80",
          1128 => x"c8",
          1129 => x"d7",
          1130 => x"79",
          1131 => x"79",
          1132 => x"65",
          1133 => x"ff",
          1134 => x"e8",
          1135 => x"2e",
          1136 => x"11",
          1137 => x"3f",
          1138 => x"70",
          1139 => x"cc",
          1140 => x"80",
          1141 => x"7e",
          1142 => x"f6",
          1143 => x"38",
          1144 => x"59",
          1145 => x"68",
          1146 => x"11",
          1147 => x"3f",
          1148 => x"dd",
          1149 => x"33",
          1150 => x"3d",
          1151 => x"51",
          1152 => x"ff",
          1153 => x"ff",
          1154 => x"e6",
          1155 => x"2e",
          1156 => x"11",
          1157 => x"3f",
          1158 => x"8d",
          1159 => x"ff",
          1160 => x"b9",
          1161 => x"08",
          1162 => x"3f",
          1163 => x"8f",
          1164 => x"05",
          1165 => x"8a",
          1166 => x"b8",
          1167 => x"3f",
          1168 => x"80",
          1169 => x"53",
          1170 => x"ea",
          1171 => x"2e",
          1172 => x"51",
          1173 => x"3d",
          1174 => x"51",
          1175 => x"91",
          1176 => x"80",
          1177 => x"08",
          1178 => x"ff",
          1179 => x"b9",
          1180 => x"33",
          1181 => x"83",
          1182 => x"f8",
          1183 => x"8c",
          1184 => x"a5",
          1185 => x"2e",
          1186 => x"70",
          1187 => x"06",
          1188 => x"38",
          1189 => x"83",
          1190 => x"55",
          1191 => x"51",
          1192 => x"d6",
          1193 => x"71",
          1194 => x"3d",
          1195 => x"51",
          1196 => x"80",
          1197 => x"0c",
          1198 => x"fe",
          1199 => x"e2",
          1200 => x"38",
          1201 => x"ce",
          1202 => x"23",
          1203 => x"53",
          1204 => x"84",
          1205 => x"38",
          1206 => x"7e",
          1207 => x"b8",
          1208 => x"05",
          1209 => x"08",
          1210 => x"3d",
          1211 => x"51",
          1212 => x"80",
          1213 => x"80",
          1214 => x"05",
          1215 => x"f0",
          1216 => x"80",
          1217 => x"81",
          1218 => x"64",
          1219 => x"39",
          1220 => x"9d",
          1221 => x"80",
          1222 => x"c8",
          1223 => x"7c",
          1224 => x"83",
          1225 => x"f5",
          1226 => x"ff",
          1227 => x"b9",
          1228 => x"59",
          1229 => x"82",
          1230 => x"39",
          1231 => x"2e",
          1232 => x"47",
          1233 => x"5c",
          1234 => x"8c",
          1235 => x"e8",
          1236 => x"b6",
          1237 => x"3f",
          1238 => x"ce",
          1239 => x"83",
          1240 => x"83",
          1241 => x"c6",
          1242 => x"80",
          1243 => x"47",
          1244 => x"5e",
          1245 => x"9c",
          1246 => x"cf",
          1247 => x"83",
          1248 => x"83",
          1249 => x"9b",
          1250 => x"b9",
          1251 => x"80",
          1252 => x"47",
          1253 => x"fc",
          1254 => x"f2",
          1255 => x"39",
          1256 => x"f8",
          1257 => x"56",
          1258 => x"da",
          1259 => x"2b",
          1260 => x"52",
          1261 => x"b9",
          1262 => x"94",
          1263 => x"80",
          1264 => x"b9",
          1265 => x"55",
          1266 => x"93",
          1267 => x"77",
          1268 => x"94",
          1269 => x"c0",
          1270 => x"81",
          1271 => x"a1",
          1272 => x"0b",
          1273 => x"72",
          1274 => x"85",
          1275 => x"ba",
          1276 => x"b0",
          1277 => x"3f",
          1278 => x"94",
          1279 => x"d2",
          1280 => x"d2",
          1281 => x"3f",
          1282 => x"80",
          1283 => x"3f",
          1284 => x"51",
          1285 => x"04",
          1286 => x"56",
          1287 => x"81",
          1288 => x"06",
          1289 => x"06",
          1290 => x"81",
          1291 => x"2e",
          1292 => x"73",
          1293 => x"72",
          1294 => x"33",
          1295 => x"70",
          1296 => x"80",
          1297 => x"38",
          1298 => x"81",
          1299 => x"09",
          1300 => x"a2",
          1301 => x"07",
          1302 => x"38",
          1303 => x"71",
          1304 => x"c8",
          1305 => x"2e",
          1306 => x"38",
          1307 => x"81",
          1308 => x"2e",
          1309 => x"15",
          1310 => x"2e",
          1311 => x"39",
          1312 => x"8b",
          1313 => x"86",
          1314 => x"52",
          1315 => x"c8",
          1316 => x"b9",
          1317 => x"3d",
          1318 => x"52",
          1319 => x"98",
          1320 => x"82",
          1321 => x"84",
          1322 => x"26",
          1323 => x"84",
          1324 => x"86",
          1325 => x"26",
          1326 => x"86",
          1327 => x"38",
          1328 => x"87",
          1329 => x"87",
          1330 => x"c0",
          1331 => x"c0",
          1332 => x"c0",
          1333 => x"c0",
          1334 => x"c0",
          1335 => x"c0",
          1336 => x"a4",
          1337 => x"80",
          1338 => x"52",
          1339 => x"0d",
          1340 => x"c0",
          1341 => x"c0",
          1342 => x"87",
          1343 => x"1c",
          1344 => x"79",
          1345 => x"08",
          1346 => x"98",
          1347 => x"87",
          1348 => x"1c",
          1349 => x"7b",
          1350 => x"08",
          1351 => x"0c",
          1352 => x"83",
          1353 => x"57",
          1354 => x"55",
          1355 => x"53",
          1356 => x"d8",
          1357 => x"3d",
          1358 => x"05",
          1359 => x"72",
          1360 => x"c8",
          1361 => x"52",
          1362 => x"38",
          1363 => x"b9",
          1364 => x"51",
          1365 => x"08",
          1366 => x"71",
          1367 => x"72",
          1368 => x"c8",
          1369 => x"52",
          1370 => x"fd",
          1371 => x"88",
          1372 => x"3f",
          1373 => x"98",
          1374 => x"38",
          1375 => x"83",
          1376 => x"c8",
          1377 => x"0d",
          1378 => x"33",
          1379 => x"70",
          1380 => x"94",
          1381 => x"06",
          1382 => x"38",
          1383 => x"51",
          1384 => x"06",
          1385 => x"93",
          1386 => x"73",
          1387 => x"80",
          1388 => x"c0",
          1389 => x"84",
          1390 => x"71",
          1391 => x"70",
          1392 => x"53",
          1393 => x"2a",
          1394 => x"38",
          1395 => x"2a",
          1396 => x"cf",
          1397 => x"8f",
          1398 => x"51",
          1399 => x"83",
          1400 => x"55",
          1401 => x"70",
          1402 => x"83",
          1403 => x"54",
          1404 => x"38",
          1405 => x"2a",
          1406 => x"80",
          1407 => x"81",
          1408 => x"81",
          1409 => x"8a",
          1410 => x"71",
          1411 => x"87",
          1412 => x"86",
          1413 => x"72",
          1414 => x"73",
          1415 => x"0c",
          1416 => x"70",
          1417 => x"72",
          1418 => x"2e",
          1419 => x"52",
          1420 => x"c0",
          1421 => x"81",
          1422 => x"d7",
          1423 => x"80",
          1424 => x"52",
          1425 => x"c0",
          1426 => x"87",
          1427 => x"0c",
          1428 => x"8c",
          1429 => x"f2",
          1430 => x"83",
          1431 => x"08",
          1432 => x"ac",
          1433 => x"9e",
          1434 => x"c0",
          1435 => x"87",
          1436 => x"0c",
          1437 => x"ac",
          1438 => x"f2",
          1439 => x"83",
          1440 => x"08",
          1441 => x"c0",
          1442 => x"87",
          1443 => x"0c",
          1444 => x"c4",
          1445 => x"80",
          1446 => x"84",
          1447 => x"82",
          1448 => x"80",
          1449 => x"88",
          1450 => x"80",
          1451 => x"f2",
          1452 => x"90",
          1453 => x"52",
          1454 => x"52",
          1455 => x"87",
          1456 => x"80",
          1457 => x"83",
          1458 => x"34",
          1459 => x"70",
          1460 => x"70",
          1461 => x"83",
          1462 => x"9e",
          1463 => x"51",
          1464 => x"81",
          1465 => x"0b",
          1466 => x"80",
          1467 => x"2e",
          1468 => x"cf",
          1469 => x"08",
          1470 => x"52",
          1471 => x"71",
          1472 => x"c0",
          1473 => x"06",
          1474 => x"38",
          1475 => x"80",
          1476 => x"80",
          1477 => x"80",
          1478 => x"f2",
          1479 => x"90",
          1480 => x"52",
          1481 => x"71",
          1482 => x"90",
          1483 => x"53",
          1484 => x"0b",
          1485 => x"80",
          1486 => x"83",
          1487 => x"34",
          1488 => x"06",
          1489 => x"f2",
          1490 => x"90",
          1491 => x"70",
          1492 => x"83",
          1493 => x"08",
          1494 => x"34",
          1495 => x"82",
          1496 => x"51",
          1497 => x"33",
          1498 => x"98",
          1499 => x"33",
          1500 => x"cf",
          1501 => x"f2",
          1502 => x"83",
          1503 => x"38",
          1504 => x"cb",
          1505 => x"84",
          1506 => x"73",
          1507 => x"55",
          1508 => x"33",
          1509 => x"cb",
          1510 => x"f2",
          1511 => x"83",
          1512 => x"38",
          1513 => x"e1",
          1514 => x"3f",
          1515 => x"bc",
          1516 => x"b0",
          1517 => x"b5",
          1518 => x"83",
          1519 => x"83",
          1520 => x"f2",
          1521 => x"ff",
          1522 => x"56",
          1523 => x"8b",
          1524 => x"c0",
          1525 => x"b9",
          1526 => x"ff",
          1527 => x"55",
          1528 => x"55",
          1529 => x"83",
          1530 => x"52",
          1531 => x"c8",
          1532 => x"31",
          1533 => x"83",
          1534 => x"87",
          1535 => x"56",
          1536 => x"a3",
          1537 => x"c0",
          1538 => x"b9",
          1539 => x"ff",
          1540 => x"55",
          1541 => x"9f",
          1542 => x"3f",
          1543 => x"83",
          1544 => x"51",
          1545 => x"08",
          1546 => x"b6",
          1547 => x"da",
          1548 => x"da",
          1549 => x"b8",
          1550 => x"b3",
          1551 => x"bd",
          1552 => x"3f",
          1553 => x"29",
          1554 => x"c8",
          1555 => x"b2",
          1556 => x"74",
          1557 => x"39",
          1558 => x"3f",
          1559 => x"2e",
          1560 => x"db",
          1561 => x"f2",
          1562 => x"f0",
          1563 => x"ff",
          1564 => x"55",
          1565 => x"39",
          1566 => x"3f",
          1567 => x"2e",
          1568 => x"d6",
          1569 => x"b1",
          1570 => x"75",
          1571 => x"83",
          1572 => x"51",
          1573 => x"33",
          1574 => x"cd",
          1575 => x"dc",
          1576 => x"f2",
          1577 => x"cb",
          1578 => x"83",
          1579 => x"dd",
          1580 => x"f2",
          1581 => x"a2",
          1582 => x"83",
          1583 => x"dd",
          1584 => x"f2",
          1585 => x"f9",
          1586 => x"83",
          1587 => x"dd",
          1588 => x"f2",
          1589 => x"d0",
          1590 => x"83",
          1591 => x"dd",
          1592 => x"f2",
          1593 => x"a7",
          1594 => x"83",
          1595 => x"dd",
          1596 => x"f2",
          1597 => x"fe",
          1598 => x"ff",
          1599 => x"ff",
          1600 => x"55",
          1601 => x"39",
          1602 => x"52",
          1603 => x"10",
          1604 => x"04",
          1605 => x"3f",
          1606 => x"51",
          1607 => x"04",
          1608 => x"3f",
          1609 => x"51",
          1610 => x"04",
          1611 => x"3f",
          1612 => x"51",
          1613 => x"04",
          1614 => x"87",
          1615 => x"dc",
          1616 => x"d9",
          1617 => x"08",
          1618 => x"52",
          1619 => x"83",
          1620 => x"38",
          1621 => x"b4",
          1622 => x"51",
          1623 => x"08",
          1624 => x"e6",
          1625 => x"57",
          1626 => x"25",
          1627 => x"05",
          1628 => x"74",
          1629 => x"2a",
          1630 => x"38",
          1631 => x"08",
          1632 => x"9b",
          1633 => x"78",
          1634 => x"c8",
          1635 => x"fc",
          1636 => x"2e",
          1637 => x"79",
          1638 => x"bf",
          1639 => x"b9",
          1640 => x"e2",
          1641 => x"0b",
          1642 => x"04",
          1643 => x"3d",
          1644 => x"57",
          1645 => x"38",
          1646 => x"10",
          1647 => x"08",
          1648 => x"b9",
          1649 => x"51",
          1650 => x"90",
          1651 => x"2e",
          1652 => x"38",
          1653 => x"54",
          1654 => x"73",
          1655 => x"04",
          1656 => x"11",
          1657 => x"3f",
          1658 => x"38",
          1659 => x"fd",
          1660 => x"ff",
          1661 => x"81",
          1662 => x"82",
          1663 => x"39",
          1664 => x"27",
          1665 => x"70",
          1666 => x"81",
          1667 => x"eb",
          1668 => x"fe",
          1669 => x"53",
          1670 => x"84",
          1671 => x"d0",
          1672 => x"f8",
          1673 => x"84",
          1674 => x"77",
          1675 => x"c8",
          1676 => x"08",
          1677 => x"ff",
          1678 => x"34",
          1679 => x"e1",
          1680 => x"74",
          1681 => x"38",
          1682 => x"3d",
          1683 => x"08",
          1684 => x"41",
          1685 => x"f3",
          1686 => x"5d",
          1687 => x"33",
          1688 => x"38",
          1689 => x"70",
          1690 => x"38",
          1691 => x"3d",
          1692 => x"8a",
          1693 => x"70",
          1694 => x"ec",
          1695 => x"84",
          1696 => x"84",
          1697 => x"97",
          1698 => x"10",
          1699 => x"70",
          1700 => x"5b",
          1701 => x"2e",
          1702 => x"87",
          1703 => x"ff",
          1704 => x"80",
          1705 => x"16",
          1706 => x"83",
          1707 => x"61",
          1708 => x"08",
          1709 => x"2e",
          1710 => x"38",
          1711 => x"76",
          1712 => x"70",
          1713 => x"80",
          1714 => x"71",
          1715 => x"de",
          1716 => x"58",
          1717 => x"90",
          1718 => x"ac",
          1719 => x"75",
          1720 => x"05",
          1721 => x"59",
          1722 => x"38",
          1723 => x"55",
          1724 => x"42",
          1725 => x"de",
          1726 => x"55",
          1727 => x"80",
          1728 => x"81",
          1729 => x"fe",
          1730 => x"80",
          1731 => x"d1",
          1732 => x"79",
          1733 => x"74",
          1734 => x"10",
          1735 => x"04",
          1736 => x"80",
          1737 => x"84",
          1738 => x"8c",
          1739 => x"38",
          1740 => x"ff",
          1741 => x"ff",
          1742 => x"fc",
          1743 => x"81",
          1744 => x"57",
          1745 => x"84",
          1746 => x"77",
          1747 => x"33",
          1748 => x"bc",
          1749 => x"7c",
          1750 => x"08",
          1751 => x"84",
          1752 => x"d1",
          1753 => x"56",
          1754 => x"ac",
          1755 => x"3f",
          1756 => x"ff",
          1757 => x"52",
          1758 => x"d1",
          1759 => x"d1",
          1760 => x"74",
          1761 => x"3f",
          1762 => x"39",
          1763 => x"56",
          1764 => x"83",
          1765 => x"55",
          1766 => x"75",
          1767 => x"ff",
          1768 => x"84",
          1769 => x"81",
          1770 => x"7b",
          1771 => x"88",
          1772 => x"74",
          1773 => x"ac",
          1774 => x"3f",
          1775 => x"ff",
          1776 => x"52",
          1777 => x"d1",
          1778 => x"d1",
          1779 => x"c7",
          1780 => x"ff",
          1781 => x"55",
          1782 => x"d5",
          1783 => x"84",
          1784 => x"52",
          1785 => x"8c",
          1786 => x"88",
          1787 => x"fa",
          1788 => x"81",
          1789 => x"7b",
          1790 => x"fc",
          1791 => x"ff",
          1792 => x"55",
          1793 => x"d4",
          1794 => x"88",
          1795 => x"c4",
          1796 => x"88",
          1797 => x"7c",
          1798 => x"76",
          1799 => x"08",
          1800 => x"84",
          1801 => x"98",
          1802 => x"57",
          1803 => x"84",
          1804 => x"b2",
          1805 => x"81",
          1806 => x"d1",
          1807 => x"24",
          1808 => x"52",
          1809 => x"81",
          1810 => x"70",
          1811 => x"56",
          1812 => x"f8",
          1813 => x"33",
          1814 => x"77",
          1815 => x"81",
          1816 => x"70",
          1817 => x"57",
          1818 => x"7b",
          1819 => x"84",
          1820 => x"ff",
          1821 => x"29",
          1822 => x"84",
          1823 => x"76",
          1824 => x"84",
          1825 => x"f7",
          1826 => x"88",
          1827 => x"8c",
          1828 => x"8c",
          1829 => x"39",
          1830 => x"80",
          1831 => x"8a",
          1832 => x"88",
          1833 => x"b9",
          1834 => x"89",
          1835 => x"76",
          1836 => x"b8",
          1837 => x"05",
          1838 => x"a0",
          1839 => x"83",
          1840 => x"57",
          1841 => x"c8",
          1842 => x"70",
          1843 => x"08",
          1844 => x"83",
          1845 => x"8c",
          1846 => x"80",
          1847 => x"d1",
          1848 => x"34",
          1849 => x"0d",
          1850 => x"80",
          1851 => x"52",
          1852 => x"d5",
          1853 => x"84",
          1854 => x"51",
          1855 => x"33",
          1856 => x"34",
          1857 => x"38",
          1858 => x"3f",
          1859 => x"0b",
          1860 => x"83",
          1861 => x"84",
          1862 => x"b6",
          1863 => x"51",
          1864 => x"08",
          1865 => x"84",
          1866 => x"ae",
          1867 => x"05",
          1868 => x"81",
          1869 => x"d1",
          1870 => x"0b",
          1871 => x"d1",
          1872 => x"b4",
          1873 => x"70",
          1874 => x"2e",
          1875 => x"ff",
          1876 => x"ff",
          1877 => x"84",
          1878 => x"ad",
          1879 => x"98",
          1880 => x"33",
          1881 => x"80",
          1882 => x"a0",
          1883 => x"8c",
          1884 => x"84",
          1885 => x"74",
          1886 => x"ac",
          1887 => x"3f",
          1888 => x"0a",
          1889 => x"33",
          1890 => x"cc",
          1891 => x"51",
          1892 => x"0a",
          1893 => x"2c",
          1894 => x"78",
          1895 => x"39",
          1896 => x"34",
          1897 => x"51",
          1898 => x"0a",
          1899 => x"2c",
          1900 => x"75",
          1901 => x"57",
          1902 => x"ac",
          1903 => x"f4",
          1904 => x"80",
          1905 => x"88",
          1906 => x"ff",
          1907 => x"8c",
          1908 => x"76",
          1909 => x"88",
          1910 => x"74",
          1911 => x"76",
          1912 => x"7a",
          1913 => x"0a",
          1914 => x"2c",
          1915 => x"75",
          1916 => x"74",
          1917 => x"06",
          1918 => x"34",
          1919 => x"25",
          1920 => x"d1",
          1921 => x"33",
          1922 => x"0a",
          1923 => x"06",
          1924 => x"81",
          1925 => x"2c",
          1926 => x"75",
          1927 => x"ac",
          1928 => x"3f",
          1929 => x"0a",
          1930 => x"33",
          1931 => x"84",
          1932 => x"51",
          1933 => x"0a",
          1934 => x"2c",
          1935 => x"74",
          1936 => x"39",
          1937 => x"2e",
          1938 => x"96",
          1939 => x"88",
          1940 => x"06",
          1941 => x"ff",
          1942 => x"84",
          1943 => x"2e",
          1944 => x"52",
          1945 => x"d5",
          1946 => x"9c",
          1947 => x"51",
          1948 => x"33",
          1949 => x"34",
          1950 => x"a8",
          1951 => x"c8",
          1952 => x"c8",
          1953 => x"b0",
          1954 => x"39",
          1955 => x"70",
          1956 => x"75",
          1957 => x"05",
          1958 => x"52",
          1959 => x"84",
          1960 => x"98",
          1961 => x"5a",
          1962 => x"fd",
          1963 => x"2e",
          1964 => x"93",
          1965 => x"ff",
          1966 => x"25",
          1967 => x"34",
          1968 => x"2e",
          1969 => x"f6",
          1970 => x"d9",
          1971 => x"0c",
          1972 => x"bc",
          1973 => x"80",
          1974 => x"56",
          1975 => x"ba",
          1976 => x"84",
          1977 => x"84",
          1978 => x"05",
          1979 => x"90",
          1980 => x"84",
          1981 => x"80",
          1982 => x"08",
          1983 => x"84",
          1984 => x"a6",
          1985 => x"88",
          1986 => x"8c",
          1987 => x"8c",
          1988 => x"39",
          1989 => x"8c",
          1990 => x"7b",
          1991 => x"04",
          1992 => x"b9",
          1993 => x"b9",
          1994 => x"53",
          1995 => x"3f",
          1996 => x"d1",
          1997 => x"52",
          1998 => x"38",
          1999 => x"ff",
          2000 => x"52",
          2001 => x"d5",
          2002 => x"dc",
          2003 => x"57",
          2004 => x"ff",
          2005 => x"a8",
          2006 => x"d1",
          2007 => x"ff",
          2008 => x"51",
          2009 => x"81",
          2010 => x"d1",
          2011 => x"80",
          2012 => x"08",
          2013 => x"84",
          2014 => x"a4",
          2015 => x"88",
          2016 => x"8c",
          2017 => x"8c",
          2018 => x"39",
          2019 => x"f3",
          2020 => x"06",
          2021 => x"54",
          2022 => x"84",
          2023 => x"b8",
          2024 => x"05",
          2025 => x"2e",
          2026 => x"74",
          2027 => x"b8",
          2028 => x"5a",
          2029 => x"77",
          2030 => x"b4",
          2031 => x"7b",
          2032 => x"83",
          2033 => x"ba",
          2034 => x"81",
          2035 => x"8c",
          2036 => x"7b",
          2037 => x"04",
          2038 => x"08",
          2039 => x"c8",
          2040 => x"08",
          2041 => x"08",
          2042 => x"b7",
          2043 => x"84",
          2044 => x"06",
          2045 => x"51",
          2046 => x"08",
          2047 => x"25",
          2048 => x"ff",
          2049 => x"34",
          2050 => x"33",
          2051 => x"70",
          2052 => x"f2",
          2053 => x"83",
          2054 => x"58",
          2055 => x"c8",
          2056 => x"70",
          2057 => x"08",
          2058 => x"1d",
          2059 => x"7d",
          2060 => x"2e",
          2061 => x"e8",
          2062 => x"79",
          2063 => x"83",
          2064 => x"ff",
          2065 => x"c8",
          2066 => x"ff",
          2067 => x"3f",
          2068 => x"87",
          2069 => x"1b",
          2070 => x"cf",
          2071 => x"83",
          2072 => x"f2",
          2073 => x"74",
          2074 => x"39",
          2075 => x"39",
          2076 => x"39",
          2077 => x"3f",
          2078 => x"f2",
          2079 => x"02",
          2080 => x"53",
          2081 => x"81",
          2082 => x"83",
          2083 => x"38",
          2084 => x"b0",
          2085 => x"a0",
          2086 => x"83",
          2087 => x"34",
          2088 => x"f4",
          2089 => x"07",
          2090 => x"7f",
          2091 => x"94",
          2092 => x"0c",
          2093 => x"76",
          2094 => x"a2",
          2095 => x"9a",
          2096 => x"a0",
          2097 => x"70",
          2098 => x"72",
          2099 => x"a7",
          2100 => x"70",
          2101 => x"71",
          2102 => x"58",
          2103 => x"84",
          2104 => x"84",
          2105 => x"83",
          2106 => x"06",
          2107 => x"5e",
          2108 => x"38",
          2109 => x"81",
          2110 => x"81",
          2111 => x"62",
          2112 => x"5d",
          2113 => x"26",
          2114 => x"76",
          2115 => x"5f",
          2116 => x"fe",
          2117 => x"77",
          2118 => x"81",
          2119 => x"74",
          2120 => x"86",
          2121 => x"80",
          2122 => x"ff",
          2123 => x"ff",
          2124 => x"29",
          2125 => x"57",
          2126 => x"81",
          2127 => x"71",
          2128 => x"2e",
          2129 => x"f8",
          2130 => x"83",
          2131 => x"90",
          2132 => x"07",
          2133 => x"79",
          2134 => x"72",
          2135 => x"70",
          2136 => x"83",
          2137 => x"86",
          2138 => x"56",
          2139 => x"14",
          2140 => x"06",
          2141 => x"06",
          2142 => x"ff",
          2143 => x"5a",
          2144 => x"79",
          2145 => x"15",
          2146 => x"81",
          2147 => x"71",
          2148 => x"81",
          2149 => x"5b",
          2150 => x"38",
          2151 => x"16",
          2152 => x"e2",
          2153 => x"da",
          2154 => x"7b",
          2155 => x"0d",
          2156 => x"73",
          2157 => x"81",
          2158 => x"80",
          2159 => x"86",
          2160 => x"80",
          2161 => x"8a",
          2162 => x"75",
          2163 => x"3f",
          2164 => x"54",
          2165 => x"73",
          2166 => x"75",
          2167 => x"80",
          2168 => x"86",
          2169 => x"81",
          2170 => x"f3",
          2171 => x"07",
          2172 => x"84",
          2173 => x"c8",
          2174 => x"bc",
          2175 => x"3d",
          2176 => x"05",
          2177 => x"5b",
          2178 => x"82",
          2179 => x"f8",
          2180 => x"71",
          2181 => x"83",
          2182 => x"71",
          2183 => x"06",
          2184 => x"53",
          2185 => x"f8",
          2186 => x"f8",
          2187 => x"05",
          2188 => x"06",
          2189 => x"8c",
          2190 => x"f8",
          2191 => x"ff",
          2192 => x"55",
          2193 => x"84",
          2194 => x"58",
          2195 => x"38",
          2196 => x"e0",
          2197 => x"72",
          2198 => x"81",
          2199 => x"b7",
          2200 => x"9f",
          2201 => x"84",
          2202 => x"e0",
          2203 => x"05",
          2204 => x"74",
          2205 => x"ff",
          2206 => x"75",
          2207 => x"ff",
          2208 => x"81",
          2209 => x"84",
          2210 => x"55",
          2211 => x"58",
          2212 => x"06",
          2213 => x"19",
          2214 => x"b9",
          2215 => x"e0",
          2216 => x"33",
          2217 => x"70",
          2218 => x"05",
          2219 => x"33",
          2220 => x"19",
          2221 => x"ce",
          2222 => x"0c",
          2223 => x"f8",
          2224 => x"ff",
          2225 => x"55",
          2226 => x"77",
          2227 => x"ff",
          2228 => x"56",
          2229 => x"fe",
          2230 => x"84",
          2231 => x"72",
          2232 => x"73",
          2233 => x"33",
          2234 => x"55",
          2235 => x"34",
          2236 => x"ff",
          2237 => x"38",
          2238 => x"75",
          2239 => x"53",
          2240 => x"0b",
          2241 => x"89",
          2242 => x"84",
          2243 => x"b7",
          2244 => x"3d",
          2245 => x"33",
          2246 => x"70",
          2247 => x"70",
          2248 => x"71",
          2249 => x"f9",
          2250 => x"86",
          2251 => x"f9",
          2252 => x"ff",
          2253 => x"38",
          2254 => x"34",
          2255 => x"3d",
          2256 => x"73",
          2257 => x"06",
          2258 => x"f8",
          2259 => x"72",
          2260 => x"55",
          2261 => x"70",
          2262 => x"0b",
          2263 => x"04",
          2264 => x"70",
          2265 => x"56",
          2266 => x"80",
          2267 => x"0d",
          2268 => x"84",
          2269 => x"51",
          2270 => x"72",
          2271 => x"b9",
          2272 => x"0b",
          2273 => x"33",
          2274 => x"52",
          2275 => x"12",
          2276 => x"d0",
          2277 => x"33",
          2278 => x"10",
          2279 => x"08",
          2280 => x"f0",
          2281 => x"70",
          2282 => x"51",
          2283 => x"9c",
          2284 => x"34",
          2285 => x"3d",
          2286 => x"9f",
          2287 => x"f4",
          2288 => x"83",
          2289 => x"80",
          2290 => x"34",
          2291 => x"fe",
          2292 => x"f4",
          2293 => x"f8",
          2294 => x"0c",
          2295 => x"33",
          2296 => x"83",
          2297 => x"f8",
          2298 => x"f8",
          2299 => x"f4",
          2300 => x"70",
          2301 => x"83",
          2302 => x"07",
          2303 => x"81",
          2304 => x"06",
          2305 => x"34",
          2306 => x"81",
          2307 => x"34",
          2308 => x"81",
          2309 => x"83",
          2310 => x"f8",
          2311 => x"51",
          2312 => x"39",
          2313 => x"80",
          2314 => x"34",
          2315 => x"81",
          2316 => x"83",
          2317 => x"f8",
          2318 => x"51",
          2319 => x"39",
          2320 => x"51",
          2321 => x"39",
          2322 => x"82",
          2323 => x"fd",
          2324 => x"05",
          2325 => x"33",
          2326 => x"33",
          2327 => x"33",
          2328 => x"82",
          2329 => x"a5",
          2330 => x"7d",
          2331 => x"b7",
          2332 => x"7b",
          2333 => x"f9",
          2334 => x"2e",
          2335 => x"84",
          2336 => x"c0",
          2337 => x"a8",
          2338 => x"83",
          2339 => x"bc",
          2340 => x"84",
          2341 => x"53",
          2342 => x"81",
          2343 => x"80",
          2344 => x"f8",
          2345 => x"7c",
          2346 => x"04",
          2347 => x"0b",
          2348 => x"f8",
          2349 => x"34",
          2350 => x"b8",
          2351 => x"57",
          2352 => x"7b",
          2353 => x"d8",
          2354 => x"84",
          2355 => x"27",
          2356 => x"05",
          2357 => x"51",
          2358 => x"81",
          2359 => x"5b",
          2360 => x"d2",
          2361 => x"84",
          2362 => x"c0",
          2363 => x"83",
          2364 => x"34",
          2365 => x"b7",
          2366 => x"34",
          2367 => x"0b",
          2368 => x"f8",
          2369 => x"92",
          2370 => x"83",
          2371 => x"80",
          2372 => x"86",
          2373 => x"fd",
          2374 => x"52",
          2375 => x"3f",
          2376 => x"5a",
          2377 => x"84",
          2378 => x"33",
          2379 => x"33",
          2380 => x"80",
          2381 => x"59",
          2382 => x"ff",
          2383 => x"59",
          2384 => x"81",
          2385 => x"38",
          2386 => x"81",
          2387 => x"82",
          2388 => x"f8",
          2389 => x"72",
          2390 => x"c4",
          2391 => x"34",
          2392 => x"33",
          2393 => x"12",
          2394 => x"fa",
          2395 => x"71",
          2396 => x"33",
          2397 => x"b7",
          2398 => x"f8",
          2399 => x"72",
          2400 => x"83",
          2401 => x"34",
          2402 => x"55",
          2403 => x"b7",
          2404 => x"ff",
          2405 => x"84",
          2406 => x"8c",
          2407 => x"80",
          2408 => x"b9",
          2409 => x"8d",
          2410 => x"f7",
          2411 => x"fe",
          2412 => x"96",
          2413 => x"ff",
          2414 => x"53",
          2415 => x"75",
          2416 => x"38",
          2417 => x"ba",
          2418 => x"54",
          2419 => x"76",
          2420 => x"13",
          2421 => x"73",
          2422 => x"83",
          2423 => x"52",
          2424 => x"84",
          2425 => x"75",
          2426 => x"ca",
          2427 => x"ff",
          2428 => x"38",
          2429 => x"76",
          2430 => x"f8",
          2431 => x"ff",
          2432 => x"53",
          2433 => x"39",
          2434 => x"52",
          2435 => x"39",
          2436 => x"fe",
          2437 => x"f3",
          2438 => x"59",
          2439 => x"82",
          2440 => x"84",
          2441 => x"38",
          2442 => x"89",
          2443 => x"33",
          2444 => x"33",
          2445 => x"84",
          2446 => x"80",
          2447 => x"f8",
          2448 => x"71",
          2449 => x"83",
          2450 => x"33",
          2451 => x"83",
          2452 => x"80",
          2453 => x"81",
          2454 => x"f8",
          2455 => x"40",
          2456 => x"84",
          2457 => x"81",
          2458 => x"81",
          2459 => x"79",
          2460 => x"83",
          2461 => x"c8",
          2462 => x"2e",
          2463 => x"fd",
          2464 => x"78",
          2465 => x"0b",
          2466 => x"33",
          2467 => x"33",
          2468 => x"84",
          2469 => x"80",
          2470 => x"f8",
          2471 => x"71",
          2472 => x"83",
          2473 => x"33",
          2474 => x"f8",
          2475 => x"34",
          2476 => x"06",
          2477 => x"33",
          2478 => x"58",
          2479 => x"98",
          2480 => x"81",
          2481 => x"ca",
          2482 => x"0b",
          2483 => x"04",
          2484 => x"9b",
          2485 => x"09",
          2486 => x"83",
          2487 => x"c8",
          2488 => x"2e",
          2489 => x"89",
          2490 => x"33",
          2491 => x"c8",
          2492 => x"77",
          2493 => x"b8",
          2494 => x"c8",
          2495 => x"2e",
          2496 => x"c4",
          2497 => x"f8",
          2498 => x"29",
          2499 => x"19",
          2500 => x"84",
          2501 => x"83",
          2502 => x"41",
          2503 => x"1f",
          2504 => x"29",
          2505 => x"86",
          2506 => x"bc",
          2507 => x"f6",
          2508 => x"29",
          2509 => x"f8",
          2510 => x"34",
          2511 => x"52",
          2512 => x"83",
          2513 => x"b7",
          2514 => x"81",
          2515 => x"71",
          2516 => x"83",
          2517 => x"7e",
          2518 => x"83",
          2519 => x"5c",
          2520 => x"81",
          2521 => x"fc",
          2522 => x"f9",
          2523 => x"b8",
          2524 => x"34",
          2525 => x"0b",
          2526 => x"b8",
          2527 => x"0c",
          2528 => x"33",
          2529 => x"33",
          2530 => x"33",
          2531 => x"b8",
          2532 => x"0c",
          2533 => x"2e",
          2534 => x"f8",
          2535 => x"81",
          2536 => x"81",
          2537 => x"a7",
          2538 => x"5c",
          2539 => x"ff",
          2540 => x"5c",
          2541 => x"2e",
          2542 => x"ff",
          2543 => x"57",
          2544 => x"ff",
          2545 => x"ff",
          2546 => x"5b",
          2547 => x"80",
          2548 => x"f8",
          2549 => x"71",
          2550 => x"0b",
          2551 => x"f8",
          2552 => x"56",
          2553 => x"80",
          2554 => x"81",
          2555 => x"f8",
          2556 => x"5d",
          2557 => x"7f",
          2558 => x"70",
          2559 => x"26",
          2560 => x"5a",
          2561 => x"77",
          2562 => x"33",
          2563 => x"56",
          2564 => x"d8",
          2565 => x"78",
          2566 => x"c8",
          2567 => x"bf",
          2568 => x"38",
          2569 => x"58",
          2570 => x"f9",
          2571 => x"3f",
          2572 => x"3d",
          2573 => x"b7",
          2574 => x"f8",
          2575 => x"75",
          2576 => x"83",
          2577 => x"29",
          2578 => x"f7",
          2579 => x"5b",
          2580 => x"80",
          2581 => x"ff",
          2582 => x"29",
          2583 => x"33",
          2584 => x"b7",
          2585 => x"f8",
          2586 => x"41",
          2587 => x"1c",
          2588 => x"29",
          2589 => x"86",
          2590 => x"bc",
          2591 => x"f6",
          2592 => x"29",
          2593 => x"f8",
          2594 => x"60",
          2595 => x"58",
          2596 => x"b7",
          2597 => x"ff",
          2598 => x"81",
          2599 => x"7b",
          2600 => x"f8",
          2601 => x"f9",
          2602 => x"ff",
          2603 => x"29",
          2604 => x"84",
          2605 => x"1b",
          2606 => x"f9",
          2607 => x"29",
          2608 => x"83",
          2609 => x"33",
          2610 => x"f8",
          2611 => x"34",
          2612 => x"06",
          2613 => x"33",
          2614 => x"40",
          2615 => x"9a",
          2616 => x"ff",
          2617 => x"d6",
          2618 => x"df",
          2619 => x"80",
          2620 => x"0d",
          2621 => x"84",
          2622 => x"f8",
          2623 => x"ff",
          2624 => x"84",
          2625 => x"c8",
          2626 => x"fa",
          2627 => x"33",
          2628 => x"b7",
          2629 => x"5b",
          2630 => x"b8",
          2631 => x"d8",
          2632 => x"b9",
          2633 => x"84",
          2634 => x"75",
          2635 => x"fe",
          2636 => x"61",
          2637 => x"39",
          2638 => x"b7",
          2639 => x"f8",
          2640 => x"f9",
          2641 => x"84",
          2642 => x"83",
          2643 => x"41",
          2644 => x"7f",
          2645 => x"b7",
          2646 => x"f8",
          2647 => x"43",
          2648 => x"34",
          2649 => x"1b",
          2650 => x"86",
          2651 => x"bc",
          2652 => x"f6",
          2653 => x"29",
          2654 => x"f8",
          2655 => x"81",
          2656 => x"60",
          2657 => x"bd",
          2658 => x"1a",
          2659 => x"0b",
          2660 => x"33",
          2661 => x"84",
          2662 => x"38",
          2663 => x"80",
          2664 => x"0d",
          2665 => x"f8",
          2666 => x"f9",
          2667 => x"83",
          2668 => x"f8",
          2669 => x"f8",
          2670 => x"f8",
          2671 => x"9e",
          2672 => x"80",
          2673 => x"22",
          2674 => x"ff",
          2675 => x"05",
          2676 => x"54",
          2677 => x"3d",
          2678 => x"76",
          2679 => x"c8",
          2680 => x"33",
          2681 => x"fe",
          2682 => x"51",
          2683 => x"80",
          2684 => x"79",
          2685 => x"fe",
          2686 => x"05",
          2687 => x"26",
          2688 => x"c7",
          2689 => x"b8",
          2690 => x"a4",
          2691 => x"9d",
          2692 => x"9f",
          2693 => x"5c",
          2694 => x"39",
          2695 => x"2e",
          2696 => x"ff",
          2697 => x"bc",
          2698 => x"fd",
          2699 => x"fd",
          2700 => x"34",
          2701 => x"06",
          2702 => x"38",
          2703 => x"34",
          2704 => x"f9",
          2705 => x"bb",
          2706 => x"25",
          2707 => x"83",
          2708 => x"b8",
          2709 => x"e0",
          2710 => x"9d",
          2711 => x"9f",
          2712 => x"5a",
          2713 => x"39",
          2714 => x"2e",
          2715 => x"41",
          2716 => x"b6",
          2717 => x"f9",
          2718 => x"29",
          2719 => x"f8",
          2720 => x"60",
          2721 => x"83",
          2722 => x"06",
          2723 => x"80",
          2724 => x"f7",
          2725 => x"c9",
          2726 => x"38",
          2727 => x"2e",
          2728 => x"0b",
          2729 => x"84",
          2730 => x"90",
          2731 => x"f8",
          2732 => x"bc",
          2733 => x"7d",
          2734 => x"f8",
          2735 => x"c9",
          2736 => x"38",
          2737 => x"33",
          2738 => x"ff",
          2739 => x"83",
          2740 => x"34",
          2741 => x"fe",
          2742 => x"c9",
          2743 => x"c7",
          2744 => x"70",
          2745 => x"fe",
          2746 => x"ff",
          2747 => x"58",
          2748 => x"33",
          2749 => x"84",
          2750 => x"83",
          2751 => x"ff",
          2752 => x"39",
          2753 => x"27",
          2754 => x"ff",
          2755 => x"9d",
          2756 => x"84",
          2757 => x"ff",
          2758 => x"5c",
          2759 => x"79",
          2760 => x"06",
          2761 => x"83",
          2762 => x"34",
          2763 => x"40",
          2764 => x"56",
          2765 => x"39",
          2766 => x"2e",
          2767 => x"84",
          2768 => x"26",
          2769 => x"84",
          2770 => x"83",
          2771 => x"86",
          2772 => x"22",
          2773 => x"83",
          2774 => x"46",
          2775 => x"2e",
          2776 => x"06",
          2777 => x"24",
          2778 => x"56",
          2779 => x"16",
          2780 => x"81",
          2781 => x"80",
          2782 => x"bb",
          2783 => x"38",
          2784 => x"34",
          2785 => x"22",
          2786 => x"90",
          2787 => x"81",
          2788 => x"5b",
          2789 => x"86",
          2790 => x"7f",
          2791 => x"42",
          2792 => x"d6",
          2793 => x"e0",
          2794 => x"33",
          2795 => x"70",
          2796 => x"05",
          2797 => x"33",
          2798 => x"1d",
          2799 => x"f7",
          2800 => x"84",
          2801 => x"05",
          2802 => x"33",
          2803 => x"18",
          2804 => x"33",
          2805 => x"58",
          2806 => x"e6",
          2807 => x"80",
          2808 => x"b9",
          2809 => x"ce",
          2810 => x"ff",
          2811 => x"40",
          2812 => x"b9",
          2813 => x"81",
          2814 => x"33",
          2815 => x"f8",
          2816 => x"2e",
          2817 => x"40",
          2818 => x"81",
          2819 => x"fe",
          2820 => x"07",
          2821 => x"10",
          2822 => x"a7",
          2823 => x"86",
          2824 => x"58",
          2825 => x"83",
          2826 => x"f8",
          2827 => x"2b",
          2828 => x"79",
          2829 => x"27",
          2830 => x"59",
          2831 => x"0c",
          2832 => x"bc",
          2833 => x"7e",
          2834 => x"83",
          2835 => x"05",
          2836 => x"8c",
          2837 => x"29",
          2838 => x"57",
          2839 => x"83",
          2840 => x"59",
          2841 => x"79",
          2842 => x"17",
          2843 => x"a0",
          2844 => x"70",
          2845 => x"75",
          2846 => x"ff",
          2847 => x"fe",
          2848 => x"80",
          2849 => x"06",
          2850 => x"7b",
          2851 => x"38",
          2852 => x"81",
          2853 => x"f5",
          2854 => x"5e",
          2855 => x"83",
          2856 => x"83",
          2857 => x"42",
          2858 => x"f8",
          2859 => x"f8",
          2860 => x"06",
          2861 => x"f4",
          2862 => x"75",
          2863 => x"f8",
          2864 => x"56",
          2865 => x"83",
          2866 => x"07",
          2867 => x"39",
          2868 => x"90",
          2869 => x"ff",
          2870 => x"f4",
          2871 => x"59",
          2872 => x"33",
          2873 => x"f4",
          2874 => x"33",
          2875 => x"83",
          2876 => x"f8",
          2877 => x"07",
          2878 => x"ea",
          2879 => x"06",
          2880 => x"f4",
          2881 => x"33",
          2882 => x"83",
          2883 => x"f8",
          2884 => x"56",
          2885 => x"39",
          2886 => x"84",
          2887 => x"fe",
          2888 => x"fa",
          2889 => x"f4",
          2890 => x"33",
          2891 => x"f4",
          2892 => x"33",
          2893 => x"f4",
          2894 => x"33",
          2895 => x"f4",
          2896 => x"33",
          2897 => x"75",
          2898 => x"83",
          2899 => x"07",
          2900 => x"ba",
          2901 => x"80",
          2902 => x"ff",
          2903 => x"f8",
          2904 => x"f9",
          2905 => x"83",
          2906 => x"c4",
          2907 => x"b8",
          2908 => x"0c",
          2909 => x"f9",
          2910 => x"ff",
          2911 => x"39",
          2912 => x"11",
          2913 => x"3f",
          2914 => x"b9",
          2915 => x"0b",
          2916 => x"b9",
          2917 => x"83",
          2918 => x"b8",
          2919 => x"84",
          2920 => x"06",
          2921 => x"b9",
          2922 => x"c8",
          2923 => x"f9",
          2924 => x"3f",
          2925 => x"06",
          2926 => x"80",
          2927 => x"81",
          2928 => x"8a",
          2929 => x"39",
          2930 => x"09",
          2931 => x"57",
          2932 => x"d9",
          2933 => x"60",
          2934 => x"f9",
          2935 => x"33",
          2936 => x"72",
          2937 => x"83",
          2938 => x"bb",
          2939 => x"78",
          2940 => x"bb",
          2941 => x"ff",
          2942 => x"a6",
          2943 => x"bc",
          2944 => x"f9",
          2945 => x"a0",
          2946 => x"5f",
          2947 => x"ff",
          2948 => x"44",
          2949 => x"f5",
          2950 => x"11",
          2951 => x"38",
          2952 => x"27",
          2953 => x"83",
          2954 => x"ff",
          2955 => x"df",
          2956 => x"76",
          2957 => x"75",
          2958 => x"06",
          2959 => x"5a",
          2960 => x"31",
          2961 => x"71",
          2962 => x"a7",
          2963 => x"7c",
          2964 => x"71",
          2965 => x"79",
          2966 => x"9a",
          2967 => x"84",
          2968 => x"05",
          2969 => x"33",
          2970 => x"18",
          2971 => x"33",
          2972 => x"58",
          2973 => x"e0",
          2974 => x"33",
          2975 => x"70",
          2976 => x"05",
          2977 => x"33",
          2978 => x"1d",
          2979 => x"ff",
          2980 => x"fa",
          2981 => x"33",
          2982 => x"b7",
          2983 => x"b7",
          2984 => x"e9",
          2985 => x"bb",
          2986 => x"5c",
          2987 => x"76",
          2988 => x"81",
          2989 => x"7a",
          2990 => x"f8",
          2991 => x"81",
          2992 => x"80",
          2993 => x"75",
          2994 => x"83",
          2995 => x"bc",
          2996 => x"7f",
          2997 => x"c5",
          2998 => x"f4",
          2999 => x"81",
          3000 => x"44",
          3001 => x"81",
          3002 => x"ff",
          3003 => x"fd",
          3004 => x"f8",
          3005 => x"31",
          3006 => x"90",
          3007 => x"26",
          3008 => x"05",
          3009 => x"70",
          3010 => x"f4",
          3011 => x"58",
          3012 => x"81",
          3013 => x"38",
          3014 => x"75",
          3015 => x"80",
          3016 => x"39",
          3017 => x"39",
          3018 => x"8e",
          3019 => x"f1",
          3020 => x"5a",
          3021 => x"80",
          3022 => x"39",
          3023 => x"84",
          3024 => x"2e",
          3025 => x"80",
          3026 => x"0d",
          3027 => x"3f",
          3028 => x"3d",
          3029 => x"05",
          3030 => x"33",
          3031 => x"11",
          3032 => x"2e",
          3033 => x"83",
          3034 => x"b9",
          3035 => x"f7",
          3036 => x"2e",
          3037 => x"71",
          3038 => x"5d",
          3039 => x"ff",
          3040 => x"81",
          3041 => x"32",
          3042 => x"5c",
          3043 => x"38",
          3044 => x"33",
          3045 => x"12",
          3046 => x"f6",
          3047 => x"05",
          3048 => x"cd",
          3049 => x"2e",
          3050 => x"86",
          3051 => x"c0",
          3052 => x"08",
          3053 => x"ee",
          3054 => x"f8",
          3055 => x"06",
          3056 => x"38",
          3057 => x"70",
          3058 => x"33",
          3059 => x"c1",
          3060 => x"38",
          3061 => x"81",
          3062 => x"85",
          3063 => x"34",
          3064 => x"f2",
          3065 => x"06",
          3066 => x"38",
          3067 => x"70",
          3068 => x"f7",
          3069 => x"86",
          3070 => x"54",
          3071 => x"81",
          3072 => x"81",
          3073 => x"38",
          3074 => x"0b",
          3075 => x"08",
          3076 => x"a4",
          3077 => x"42",
          3078 => x"16",
          3079 => x"38",
          3080 => x"80",
          3081 => x"16",
          3082 => x"38",
          3083 => x"81",
          3084 => x"73",
          3085 => x"90",
          3086 => x"da",
          3087 => x"81",
          3088 => x"90",
          3089 => x"80",
          3090 => x"05",
          3091 => x"73",
          3092 => x"87",
          3093 => x"0c",
          3094 => x"57",
          3095 => x"76",
          3096 => x"a4",
          3097 => x"26",
          3098 => x"c8",
          3099 => x"f7",
          3100 => x"38",
          3101 => x"08",
          3102 => x"38",
          3103 => x"54",
          3104 => x"73",
          3105 => x"9c",
          3106 => x"ff",
          3107 => x"83",
          3108 => x"c4",
          3109 => x"fc",
          3110 => x"72",
          3111 => x"2e",
          3112 => x"81",
          3113 => x"fe",
          3114 => x"59",
          3115 => x"2e",
          3116 => x"81",
          3117 => x"80",
          3118 => x"87",
          3119 => x"72",
          3120 => x"9c",
          3121 => x"76",
          3122 => x"71",
          3123 => x"80",
          3124 => x"10",
          3125 => x"78",
          3126 => x"5b",
          3127 => x"08",
          3128 => x"39",
          3129 => x"38",
          3130 => x"39",
          3131 => x"2e",
          3132 => x"be",
          3133 => x"e8",
          3134 => x"80",
          3135 => x"8a",
          3136 => x"f9",
          3137 => x"38",
          3138 => x"f7",
          3139 => x"7c",
          3140 => x"81",
          3141 => x"e2",
          3142 => x"80",
          3143 => x"33",
          3144 => x"ff",
          3145 => x"78",
          3146 => x"04",
          3147 => x"f6",
          3148 => x"83",
          3149 => x"7a",
          3150 => x"39",
          3151 => x"ff",
          3152 => x"0b",
          3153 => x"39",
          3154 => x"ff",
          3155 => x"16",
          3156 => x"38",
          3157 => x"2e",
          3158 => x"f7",
          3159 => x"98",
          3160 => x"fb",
          3161 => x"83",
          3162 => x"59",
          3163 => x"fc",
          3164 => x"f7",
          3165 => x"72",
          3166 => x"34",
          3167 => x"f7",
          3168 => x"83",
          3169 => x"5d",
          3170 => x"9c",
          3171 => x"fc",
          3172 => x"fc",
          3173 => x"06",
          3174 => x"76",
          3175 => x"80",
          3176 => x"75",
          3177 => x"bf",
          3178 => x"0b",
          3179 => x"83",
          3180 => x"34",
          3181 => x"83",
          3182 => x"38",
          3183 => x"ff",
          3184 => x"ff",
          3185 => x"79",
          3186 => x"f8",
          3187 => x"15",
          3188 => x"80",
          3189 => x"b7",
          3190 => x"ff",
          3191 => x"80",
          3192 => x"59",
          3193 => x"ff",
          3194 => x"39",
          3195 => x"08",
          3196 => x"e5",
          3197 => x"83",
          3198 => x"80",
          3199 => x"82",
          3200 => x"0b",
          3201 => x"a3",
          3202 => x"d4",
          3203 => x"0b",
          3204 => x"0b",
          3205 => x"80",
          3206 => x"83",
          3207 => x"05",
          3208 => x"87",
          3209 => x"2e",
          3210 => x"98",
          3211 => x"87",
          3212 => x"87",
          3213 => x"70",
          3214 => x"71",
          3215 => x"98",
          3216 => x"87",
          3217 => x"98",
          3218 => x"38",
          3219 => x"08",
          3220 => x"71",
          3221 => x"98",
          3222 => x"38",
          3223 => x"81",
          3224 => x"98",
          3225 => x"fe",
          3226 => x"76",
          3227 => x"04",
          3228 => x"3d",
          3229 => x"84",
          3230 => x"0b",
          3231 => x"87",
          3232 => x"2a",
          3233 => x"15",
          3234 => x"15",
          3235 => x"15",
          3236 => x"d4",
          3237 => x"f3",
          3238 => x"85",
          3239 => x"fe",
          3240 => x"f0",
          3241 => x"08",
          3242 => x"90",
          3243 => x"52",
          3244 => x"72",
          3245 => x"c0",
          3246 => x"27",
          3247 => x"38",
          3248 => x"55",
          3249 => x"55",
          3250 => x"c0",
          3251 => x"53",
          3252 => x"c0",
          3253 => x"f6",
          3254 => x"9c",
          3255 => x"38",
          3256 => x"c0",
          3257 => x"83",
          3258 => x"70",
          3259 => x"2e",
          3260 => x"52",
          3261 => x"81",
          3262 => x"c6",
          3263 => x"52",
          3264 => x"81",
          3265 => x"53",
          3266 => x"84",
          3267 => x"81",
          3268 => x"0d",
          3269 => x"0d",
          3270 => x"56",
          3271 => x"77",
          3272 => x"70",
          3273 => x"57",
          3274 => x"51",
          3275 => x"52",
          3276 => x"34",
          3277 => x"11",
          3278 => x"70",
          3279 => x"05",
          3280 => x"34",
          3281 => x"d4",
          3282 => x"f3",
          3283 => x"85",
          3284 => x"fe",
          3285 => x"f0",
          3286 => x"08",
          3287 => x"90",
          3288 => x"52",
          3289 => x"72",
          3290 => x"c0",
          3291 => x"27",
          3292 => x"38",
          3293 => x"55",
          3294 => x"55",
          3295 => x"c0",
          3296 => x"53",
          3297 => x"c0",
          3298 => x"f6",
          3299 => x"9c",
          3300 => x"38",
          3301 => x"c0",
          3302 => x"83",
          3303 => x"70",
          3304 => x"2e",
          3305 => x"71",
          3306 => x"ff",
          3307 => x"81",
          3308 => x"3d",
          3309 => x"3d",
          3310 => x"d0",
          3311 => x"08",
          3312 => x"80",
          3313 => x"c0",
          3314 => x"56",
          3315 => x"98",
          3316 => x"08",
          3317 => x"15",
          3318 => x"52",
          3319 => x"fe",
          3320 => x"08",
          3321 => x"c8",
          3322 => x"c0",
          3323 => x"ce",
          3324 => x"08",
          3325 => x"70",
          3326 => x"87",
          3327 => x"73",
          3328 => x"db",
          3329 => x"72",
          3330 => x"53",
          3331 => x"52",
          3332 => x"ff",
          3333 => x"39",
          3334 => x"fe",
          3335 => x"f9",
          3336 => x"71",
          3337 => x"06",
          3338 => x"81",
          3339 => x"2b",
          3340 => x"33",
          3341 => x"5c",
          3342 => x"52",
          3343 => x"af",
          3344 => x"12",
          3345 => x"07",
          3346 => x"71",
          3347 => x"53",
          3348 => x"24",
          3349 => x"14",
          3350 => x"07",
          3351 => x"56",
          3352 => x"ff",
          3353 => x"b9",
          3354 => x"85",
          3355 => x"88",
          3356 => x"84",
          3357 => x"b9",
          3358 => x"13",
          3359 => x"b9",
          3360 => x"73",
          3361 => x"16",
          3362 => x"2b",
          3363 => x"2a",
          3364 => x"75",
          3365 => x"86",
          3366 => x"2b",
          3367 => x"16",
          3368 => x"07",
          3369 => x"53",
          3370 => x"85",
          3371 => x"16",
          3372 => x"8b",
          3373 => x"5a",
          3374 => x"13",
          3375 => x"2a",
          3376 => x"34",
          3377 => x"08",
          3378 => x"88",
          3379 => x"88",
          3380 => x"34",
          3381 => x"08",
          3382 => x"71",
          3383 => x"05",
          3384 => x"2b",
          3385 => x"06",
          3386 => x"53",
          3387 => x"82",
          3388 => x"b9",
          3389 => x"12",
          3390 => x"07",
          3391 => x"71",
          3392 => x"70",
          3393 => x"57",
          3394 => x"14",
          3395 => x"82",
          3396 => x"2b",
          3397 => x"33",
          3398 => x"90",
          3399 => x"57",
          3400 => x"38",
          3401 => x"2b",
          3402 => x"2a",
          3403 => x"81",
          3404 => x"17",
          3405 => x"2b",
          3406 => x"14",
          3407 => x"07",
          3408 => x"58",
          3409 => x"75",
          3410 => x"f9",
          3411 => x"58",
          3412 => x"80",
          3413 => x"3f",
          3414 => x"0b",
          3415 => x"84",
          3416 => x"76",
          3417 => x"b5",
          3418 => x"75",
          3419 => x"b9",
          3420 => x"81",
          3421 => x"08",
          3422 => x"87",
          3423 => x"b9",
          3424 => x"07",
          3425 => x"2a",
          3426 => x"34",
          3427 => x"22",
          3428 => x"08",
          3429 => x"15",
          3430 => x"ee",
          3431 => x"53",
          3432 => x"fb",
          3433 => x"ff",
          3434 => x"ff",
          3435 => x"33",
          3436 => x"70",
          3437 => x"ff",
          3438 => x"75",
          3439 => x"12",
          3440 => x"ff",
          3441 => x"ff",
          3442 => x"5c",
          3443 => x"70",
          3444 => x"58",
          3445 => x"88",
          3446 => x"73",
          3447 => x"74",
          3448 => x"11",
          3449 => x"2b",
          3450 => x"56",
          3451 => x"83",
          3452 => x"26",
          3453 => x"2e",
          3454 => x"88",
          3455 => x"11",
          3456 => x"2a",
          3457 => x"34",
          3458 => x"08",
          3459 => x"82",
          3460 => x"b9",
          3461 => x"12",
          3462 => x"2b",
          3463 => x"83",
          3464 => x"58",
          3465 => x"12",
          3466 => x"83",
          3467 => x"54",
          3468 => x"84",
          3469 => x"33",
          3470 => x"83",
          3471 => x"53",
          3472 => x"15",
          3473 => x"55",
          3474 => x"33",
          3475 => x"54",
          3476 => x"71",
          3477 => x"70",
          3478 => x"71",
          3479 => x"05",
          3480 => x"15",
          3481 => x"b8",
          3482 => x"11",
          3483 => x"07",
          3484 => x"70",
          3485 => x"84",
          3486 => x"70",
          3487 => x"04",
          3488 => x"8b",
          3489 => x"84",
          3490 => x"2b",
          3491 => x"53",
          3492 => x"85",
          3493 => x"19",
          3494 => x"8b",
          3495 => x"86",
          3496 => x"2b",
          3497 => x"52",
          3498 => x"34",
          3499 => x"08",
          3500 => x"88",
          3501 => x"88",
          3502 => x"34",
          3503 => x"08",
          3504 => x"f9",
          3505 => x"58",
          3506 => x"54",
          3507 => x"0c",
          3508 => x"91",
          3509 => x"c8",
          3510 => x"f4",
          3511 => x"0b",
          3512 => x"53",
          3513 => x"cd",
          3514 => x"76",
          3515 => x"84",
          3516 => x"34",
          3517 => x"b8",
          3518 => x"0b",
          3519 => x"84",
          3520 => x"80",
          3521 => x"88",
          3522 => x"17",
          3523 => x"b4",
          3524 => x"b8",
          3525 => x"82",
          3526 => x"77",
          3527 => x"fe",
          3528 => x"41",
          3529 => x"59",
          3530 => x"38",
          3531 => x"80",
          3532 => x"60",
          3533 => x"2a",
          3534 => x"55",
          3535 => x"78",
          3536 => x"06",
          3537 => x"81",
          3538 => x"75",
          3539 => x"10",
          3540 => x"61",
          3541 => x"88",
          3542 => x"2c",
          3543 => x"43",
          3544 => x"42",
          3545 => x"15",
          3546 => x"07",
          3547 => x"81",
          3548 => x"2b",
          3549 => x"80",
          3550 => x"27",
          3551 => x"62",
          3552 => x"85",
          3553 => x"25",
          3554 => x"79",
          3555 => x"33",
          3556 => x"83",
          3557 => x"12",
          3558 => x"07",
          3559 => x"58",
          3560 => x"1e",
          3561 => x"8b",
          3562 => x"86",
          3563 => x"2b",
          3564 => x"14",
          3565 => x"07",
          3566 => x"5b",
          3567 => x"84",
          3568 => x"b9",
          3569 => x"85",
          3570 => x"2b",
          3571 => x"15",
          3572 => x"2a",
          3573 => x"57",
          3574 => x"34",
          3575 => x"81",
          3576 => x"ff",
          3577 => x"5e",
          3578 => x"34",
          3579 => x"11",
          3580 => x"71",
          3581 => x"81",
          3582 => x"88",
          3583 => x"55",
          3584 => x"34",
          3585 => x"33",
          3586 => x"83",
          3587 => x"83",
          3588 => x"88",
          3589 => x"55",
          3590 => x"1a",
          3591 => x"82",
          3592 => x"2b",
          3593 => x"2b",
          3594 => x"05",
          3595 => x"b8",
          3596 => x"1c",
          3597 => x"5f",
          3598 => x"54",
          3599 => x"0d",
          3600 => x"b8",
          3601 => x"23",
          3602 => x"ff",
          3603 => x"b9",
          3604 => x"0b",
          3605 => x"5d",
          3606 => x"1e",
          3607 => x"86",
          3608 => x"84",
          3609 => x"ff",
          3610 => x"ff",
          3611 => x"5b",
          3612 => x"18",
          3613 => x"10",
          3614 => x"05",
          3615 => x"0b",
          3616 => x"57",
          3617 => x"82",
          3618 => x"fe",
          3619 => x"84",
          3620 => x"95",
          3621 => x"b8",
          3622 => x"44",
          3623 => x"71",
          3624 => x"70",
          3625 => x"63",
          3626 => x"84",
          3627 => x"57",
          3628 => x"19",
          3629 => x"70",
          3630 => x"07",
          3631 => x"74",
          3632 => x"88",
          3633 => x"5d",
          3634 => x"ff",
          3635 => x"84",
          3636 => x"34",
          3637 => x"b8",
          3638 => x"3f",
          3639 => x"31",
          3640 => x"fa",
          3641 => x"76",
          3642 => x"17",
          3643 => x"07",
          3644 => x"81",
          3645 => x"2b",
          3646 => x"45",
          3647 => x"ff",
          3648 => x"38",
          3649 => x"83",
          3650 => x"fc",
          3651 => x"f4",
          3652 => x"0b",
          3653 => x"53",
          3654 => x"c4",
          3655 => x"7e",
          3656 => x"84",
          3657 => x"34",
          3658 => x"b8",
          3659 => x"0b",
          3660 => x"84",
          3661 => x"80",
          3662 => x"88",
          3663 => x"88",
          3664 => x"84",
          3665 => x"84",
          3666 => x"43",
          3667 => x"83",
          3668 => x"24",
          3669 => x"06",
          3670 => x"fc",
          3671 => x"38",
          3672 => x"73",
          3673 => x"04",
          3674 => x"33",
          3675 => x"7a",
          3676 => x"71",
          3677 => x"05",
          3678 => x"88",
          3679 => x"45",
          3680 => x"56",
          3681 => x"85",
          3682 => x"17",
          3683 => x"8b",
          3684 => x"86",
          3685 => x"2b",
          3686 => x"48",
          3687 => x"05",
          3688 => x"b9",
          3689 => x"33",
          3690 => x"06",
          3691 => x"7b",
          3692 => x"b9",
          3693 => x"83",
          3694 => x"2b",
          3695 => x"33",
          3696 => x"5e",
          3697 => x"76",
          3698 => x"b9",
          3699 => x"12",
          3700 => x"07",
          3701 => x"33",
          3702 => x"40",
          3703 => x"78",
          3704 => x"84",
          3705 => x"33",
          3706 => x"66",
          3707 => x"52",
          3708 => x"fe",
          3709 => x"1e",
          3710 => x"5c",
          3711 => x"0b",
          3712 => x"84",
          3713 => x"7f",
          3714 => x"ed",
          3715 => x"76",
          3716 => x"b9",
          3717 => x"81",
          3718 => x"08",
          3719 => x"87",
          3720 => x"b9",
          3721 => x"07",
          3722 => x"2a",
          3723 => x"34",
          3724 => x"22",
          3725 => x"08",
          3726 => x"1c",
          3727 => x"51",
          3728 => x"39",
          3729 => x"8b",
          3730 => x"84",
          3731 => x"2b",
          3732 => x"43",
          3733 => x"63",
          3734 => x"08",
          3735 => x"33",
          3736 => x"74",
          3737 => x"71",
          3738 => x"5f",
          3739 => x"64",
          3740 => x"34",
          3741 => x"81",
          3742 => x"ff",
          3743 => x"58",
          3744 => x"34",
          3745 => x"33",
          3746 => x"83",
          3747 => x"12",
          3748 => x"2b",
          3749 => x"88",
          3750 => x"5d",
          3751 => x"83",
          3752 => x"1f",
          3753 => x"2b",
          3754 => x"33",
          3755 => x"81",
          3756 => x"5d",
          3757 => x"60",
          3758 => x"83",
          3759 => x"86",
          3760 => x"2b",
          3761 => x"18",
          3762 => x"07",
          3763 => x"41",
          3764 => x"1e",
          3765 => x"84",
          3766 => x"2b",
          3767 => x"14",
          3768 => x"07",
          3769 => x"5a",
          3770 => x"34",
          3771 => x"b8",
          3772 => x"71",
          3773 => x"70",
          3774 => x"75",
          3775 => x"b8",
          3776 => x"33",
          3777 => x"74",
          3778 => x"88",
          3779 => x"f8",
          3780 => x"54",
          3781 => x"7f",
          3782 => x"84",
          3783 => x"81",
          3784 => x"2b",
          3785 => x"33",
          3786 => x"06",
          3787 => x"5b",
          3788 => x"81",
          3789 => x"1f",
          3790 => x"8b",
          3791 => x"86",
          3792 => x"2b",
          3793 => x"14",
          3794 => x"07",
          3795 => x"5c",
          3796 => x"77",
          3797 => x"84",
          3798 => x"33",
          3799 => x"83",
          3800 => x"87",
          3801 => x"88",
          3802 => x"41",
          3803 => x"16",
          3804 => x"33",
          3805 => x"81",
          3806 => x"5c",
          3807 => x"1a",
          3808 => x"82",
          3809 => x"2b",
          3810 => x"33",
          3811 => x"70",
          3812 => x"5a",
          3813 => x"1a",
          3814 => x"70",
          3815 => x"71",
          3816 => x"33",
          3817 => x"70",
          3818 => x"5a",
          3819 => x"83",
          3820 => x"1f",
          3821 => x"88",
          3822 => x"83",
          3823 => x"84",
          3824 => x"b9",
          3825 => x"05",
          3826 => x"44",
          3827 => x"87",
          3828 => x"2b",
          3829 => x"1d",
          3830 => x"2a",
          3831 => x"61",
          3832 => x"34",
          3833 => x"11",
          3834 => x"71",
          3835 => x"33",
          3836 => x"70",
          3837 => x"59",
          3838 => x"7a",
          3839 => x"08",
          3840 => x"88",
          3841 => x"88",
          3842 => x"34",
          3843 => x"08",
          3844 => x"71",
          3845 => x"05",
          3846 => x"2b",
          3847 => x"06",
          3848 => x"5c",
          3849 => x"82",
          3850 => x"b9",
          3851 => x"12",
          3852 => x"07",
          3853 => x"71",
          3854 => x"70",
          3855 => x"59",
          3856 => x"1e",
          3857 => x"f3",
          3858 => x"a1",
          3859 => x"b9",
          3860 => x"53",
          3861 => x"fe",
          3862 => x"3f",
          3863 => x"38",
          3864 => x"7a",
          3865 => x"76",
          3866 => x"8a",
          3867 => x"3d",
          3868 => x"84",
          3869 => x"08",
          3870 => x"52",
          3871 => x"85",
          3872 => x"3d",
          3873 => x"b9",
          3874 => x"b4",
          3875 => x"84",
          3876 => x"84",
          3877 => x"81",
          3878 => x"08",
          3879 => x"85",
          3880 => x"76",
          3881 => x"34",
          3882 => x"22",
          3883 => x"83",
          3884 => x"51",
          3885 => x"89",
          3886 => x"10",
          3887 => x"f8",
          3888 => x"81",
          3889 => x"80",
          3890 => x"ff",
          3891 => x"81",
          3892 => x"b9",
          3893 => x"c8",
          3894 => x"0d",
          3895 => x"71",
          3896 => x"bb",
          3897 => x"06",
          3898 => x"c4",
          3899 => x"53",
          3900 => x"0d",
          3901 => x"02",
          3902 => x"57",
          3903 => x"38",
          3904 => x"81",
          3905 => x"73",
          3906 => x"0c",
          3907 => x"ca",
          3908 => x"06",
          3909 => x"c0",
          3910 => x"79",
          3911 => x"80",
          3912 => x"81",
          3913 => x"0c",
          3914 => x"81",
          3915 => x"56",
          3916 => x"39",
          3917 => x"8c",
          3918 => x"59",
          3919 => x"84",
          3920 => x"06",
          3921 => x"58",
          3922 => x"78",
          3923 => x"3f",
          3924 => x"55",
          3925 => x"98",
          3926 => x"78",
          3927 => x"06",
          3928 => x"54",
          3929 => x"8b",
          3930 => x"19",
          3931 => x"79",
          3932 => x"fc",
          3933 => x"05",
          3934 => x"53",
          3935 => x"87",
          3936 => x"72",
          3937 => x"38",
          3938 => x"81",
          3939 => x"71",
          3940 => x"38",
          3941 => x"86",
          3942 => x"0c",
          3943 => x"0d",
          3944 => x"84",
          3945 => x"71",
          3946 => x"53",
          3947 => x"81",
          3948 => x"2e",
          3949 => x"55",
          3950 => x"08",
          3951 => x"87",
          3952 => x"82",
          3953 => x"38",
          3954 => x"38",
          3955 => x"58",
          3956 => x"56",
          3957 => x"a8",
          3958 => x"81",
          3959 => x"18",
          3960 => x"c8",
          3961 => x"78",
          3962 => x"04",
          3963 => x"18",
          3964 => x"fc",
          3965 => x"08",
          3966 => x"84",
          3967 => x"18",
          3968 => x"1a",
          3969 => x"56",
          3970 => x"82",
          3971 => x"81",
          3972 => x"1b",
          3973 => x"fc",
          3974 => x"75",
          3975 => x"38",
          3976 => x"09",
          3977 => x"5a",
          3978 => x"70",
          3979 => x"76",
          3980 => x"19",
          3981 => x"34",
          3982 => x"b9",
          3983 => x"34",
          3984 => x"f2",
          3985 => x"0b",
          3986 => x"84",
          3987 => x"9f",
          3988 => x"84",
          3989 => x"7a",
          3990 => x"56",
          3991 => x"2a",
          3992 => x"18",
          3993 => x"7a",
          3994 => x"34",
          3995 => x"19",
          3996 => x"a7",
          3997 => x"70",
          3998 => x"53",
          3999 => x"e8",
          4000 => x"80",
          4001 => x"3f",
          4002 => x"b7",
          4003 => x"60",
          4004 => x"76",
          4005 => x"26",
          4006 => x"c8",
          4007 => x"33",
          4008 => x"38",
          4009 => x"81",
          4010 => x"81",
          4011 => x"08",
          4012 => x"08",
          4013 => x"5c",
          4014 => x"de",
          4015 => x"52",
          4016 => x"84",
          4017 => x"ff",
          4018 => x"7a",
          4019 => x"17",
          4020 => x"2a",
          4021 => x"59",
          4022 => x"80",
          4023 => x"5d",
          4024 => x"b5",
          4025 => x"52",
          4026 => x"84",
          4027 => x"ff",
          4028 => x"79",
          4029 => x"17",
          4030 => x"07",
          4031 => x"5d",
          4032 => x"76",
          4033 => x"8f",
          4034 => x"18",
          4035 => x"2e",
          4036 => x"71",
          4037 => x"81",
          4038 => x"53",
          4039 => x"f7",
          4040 => x"2e",
          4041 => x"b4",
          4042 => x"10",
          4043 => x"81",
          4044 => x"07",
          4045 => x"3d",
          4046 => x"06",
          4047 => x"18",
          4048 => x"2e",
          4049 => x"71",
          4050 => x"81",
          4051 => x"53",
          4052 => x"f6",
          4053 => x"2e",
          4054 => x"b4",
          4055 => x"82",
          4056 => x"05",
          4057 => x"90",
          4058 => x"33",
          4059 => x"71",
          4060 => x"84",
          4061 => x"5a",
          4062 => x"b4",
          4063 => x"81",
          4064 => x"81",
          4065 => x"09",
          4066 => x"c8",
          4067 => x"a8",
          4068 => x"5b",
          4069 => x"84",
          4070 => x"2e",
          4071 => x"54",
          4072 => x"53",
          4073 => x"98",
          4074 => x"54",
          4075 => x"53",
          4076 => x"3f",
          4077 => x"81",
          4078 => x"08",
          4079 => x"18",
          4080 => x"27",
          4081 => x"82",
          4082 => x"08",
          4083 => x"17",
          4084 => x"18",
          4085 => x"5a",
          4086 => x"81",
          4087 => x"08",
          4088 => x"18",
          4089 => x"5e",
          4090 => x"38",
          4091 => x"09",
          4092 => x"b4",
          4093 => x"7b",
          4094 => x"3f",
          4095 => x"b4",
          4096 => x"81",
          4097 => x"81",
          4098 => x"09",
          4099 => x"c8",
          4100 => x"a8",
          4101 => x"5b",
          4102 => x"91",
          4103 => x"2e",
          4104 => x"54",
          4105 => x"53",
          4106 => x"90",
          4107 => x"54",
          4108 => x"53",
          4109 => x"f8",
          4110 => x"f9",
          4111 => x"0d",
          4112 => x"58",
          4113 => x"1a",
          4114 => x"74",
          4115 => x"81",
          4116 => x"38",
          4117 => x"0d",
          4118 => x"05",
          4119 => x"5c",
          4120 => x"19",
          4121 => x"09",
          4122 => x"77",
          4123 => x"51",
          4124 => x"80",
          4125 => x"77",
          4126 => x"b0",
          4127 => x"05",
          4128 => x"76",
          4129 => x"79",
          4130 => x"34",
          4131 => x"0d",
          4132 => x"fe",
          4133 => x"08",
          4134 => x"58",
          4135 => x"83",
          4136 => x"2e",
          4137 => x"54",
          4138 => x"33",
          4139 => x"08",
          4140 => x"5a",
          4141 => x"fe",
          4142 => x"06",
          4143 => x"70",
          4144 => x"0a",
          4145 => x"7d",
          4146 => x"1d",
          4147 => x"1d",
          4148 => x"1d",
          4149 => x"e8",
          4150 => x"2a",
          4151 => x"59",
          4152 => x"80",
          4153 => x"5d",
          4154 => x"d4",
          4155 => x"52",
          4156 => x"84",
          4157 => x"ff",
          4158 => x"7b",
          4159 => x"ff",
          4160 => x"81",
          4161 => x"80",
          4162 => x"f0",
          4163 => x"56",
          4164 => x"1a",
          4165 => x"05",
          4166 => x"5f",
          4167 => x"54",
          4168 => x"1a",
          4169 => x"58",
          4170 => x"81",
          4171 => x"08",
          4172 => x"a8",
          4173 => x"b9",
          4174 => x"7a",
          4175 => x"74",
          4176 => x"75",
          4177 => x"ee",
          4178 => x"2e",
          4179 => x"b4",
          4180 => x"83",
          4181 => x"2a",
          4182 => x"2a",
          4183 => x"06",
          4184 => x"0b",
          4185 => x"54",
          4186 => x"1a",
          4187 => x"5a",
          4188 => x"81",
          4189 => x"08",
          4190 => x"a8",
          4191 => x"b9",
          4192 => x"77",
          4193 => x"55",
          4194 => x"bd",
          4195 => x"52",
          4196 => x"7b",
          4197 => x"53",
          4198 => x"52",
          4199 => x"b9",
          4200 => x"fd",
          4201 => x"1a",
          4202 => x"08",
          4203 => x"08",
          4204 => x"fc",
          4205 => x"82",
          4206 => x"81",
          4207 => x"19",
          4208 => x"fc",
          4209 => x"19",
          4210 => x"ed",
          4211 => x"08",
          4212 => x"38",
          4213 => x"b4",
          4214 => x"a0",
          4215 => x"5f",
          4216 => x"38",
          4217 => x"09",
          4218 => x"7c",
          4219 => x"51",
          4220 => x"39",
          4221 => x"81",
          4222 => x"58",
          4223 => x"fe",
          4224 => x"06",
          4225 => x"76",
          4226 => x"f9",
          4227 => x"7b",
          4228 => x"05",
          4229 => x"2b",
          4230 => x"07",
          4231 => x"34",
          4232 => x"34",
          4233 => x"34",
          4234 => x"34",
          4235 => x"7e",
          4236 => x"8a",
          4237 => x"2e",
          4238 => x"27",
          4239 => x"56",
          4240 => x"76",
          4241 => x"81",
          4242 => x"89",
          4243 => x"b2",
          4244 => x"3f",
          4245 => x"d0",
          4246 => x"81",
          4247 => x"09",
          4248 => x"70",
          4249 => x"82",
          4250 => x"06",
          4251 => x"b9",
          4252 => x"57",
          4253 => x"58",
          4254 => x"a4",
          4255 => x"08",
          4256 => x"55",
          4257 => x"38",
          4258 => x"26",
          4259 => x"81",
          4260 => x"83",
          4261 => x"ef",
          4262 => x"08",
          4263 => x"c8",
          4264 => x"80",
          4265 => x"08",
          4266 => x"85",
          4267 => x"9a",
          4268 => x"27",
          4269 => x"27",
          4270 => x"fe",
          4271 => x"38",
          4272 => x"f5",
          4273 => x"c8",
          4274 => x"07",
          4275 => x"c4",
          4276 => x"1a",
          4277 => x"1a",
          4278 => x"38",
          4279 => x"33",
          4280 => x"75",
          4281 => x"3d",
          4282 => x"0c",
          4283 => x"08",
          4284 => x"ff",
          4285 => x"51",
          4286 => x"55",
          4287 => x"84",
          4288 => x"ff",
          4289 => x"81",
          4290 => x"7a",
          4291 => x"f0",
          4292 => x"9f",
          4293 => x"90",
          4294 => x"80",
          4295 => x"26",
          4296 => x"82",
          4297 => x"79",
          4298 => x"19",
          4299 => x"08",
          4300 => x"38",
          4301 => x"73",
          4302 => x"19",
          4303 => x"0c",
          4304 => x"b9",
          4305 => x"17",
          4306 => x"38",
          4307 => x"59",
          4308 => x"08",
          4309 => x"80",
          4310 => x"17",
          4311 => x"05",
          4312 => x"91",
          4313 => x"3f",
          4314 => x"c8",
          4315 => x"84",
          4316 => x"9c",
          4317 => x"73",
          4318 => x"54",
          4319 => x"39",
          4320 => x"3d",
          4321 => x"08",
          4322 => x"57",
          4323 => x"80",
          4324 => x"55",
          4325 => x"79",
          4326 => x"81",
          4327 => x"a9",
          4328 => x"57",
          4329 => x"77",
          4330 => x"78",
          4331 => x"56",
          4332 => x"0d",
          4333 => x"22",
          4334 => x"7b",
          4335 => x"9c",
          4336 => x"56",
          4337 => x"d0",
          4338 => x"ff",
          4339 => x"b9",
          4340 => x"80",
          4341 => x"52",
          4342 => x"c8",
          4343 => x"08",
          4344 => x"84",
          4345 => x"38",
          4346 => x"2e",
          4347 => x"83",
          4348 => x"38",
          4349 => x"59",
          4350 => x"38",
          4351 => x"1b",
          4352 => x"0c",
          4353 => x"55",
          4354 => x"ff",
          4355 => x"8a",
          4356 => x"80",
          4357 => x"52",
          4358 => x"84",
          4359 => x"16",
          4360 => x"84",
          4361 => x"0d",
          4362 => x"b8",
          4363 => x"56",
          4364 => x"80",
          4365 => x"1a",
          4366 => x"31",
          4367 => x"e8",
          4368 => x"2e",
          4369 => x"54",
          4370 => x"53",
          4371 => x"c8",
          4372 => x"55",
          4373 => x"76",
          4374 => x"94",
          4375 => x"fe",
          4376 => x"27",
          4377 => x"71",
          4378 => x"0c",
          4379 => x"b9",
          4380 => x"3d",
          4381 => x"08",
          4382 => x"08",
          4383 => x"d2",
          4384 => x"58",
          4385 => x"38",
          4386 => x"78",
          4387 => x"81",
          4388 => x"19",
          4389 => x"c8",
          4390 => x"81",
          4391 => x"76",
          4392 => x"33",
          4393 => x"38",
          4394 => x"ff",
          4395 => x"76",
          4396 => x"32",
          4397 => x"25",
          4398 => x"93",
          4399 => x"61",
          4400 => x"2e",
          4401 => x"52",
          4402 => x"c8",
          4403 => x"b2",
          4404 => x"dc",
          4405 => x"3d",
          4406 => x"53",
          4407 => x"a8",
          4408 => x"78",
          4409 => x"84",
          4410 => x"19",
          4411 => x"c8",
          4412 => x"27",
          4413 => x"60",
          4414 => x"38",
          4415 => x"08",
          4416 => x"51",
          4417 => x"39",
          4418 => x"e7",
          4419 => x"7a",
          4420 => x"77",
          4421 => x"7f",
          4422 => x"7d",
          4423 => x"5d",
          4424 => x"2e",
          4425 => x"39",
          4426 => x"7a",
          4427 => x"04",
          4428 => x"33",
          4429 => x"cb",
          4430 => x"9a",
          4431 => x"56",
          4432 => x"70",
          4433 => x"51",
          4434 => x"c8",
          4435 => x"71",
          4436 => x"56",
          4437 => x"81",
          4438 => x"61",
          4439 => x"81",
          4440 => x"27",
          4441 => x"81",
          4442 => x"38",
          4443 => x"79",
          4444 => x"ff",
          4445 => x"fd",
          4446 => x"ca",
          4447 => x"7c",
          4448 => x"81",
          4449 => x"70",
          4450 => x"70",
          4451 => x"59",
          4452 => x"81",
          4453 => x"84",
          4454 => x"ef",
          4455 => x"80",
          4456 => x"b9",
          4457 => x"82",
          4458 => x"ff",
          4459 => x"98",
          4460 => x"08",
          4461 => x"33",
          4462 => x"81",
          4463 => x"53",
          4464 => x"dc",
          4465 => x"2e",
          4466 => x"b4",
          4467 => x"38",
          4468 => x"76",
          4469 => x"33",
          4470 => x"58",
          4471 => x"2e",
          4472 => x"06",
          4473 => x"74",
          4474 => x"e5",
          4475 => x"58",
          4476 => x"80",
          4477 => x"33",
          4478 => x"ff",
          4479 => x"74",
          4480 => x"33",
          4481 => x"0b",
          4482 => x"05",
          4483 => x"33",
          4484 => x"42",
          4485 => x"75",
          4486 => x"ff",
          4487 => x"51",
          4488 => x"5a",
          4489 => x"8f",
          4490 => x"3d",
          4491 => x"53",
          4492 => x"80",
          4493 => x"78",
          4494 => x"84",
          4495 => x"1b",
          4496 => x"c8",
          4497 => x"27",
          4498 => x"79",
          4499 => x"38",
          4500 => x"08",
          4501 => x"51",
          4502 => x"39",
          4503 => x"33",
          4504 => x"60",
          4505 => x"06",
          4506 => x"19",
          4507 => x"1f",
          4508 => x"5f",
          4509 => x"55",
          4510 => x"92",
          4511 => x"b9",
          4512 => x"fe",
          4513 => x"38",
          4514 => x"0c",
          4515 => x"7e",
          4516 => x"8c",
          4517 => x"33",
          4518 => x"76",
          4519 => x"06",
          4520 => x"77",
          4521 => x"79",
          4522 => x"88",
          4523 => x"2e",
          4524 => x"ff",
          4525 => x"3f",
          4526 => x"05",
          4527 => x"56",
          4528 => x"c8",
          4529 => x"38",
          4530 => x"27",
          4531 => x"2a",
          4532 => x"92",
          4533 => x"10",
          4534 => x"fe",
          4535 => x"06",
          4536 => x"84",
          4537 => x"76",
          4538 => x"81",
          4539 => x"0d",
          4540 => x"81",
          4541 => x"56",
          4542 => x"08",
          4543 => x"2e",
          4544 => x"70",
          4545 => x"95",
          4546 => x"7b",
          4547 => x"57",
          4548 => x"ff",
          4549 => x"db",
          4550 => x"76",
          4551 => x"0b",
          4552 => x"40",
          4553 => x"8b",
          4554 => x"81",
          4555 => x"58",
          4556 => x"85",
          4557 => x"22",
          4558 => x"74",
          4559 => x"81",
          4560 => x"70",
          4561 => x"81",
          4562 => x"2e",
          4563 => x"57",
          4564 => x"38",
          4565 => x"02",
          4566 => x"76",
          4567 => x"27",
          4568 => x"34",
          4569 => x"59",
          4570 => x"59",
          4571 => x"56",
          4572 => x"55",
          4573 => x"56",
          4574 => x"1a",
          4575 => x"09",
          4576 => x"a0",
          4577 => x"3d",
          4578 => x"33",
          4579 => x"76",
          4580 => x"8f",
          4581 => x"81",
          4582 => x"91",
          4583 => x"82",
          4584 => x"84",
          4585 => x"06",
          4586 => x"33",
          4587 => x"05",
          4588 => x"81",
          4589 => x"80",
          4590 => x"51",
          4591 => x"08",
          4592 => x"8c",
          4593 => x"b9",
          4594 => x"c8",
          4595 => x"08",
          4596 => x"2e",
          4597 => x"7f",
          4598 => x"38",
          4599 => x"81",
          4600 => x"b9",
          4601 => x"56",
          4602 => x"56",
          4603 => x"33",
          4604 => x"c9",
          4605 => x"07",
          4606 => x"38",
          4607 => x"89",
          4608 => x"3f",
          4609 => x"c8",
          4610 => x"58",
          4611 => x"58",
          4612 => x"7f",
          4613 => x"b4",
          4614 => x"1c",
          4615 => x"38",
          4616 => x"81",
          4617 => x"b9",
          4618 => x"57",
          4619 => x"58",
          4620 => x"1f",
          4621 => x"05",
          4622 => x"38",
          4623 => x"58",
          4624 => x"77",
          4625 => x"55",
          4626 => x"1f",
          4627 => x"1b",
          4628 => x"56",
          4629 => x"0d",
          4630 => x"72",
          4631 => x"38",
          4632 => x"c2",
          4633 => x"b9",
          4634 => x"fe",
          4635 => x"53",
          4636 => x"80",
          4637 => x"09",
          4638 => x"c8",
          4639 => x"a8",
          4640 => x"08",
          4641 => x"60",
          4642 => x"c8",
          4643 => x"2b",
          4644 => x"7d",
          4645 => x"08",
          4646 => x"38",
          4647 => x"8b",
          4648 => x"29",
          4649 => x"57",
          4650 => x"19",
          4651 => x"81",
          4652 => x"1e",
          4653 => x"77",
          4654 => x"7a",
          4655 => x"38",
          4656 => x"81",
          4657 => x"b9",
          4658 => x"57",
          4659 => x"58",
          4660 => x"9c",
          4661 => x"5c",
          4662 => x"8b",
          4663 => x"9a",
          4664 => x"8d",
          4665 => x"59",
          4666 => x"78",
          4667 => x"58",
          4668 => x"05",
          4669 => x"34",
          4670 => x"76",
          4671 => x"18",
          4672 => x"83",
          4673 => x"10",
          4674 => x"2e",
          4675 => x"0b",
          4676 => x"e9",
          4677 => x"84",
          4678 => x"ff",
          4679 => x"eb",
          4680 => x"b8",
          4681 => x"59",
          4682 => x"c8",
          4683 => x"08",
          4684 => x"1d",
          4685 => x"41",
          4686 => x"38",
          4687 => x"09",
          4688 => x"b4",
          4689 => x"78",
          4690 => x"3f",
          4691 => x"1f",
          4692 => x"81",
          4693 => x"38",
          4694 => x"76",
          4695 => x"39",
          4696 => x"39",
          4697 => x"52",
          4698 => x"84",
          4699 => x"06",
          4700 => x"1d",
          4701 => x"31",
          4702 => x"38",
          4703 => x"aa",
          4704 => x"f8",
          4705 => x"80",
          4706 => x"75",
          4707 => x"59",
          4708 => x"fa",
          4709 => x"a0",
          4710 => x"1c",
          4711 => x"39",
          4712 => x"08",
          4713 => x"51",
          4714 => x"3d",
          4715 => x"5c",
          4716 => x"08",
          4717 => x"08",
          4718 => x"71",
          4719 => x"58",
          4720 => x"38",
          4721 => x"1b",
          4722 => x"80",
          4723 => x"06",
          4724 => x"83",
          4725 => x"22",
          4726 => x"7a",
          4727 => x"06",
          4728 => x"57",
          4729 => x"89",
          4730 => x"16",
          4731 => x"74",
          4732 => x"81",
          4733 => x"70",
          4734 => x"77",
          4735 => x"8b",
          4736 => x"34",
          4737 => x"05",
          4738 => x"27",
          4739 => x"55",
          4740 => x"33",
          4741 => x"38",
          4742 => x"7c",
          4743 => x"17",
          4744 => x"55",
          4745 => x"34",
          4746 => x"88",
          4747 => x"83",
          4748 => x"2b",
          4749 => x"70",
          4750 => x"07",
          4751 => x"17",
          4752 => x"5b",
          4753 => x"1e",
          4754 => x"71",
          4755 => x"1e",
          4756 => x"55",
          4757 => x"81",
          4758 => x"b5",
          4759 => x"81",
          4760 => x"83",
          4761 => x"27",
          4762 => x"38",
          4763 => x"74",
          4764 => x"80",
          4765 => x"19",
          4766 => x"79",
          4767 => x"30",
          4768 => x"72",
          4769 => x"80",
          4770 => x"05",
          4771 => x"5b",
          4772 => x"5a",
          4773 => x"38",
          4774 => x"89",
          4775 => x"78",
          4776 => x"8c",
          4777 => x"b4",
          4778 => x"06",
          4779 => x"14",
          4780 => x"73",
          4781 => x"16",
          4782 => x"33",
          4783 => x"b7",
          4784 => x"53",
          4785 => x"25",
          4786 => x"58",
          4787 => x"70",
          4788 => x"70",
          4789 => x"83",
          4790 => x"81",
          4791 => x"38",
          4792 => x"33",
          4793 => x"9f",
          4794 => x"8c",
          4795 => x"70",
          4796 => x"81",
          4797 => x"2e",
          4798 => x"27",
          4799 => x"76",
          4800 => x"ff",
          4801 => x"73",
          4802 => x"5b",
          4803 => x"dc",
          4804 => x"26",
          4805 => x"e4",
          4806 => x"54",
          4807 => x"73",
          4808 => x"33",
          4809 => x"73",
          4810 => x"7a",
          4811 => x"80",
          4812 => x"7d",
          4813 => x"05",
          4814 => x"2e",
          4815 => x"73",
          4816 => x"25",
          4817 => x"80",
          4818 => x"54",
          4819 => x"2e",
          4820 => x"30",
          4821 => x"57",
          4822 => x"73",
          4823 => x"55",
          4824 => x"39",
          4825 => x"e7",
          4826 => x"ff",
          4827 => x"54",
          4828 => x"0d",
          4829 => x"ff",
          4830 => x"e3",
          4831 => x"1d",
          4832 => x"3f",
          4833 => x"0c",
          4834 => x"dc",
          4835 => x"07",
          4836 => x"a1",
          4837 => x"33",
          4838 => x"38",
          4839 => x"80",
          4840 => x"e1",
          4841 => x"82",
          4842 => x"38",
          4843 => x"17",
          4844 => x"17",
          4845 => x"a0",
          4846 => x"42",
          4847 => x"84",
          4848 => x"76",
          4849 => x"80",
          4850 => x"38",
          4851 => x"06",
          4852 => x"2e",
          4853 => x"06",
          4854 => x"76",
          4855 => x"05",
          4856 => x"9d",
          4857 => x"ff",
          4858 => x"fe",
          4859 => x"2e",
          4860 => x"a0",
          4861 => x"05",
          4862 => x"38",
          4863 => x"70",
          4864 => x"74",
          4865 => x"2e",
          4866 => x"30",
          4867 => x"77",
          4868 => x"38",
          4869 => x"81",
          4870 => x"72",
          4871 => x"51",
          4872 => x"38",
          4873 => x"77",
          4874 => x"75",
          4875 => x"5b",
          4876 => x"77",
          4877 => x"22",
          4878 => x"95",
          4879 => x"e5",
          4880 => x"82",
          4881 => x"8c",
          4882 => x"55",
          4883 => x"81",
          4884 => x"7d",
          4885 => x"38",
          4886 => x"81",
          4887 => x"79",
          4888 => x"7b",
          4889 => x"08",
          4890 => x"c8",
          4891 => x"b9",
          4892 => x"fb",
          4893 => x"5a",
          4894 => x"82",
          4895 => x"38",
          4896 => x"8c",
          4897 => x"39",
          4898 => x"22",
          4899 => x"f0",
          4900 => x"79",
          4901 => x"18",
          4902 => x"06",
          4903 => x"ae",
          4904 => x"76",
          4905 => x"0b",
          4906 => x"73",
          4907 => x"70",
          4908 => x"8a",
          4909 => x"58",
          4910 => x"bf",
          4911 => x"33",
          4912 => x"d6",
          4913 => x"77",
          4914 => x"84",
          4915 => x"2e",
          4916 => x"ff",
          4917 => x"80",
          4918 => x"62",
          4919 => x"2e",
          4920 => x"7b",
          4921 => x"77",
          4922 => x"38",
          4923 => x"fb",
          4924 => x"56",
          4925 => x"81",
          4926 => x"77",
          4927 => x"38",
          4928 => x"85",
          4929 => x"09",
          4930 => x"ff",
          4931 => x"84",
          4932 => x"74",
          4933 => x"75",
          4934 => x"78",
          4935 => x"07",
          4936 => x"a4",
          4937 => x"52",
          4938 => x"b9",
          4939 => x"87",
          4940 => x"2e",
          4941 => x"e5",
          4942 => x"ff",
          4943 => x"81",
          4944 => x"e4",
          4945 => x"54",
          4946 => x"73",
          4947 => x"33",
          4948 => x"73",
          4949 => x"78",
          4950 => x"73",
          4951 => x"70",
          4952 => x"15",
          4953 => x"81",
          4954 => x"70",
          4955 => x"53",
          4956 => x"34",
          4957 => x"fc",
          4958 => x"e4",
          4959 => x"53",
          4960 => x"df",
          4961 => x"5b",
          4962 => x"5b",
          4963 => x"cc",
          4964 => x"2b",
          4965 => x"57",
          4966 => x"75",
          4967 => x"81",
          4968 => x"74",
          4969 => x"39",
          4970 => x"5a",
          4971 => x"fa",
          4972 => x"2a",
          4973 => x"85",
          4974 => x"0d",
          4975 => x"88",
          4976 => x"5e",
          4977 => x"59",
          4978 => x"38",
          4979 => x"9f",
          4980 => x"d0",
          4981 => x"85",
          4982 => x"80",
          4983 => x"10",
          4984 => x"5a",
          4985 => x"38",
          4986 => x"77",
          4987 => x"38",
          4988 => x"3f",
          4989 => x"70",
          4990 => x"86",
          4991 => x"5d",
          4992 => x"34",
          4993 => x"bb",
          4994 => x"ff",
          4995 => x"58",
          4996 => x"8d",
          4997 => x"8a",
          4998 => x"7a",
          4999 => x"0c",
          5000 => x"53",
          5001 => x"52",
          5002 => x"c8",
          5003 => x"81",
          5004 => x"78",
          5005 => x"b6",
          5006 => x"56",
          5007 => x"85",
          5008 => x"84",
          5009 => x"bf",
          5010 => x"cd",
          5011 => x"c5",
          5012 => x"18",
          5013 => x"7c",
          5014 => x"ad",
          5015 => x"18",
          5016 => x"75",
          5017 => x"33",
          5018 => x"88",
          5019 => x"07",
          5020 => x"5a",
          5021 => x"18",
          5022 => x"34",
          5023 => x"81",
          5024 => x"7c",
          5025 => x"ff",
          5026 => x"33",
          5027 => x"77",
          5028 => x"ff",
          5029 => x"38",
          5030 => x"33",
          5031 => x"88",
          5032 => x"5a",
          5033 => x"cc",
          5034 => x"88",
          5035 => x"80",
          5036 => x"33",
          5037 => x"81",
          5038 => x"75",
          5039 => x"42",
          5040 => x"c6",
          5041 => x"58",
          5042 => x"38",
          5043 => x"79",
          5044 => x"74",
          5045 => x"84",
          5046 => x"08",
          5047 => x"c8",
          5048 => x"83",
          5049 => x"26",
          5050 => x"26",
          5051 => x"70",
          5052 => x"7b",
          5053 => x"b0",
          5054 => x"8a",
          5055 => x"58",
          5056 => x"16",
          5057 => x"82",
          5058 => x"81",
          5059 => x"83",
          5060 => x"78",
          5061 => x"0b",
          5062 => x"0c",
          5063 => x"83",
          5064 => x"84",
          5065 => x"84",
          5066 => x"84",
          5067 => x"0b",
          5068 => x"b9",
          5069 => x"0b",
          5070 => x"04",
          5071 => x"06",
          5072 => x"38",
          5073 => x"05",
          5074 => x"38",
          5075 => x"40",
          5076 => x"70",
          5077 => x"05",
          5078 => x"56",
          5079 => x"70",
          5080 => x"17",
          5081 => x"17",
          5082 => x"30",
          5083 => x"2e",
          5084 => x"be",
          5085 => x"72",
          5086 => x"55",
          5087 => x"1c",
          5088 => x"ff",
          5089 => x"78",
          5090 => x"2a",
          5091 => x"c5",
          5092 => x"78",
          5093 => x"09",
          5094 => x"81",
          5095 => x"7b",
          5096 => x"38",
          5097 => x"93",
          5098 => x"fa",
          5099 => x"2e",
          5100 => x"80",
          5101 => x"2b",
          5102 => x"07",
          5103 => x"07",
          5104 => x"7a",
          5105 => x"90",
          5106 => x"be",
          5107 => x"30",
          5108 => x"3d",
          5109 => x"b6",
          5110 => x"78",
          5111 => x"80",
          5112 => x"ff",
          5113 => x"56",
          5114 => x"7a",
          5115 => x"51",
          5116 => x"08",
          5117 => x"56",
          5118 => x"bf",
          5119 => x"88",
          5120 => x"82",
          5121 => x"38",
          5122 => x"75",
          5123 => x"81",
          5124 => x"7a",
          5125 => x"75",
          5126 => x"77",
          5127 => x"b9",
          5128 => x"2e",
          5129 => x"81",
          5130 => x"2e",
          5131 => x"5a",
          5132 => x"f8",
          5133 => x"83",
          5134 => x"81",
          5135 => x"40",
          5136 => x"52",
          5137 => x"38",
          5138 => x"81",
          5139 => x"58",
          5140 => x"70",
          5141 => x"ff",
          5142 => x"2e",
          5143 => x"38",
          5144 => x"7c",
          5145 => x"0c",
          5146 => x"80",
          5147 => x"8a",
          5148 => x"ff",
          5149 => x"0c",
          5150 => x"ee",
          5151 => x"78",
          5152 => x"81",
          5153 => x"1b",
          5154 => x"83",
          5155 => x"85",
          5156 => x"5c",
          5157 => x"33",
          5158 => x"71",
          5159 => x"77",
          5160 => x"2e",
          5161 => x"83",
          5162 => x"c6",
          5163 => x"18",
          5164 => x"75",
          5165 => x"38",
          5166 => x"08",
          5167 => x"5b",
          5168 => x"9b",
          5169 => x"52",
          5170 => x"3f",
          5171 => x"38",
          5172 => x"0c",
          5173 => x"34",
          5174 => x"33",
          5175 => x"82",
          5176 => x"fc",
          5177 => x"12",
          5178 => x"07",
          5179 => x"2b",
          5180 => x"45",
          5181 => x"a4",
          5182 => x"38",
          5183 => x"12",
          5184 => x"07",
          5185 => x"2b",
          5186 => x"5b",
          5187 => x"e4",
          5188 => x"38",
          5189 => x"12",
          5190 => x"07",
          5191 => x"2b",
          5192 => x"5d",
          5193 => x"12",
          5194 => x"07",
          5195 => x"2b",
          5196 => x"0c",
          5197 => x"45",
          5198 => x"d1",
          5199 => x"d1",
          5200 => x"d1",
          5201 => x"98",
          5202 => x"24",
          5203 => x"56",
          5204 => x"08",
          5205 => x"33",
          5206 => x"b9",
          5207 => x"81",
          5208 => x"18",
          5209 => x"31",
          5210 => x"38",
          5211 => x"81",
          5212 => x"fd",
          5213 => x"f3",
          5214 => x"83",
          5215 => x"39",
          5216 => x"33",
          5217 => x"58",
          5218 => x"42",
          5219 => x"83",
          5220 => x"2b",
          5221 => x"70",
          5222 => x"07",
          5223 => x"5a",
          5224 => x"39",
          5225 => x"38",
          5226 => x"2e",
          5227 => x"5a",
          5228 => x"79",
          5229 => x"54",
          5230 => x"53",
          5231 => x"ad",
          5232 => x"0d",
          5233 => x"43",
          5234 => x"5a",
          5235 => x"78",
          5236 => x"26",
          5237 => x"38",
          5238 => x"d9",
          5239 => x"74",
          5240 => x"84",
          5241 => x"73",
          5242 => x"62",
          5243 => x"74",
          5244 => x"54",
          5245 => x"93",
          5246 => x"81",
          5247 => x"84",
          5248 => x"8b",
          5249 => x"0d",
          5250 => x"ff",
          5251 => x"91",
          5252 => x"d0",
          5253 => x"f7",
          5254 => x"5e",
          5255 => x"79",
          5256 => x"81",
          5257 => x"57",
          5258 => x"15",
          5259 => x"9f",
          5260 => x"e0",
          5261 => x"74",
          5262 => x"76",
          5263 => x"ff",
          5264 => x"70",
          5265 => x"57",
          5266 => x"1b",
          5267 => x"ff",
          5268 => x"7a",
          5269 => x"0c",
          5270 => x"6c",
          5271 => x"56",
          5272 => x"38",
          5273 => x"cc",
          5274 => x"58",
          5275 => x"57",
          5276 => x"38",
          5277 => x"b9",
          5278 => x"40",
          5279 => x"e1",
          5280 => x"84",
          5281 => x"38",
          5282 => x"81",
          5283 => x"38",
          5284 => x"88",
          5285 => x"83",
          5286 => x"81",
          5287 => x"12",
          5288 => x"33",
          5289 => x"2e",
          5290 => x"34",
          5291 => x"90",
          5292 => x"34",
          5293 => x"7e",
          5294 => x"34",
          5295 => x"5d",
          5296 => x"5b",
          5297 => x"9d",
          5298 => x"80",
          5299 => x"0b",
          5300 => x"e2",
          5301 => x"08",
          5302 => x"89",
          5303 => x"8a",
          5304 => x"a3",
          5305 => x"98",
          5306 => x"b8",
          5307 => x"7c",
          5308 => x"02",
          5309 => x"81",
          5310 => x"77",
          5311 => x"2e",
          5312 => x"81",
          5313 => x"56",
          5314 => x"c0",
          5315 => x"1b",
          5316 => x"11",
          5317 => x"07",
          5318 => x"7b",
          5319 => x"1a",
          5320 => x"12",
          5321 => x"07",
          5322 => x"2b",
          5323 => x"05",
          5324 => x"59",
          5325 => x"1a",
          5326 => x"91",
          5327 => x"77",
          5328 => x"2e",
          5329 => x"f1",
          5330 => x"22",
          5331 => x"76",
          5332 => x"5b",
          5333 => x"70",
          5334 => x"84",
          5335 => x"ac",
          5336 => x"84",
          5337 => x"82",
          5338 => x"80",
          5339 => x"39",
          5340 => x"5e",
          5341 => x"06",
          5342 => x"88",
          5343 => x"87",
          5344 => x"84",
          5345 => x"79",
          5346 => x"08",
          5347 => x"c8",
          5348 => x"31",
          5349 => x"33",
          5350 => x"90",
          5351 => x"fd",
          5352 => x"81",
          5353 => x"ab",
          5354 => x"84",
          5355 => x"38",
          5356 => x"d9",
          5357 => x"83",
          5358 => x"51",
          5359 => x"08",
          5360 => x"11",
          5361 => x"75",
          5362 => x"18",
          5363 => x"74",
          5364 => x"26",
          5365 => x"0b",
          5366 => x"34",
          5367 => x"17",
          5368 => x"07",
          5369 => x"8e",
          5370 => x"a1",
          5371 => x"91",
          5372 => x"17",
          5373 => x"9a",
          5374 => x"7d",
          5375 => x"06",
          5376 => x"7f",
          5377 => x"16",
          5378 => x"33",
          5379 => x"b5",
          5380 => x"52",
          5381 => x"3f",
          5382 => x"38",
          5383 => x"0c",
          5384 => x"0c",
          5385 => x"80",
          5386 => x"b4",
          5387 => x"81",
          5388 => x"3f",
          5389 => x"81",
          5390 => x"08",
          5391 => x"17",
          5392 => x"55",
          5393 => x"38",
          5394 => x"09",
          5395 => x"b4",
          5396 => x"79",
          5397 => x"b8",
          5398 => x"94",
          5399 => x"77",
          5400 => x"75",
          5401 => x"f8",
          5402 => x"08",
          5403 => x"27",
          5404 => x"71",
          5405 => x"74",
          5406 => x"2a",
          5407 => x"ed",
          5408 => x"f7",
          5409 => x"f7",
          5410 => x"80",
          5411 => x"57",
          5412 => x"62",
          5413 => x"80",
          5414 => x"9f",
          5415 => x"97",
          5416 => x"8f",
          5417 => x"59",
          5418 => x"80",
          5419 => x"8c",
          5420 => x"84",
          5421 => x"87",
          5422 => x"94",
          5423 => x"56",
          5424 => x"7b",
          5425 => x"75",
          5426 => x"38",
          5427 => x"2a",
          5428 => x"d3",
          5429 => x"27",
          5430 => x"f0",
          5431 => x"98",
          5432 => x"fe",
          5433 => x"e7",
          5434 => x"b0",
          5435 => x"2e",
          5436 => x"2a",
          5437 => x"38",
          5438 => x"38",
          5439 => x"53",
          5440 => x"9f",
          5441 => x"98",
          5442 => x"75",
          5443 => x"77",
          5444 => x"84",
          5445 => x"58",
          5446 => x"33",
          5447 => x"15",
          5448 => x"58",
          5449 => x"0c",
          5450 => x"59",
          5451 => x"af",
          5452 => x"0c",
          5453 => x"c8",
          5454 => x"fe",
          5455 => x"83",
          5456 => x"5b",
          5457 => x"76",
          5458 => x"38",
          5459 => x"41",
          5460 => x"80",
          5461 => x"19",
          5462 => x"b1",
          5463 => x"85",
          5464 => x"1a",
          5465 => x"1b",
          5466 => x"5a",
          5467 => x"2e",
          5468 => x"56",
          5469 => x"ff",
          5470 => x"38",
          5471 => x"70",
          5472 => x"75",
          5473 => x"b4",
          5474 => x"81",
          5475 => x"3f",
          5476 => x"2e",
          5477 => x"b9",
          5478 => x"08",
          5479 => x"08",
          5480 => x"fe",
          5481 => x"82",
          5482 => x"81",
          5483 => x"05",
          5484 => x"ff",
          5485 => x"39",
          5486 => x"56",
          5487 => x"79",
          5488 => x"c8",
          5489 => x"33",
          5490 => x"c8",
          5491 => x"38",
          5492 => x"39",
          5493 => x"84",
          5494 => x"82",
          5495 => x"b9",
          5496 => x"3d",
          5497 => x"5c",
          5498 => x"80",
          5499 => x"80",
          5500 => x"80",
          5501 => x"1b",
          5502 => x"fd",
          5503 => x"76",
          5504 => x"74",
          5505 => x"81",
          5506 => x"76",
          5507 => x"08",
          5508 => x"84",
          5509 => x"82",
          5510 => x"7e",
          5511 => x"ff",
          5512 => x"78",
          5513 => x"1a",
          5514 => x"38",
          5515 => x"ff",
          5516 => x"0c",
          5517 => x"1b",
          5518 => x"1b",
          5519 => x"08",
          5520 => x"58",
          5521 => x"8a",
          5522 => x"08",
          5523 => x"de",
          5524 => x"5c",
          5525 => x"19",
          5526 => x"79",
          5527 => x"52",
          5528 => x"3f",
          5529 => x"60",
          5530 => x"74",
          5531 => x"b8",
          5532 => x"56",
          5533 => x"70",
          5534 => x"75",
          5535 => x"34",
          5536 => x"7e",
          5537 => x"1c",
          5538 => x"8c",
          5539 => x"75",
          5540 => x"8c",
          5541 => x"1a",
          5542 => x"7a",
          5543 => x"b9",
          5544 => x"84",
          5545 => x"83",
          5546 => x"60",
          5547 => x"08",
          5548 => x"80",
          5549 => x"83",
          5550 => x"08",
          5551 => x"17",
          5552 => x"2e",
          5553 => x"54",
          5554 => x"33",
          5555 => x"c8",
          5556 => x"81",
          5557 => x"bf",
          5558 => x"06",
          5559 => x"56",
          5560 => x"70",
          5561 => x"05",
          5562 => x"38",
          5563 => x"fe",
          5564 => x"53",
          5565 => x"52",
          5566 => x"84",
          5567 => x"06",
          5568 => x"83",
          5569 => x"08",
          5570 => x"74",
          5571 => x"82",
          5572 => x"81",
          5573 => x"16",
          5574 => x"52",
          5575 => x"3f",
          5576 => x"08",
          5577 => x"38",
          5578 => x"38",
          5579 => x"08",
          5580 => x"58",
          5581 => x"79",
          5582 => x"c8",
          5583 => x"d8",
          5584 => x"39",
          5585 => x"3f",
          5586 => x"c8",
          5587 => x"54",
          5588 => x"53",
          5589 => x"b8",
          5590 => x"38",
          5591 => x"b4",
          5592 => x"77",
          5593 => x"82",
          5594 => x"81",
          5595 => x"16",
          5596 => x"52",
          5597 => x"3f",
          5598 => x"33",
          5599 => x"c8",
          5600 => x"38",
          5601 => x"39",
          5602 => x"16",
          5603 => x"ff",
          5604 => x"80",
          5605 => x"17",
          5606 => x"31",
          5607 => x"98",
          5608 => x"2e",
          5609 => x"54",
          5610 => x"53",
          5611 => x"96",
          5612 => x"94",
          5613 => x"81",
          5614 => x"b9",
          5615 => x"0b",
          5616 => x"c8",
          5617 => x"0d",
          5618 => x"9f",
          5619 => x"97",
          5620 => x"8f",
          5621 => x"58",
          5622 => x"80",
          5623 => x"d8",
          5624 => x"81",
          5625 => x"c8",
          5626 => x"b4",
          5627 => x"17",
          5628 => x"54",
          5629 => x"33",
          5630 => x"c8",
          5631 => x"81",
          5632 => x"90",
          5633 => x"a0",
          5634 => x"77",
          5635 => x"ff",
          5636 => x"34",
          5637 => x"34",
          5638 => x"56",
          5639 => x"8c",
          5640 => x"88",
          5641 => x"90",
          5642 => x"98",
          5643 => x"7a",
          5644 => x"0b",
          5645 => x"18",
          5646 => x"0b",
          5647 => x"83",
          5648 => x"3f",
          5649 => x"81",
          5650 => x"34",
          5651 => x"0d",
          5652 => x"b8",
          5653 => x"5b",
          5654 => x"b9",
          5655 => x"c8",
          5656 => x"a8",
          5657 => x"57",
          5658 => x"8e",
          5659 => x"2e",
          5660 => x"54",
          5661 => x"53",
          5662 => x"92",
          5663 => x"78",
          5664 => x"74",
          5665 => x"8c",
          5666 => x"88",
          5667 => x"90",
          5668 => x"98",
          5669 => x"7a",
          5670 => x"0b",
          5671 => x"18",
          5672 => x"0b",
          5673 => x"83",
          5674 => x"3f",
          5675 => x"81",
          5676 => x"34",
          5677 => x"ff",
          5678 => x"81",
          5679 => x"78",
          5680 => x"3d",
          5681 => x"3f",
          5682 => x"c8",
          5683 => x"2e",
          5684 => x"2e",
          5685 => x"2e",
          5686 => x"22",
          5687 => x"80",
          5688 => x"38",
          5689 => x"0c",
          5690 => x"51",
          5691 => x"08",
          5692 => x"75",
          5693 => x"0d",
          5694 => x"80",
          5695 => x"57",
          5696 => x"ba",
          5697 => x"ba",
          5698 => x"51",
          5699 => x"d1",
          5700 => x"0c",
          5701 => x"b9",
          5702 => x"33",
          5703 => x"53",
          5704 => x"19",
          5705 => x"54",
          5706 => x"0b",
          5707 => x"79",
          5708 => x"33",
          5709 => x"9f",
          5710 => x"89",
          5711 => x"53",
          5712 => x"26",
          5713 => x"06",
          5714 => x"55",
          5715 => x"85",
          5716 => x"32",
          5717 => x"76",
          5718 => x"92",
          5719 => x"83",
          5720 => x"fe",
          5721 => x"77",
          5722 => x"3d",
          5723 => x"52",
          5724 => x"b9",
          5725 => x"80",
          5726 => x"0c",
          5727 => x"52",
          5728 => x"3f",
          5729 => x"c8",
          5730 => x"05",
          5731 => x"77",
          5732 => x"33",
          5733 => x"75",
          5734 => x"11",
          5735 => x"07",
          5736 => x"79",
          5737 => x"0c",
          5738 => x"0d",
          5739 => x"09",
          5740 => x"84",
          5741 => x"95",
          5742 => x"2b",
          5743 => x"1b",
          5744 => x"98",
          5745 => x"0c",
          5746 => x"0d",
          5747 => x"08",
          5748 => x"80",
          5749 => x"e5",
          5750 => x"c8",
          5751 => x"c8",
          5752 => x"61",
          5753 => x"58",
          5754 => x"80",
          5755 => x"98",
          5756 => x"ff",
          5757 => x"59",
          5758 => x"60",
          5759 => x"16",
          5760 => x"c8",
          5761 => x"83",
          5762 => x"16",
          5763 => x"c9",
          5764 => x"85",
          5765 => x"17",
          5766 => x"3d",
          5767 => x"71",
          5768 => x"40",
          5769 => x"da",
          5770 => x"52",
          5771 => x"b9",
          5772 => x"82",
          5773 => x"a8",
          5774 => x"84",
          5775 => x"3d",
          5776 => x"71",
          5777 => x"58",
          5778 => x"fd",
          5779 => x"b9",
          5780 => x"e2",
          5781 => x"b9",
          5782 => x"78",
          5783 => x"c8",
          5784 => x"52",
          5785 => x"7f",
          5786 => x"2e",
          5787 => x"81",
          5788 => x"f5",
          5789 => x"81",
          5790 => x"7e",
          5791 => x"e6",
          5792 => x"59",
          5793 => x"76",
          5794 => x"08",
          5795 => x"da",
          5796 => x"77",
          5797 => x"84",
          5798 => x"e5",
          5799 => x"59",
          5800 => x"38",
          5801 => x"5f",
          5802 => x"7a",
          5803 => x"7a",
          5804 => x"33",
          5805 => x"17",
          5806 => x"7c",
          5807 => x"2e",
          5808 => x"59",
          5809 => x"0c",
          5810 => x"33",
          5811 => x"90",
          5812 => x"fd",
          5813 => x"33",
          5814 => x"79",
          5815 => x"80",
          5816 => x"84",
          5817 => x"08",
          5818 => x"39",
          5819 => x"16",
          5820 => x"ff",
          5821 => x"c8",
          5822 => x"08",
          5823 => x"17",
          5824 => x"55",
          5825 => x"38",
          5826 => x"09",
          5827 => x"b4",
          5828 => x"7d",
          5829 => x"b8",
          5830 => x"18",
          5831 => x"af",
          5832 => x"33",
          5833 => x"70",
          5834 => x"5a",
          5835 => x"e8",
          5836 => x"08",
          5837 => x"7c",
          5838 => x"27",
          5839 => x"18",
          5840 => x"70",
          5841 => x"d4",
          5842 => x"7c",
          5843 => x"e4",
          5844 => x"7d",
          5845 => x"9f",
          5846 => x"97",
          5847 => x"8f",
          5848 => x"59",
          5849 => x"80",
          5850 => x"c2",
          5851 => x"ba",
          5852 => x"26",
          5853 => x"80",
          5854 => x"79",
          5855 => x"5a",
          5856 => x"75",
          5857 => x"3f",
          5858 => x"54",
          5859 => x"3f",
          5860 => x"d5",
          5861 => x"17",
          5862 => x"56",
          5863 => x"38",
          5864 => x"76",
          5865 => x"0c",
          5866 => x"06",
          5867 => x"fe",
          5868 => x"f3",
          5869 => x"b9",
          5870 => x"73",
          5871 => x"82",
          5872 => x"08",
          5873 => x"0c",
          5874 => x"34",
          5875 => x"8b",
          5876 => x"81",
          5877 => x"bb",
          5878 => x"80",
          5879 => x"fe",
          5880 => x"15",
          5881 => x"73",
          5882 => x"c0",
          5883 => x"83",
          5884 => x"38",
          5885 => x"77",
          5886 => x"c8",
          5887 => x"94",
          5888 => x"80",
          5889 => x"0c",
          5890 => x"a8",
          5891 => x"15",
          5892 => x"ff",
          5893 => x"79",
          5894 => x"5a",
          5895 => x"38",
          5896 => x"18",
          5897 => x"5a",
          5898 => x"8c",
          5899 => x"52",
          5900 => x"b9",
          5901 => x"14",
          5902 => x"b9",
          5903 => x"cf",
          5904 => x"c9",
          5905 => x"cb",
          5906 => x"b9",
          5907 => x"b9",
          5908 => x"84",
          5909 => x"98",
          5910 => x"91",
          5911 => x"0c",
          5912 => x"7c",
          5913 => x"38",
          5914 => x"8d",
          5915 => x"84",
          5916 => x"08",
          5917 => x"74",
          5918 => x"3d",
          5919 => x"75",
          5920 => x"c8",
          5921 => x"d1",
          5922 => x"59",
          5923 => x"16",
          5924 => x"54",
          5925 => x"16",
          5926 => x"71",
          5927 => x"5d",
          5928 => x"38",
          5929 => x"18",
          5930 => x"51",
          5931 => x"08",
          5932 => x"80",
          5933 => x"fe",
          5934 => x"fe",
          5935 => x"33",
          5936 => x"7a",
          5937 => x"bc",
          5938 => x"54",
          5939 => x"53",
          5940 => x"52",
          5941 => x"22",
          5942 => x"2e",
          5943 => x"84",
          5944 => x"c8",
          5945 => x"33",
          5946 => x"c8",
          5947 => x"71",
          5948 => x"3d",
          5949 => x"74",
          5950 => x"73",
          5951 => x"72",
          5952 => x"84",
          5953 => x"81",
          5954 => x"53",
          5955 => x"80",
          5956 => x"9d",
          5957 => x"84",
          5958 => x"84",
          5959 => x"74",
          5960 => x"74",
          5961 => x"c8",
          5962 => x"07",
          5963 => x"55",
          5964 => x"8a",
          5965 => x"52",
          5966 => x"74",
          5967 => x"c8",
          5968 => x"07",
          5969 => x"55",
          5970 => x"51",
          5971 => x"08",
          5972 => x"04",
          5973 => x"3f",
          5974 => x"72",
          5975 => x"56",
          5976 => x"57",
          5977 => x"3d",
          5978 => x"c8",
          5979 => x"2e",
          5980 => x"95",
          5981 => x"ff",
          5982 => x"55",
          5983 => x"80",
          5984 => x"58",
          5985 => x"2e",
          5986 => x"b0",
          5987 => x"95",
          5988 => x"c8",
          5989 => x"0d",
          5990 => x"3d",
          5991 => x"b9",
          5992 => x"b9",
          5993 => x"74",
          5994 => x"13",
          5995 => x"26",
          5996 => x"b9",
          5997 => x"b9",
          5998 => x"81",
          5999 => x"08",
          6000 => x"77",
          6001 => x"5c",
          6002 => x"82",
          6003 => x"5d",
          6004 => x"53",
          6005 => x"fe",
          6006 => x"80",
          6007 => x"79",
          6008 => x"7d",
          6009 => x"82",
          6010 => x"05",
          6011 => x"90",
          6012 => x"33",
          6013 => x"71",
          6014 => x"70",
          6015 => x"84",
          6016 => x"43",
          6017 => x"40",
          6018 => x"7f",
          6019 => x"33",
          6020 => x"79",
          6021 => x"04",
          6022 => x"17",
          6023 => x"fe",
          6024 => x"c8",
          6025 => x"08",
          6026 => x"18",
          6027 => x"55",
          6028 => x"38",
          6029 => x"09",
          6030 => x"b4",
          6031 => x"7c",
          6032 => x"e0",
          6033 => x"77",
          6034 => x"77",
          6035 => x"c8",
          6036 => x"b9",
          6037 => x"84",
          6038 => x"c8",
          6039 => x"18",
          6040 => x"08",
          6041 => x"7a",
          6042 => x"07",
          6043 => x"39",
          6044 => x"71",
          6045 => x"70",
          6046 => x"06",
          6047 => x"5f",
          6048 => x"39",
          6049 => x"58",
          6050 => x"0c",
          6051 => x"84",
          6052 => x"58",
          6053 => x"57",
          6054 => x"76",
          6055 => x"74",
          6056 => x"86",
          6057 => x"78",
          6058 => x"73",
          6059 => x"33",
          6060 => x"33",
          6061 => x"87",
          6062 => x"94",
          6063 => x"27",
          6064 => x"17",
          6065 => x"27",
          6066 => x"b3",
          6067 => x"0c",
          6068 => x"80",
          6069 => x"75",
          6070 => x"34",
          6071 => x"8b",
          6072 => x"27",
          6073 => x"fe",
          6074 => x"59",
          6075 => x"e9",
          6076 => x"82",
          6077 => x"2e",
          6078 => x"75",
          6079 => x"c8",
          6080 => x"fe",
          6081 => x"74",
          6082 => x"94",
          6083 => x"54",
          6084 => x"79",
          6085 => x"15",
          6086 => x"b9",
          6087 => x"95",
          6088 => x"8f",
          6089 => x"54",
          6090 => x"fe",
          6091 => x"51",
          6092 => x"08",
          6093 => x"c8",
          6094 => x"81",
          6095 => x"08",
          6096 => x"84",
          6097 => x"08",
          6098 => x"c8",
          6099 => x"c8",
          6100 => x"38",
          6101 => x"74",
          6102 => x"84",
          6103 => x"08",
          6104 => x"fe",
          6105 => x"59",
          6106 => x"cb",
          6107 => x"80",
          6108 => x"2e",
          6109 => x"75",
          6110 => x"c8",
          6111 => x"fe",
          6112 => x"74",
          6113 => x"17",
          6114 => x"73",
          6115 => x"26",
          6116 => x"90",
          6117 => x"56",
          6118 => x"33",
          6119 => x"e7",
          6120 => x"54",
          6121 => x"90",
          6122 => x"81",
          6123 => x"f0",
          6124 => x"39",
          6125 => x"0d",
          6126 => x"52",
          6127 => x"84",
          6128 => x"08",
          6129 => x"c8",
          6130 => x"a8",
          6131 => x"59",
          6132 => x"08",
          6133 => x"02",
          6134 => x"81",
          6135 => x"38",
          6136 => x"c4",
          6137 => x"81",
          6138 => x"b4",
          6139 => x"33",
          6140 => x"73",
          6141 => x"83",
          6142 => x"81",
          6143 => x"38",
          6144 => x"ff",
          6145 => x"b9",
          6146 => x"55",
          6147 => x"08",
          6148 => x"38",
          6149 => x"ff",
          6150 => x"56",
          6151 => x"0b",
          6152 => x"04",
          6153 => x"98",
          6154 => x"5d",
          6155 => x"c8",
          6156 => x"c8",
          6157 => x"a8",
          6158 => x"2e",
          6159 => x"ff",
          6160 => x"56",
          6161 => x"38",
          6162 => x"56",
          6163 => x"80",
          6164 => x"55",
          6165 => x"08",
          6166 => x"75",
          6167 => x"db",
          6168 => x"c8",
          6169 => x"5d",
          6170 => x"17",
          6171 => x"17",
          6172 => x"09",
          6173 => x"75",
          6174 => x"51",
          6175 => x"08",
          6176 => x"58",
          6177 => x"ab",
          6178 => x"34",
          6179 => x"08",
          6180 => x"78",
          6181 => x"c8",
          6182 => x"2e",
          6183 => x"81",
          6184 => x"c8",
          6185 => x"7c",
          6186 => x"90",
          6187 => x"7a",
          6188 => x"84",
          6189 => x"17",
          6190 => x"c8",
          6191 => x"27",
          6192 => x"74",
          6193 => x"38",
          6194 => x"08",
          6195 => x"51",
          6196 => x"c5",
          6197 => x"e1",
          6198 => x"e4",
          6199 => x"b9",
          6200 => x"84",
          6201 => x"38",
          6202 => x"cb",
          6203 => x"fe",
          6204 => x"b3",
          6205 => x"19",
          6206 => x"ff",
          6207 => x"84",
          6208 => x"18",
          6209 => x"a1",
          6210 => x"56",
          6211 => x"56",
          6212 => x"39",
          6213 => x"ff",
          6214 => x"b2",
          6215 => x"84",
          6216 => x"75",
          6217 => x"04",
          6218 => x"52",
          6219 => x"c8",
          6220 => x"38",
          6221 => x"3d",
          6222 => x"2e",
          6223 => x"f3",
          6224 => x"56",
          6225 => x"7d",
          6226 => x"5d",
          6227 => x"08",
          6228 => x"83",
          6229 => x"81",
          6230 => x"08",
          6231 => x"c9",
          6232 => x"12",
          6233 => x"38",
          6234 => x"5a",
          6235 => x"38",
          6236 => x"19",
          6237 => x"0c",
          6238 => x"55",
          6239 => x"ff",
          6240 => x"8a",
          6241 => x"f9",
          6242 => x"52",
          6243 => x"3f",
          6244 => x"81",
          6245 => x"84",
          6246 => x"b8",
          6247 => x"58",
          6248 => x"b9",
          6249 => x"08",
          6250 => x"18",
          6251 => x"27",
          6252 => x"7a",
          6253 => x"38",
          6254 => x"08",
          6255 => x"51",
          6256 => x"81",
          6257 => x"7c",
          6258 => x"08",
          6259 => x"51",
          6260 => x"08",
          6261 => x"fd",
          6262 => x"2e",
          6263 => x"ff",
          6264 => x"52",
          6265 => x"b9",
          6266 => x"08",
          6267 => x"59",
          6268 => x"94",
          6269 => x"5c",
          6270 => x"7a",
          6271 => x"c8",
          6272 => x"22",
          6273 => x"81",
          6274 => x"fe",
          6275 => x"56",
          6276 => x"ff",
          6277 => x"ae",
          6278 => x"0b",
          6279 => x"80",
          6280 => x"34",
          6281 => x"cc",
          6282 => x"83",
          6283 => x"d2",
          6284 => x"80",
          6285 => x"83",
          6286 => x"0b",
          6287 => x"56",
          6288 => x"70",
          6289 => x"75",
          6290 => x"d9",
          6291 => x"ff",
          6292 => x"17",
          6293 => x"f3",
          6294 => x"2e",
          6295 => x"83",
          6296 => x"3f",
          6297 => x"c8",
          6298 => x"b9",
          6299 => x"c8",
          6300 => x"17",
          6301 => x"7d",
          6302 => x"77",
          6303 => x"7c",
          6304 => x"38",
          6305 => x"7d",
          6306 => x"51",
          6307 => x"08",
          6308 => x"3d",
          6309 => x"80",
          6310 => x"76",
          6311 => x"7b",
          6312 => x"34",
          6313 => x"17",
          6314 => x"1a",
          6315 => x"39",
          6316 => x"34",
          6317 => x"34",
          6318 => x"7d",
          6319 => x"51",
          6320 => x"08",
          6321 => x"b3",
          6322 => x"5f",
          6323 => x"81",
          6324 => x"56",
          6325 => x"ed",
          6326 => x"82",
          6327 => x"b2",
          6328 => x"b9",
          6329 => x"80",
          6330 => x"0c",
          6331 => x"0c",
          6332 => x"52",
          6333 => x"c8",
          6334 => x"38",
          6335 => x"06",
          6336 => x"0b",
          6337 => x"55",
          6338 => x"70",
          6339 => x"74",
          6340 => x"7a",
          6341 => x"57",
          6342 => x"ff",
          6343 => x"08",
          6344 => x"84",
          6345 => x"08",
          6346 => x"2e",
          6347 => x"c8",
          6348 => x"d0",
          6349 => x"58",
          6350 => x"78",
          6351 => x"78",
          6352 => x"08",
          6353 => x"5e",
          6354 => x"5c",
          6355 => x"ff",
          6356 => x"26",
          6357 => x"06",
          6358 => x"99",
          6359 => x"ff",
          6360 => x"2a",
          6361 => x"06",
          6362 => x"7a",
          6363 => x"2a",
          6364 => x"2e",
          6365 => x"5c",
          6366 => x"08",
          6367 => x"83",
          6368 => x"82",
          6369 => x"b2",
          6370 => x"b9",
          6371 => x"fd",
          6372 => x"3d",
          6373 => x"38",
          6374 => x"b9",
          6375 => x"fd",
          6376 => x"19",
          6377 => x"56",
          6378 => x"75",
          6379 => x"5a",
          6380 => x"33",
          6381 => x"84",
          6382 => x"38",
          6383 => x"34",
          6384 => x"8b",
          6385 => x"57",
          6386 => x"a7",
          6387 => x"7f",
          6388 => x"88",
          6389 => x"57",
          6390 => x"16",
          6391 => x"75",
          6392 => x"22",
          6393 => x"57",
          6394 => x"75",
          6395 => x"2e",
          6396 => x"83",
          6397 => x"17",
          6398 => x"f1",
          6399 => x"85",
          6400 => x"18",
          6401 => x"56",
          6402 => x"33",
          6403 => x"bb",
          6404 => x"5d",
          6405 => x"88",
          6406 => x"76",
          6407 => x"06",
          6408 => x"80",
          6409 => x"75",
          6410 => x"0b",
          6411 => x"08",
          6412 => x"ff",
          6413 => x"fe",
          6414 => x"55",
          6415 => x"b8",
          6416 => x"5a",
          6417 => x"83",
          6418 => x"2e",
          6419 => x"54",
          6420 => x"33",
          6421 => x"c8",
          6422 => x"81",
          6423 => x"77",
          6424 => x"7a",
          6425 => x"19",
          6426 => x"78",
          6427 => x"c8",
          6428 => x"2e",
          6429 => x"2e",
          6430 => x"db",
          6431 => x"84",
          6432 => x"b1",
          6433 => x"c8",
          6434 => x"33",
          6435 => x"90",
          6436 => x"fd",
          6437 => x"2e",
          6438 => x"80",
          6439 => x"c8",
          6440 => x"b4",
          6441 => x"33",
          6442 => x"84",
          6443 => x"06",
          6444 => x"83",
          6445 => x"08",
          6446 => x"74",
          6447 => x"82",
          6448 => x"81",
          6449 => x"16",
          6450 => x"52",
          6451 => x"3f",
          6452 => x"b4",
          6453 => x"81",
          6454 => x"3f",
          6455 => x"c9",
          6456 => x"34",
          6457 => x"84",
          6458 => x"18",
          6459 => x"33",
          6460 => x"fc",
          6461 => x"a0",
          6462 => x"17",
          6463 => x"5c",
          6464 => x"80",
          6465 => x"e3",
          6466 => x"3d",
          6467 => x"a2",
          6468 => x"84",
          6469 => x"75",
          6470 => x"04",
          6471 => x"05",
          6472 => x"c8",
          6473 => x"38",
          6474 => x"06",
          6475 => x"a7",
          6476 => x"71",
          6477 => x"57",
          6478 => x"81",
          6479 => x"e2",
          6480 => x"b9",
          6481 => x"3d",
          6482 => x"cc",
          6483 => x"d9",
          6484 => x"b9",
          6485 => x"84",
          6486 => x"78",
          6487 => x"51",
          6488 => x"08",
          6489 => x"02",
          6490 => x"56",
          6491 => x"18",
          6492 => x"07",
          6493 => x"76",
          6494 => x"76",
          6495 => x"76",
          6496 => x"78",
          6497 => x"51",
          6498 => x"08",
          6499 => x"04",
          6500 => x"80",
          6501 => x"3d",
          6502 => x"c8",
          6503 => x"84",
          6504 => x"56",
          6505 => x"70",
          6506 => x"38",
          6507 => x"56",
          6508 => x"81",
          6509 => x"2e",
          6510 => x"58",
          6511 => x"2e",
          6512 => x"5a",
          6513 => x"81",
          6514 => x"16",
          6515 => x"c9",
          6516 => x"85",
          6517 => x"17",
          6518 => x"70",
          6519 => x"83",
          6520 => x"84",
          6521 => x"b8",
          6522 => x"71",
          6523 => x"14",
          6524 => x"33",
          6525 => x"57",
          6526 => x"9a",
          6527 => x"80",
          6528 => x"f4",
          6529 => x"84",
          6530 => x"38",
          6531 => x"b8",
          6532 => x"b0",
          6533 => x"b8",
          6534 => x"5b",
          6535 => x"b9",
          6536 => x"fe",
          6537 => x"17",
          6538 => x"31",
          6539 => x"a0",
          6540 => x"16",
          6541 => x"06",
          6542 => x"08",
          6543 => x"81",
          6544 => x"79",
          6545 => x"52",
          6546 => x"3f",
          6547 => x"8d",
          6548 => x"51",
          6549 => x"08",
          6550 => x"38",
          6551 => x"08",
          6552 => x"19",
          6553 => x"75",
          6554 => x"ec",
          6555 => x"76",
          6556 => x"ff",
          6557 => x"58",
          6558 => x"39",
          6559 => x"0d",
          6560 => x"52",
          6561 => x"84",
          6562 => x"08",
          6563 => x"7d",
          6564 => x"58",
          6565 => x"74",
          6566 => x"ff",
          6567 => x"27",
          6568 => x"5c",
          6569 => x"57",
          6570 => x"0c",
          6571 => x"38",
          6572 => x"52",
          6573 => x"3f",
          6574 => x"06",
          6575 => x"83",
          6576 => x"70",
          6577 => x"80",
          6578 => x"77",
          6579 => x"70",
          6580 => x"80",
          6581 => x"81",
          6582 => x"59",
          6583 => x"27",
          6584 => x"96",
          6585 => x"76",
          6586 => x"05",
          6587 => x"70",
          6588 => x"3d",
          6589 => x"5b",
          6590 => x"d1",
          6591 => x"76",
          6592 => x"2e",
          6593 => x"16",
          6594 => x"09",
          6595 => x"79",
          6596 => x"52",
          6597 => x"e4",
          6598 => x"b9",
          6599 => x"56",
          6600 => x"0d",
          6601 => x"e7",
          6602 => x"ff",
          6603 => x"56",
          6604 => x"0d",
          6605 => x"c3",
          6606 => x"ee",
          6607 => x"b9",
          6608 => x"2e",
          6609 => x"57",
          6610 => x"76",
          6611 => x"55",
          6612 => x"83",
          6613 => x"3f",
          6614 => x"ff",
          6615 => x"38",
          6616 => x"c8",
          6617 => x"ee",
          6618 => x"e6",
          6619 => x"58",
          6620 => x"08",
          6621 => x"09",
          6622 => x"c8",
          6623 => x"08",
          6624 => x"2e",
          6625 => x"79",
          6626 => x"81",
          6627 => x"18",
          6628 => x"b9",
          6629 => x"57",
          6630 => x"57",
          6631 => x"70",
          6632 => x"2e",
          6633 => x"25",
          6634 => x"81",
          6635 => x"2e",
          6636 => x"ef",
          6637 => x"84",
          6638 => x"38",
          6639 => x"38",
          6640 => x"6c",
          6641 => x"58",
          6642 => x"6b",
          6643 => x"6c",
          6644 => x"05",
          6645 => x"34",
          6646 => x"eb",
          6647 => x"76",
          6648 => x"55",
          6649 => x"5a",
          6650 => x"83",
          6651 => x"3f",
          6652 => x"39",
          6653 => x"b4",
          6654 => x"33",
          6655 => x"c8",
          6656 => x"c3",
          6657 => x"34",
          6658 => x"5c",
          6659 => x"82",
          6660 => x"38",
          6661 => x"39",
          6662 => x"ed",
          6663 => x"84",
          6664 => x"38",
          6665 => x"78",
          6666 => x"39",
          6667 => x"08",
          6668 => x"51",
          6669 => x"f2",
          6670 => x"80",
          6671 => x"56",
          6672 => x"55",
          6673 => x"54",
          6674 => x"22",
          6675 => x"2e",
          6676 => x"75",
          6677 => x"75",
          6678 => x"a2",
          6679 => x"90",
          6680 => x"56",
          6681 => x"7e",
          6682 => x"55",
          6683 => x"cb",
          6684 => x"70",
          6685 => x"08",
          6686 => x"5f",
          6687 => x"9c",
          6688 => x"58",
          6689 => x"52",
          6690 => x"15",
          6691 => x"26",
          6692 => x"08",
          6693 => x"c8",
          6694 => x"b9",
          6695 => x"59",
          6696 => x"2e",
          6697 => x"75",
          6698 => x"3d",
          6699 => x"0c",
          6700 => x"51",
          6701 => x"08",
          6702 => x"73",
          6703 => x"7b",
          6704 => x"56",
          6705 => x"18",
          6706 => x"73",
          6707 => x"dd",
          6708 => x"b9",
          6709 => x"19",
          6710 => x"38",
          6711 => x"80",
          6712 => x"0c",
          6713 => x"80",
          6714 => x"9c",
          6715 => x"58",
          6716 => x"76",
          6717 => x"33",
          6718 => x"75",
          6719 => x"97",
          6720 => x"39",
          6721 => x"fe",
          6722 => x"39",
          6723 => x"a3",
          6724 => x"05",
          6725 => x"ff",
          6726 => x"40",
          6727 => x"70",
          6728 => x"56",
          6729 => x"74",
          6730 => x"38",
          6731 => x"24",
          6732 => x"d1",
          6733 => x"80",
          6734 => x"16",
          6735 => x"bd",
          6736 => x"79",
          6737 => x"c8",
          6738 => x"5d",
          6739 => x"75",
          6740 => x"7f",
          6741 => x"53",
          6742 => x"3f",
          6743 => x"6d",
          6744 => x"74",
          6745 => x"ff",
          6746 => x"38",
          6747 => x"7f",
          6748 => x"0a",
          6749 => x"06",
          6750 => x"2a",
          6751 => x"2b",
          6752 => x"2e",
          6753 => x"25",
          6754 => x"83",
          6755 => x"38",
          6756 => x"51",
          6757 => x"b9",
          6758 => x"ff",
          6759 => x"71",
          6760 => x"77",
          6761 => x"82",
          6762 => x"83",
          6763 => x"2e",
          6764 => x"11",
          6765 => x"71",
          6766 => x"72",
          6767 => x"83",
          6768 => x"33",
          6769 => x"81",
          6770 => x"75",
          6771 => x"42",
          6772 => x"4e",
          6773 => x"78",
          6774 => x"82",
          6775 => x"26",
          6776 => x"81",
          6777 => x"f9",
          6778 => x"2e",
          6779 => x"83",
          6780 => x"46",
          6781 => x"c2",
          6782 => x"57",
          6783 => x"58",
          6784 => x"26",
          6785 => x"10",
          6786 => x"74",
          6787 => x"ee",
          6788 => x"83",
          6789 => x"05",
          6790 => x"26",
          6791 => x"08",
          6792 => x"11",
          6793 => x"83",
          6794 => x"a0",
          6795 => x"66",
          6796 => x"31",
          6797 => x"89",
          6798 => x"29",
          6799 => x"79",
          6800 => x"7d",
          6801 => x"56",
          6802 => x"08",
          6803 => x"62",
          6804 => x"38",
          6805 => x"08",
          6806 => x"38",
          6807 => x"89",
          6808 => x"8b",
          6809 => x"3d",
          6810 => x"4e",
          6811 => x"c8",
          6812 => x"0c",
          6813 => x"ff",
          6814 => x"91",
          6815 => x"d0",
          6816 => x"b2",
          6817 => x"5c",
          6818 => x"81",
          6819 => x"58",
          6820 => x"62",
          6821 => x"81",
          6822 => x"45",
          6823 => x"70",
          6824 => x"70",
          6825 => x"09",
          6826 => x"38",
          6827 => x"07",
          6828 => x"7a",
          6829 => x"84",
          6830 => x"98",
          6831 => x"3d",
          6832 => x"fe",
          6833 => x"c8",
          6834 => x"77",
          6835 => x"75",
          6836 => x"57",
          6837 => x"7f",
          6838 => x"fa",
          6839 => x"38",
          6840 => x"95",
          6841 => x"67",
          6842 => x"70",
          6843 => x"84",
          6844 => x"38",
          6845 => x"80",
          6846 => x"76",
          6847 => x"84",
          6848 => x"81",
          6849 => x"27",
          6850 => x"57",
          6851 => x"57",
          6852 => x"34",
          6853 => x"61",
          6854 => x"70",
          6855 => x"05",
          6856 => x"38",
          6857 => x"82",
          6858 => x"05",
          6859 => x"6a",
          6860 => x"5c",
          6861 => x"90",
          6862 => x"5a",
          6863 => x"9e",
          6864 => x"05",
          6865 => x"26",
          6866 => x"06",
          6867 => x"88",
          6868 => x"f8",
          6869 => x"05",
          6870 => x"61",
          6871 => x"34",
          6872 => x"2a",
          6873 => x"90",
          6874 => x"7e",
          6875 => x"b9",
          6876 => x"83",
          6877 => x"05",
          6878 => x"61",
          6879 => x"05",
          6880 => x"74",
          6881 => x"4b",
          6882 => x"61",
          6883 => x"34",
          6884 => x"59",
          6885 => x"33",
          6886 => x"15",
          6887 => x"05",
          6888 => x"ff",
          6889 => x"54",
          6890 => x"c6",
          6891 => x"08",
          6892 => x"83",
          6893 => x"55",
          6894 => x"ff",
          6895 => x"41",
          6896 => x"87",
          6897 => x"83",
          6898 => x"88",
          6899 => x"81",
          6900 => x"78",
          6901 => x"98",
          6902 => x"65",
          6903 => x"59",
          6904 => x"51",
          6905 => x"08",
          6906 => x"55",
          6907 => x"ff",
          6908 => x"77",
          6909 => x"7f",
          6910 => x"89",
          6911 => x"38",
          6912 => x"83",
          6913 => x"60",
          6914 => x"84",
          6915 => x"1b",
          6916 => x"38",
          6917 => x"86",
          6918 => x"38",
          6919 => x"81",
          6920 => x"2a",
          6921 => x"84",
          6922 => x"81",
          6923 => x"f4",
          6924 => x"6b",
          6925 => x"67",
          6926 => x"67",
          6927 => x"34",
          6928 => x"80",
          6929 => x"f8",
          6930 => x"84",
          6931 => x"57",
          6932 => x"c8",
          6933 => x"83",
          6934 => x"05",
          6935 => x"84",
          6936 => x"34",
          6937 => x"88",
          6938 => x"34",
          6939 => x"cc",
          6940 => x"61",
          6941 => x"53",
          6942 => x"3f",
          6943 => x"c9",
          6944 => x"fe",
          6945 => x"c8",
          6946 => x"08",
          6947 => x"84",
          6948 => x"e4",
          6949 => x"f6",
          6950 => x"2a",
          6951 => x"56",
          6952 => x"77",
          6953 => x"77",
          6954 => x"58",
          6955 => x"27",
          6956 => x"f6",
          6957 => x"10",
          6958 => x"5c",
          6959 => x"08",
          6960 => x"ff",
          6961 => x"8e",
          6962 => x"08",
          6963 => x"7a",
          6964 => x"7a",
          6965 => x"39",
          6966 => x"f8",
          6967 => x"75",
          6968 => x"49",
          6969 => x"2a",
          6970 => x"98",
          6971 => x"f9",
          6972 => x"34",
          6973 => x"61",
          6974 => x"80",
          6975 => x"34",
          6976 => x"05",
          6977 => x"a6",
          6978 => x"61",
          6979 => x"34",
          6980 => x"ae",
          6981 => x"81",
          6982 => x"05",
          6983 => x"61",
          6984 => x"c0",
          6985 => x"34",
          6986 => x"a4",
          6987 => x"58",
          6988 => x"ff",
          6989 => x"38",
          6990 => x"70",
          6991 => x"74",
          6992 => x"80",
          6993 => x"d9",
          6994 => x"f4",
          6995 => x"42",
          6996 => x"54",
          6997 => x"79",
          6998 => x"39",
          6999 => x"3d",
          7000 => x"61",
          7001 => x"05",
          7002 => x"4c",
          7003 => x"05",
          7004 => x"61",
          7005 => x"34",
          7006 => x"89",
          7007 => x"8f",
          7008 => x"76",
          7009 => x"51",
          7010 => x"56",
          7011 => x"34",
          7012 => x"5c",
          7013 => x"34",
          7014 => x"05",
          7015 => x"05",
          7016 => x"f2",
          7017 => x"61",
          7018 => x"83",
          7019 => x"e7",
          7020 => x"61",
          7021 => x"59",
          7022 => x"90",
          7023 => x"34",
          7024 => x"eb",
          7025 => x"34",
          7026 => x"61",
          7027 => x"ef",
          7028 => x"aa",
          7029 => x"60",
          7030 => x"81",
          7031 => x"51",
          7032 => x"55",
          7033 => x"61",
          7034 => x"5a",
          7035 => x"8d",
          7036 => x"81",
          7037 => x"b4",
          7038 => x"9e",
          7039 => x"2e",
          7040 => x"58",
          7041 => x"86",
          7042 => x"76",
          7043 => x"55",
          7044 => x"0d",
          7045 => x"05",
          7046 => x"2e",
          7047 => x"80",
          7048 => x"77",
          7049 => x"34",
          7050 => x"38",
          7051 => x"18",
          7052 => x"fc",
          7053 => x"76",
          7054 => x"7a",
          7055 => x"2a",
          7056 => x"88",
          7057 => x"8d",
          7058 => x"a3",
          7059 => x"05",
          7060 => x"77",
          7061 => x"58",
          7062 => x"a1",
          7063 => x"80",
          7064 => x"80",
          7065 => x"56",
          7066 => x"74",
          7067 => x"0c",
          7068 => x"80",
          7069 => x"ac",
          7070 => x"76",
          7071 => x"b9",
          7072 => x"ba",
          7073 => x"9f",
          7074 => x"11",
          7075 => x"08",
          7076 => x"32",
          7077 => x"70",
          7078 => x"39",
          7079 => x"ff",
          7080 => x"9f",
          7081 => x"02",
          7082 => x"80",
          7083 => x"72",
          7084 => x"b9",
          7085 => x"ff",
          7086 => x"2e",
          7087 => x"2e",
          7088 => x"72",
          7089 => x"83",
          7090 => x"ff",
          7091 => x"8c",
          7092 => x"81",
          7093 => x"b9",
          7094 => x"fe",
          7095 => x"84",
          7096 => x"53",
          7097 => x"53",
          7098 => x"0d",
          7099 => x"06",
          7100 => x"38",
          7101 => x"22",
          7102 => x"0d",
          7103 => x"83",
          7104 => x"83",
          7105 => x"56",
          7106 => x"74",
          7107 => x"30",
          7108 => x"54",
          7109 => x"70",
          7110 => x"2a",
          7111 => x"52",
          7112 => x"cf",
          7113 => x"05",
          7114 => x"25",
          7115 => x"70",
          7116 => x"84",
          7117 => x"83",
          7118 => x"88",
          7119 => x"c9",
          7120 => x"a0",
          7121 => x"51",
          7122 => x"70",
          7123 => x"39",
          7124 => x"57",
          7125 => x"ff",
          7126 => x"16",
          7127 => x"d0",
          7128 => x"06",
          7129 => x"83",
          7130 => x"39",
          7131 => x"31",
          7132 => x"55",
          7133 => x"75",
          7134 => x"39",
          7135 => x"00",
          7136 => x"ff",
          7137 => x"00",
          7138 => x"00",
          7139 => x"00",
          7140 => x"00",
          7141 => x"00",
          7142 => x"00",
          7143 => x"00",
          7144 => x"00",
          7145 => x"00",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"69",
          7374 => x"69",
          7375 => x"69",
          7376 => x"6c",
          7377 => x"65",
          7378 => x"63",
          7379 => x"63",
          7380 => x"64",
          7381 => x"64",
          7382 => x"65",
          7383 => x"65",
          7384 => x"69",
          7385 => x"66",
          7386 => x"00",
          7387 => x"65",
          7388 => x"65",
          7389 => x"6e",
          7390 => x"65",
          7391 => x"6c",
          7392 => x"62",
          7393 => x"62",
          7394 => x"69",
          7395 => x"64",
          7396 => x"77",
          7397 => x"2e",
          7398 => x"65",
          7399 => x"63",
          7400 => x"00",
          7401 => x"61",
          7402 => x"20",
          7403 => x"00",
          7404 => x"66",
          7405 => x"6d",
          7406 => x"00",
          7407 => x"69",
          7408 => x"64",
          7409 => x"75",
          7410 => x"61",
          7411 => x"6e",
          7412 => x"00",
          7413 => x"74",
          7414 => x"64",
          7415 => x"6d",
          7416 => x"20",
          7417 => x"74",
          7418 => x"64",
          7419 => x"6b",
          7420 => x"6e",
          7421 => x"6c",
          7422 => x"72",
          7423 => x"62",
          7424 => x"6e",
          7425 => x"00",
          7426 => x"20",
          7427 => x"72",
          7428 => x"2e",
          7429 => x"68",
          7430 => x"6e",
          7431 => x"00",
          7432 => x"61",
          7433 => x"65",
          7434 => x"00",
          7435 => x"73",
          7436 => x"2e",
          7437 => x"69",
          7438 => x"61",
          7439 => x"6f",
          7440 => x"6f",
          7441 => x"6f",
          7442 => x"6f",
          7443 => x"69",
          7444 => x"72",
          7445 => x"6e",
          7446 => x"65",
          7447 => x"69",
          7448 => x"72",
          7449 => x"73",
          7450 => x"25",
          7451 => x"73",
          7452 => x"25",
          7453 => x"73",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"30",
          7458 => x"7c",
          7459 => x"20",
          7460 => x"00",
          7461 => x"20",
          7462 => x"4f",
          7463 => x"20",
          7464 => x"2f",
          7465 => x"31",
          7466 => x"5a",
          7467 => x"20",
          7468 => x"73",
          7469 => x"0a",
          7470 => x"20",
          7471 => x"41",
          7472 => x"20",
          7473 => x"20",
          7474 => x"38",
          7475 => x"20",
          7476 => x"64",
          7477 => x"20",
          7478 => x"20",
          7479 => x"38",
          7480 => x"50",
          7481 => x"72",
          7482 => x"64",
          7483 => x"41",
          7484 => x"69",
          7485 => x"74",
          7486 => x"20",
          7487 => x"72",
          7488 => x"41",
          7489 => x"69",
          7490 => x"74",
          7491 => x"20",
          7492 => x"72",
          7493 => x"4f",
          7494 => x"69",
          7495 => x"74",
          7496 => x"20",
          7497 => x"72",
          7498 => x"53",
          7499 => x"72",
          7500 => x"69",
          7501 => x"65",
          7502 => x"65",
          7503 => x"70",
          7504 => x"2e",
          7505 => x"69",
          7506 => x"72",
          7507 => x"75",
          7508 => x"62",
          7509 => x"4f",
          7510 => x"73",
          7511 => x"64",
          7512 => x"74",
          7513 => x"73",
          7514 => x"30",
          7515 => x"65",
          7516 => x"61",
          7517 => x"00",
          7518 => x"64",
          7519 => x"3a",
          7520 => x"6f",
          7521 => x"00",
          7522 => x"69",
          7523 => x"73",
          7524 => x"00",
          7525 => x"72",
          7526 => x"67",
          7527 => x"65",
          7528 => x"67",
          7529 => x"61",
          7530 => x"00",
          7531 => x"6e",
          7532 => x"40",
          7533 => x"2e",
          7534 => x"61",
          7535 => x"72",
          7536 => x"65",
          7537 => x"00",
          7538 => x"74",
          7539 => x"65",
          7540 => x"78",
          7541 => x"30",
          7542 => x"6c",
          7543 => x"30",
          7544 => x"58",
          7545 => x"72",
          7546 => x"00",
          7547 => x"28",
          7548 => x"25",
          7549 => x"38",
          7550 => x"6f",
          7551 => x"2e",
          7552 => x"20",
          7553 => x"6c",
          7554 => x"2e",
          7555 => x"75",
          7556 => x"72",
          7557 => x"6c",
          7558 => x"64",
          7559 => x"00",
          7560 => x"79",
          7561 => x"74",
          7562 => x"6e",
          7563 => x"65",
          7564 => x"61",
          7565 => x"3f",
          7566 => x"2f",
          7567 => x"64",
          7568 => x"64",
          7569 => x"6f",
          7570 => x"74",
          7571 => x"0a",
          7572 => x"20",
          7573 => x"6e",
          7574 => x"64",
          7575 => x"3a",
          7576 => x"50",
          7577 => x"20",
          7578 => x"41",
          7579 => x"3d",
          7580 => x"00",
          7581 => x"50",
          7582 => x"79",
          7583 => x"41",
          7584 => x"3d",
          7585 => x"00",
          7586 => x"74",
          7587 => x"72",
          7588 => x"73",
          7589 => x"3d",
          7590 => x"00",
          7591 => x"00",
          7592 => x"50",
          7593 => x"20",
          7594 => x"20",
          7595 => x"3d",
          7596 => x"00",
          7597 => x"79",
          7598 => x"6f",
          7599 => x"20",
          7600 => x"3d",
          7601 => x"64",
          7602 => x"20",
          7603 => x"6f",
          7604 => x"4d",
          7605 => x"46",
          7606 => x"2e",
          7607 => x"0a",
          7608 => x"44",
          7609 => x"63",
          7610 => x"20",
          7611 => x"3d",
          7612 => x"64",
          7613 => x"20",
          7614 => x"20",
          7615 => x"20",
          7616 => x"00",
          7617 => x"42",
          7618 => x"20",
          7619 => x"4f",
          7620 => x"00",
          7621 => x"4e",
          7622 => x"20",
          7623 => x"6c",
          7624 => x"2e",
          7625 => x"49",
          7626 => x"20",
          7627 => x"20",
          7628 => x"2e",
          7629 => x"44",
          7630 => x"20",
          7631 => x"73",
          7632 => x"2e",
          7633 => x"41",
          7634 => x"20",
          7635 => x"30",
          7636 => x"20",
          7637 => x"20",
          7638 => x"38",
          7639 => x"2e",
          7640 => x"4e",
          7641 => x"20",
          7642 => x"30",
          7643 => x"20",
          7644 => x"20",
          7645 => x"38",
          7646 => x"2e",
          7647 => x"42",
          7648 => x"20",
          7649 => x"30",
          7650 => x"28",
          7651 => x"43",
          7652 => x"29",
          7653 => x"77",
          7654 => x"00",
          7655 => x"00",
          7656 => x"6d",
          7657 => x"00",
          7658 => x"00",
          7659 => x"00",
          7660 => x"00",
          7661 => x"00",
          7662 => x"00",
          7663 => x"00",
          7664 => x"00",
          7665 => x"00",
          7666 => x"00",
          7667 => x"00",
          7668 => x"00",
          7669 => x"00",
          7670 => x"00",
          7671 => x"00",
          7672 => x"00",
          7673 => x"00",
          7674 => x"00",
          7675 => x"00",
          7676 => x"00",
          7677 => x"00",
          7678 => x"00",
          7679 => x"00",
          7680 => x"00",
          7681 => x"00",
          7682 => x"00",
          7683 => x"00",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"00",
          7690 => x"00",
          7691 => x"5b",
          7692 => x"5b",
          7693 => x"5b",
          7694 => x"5b",
          7695 => x"5b",
          7696 => x"5b",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"61",
          7703 => x"65",
          7704 => x"65",
          7705 => x"79",
          7706 => x"64",
          7707 => x"67",
          7708 => x"72",
          7709 => x"00",
          7710 => x"30",
          7711 => x"0a",
          7712 => x"64",
          7713 => x"65",
          7714 => x"69",
          7715 => x"69",
          7716 => x"4f",
          7717 => x"25",
          7718 => x"5b",
          7719 => x"5b",
          7720 => x"5b",
          7721 => x"5b",
          7722 => x"5b",
          7723 => x"5b",
          7724 => x"5b",
          7725 => x"5b",
          7726 => x"5b",
          7727 => x"5b",
          7728 => x"5b",
          7729 => x"5b",
          7730 => x"5b",
          7731 => x"5b",
          7732 => x"5b",
          7733 => x"5b",
          7734 => x"00",
          7735 => x"00",
          7736 => x"25",
          7737 => x"2c",
          7738 => x"30",
          7739 => x"3a",
          7740 => x"64",
          7741 => x"25",
          7742 => x"64",
          7743 => x"00",
          7744 => x"00",
          7745 => x"3b",
          7746 => x"65",
          7747 => x"72",
          7748 => x"70",
          7749 => x"30",
          7750 => x"77",
          7751 => x"30",
          7752 => x"64",
          7753 => x"00",
          7754 => x"73",
          7755 => x"65",
          7756 => x"44",
          7757 => x"3f",
          7758 => x"2c",
          7759 => x"41",
          7760 => x"00",
          7761 => x"44",
          7762 => x"4f",
          7763 => x"20",
          7764 => x"20",
          7765 => x"4d",
          7766 => x"54",
          7767 => x"00",
          7768 => x"00",
          7769 => x"03",
          7770 => x"16",
          7771 => x"9a",
          7772 => x"45",
          7773 => x"92",
          7774 => x"99",
          7775 => x"49",
          7776 => x"a9",
          7777 => x"b1",
          7778 => x"b9",
          7779 => x"c1",
          7780 => x"c9",
          7781 => x"d1",
          7782 => x"d9",
          7783 => x"e1",
          7784 => x"e9",
          7785 => x"f1",
          7786 => x"f9",
          7787 => x"2e",
          7788 => x"22",
          7789 => x"00",
          7790 => x"10",
          7791 => x"00",
          7792 => x"04",
          7793 => x"00",
          7794 => x"e9",
          7795 => x"e5",
          7796 => x"e8",
          7797 => x"c4",
          7798 => x"c6",
          7799 => x"fb",
          7800 => x"dc",
          7801 => x"a7",
          7802 => x"f3",
          7803 => x"aa",
          7804 => x"ac",
          7805 => x"ab",
          7806 => x"93",
          7807 => x"62",
          7808 => x"51",
          7809 => x"5b",
          7810 => x"2c",
          7811 => x"5e",
          7812 => x"69",
          7813 => x"6c",
          7814 => x"65",
          7815 => x"53",
          7816 => x"0c",
          7817 => x"90",
          7818 => x"93",
          7819 => x"b5",
          7820 => x"a9",
          7821 => x"b5",
          7822 => x"65",
          7823 => x"f7",
          7824 => x"b7",
          7825 => x"a0",
          7826 => x"e0",
          7827 => x"ff",
          7828 => x"30",
          7829 => x"10",
          7830 => x"06",
          7831 => x"81",
          7832 => x"84",
          7833 => x"89",
          7834 => x"8d",
          7835 => x"91",
          7836 => x"f6",
          7837 => x"98",
          7838 => x"9d",
          7839 => x"a0",
          7840 => x"a4",
          7841 => x"a9",
          7842 => x"ac",
          7843 => x"b1",
          7844 => x"b5",
          7845 => x"b8",
          7846 => x"bc",
          7847 => x"c1",
          7848 => x"c5",
          7849 => x"c7",
          7850 => x"cd",
          7851 => x"8e",
          7852 => x"03",
          7853 => x"f8",
          7854 => x"3a",
          7855 => x"3b",
          7856 => x"40",
          7857 => x"0a",
          7858 => x"86",
          7859 => x"58",
          7860 => x"5c",
          7861 => x"93",
          7862 => x"64",
          7863 => x"97",
          7864 => x"6c",
          7865 => x"70",
          7866 => x"74",
          7867 => x"78",
          7868 => x"7c",
          7869 => x"a6",
          7870 => x"84",
          7871 => x"ae",
          7872 => x"45",
          7873 => x"90",
          7874 => x"03",
          7875 => x"ac",
          7876 => x"89",
          7877 => x"c2",
          7878 => x"c4",
          7879 => x"8c",
          7880 => x"18",
          7881 => x"f3",
          7882 => x"f7",
          7883 => x"fa",
          7884 => x"10",
          7885 => x"36",
          7886 => x"01",
          7887 => x"61",
          7888 => x"7d",
          7889 => x"96",
          7890 => x"08",
          7891 => x"08",
          7892 => x"06",
          7893 => x"52",
          7894 => x"56",
          7895 => x"70",
          7896 => x"c8",
          7897 => x"da",
          7898 => x"ea",
          7899 => x"80",
          7900 => x"a0",
          7901 => x"b8",
          7902 => x"cc",
          7903 => x"02",
          7904 => x"01",
          7905 => x"fc",
          7906 => x"70",
          7907 => x"83",
          7908 => x"2f",
          7909 => x"06",
          7910 => x"64",
          7911 => x"1a",
          7912 => x"00",
          7913 => x"00",
          7914 => x"00",
          7915 => x"00",
          7916 => x"00",
          7917 => x"00",
          7918 => x"00",
          7919 => x"00",
          7920 => x"00",
          7921 => x"00",
          7922 => x"00",
          7923 => x"00",
          7924 => x"00",
          7925 => x"00",
          7926 => x"00",
          7927 => x"00",
          7928 => x"00",
          7929 => x"00",
          7930 => x"00",
          7931 => x"00",
          7932 => x"00",
          7933 => x"00",
          7934 => x"00",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"00",
          7963 => x"00",
          7964 => x"00",
          7965 => x"00",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"81",
          7973 => x"7f",
          7974 => x"00",
          7975 => x"00",
          7976 => x"f5",
          7977 => x"00",
          7978 => x"01",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"00",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"fc",
          7996 => x"7a",
          7997 => x"72",
          7998 => x"6a",
          7999 => x"62",
          8000 => x"32",
          8001 => x"f3",
          8002 => x"7f",
          8003 => x"f0",
          8004 => x"81",
          8005 => x"fc",
          8006 => x"5a",
          8007 => x"52",
          8008 => x"4a",
          8009 => x"42",
          8010 => x"32",
          8011 => x"f3",
          8012 => x"7f",
          8013 => x"f0",
          8014 => x"81",
          8015 => x"fc",
          8016 => x"5a",
          8017 => x"52",
          8018 => x"4a",
          8019 => x"42",
          8020 => x"22",
          8021 => x"7e",
          8022 => x"e2",
          8023 => x"f0",
          8024 => x"86",
          8025 => x"fe",
          8026 => x"1a",
          8027 => x"12",
          8028 => x"0a",
          8029 => x"02",
          8030 => x"f0",
          8031 => x"1e",
          8032 => x"f0",
          8033 => x"f0",
          8034 => x"81",
          8035 => x"f0",
          8036 => x"77",
          8037 => x"70",
          8038 => x"5d",
          8039 => x"6e",
          8040 => x"36",
          8041 => x"9f",
          8042 => x"c5",
          8043 => x"f0",
          8044 => x"81",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"cf",
          9082 => x"fd",
          9083 => x"c5",
          9084 => x"ee",
          9085 => x"65",
          9086 => x"2a",
          9087 => x"25",
          9088 => x"2b",
          9089 => x"05",
          9090 => x"0d",
          9091 => x"15",
          9092 => x"54",
          9093 => x"85",
          9094 => x"8d",
          9095 => x"95",
          9096 => x"40",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"04",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"00",
             3 => x"00",
             4 => x"88",
             5 => x"08",
             6 => x"04",
             7 => x"00",
             8 => x"71",
             9 => x"81",
            10 => x"ff",
            11 => x"00",
            12 => x"71",
            13 => x"83",
            14 => x"2b",
            15 => x"0b",
            16 => x"72",
            17 => x"09",
            18 => x"07",
            19 => x"00",
            20 => x"72",
            21 => x"51",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"09",
            26 => x"0a",
            27 => x"51",
            28 => x"72",
            29 => x"51",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"72",
            45 => x"0b",
            46 => x"00",
            47 => x"00",
            48 => x"72",
            49 => x"09",
            50 => x"06",
            51 => x"00",
            52 => x"71",
            53 => x"06",
            54 => x"0b",
            55 => x"51",
            56 => x"72",
            57 => x"81",
            58 => x"51",
            59 => x"00",
            60 => x"72",
            61 => x"81",
            62 => x"53",
            63 => x"00",
            64 => x"71",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"72",
            69 => x"04",
            70 => x"00",
            71 => x"00",
            72 => x"72",
            73 => x"07",
            74 => x"00",
            75 => x"00",
            76 => x"71",
            77 => x"81",
            78 => x"81",
            79 => x"00",
            80 => x"71",
            81 => x"f4",
            82 => x"06",
            83 => x"00",
            84 => x"88",
            85 => x"0b",
            86 => x"88",
            87 => x"0c",
            88 => x"88",
            89 => x"0b",
            90 => x"88",
            91 => x"0c",
            92 => x"72",
            93 => x"81",
            94 => x"73",
            95 => x"07",
            96 => x"72",
            97 => x"09",
            98 => x"06",
            99 => x"06",
           100 => x"05",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"04",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"71",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"04",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"02",
           117 => x"04",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"02",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"0b",
           134 => x"96",
           135 => x"0b",
           136 => x"0b",
           137 => x"d6",
           138 => x"0b",
           139 => x"0b",
           140 => x"96",
           141 => x"0b",
           142 => x"0b",
           143 => x"d7",
           144 => x"0b",
           145 => x"0b",
           146 => x"9b",
           147 => x"0b",
           148 => x"0b",
           149 => x"df",
           150 => x"0b",
           151 => x"0b",
           152 => x"a3",
           153 => x"0b",
           154 => x"0b",
           155 => x"e7",
           156 => x"0b",
           157 => x"0b",
           158 => x"ab",
           159 => x"0b",
           160 => x"0b",
           161 => x"ef",
           162 => x"0b",
           163 => x"0b",
           164 => x"b3",
           165 => x"0b",
           166 => x"0b",
           167 => x"f7",
           168 => x"0b",
           169 => x"0b",
           170 => x"bb",
           171 => x"0b",
           172 => x"0b",
           173 => x"fe",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"04",
           193 => x"0c",
           194 => x"08",
           195 => x"d4",
           196 => x"08",
           197 => x"d4",
           198 => x"08",
           199 => x"d4",
           200 => x"08",
           201 => x"d4",
           202 => x"08",
           203 => x"d4",
           204 => x"08",
           205 => x"d4",
           206 => x"08",
           207 => x"d4",
           208 => x"08",
           209 => x"d4",
           210 => x"08",
           211 => x"d4",
           212 => x"08",
           213 => x"d4",
           214 => x"08",
           215 => x"d4",
           216 => x"08",
           217 => x"d4",
           218 => x"d4",
           219 => x"b9",
           220 => x"b9",
           221 => x"84",
           222 => x"84",
           223 => x"04",
           224 => x"2d",
           225 => x"90",
           226 => x"ae",
           227 => x"80",
           228 => x"e3",
           229 => x"c0",
           230 => x"82",
           231 => x"80",
           232 => x"0c",
           233 => x"08",
           234 => x"d4",
           235 => x"d4",
           236 => x"b9",
           237 => x"b9",
           238 => x"84",
           239 => x"84",
           240 => x"04",
           241 => x"2d",
           242 => x"90",
           243 => x"8b",
           244 => x"80",
           245 => x"f3",
           246 => x"c0",
           247 => x"83",
           248 => x"80",
           249 => x"0c",
           250 => x"08",
           251 => x"d4",
           252 => x"d4",
           253 => x"b9",
           254 => x"b9",
           255 => x"84",
           256 => x"84",
           257 => x"04",
           258 => x"2d",
           259 => x"90",
           260 => x"d0",
           261 => x"80",
           262 => x"e3",
           263 => x"c0",
           264 => x"82",
           265 => x"80",
           266 => x"0c",
           267 => x"08",
           268 => x"d4",
           269 => x"d4",
           270 => x"b9",
           271 => x"b9",
           272 => x"84",
           273 => x"84",
           274 => x"04",
           275 => x"2d",
           276 => x"90",
           277 => x"92",
           278 => x"80",
           279 => x"b9",
           280 => x"c0",
           281 => x"83",
           282 => x"80",
           283 => x"0c",
           284 => x"08",
           285 => x"d4",
           286 => x"d4",
           287 => x"b9",
           288 => x"b9",
           289 => x"84",
           290 => x"84",
           291 => x"04",
           292 => x"2d",
           293 => x"90",
           294 => x"a5",
           295 => x"80",
           296 => x"9a",
           297 => x"80",
           298 => x"db",
           299 => x"c0",
           300 => x"81",
           301 => x"80",
           302 => x"0c",
           303 => x"08",
           304 => x"d4",
           305 => x"d4",
           306 => x"04",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"53",
           311 => x"06",
           312 => x"05",
           313 => x"06",
           314 => x"72",
           315 => x"05",
           316 => x"53",
           317 => x"04",
           318 => x"27",
           319 => x"53",
           320 => x"8c",
           321 => x"fc",
           322 => x"05",
           323 => x"d5",
           324 => x"3d",
           325 => x"7c",
           326 => x"80",
           327 => x"80",
           328 => x"80",
           329 => x"32",
           330 => x"51",
           331 => x"b7",
           332 => x"51",
           333 => x"53",
           334 => x"38",
           335 => x"05",
           336 => x"70",
           337 => x"54",
           338 => x"80",
           339 => x"c8",
           340 => x"84",
           341 => x"f5",
           342 => x"05",
           343 => x"58",
           344 => x"8d",
           345 => x"19",
           346 => x"04",
           347 => x"53",
           348 => x"3d",
           349 => x"65",
           350 => x"0c",
           351 => x"32",
           352 => x"72",
           353 => x"38",
           354 => x"c5",
           355 => x"5c",
           356 => x"17",
           357 => x"76",
           358 => x"51",
           359 => x"2e",
           360 => x"32",
           361 => x"9e",
           362 => x"33",
           363 => x"08",
           364 => x"3d",
           365 => x"10",
           366 => x"2b",
           367 => x"0a",
           368 => x"52",
           369 => x"81",
           370 => x"ff",
           371 => x"76",
           372 => x"a5",
           373 => x"73",
           374 => x"58",
           375 => x"39",
           376 => x"7b",
           377 => x"8d",
           378 => x"54",
           379 => x"06",
           380 => x"53",
           381 => x"10",
           382 => x"08",
           383 => x"d8",
           384 => x"51",
           385 => x"5b",
           386 => x"80",
           387 => x"7f",
           388 => x"ff",
           389 => x"b9",
           390 => x"9a",
           391 => x"06",
           392 => x"56",
           393 => x"b9",
           394 => x"70",
           395 => x"51",
           396 => x"56",
           397 => x"84",
           398 => x"06",
           399 => x"77",
           400 => x"05",
           401 => x"2a",
           402 => x"2e",
           403 => x"f8",
           404 => x"8b",
           405 => x"80",
           406 => x"7a",
           407 => x"72",
           408 => x"70",
           409 => x"24",
           410 => x"06",
           411 => x"56",
           412 => x"2e",
           413 => x"2b",
           414 => x"56",
           415 => x"38",
           416 => x"85",
           417 => x"54",
           418 => x"81",
           419 => x"81",
           420 => x"88",
           421 => x"b2",
           422 => x"fc",
           423 => x"40",
           424 => x"52",
           425 => x"84",
           426 => x"70",
           427 => x"24",
           428 => x"80",
           429 => x"0a",
           430 => x"2c",
           431 => x"38",
           432 => x"78",
           433 => x"0a",
           434 => x"74",
           435 => x"70",
           436 => x"81",
           437 => x"d8",
           438 => x"38",
           439 => x"7d",
           440 => x"52",
           441 => x"a5",
           442 => x"81",
           443 => x"7a",
           444 => x"84",
           445 => x"70",
           446 => x"25",
           447 => x"86",
           448 => x"5b",
           449 => x"76",
           450 => x"80",
           451 => x"60",
           452 => x"ff",
           453 => x"fb",
           454 => x"fe",
           455 => x"98",
           456 => x"29",
           457 => x"5e",
           458 => x"87",
           459 => x"fe",
           460 => x"29",
           461 => x"5a",
           462 => x"38",
           463 => x"e2",
           464 => x"06",
           465 => x"fe",
           466 => x"05",
           467 => x"39",
           468 => x"5b",
           469 => x"ab",
           470 => x"57",
           471 => x"75",
           472 => x"78",
           473 => x"05",
           474 => x"e3",
           475 => x"56",
           476 => x"39",
           477 => x"53",
           478 => x"df",
           479 => x"84",
           480 => x"84",
           481 => x"89",
           482 => x"5b",
           483 => x"f9",
           484 => x"05",
           485 => x"41",
           486 => x"87",
           487 => x"ff",
           488 => x"54",
           489 => x"39",
           490 => x"5b",
           491 => x"7f",
           492 => x"06",
           493 => x"38",
           494 => x"c8",
           495 => x"31",
           496 => x"81",
           497 => x"f7",
           498 => x"84",
           499 => x"70",
           500 => x"25",
           501 => x"83",
           502 => x"51",
           503 => x"81",
           504 => x"51",
           505 => x"06",
           506 => x"fa",
           507 => x"31",
           508 => x"80",
           509 => x"90",
           510 => x"51",
           511 => x"73",
           512 => x"39",
           513 => x"e5",
           514 => x"2e",
           515 => x"74",
           516 => x"53",
           517 => x"82",
           518 => x"51",
           519 => x"52",
           520 => x"c8",
           521 => x"31",
           522 => x"7a",
           523 => x"bf",
           524 => x"fe",
           525 => x"75",
           526 => x"3d",
           527 => x"80",
           528 => x"33",
           529 => x"06",
           530 => x"72",
           531 => x"38",
           532 => x"72",
           533 => x"08",
           534 => x"72",
           535 => x"83",
           536 => x"56",
           537 => x"84",
           538 => x"d5",
           539 => x"52",
           540 => x"2d",
           541 => x"38",
           542 => x"c8",
           543 => x"0d",
           544 => x"16",
           545 => x"81",
           546 => x"72",
           547 => x"73",
           548 => x"77",
           549 => x"56",
           550 => x"0d",
           551 => x"53",
           552 => x"72",
           553 => x"84",
           554 => x"ff",
           555 => x"57",
           556 => x"0d",
           557 => x"85",
           558 => x"0d",
           559 => x"2a",
           560 => x"57",
           561 => x"2a",
           562 => x"38",
           563 => x"08",
           564 => x"76",
           565 => x"8c",
           566 => x"0c",
           567 => x"88",
           568 => x"ff",
           569 => x"2d",
           570 => x"38",
           571 => x"0c",
           572 => x"77",
           573 => x"70",
           574 => x"56",
           575 => x"2a",
           576 => x"82",
           577 => x"80",
           578 => x"53",
           579 => x"13",
           580 => x"8c",
           581 => x"73",
           582 => x"04",
           583 => x"17",
           584 => x"17",
           585 => x"0c",
           586 => x"16",
           587 => x"08",
           588 => x"ff",
           589 => x"07",
           590 => x"2e",
           591 => x"85",
           592 => x"c8",
           593 => x"07",
           594 => x"ec",
           595 => x"54",
           596 => x"33",
           597 => x"72",
           598 => x"72",
           599 => x"38",
           600 => x"0d",
           601 => x"7a",
           602 => x"9d",
           603 => x"80",
           604 => x"53",
           605 => x"ff",
           606 => x"b9",
           607 => x"12",
           608 => x"14",
           609 => x"53",
           610 => x"51",
           611 => x"ff",
           612 => x"ff",
           613 => x"fe",
           614 => x"70",
           615 => x"38",
           616 => x"c8",
           617 => x"3d",
           618 => x"72",
           619 => x"72",
           620 => x"38",
           621 => x"0d",
           622 => x"79",
           623 => x"93",
           624 => x"73",
           625 => x"51",
           626 => x"0c",
           627 => x"76",
           628 => x"2e",
           629 => x"05",
           630 => x"09",
           631 => x"71",
           632 => x"72",
           633 => x"c8",
           634 => x"2e",
           635 => x"72",
           636 => x"52",
           637 => x"72",
           638 => x"3d",
           639 => x"86",
           640 => x"79",
           641 => x"84",
           642 => x"81",
           643 => x"84",
           644 => x"08",
           645 => x"08",
           646 => x"75",
           647 => x"b1",
           648 => x"84",
           649 => x"fd",
           650 => x"55",
           651 => x"72",
           652 => x"80",
           653 => x"ff",
           654 => x"13",
           655 => x"b9",
           656 => x"3d",
           657 => x"54",
           658 => x"72",
           659 => x"51",
           660 => x"0c",
           661 => x"78",
           662 => x"2e",
           663 => x"84",
           664 => x"73",
           665 => x"e3",
           666 => x"53",
           667 => x"38",
           668 => x"38",
           669 => x"31",
           670 => x"80",
           671 => x"10",
           672 => x"07",
           673 => x"70",
           674 => x"31",
           675 => x"58",
           676 => x"76",
           677 => x"88",
           678 => x"70",
           679 => x"72",
           680 => x"71",
           681 => x"80",
           682 => x"2b",
           683 => x"81",
           684 => x"82",
           685 => x"55",
           686 => x"70",
           687 => x"31",
           688 => x"32",
           689 => x"31",
           690 => x"0c",
           691 => x"5a",
           692 => x"56",
           693 => x"3d",
           694 => x"70",
           695 => x"3f",
           696 => x"71",
           697 => x"3d",
           698 => x"58",
           699 => x"38",
           700 => x"c8",
           701 => x"2e",
           702 => x"72",
           703 => x"53",
           704 => x"53",
           705 => x"74",
           706 => x"2b",
           707 => x"76",
           708 => x"2a",
           709 => x"31",
           710 => x"7b",
           711 => x"5c",
           712 => x"74",
           713 => x"88",
           714 => x"9f",
           715 => x"7b",
           716 => x"73",
           717 => x"31",
           718 => x"b4",
           719 => x"75",
           720 => x"0d",
           721 => x"57",
           722 => x"33",
           723 => x"81",
           724 => x"0c",
           725 => x"f3",
           726 => x"73",
           727 => x"58",
           728 => x"38",
           729 => x"80",
           730 => x"38",
           731 => x"53",
           732 => x"53",
           733 => x"70",
           734 => x"27",
           735 => x"83",
           736 => x"70",
           737 => x"73",
           738 => x"2e",
           739 => x"0c",
           740 => x"8b",
           741 => x"79",
           742 => x"b0",
           743 => x"81",
           744 => x"55",
           745 => x"58",
           746 => x"56",
           747 => x"53",
           748 => x"fe",
           749 => x"8b",
           750 => x"70",
           751 => x"56",
           752 => x"c8",
           753 => x"0d",
           754 => x"0c",
           755 => x"73",
           756 => x"81",
           757 => x"55",
           758 => x"2e",
           759 => x"83",
           760 => x"89",
           761 => x"56",
           762 => x"e0",
           763 => x"81",
           764 => x"81",
           765 => x"8f",
           766 => x"54",
           767 => x"72",
           768 => x"29",
           769 => x"33",
           770 => x"be",
           771 => x"30",
           772 => x"84",
           773 => x"81",
           774 => x"56",
           775 => x"06",
           776 => x"0c",
           777 => x"2e",
           778 => x"2e",
           779 => x"c6",
           780 => x"58",
           781 => x"84",
           782 => x"82",
           783 => x"33",
           784 => x"80",
           785 => x"0d",
           786 => x"c8",
           787 => x"0c",
           788 => x"93",
           789 => x"be",
           790 => x"ce",
           791 => x"0d",
           792 => x"3f",
           793 => x"51",
           794 => x"83",
           795 => x"3d",
           796 => x"92",
           797 => x"84",
           798 => x"04",
           799 => x"83",
           800 => x"ee",
           801 => x"cf",
           802 => x"0d",
           803 => x"3f",
           804 => x"51",
           805 => x"83",
           806 => x"3d",
           807 => x"ba",
           808 => x"d4",
           809 => x"04",
           810 => x"83",
           811 => x"ee",
           812 => x"d1",
           813 => x"0d",
           814 => x"3f",
           815 => x"51",
           816 => x"83",
           817 => x"3d",
           818 => x"e2",
           819 => x"0d",
           820 => x"33",
           821 => x"7b",
           822 => x"78",
           823 => x"81",
           824 => x"06",
           825 => x"38",
           826 => x"52",
           827 => x"c8",
           828 => x"2e",
           829 => x"97",
           830 => x"25",
           831 => x"53",
           832 => x"38",
           833 => x"87",
           834 => x"78",
           835 => x"84",
           836 => x"53",
           837 => x"df",
           838 => x"3d",
           839 => x"c0",
           840 => x"59",
           841 => x"53",
           842 => x"3f",
           843 => x"c8",
           844 => x"80",
           845 => x"17",
           846 => x"74",
           847 => x"08",
           848 => x"b9",
           849 => x"78",
           850 => x"3f",
           851 => x"02",
           852 => x"ff",
           853 => x"fd",
           854 => x"38",
           855 => x"2e",
           856 => x"8a",
           857 => x"a8",
           858 => x"c8",
           859 => x"84",
           860 => x"8a",
           861 => x"61",
           862 => x"33",
           863 => x"5c",
           864 => x"82",
           865 => x"dd",
           866 => x"f7",
           867 => x"38",
           868 => x"a0",
           869 => x"72",
           870 => x"52",
           871 => x"81",
           872 => x"a0",
           873 => x"dc",
           874 => x"3f",
           875 => x"38",
           876 => x"55",
           877 => x"80",
           878 => x"53",
           879 => x"56",
           880 => x"fe",
           881 => x"ac",
           882 => x"81",
           883 => x"83",
           884 => x"18",
           885 => x"c3",
           886 => x"70",
           887 => x"81",
           888 => x"38",
           889 => x"b9",
           890 => x"8f",
           891 => x"dc",
           892 => x"08",
           893 => x"78",
           894 => x"39",
           895 => x"82",
           896 => x"a0",
           897 => x"fe",
           898 => x"27",
           899 => x"9c",
           900 => x"d5",
           901 => x"c5",
           902 => x"99",
           903 => x"3f",
           904 => x"54",
           905 => x"27",
           906 => x"7a",
           907 => x"d1",
           908 => x"84",
           909 => x"ea",
           910 => x"fd",
           911 => x"73",
           912 => x"fe",
           913 => x"b9",
           914 => x"59",
           915 => x"59",
           916 => x"fc",
           917 => x"80",
           918 => x"08",
           919 => x"32",
           920 => x"70",
           921 => x"55",
           922 => x"25",
           923 => x"3f",
           924 => x"98",
           925 => x"9b",
           926 => x"75",
           927 => x"58",
           928 => x"fd",
           929 => x"0c",
           930 => x"87",
           931 => x"3f",
           932 => x"c0",
           933 => x"fc",
           934 => x"51",
           935 => x"2a",
           936 => x"89",
           937 => x"51",
           938 => x"2a",
           939 => x"ad",
           940 => x"51",
           941 => x"2a",
           942 => x"d2",
           943 => x"51",
           944 => x"81",
           945 => x"3f",
           946 => x"94",
           947 => x"3f",
           948 => x"3f",
           949 => x"fc",
           950 => x"3f",
           951 => x"2a",
           952 => x"38",
           953 => x"83",
           954 => x"51",
           955 => x"81",
           956 => x"9c",
           957 => x"3f",
           958 => x"80",
           959 => x"70",
           960 => x"fe",
           961 => x"9b",
           962 => x"ac",
           963 => x"85",
           964 => x"80",
           965 => x"81",
           966 => x"51",
           967 => x"3f",
           968 => x"52",
           969 => x"bd",
           970 => x"d4",
           971 => x"9a",
           972 => x"06",
           973 => x"38",
           974 => x"3f",
           975 => x"80",
           976 => x"70",
           977 => x"fd",
           978 => x"0d",
           979 => x"d0",
           980 => x"81",
           981 => x"81",
           982 => x"61",
           983 => x"51",
           984 => x"d5",
           985 => x"80",
           986 => x"ae",
           987 => x"70",
           988 => x"2e",
           989 => x"88",
           990 => x"82",
           991 => x"5a",
           992 => x"33",
           993 => x"8c",
           994 => x"7b",
           995 => x"9b",
           996 => x"ee",
           997 => x"ff",
           998 => x"c8",
           999 => x"5d",
          1000 => x"8b",
          1001 => x"2e",
          1002 => x"ff",
          1003 => x"38",
          1004 => x"fe",
          1005 => x"e9",
          1006 => x"84",
          1007 => x"38",
          1008 => x"ff",
          1009 => x"b9",
          1010 => x"7a",
          1011 => x"c8",
          1012 => x"c8",
          1013 => x"0b",
          1014 => x"8d",
          1015 => x"38",
          1016 => x"54",
          1017 => x"51",
          1018 => x"84",
          1019 => x"80",
          1020 => x"0a",
          1021 => x"b9",
          1022 => x"70",
          1023 => x"5b",
          1024 => x"83",
          1025 => x"78",
          1026 => x"81",
          1027 => x"38",
          1028 => x"5d",
          1029 => x"81",
          1030 => x"3f",
          1031 => x"7e",
          1032 => x"51",
          1033 => x"bc",
          1034 => x"79",
          1035 => x"98",
          1036 => x"cd",
          1037 => x"38",
          1038 => x"34",
          1039 => x"7e",
          1040 => x"c8",
          1041 => x"c8",
          1042 => x"83",
          1043 => x"5f",
          1044 => x"fc",
          1045 => x"51",
          1046 => x"0b",
          1047 => x"53",
          1048 => x"3f",
          1049 => x"38",
          1050 => x"1b",
          1051 => x"80",
          1052 => x"05",
          1053 => x"d5",
          1054 => x"60",
          1055 => x"82",
          1056 => x"61",
          1057 => x"81",
          1058 => x"ae",
          1059 => x"3f",
          1060 => x"90",
          1061 => x"83",
          1062 => x"94",
          1063 => x"93",
          1064 => x"39",
          1065 => x"52",
          1066 => x"39",
          1067 => x"83",
          1068 => x"59",
          1069 => x"8a",
          1070 => x"b8",
          1071 => x"05",
          1072 => x"08",
          1073 => x"83",
          1074 => x"5a",
          1075 => x"2e",
          1076 => x"52",
          1077 => x"fa",
          1078 => x"53",
          1079 => x"84",
          1080 => x"38",
          1081 => x"bf",
          1082 => x"fe",
          1083 => x"e9",
          1084 => x"2e",
          1085 => x"11",
          1086 => x"3f",
          1087 => x"64",
          1088 => x"d7",
          1089 => x"a8",
          1090 => x"d0",
          1091 => x"78",
          1092 => x"26",
          1093 => x"46",
          1094 => x"11",
          1095 => x"3f",
          1096 => x"fe",
          1097 => x"ff",
          1098 => x"b9",
          1099 => x"78",
          1100 => x"51",
          1101 => x"53",
          1102 => x"3f",
          1103 => x"2e",
          1104 => x"ca",
          1105 => x"cf",
          1106 => x"ff",
          1107 => x"b9",
          1108 => x"b8",
          1109 => x"05",
          1110 => x"08",
          1111 => x"fe",
          1112 => x"e9",
          1113 => x"2e",
          1114 => x"ce",
          1115 => x"7c",
          1116 => x"7a",
          1117 => x"95",
          1118 => x"53",
          1119 => x"8f",
          1120 => x"81",
          1121 => x"ff",
          1122 => x"e8",
          1123 => x"2e",
          1124 => x"11",
          1125 => x"3f",
          1126 => x"8e",
          1127 => x"ff",
          1128 => x"b9",
          1129 => x"83",
          1130 => x"5a",
          1131 => x"5c",
          1132 => x"34",
          1133 => x"3d",
          1134 => x"51",
          1135 => x"80",
          1136 => x"fc",
          1137 => x"fd",
          1138 => x"68",
          1139 => x"51",
          1140 => x"53",
          1141 => x"3f",
          1142 => x"2e",
          1143 => x"97",
          1144 => x"68",
          1145 => x"34",
          1146 => x"fc",
          1147 => x"ad",
          1148 => x"f5",
          1149 => x"05",
          1150 => x"b8",
          1151 => x"05",
          1152 => x"08",
          1153 => x"3d",
          1154 => x"51",
          1155 => x"80",
          1156 => x"fc",
          1157 => x"dd",
          1158 => x"f5",
          1159 => x"53",
          1160 => x"84",
          1161 => x"c8",
          1162 => x"b7",
          1163 => x"27",
          1164 => x"84",
          1165 => x"38",
          1166 => x"39",
          1167 => x"b1",
          1168 => x"ff",
          1169 => x"81",
          1170 => x"51",
          1171 => x"80",
          1172 => x"08",
          1173 => x"b8",
          1174 => x"05",
          1175 => x"08",
          1176 => x"79",
          1177 => x"84",
          1178 => x"53",
          1179 => x"84",
          1180 => x"cc",
          1181 => x"38",
          1182 => x"fe",
          1183 => x"e5",
          1184 => x"2e",
          1185 => x"88",
          1186 => x"32",
          1187 => x"7e",
          1188 => x"88",
          1189 => x"46",
          1190 => x"80",
          1191 => x"68",
          1192 => x"51",
          1193 => x"64",
          1194 => x"b8",
          1195 => x"05",
          1196 => x"08",
          1197 => x"71",
          1198 => x"3d",
          1199 => x"51",
          1200 => x"c6",
          1201 => x"80",
          1202 => x"40",
          1203 => x"11",
          1204 => x"3f",
          1205 => x"96",
          1206 => x"22",
          1207 => x"45",
          1208 => x"80",
          1209 => x"c8",
          1210 => x"b8",
          1211 => x"05",
          1212 => x"08",
          1213 => x"02",
          1214 => x"81",
          1215 => x"fe",
          1216 => x"e1",
          1217 => x"2e",
          1218 => x"5d",
          1219 => x"e1",
          1220 => x"f3",
          1221 => x"54",
          1222 => x"51",
          1223 => x"52",
          1224 => x"39",
          1225 => x"f0",
          1226 => x"53",
          1227 => x"84",
          1228 => x"64",
          1229 => x"70",
          1230 => x"e7",
          1231 => x"80",
          1232 => x"08",
          1233 => x"33",
          1234 => x"f2",
          1235 => x"d8",
          1236 => x"f7",
          1237 => x"ca",
          1238 => x"f2",
          1239 => x"38",
          1240 => x"39",
          1241 => x"f9",
          1242 => x"78",
          1243 => x"08",
          1244 => x"33",
          1245 => x"f2",
          1246 => x"f2",
          1247 => x"38",
          1248 => x"39",
          1249 => x"2e",
          1250 => x"fb",
          1251 => x"7c",
          1252 => x"08",
          1253 => x"08",
          1254 => x"83",
          1255 => x"b5",
          1256 => x"b9",
          1257 => x"08",
          1258 => x"51",
          1259 => x"90",
          1260 => x"80",
          1261 => x"84",
          1262 => x"c0",
          1263 => x"84",
          1264 => x"84",
          1265 => x"57",
          1266 => x"da",
          1267 => x"07",
          1268 => x"c0",
          1269 => x"87",
          1270 => x"5c",
          1271 => x"05",
          1272 => x"a8",
          1273 => x"70",
          1274 => x"b7",
          1275 => x"3f",
          1276 => x"d2",
          1277 => x"9f",
          1278 => x"55",
          1279 => x"83",
          1280 => x"83",
          1281 => x"b2",
          1282 => x"3f",
          1283 => x"ef",
          1284 => x"98",
          1285 => x"80",
          1286 => x"56",
          1287 => x"2e",
          1288 => x"ff",
          1289 => x"81",
          1290 => x"70",
          1291 => x"a0",
          1292 => x"54",
          1293 => x"52",
          1294 => x"72",
          1295 => x"54",
          1296 => x"70",
          1297 => x"86",
          1298 => x"73",
          1299 => x"2e",
          1300 => x"70",
          1301 => x"76",
          1302 => x"88",
          1303 => x"34",
          1304 => x"b9",
          1305 => x"80",
          1306 => x"be",
          1307 => x"70",
          1308 => x"a2",
          1309 => x"81",
          1310 => x"81",
          1311 => x"dc",
          1312 => x"08",
          1313 => x"0c",
          1314 => x"05",
          1315 => x"b9",
          1316 => x"84",
          1317 => x"fc",
          1318 => x"05",
          1319 => x"81",
          1320 => x"54",
          1321 => x"38",
          1322 => x"97",
          1323 => x"54",
          1324 => x"38",
          1325 => x"bb",
          1326 => x"55",
          1327 => x"d9",
          1328 => x"73",
          1329 => x"0b",
          1330 => x"87",
          1331 => x"87",
          1332 => x"87",
          1333 => x"87",
          1334 => x"87",
          1335 => x"87",
          1336 => x"98",
          1337 => x"0c",
          1338 => x"80",
          1339 => x"3d",
          1340 => x"87",
          1341 => x"87",
          1342 => x"23",
          1343 => x"82",
          1344 => x"5a",
          1345 => x"b0",
          1346 => x"c0",
          1347 => x"34",
          1348 => x"86",
          1349 => x"5c",
          1350 => x"a0",
          1351 => x"7d",
          1352 => x"7b",
          1353 => x"33",
          1354 => x"33",
          1355 => x"33",
          1356 => x"83",
          1357 => x"8f",
          1358 => x"93",
          1359 => x"38",
          1360 => x"b9",
          1361 => x"51",
          1362 => x"86",
          1363 => x"84",
          1364 => x"72",
          1365 => x"c8",
          1366 => x"52",
          1367 => x"38",
          1368 => x"b9",
          1369 => x"51",
          1370 => x"39",
          1371 => x"71",
          1372 => x"c3",
          1373 => x"70",
          1374 => x"eb",
          1375 => x"52",
          1376 => x"b9",
          1377 => x"3d",
          1378 => x"80",
          1379 => x"55",
          1380 => x"c0",
          1381 => x"81",
          1382 => x"8c",
          1383 => x"51",
          1384 => x"81",
          1385 => x"71",
          1386 => x"38",
          1387 => x"94",
          1388 => x"87",
          1389 => x"74",
          1390 => x"04",
          1391 => x"51",
          1392 => x"06",
          1393 => x"93",
          1394 => x"c0",
          1395 => x"96",
          1396 => x"70",
          1397 => x"02",
          1398 => x"2a",
          1399 => x"34",
          1400 => x"78",
          1401 => x"57",
          1402 => x"15",
          1403 => x"06",
          1404 => x"ff",
          1405 => x"96",
          1406 => x"70",
          1407 => x"70",
          1408 => x"72",
          1409 => x"2e",
          1410 => x"52",
          1411 => x"51",
          1412 => x"2e",
          1413 => x"73",
          1414 => x"57",
          1415 => x"c8",
          1416 => x"2a",
          1417 => x"38",
          1418 => x"80",
          1419 => x"06",
          1420 => x"87",
          1421 => x"70",
          1422 => x"38",
          1423 => x"9e",
          1424 => x"52",
          1425 => x"87",
          1426 => x"0c",
          1427 => x"88",
          1428 => x"f2",
          1429 => x"83",
          1430 => x"08",
          1431 => x"a0",
          1432 => x"9e",
          1433 => x"c0",
          1434 => x"87",
          1435 => x"0c",
          1436 => x"a8",
          1437 => x"f2",
          1438 => x"83",
          1439 => x"08",
          1440 => x"80",
          1441 => x"87",
          1442 => x"0c",
          1443 => x"c0",
          1444 => x"f2",
          1445 => x"34",
          1446 => x"70",
          1447 => x"70",
          1448 => x"34",
          1449 => x"70",
          1450 => x"70",
          1451 => x"83",
          1452 => x"9e",
          1453 => x"51",
          1454 => x"81",
          1455 => x"0b",
          1456 => x"80",
          1457 => x"2e",
          1458 => x"cc",
          1459 => x"08",
          1460 => x"52",
          1461 => x"71",
          1462 => x"c0",
          1463 => x"06",
          1464 => x"38",
          1465 => x"80",
          1466 => x"84",
          1467 => x"80",
          1468 => x"f2",
          1469 => x"90",
          1470 => x"52",
          1471 => x"52",
          1472 => x"87",
          1473 => x"80",
          1474 => x"83",
          1475 => x"34",
          1476 => x"70",
          1477 => x"70",
          1478 => x"83",
          1479 => x"9e",
          1480 => x"52",
          1481 => x"52",
          1482 => x"9e",
          1483 => x"2a",
          1484 => x"80",
          1485 => x"84",
          1486 => x"2e",
          1487 => x"d5",
          1488 => x"f0",
          1489 => x"83",
          1490 => x"9e",
          1491 => x"52",
          1492 => x"71",
          1493 => x"90",
          1494 => x"d8",
          1495 => x"fd",
          1496 => x"84",
          1497 => x"c8",
          1498 => x"d9",
          1499 => x"ca",
          1500 => x"f2",
          1501 => x"83",
          1502 => x"38",
          1503 => x"f4",
          1504 => x"84",
          1505 => x"75",
          1506 => x"54",
          1507 => x"33",
          1508 => x"c9",
          1509 => x"f2",
          1510 => x"83",
          1511 => x"38",
          1512 => x"e9",
          1513 => x"81",
          1514 => x"a2",
          1515 => x"d9",
          1516 => x"f2",
          1517 => x"ff",
          1518 => x"52",
          1519 => x"3f",
          1520 => x"83",
          1521 => x"51",
          1522 => x"08",
          1523 => x"ca",
          1524 => x"84",
          1525 => x"84",
          1526 => x"51",
          1527 => x"33",
          1528 => x"33",
          1529 => x"04",
          1530 => x"c0",
          1531 => x"b9",
          1532 => x"71",
          1533 => x"52",
          1534 => x"3f",
          1535 => x"08",
          1536 => x"c9",
          1537 => x"84",
          1538 => x"84",
          1539 => x"51",
          1540 => x"33",
          1541 => x"ff",
          1542 => x"c2",
          1543 => x"3f",
          1544 => x"bc",
          1545 => x"b0",
          1546 => x"b3",
          1547 => x"83",
          1548 => x"83",
          1549 => x"f2",
          1550 => x"ff",
          1551 => x"56",
          1552 => x"a4",
          1553 => x"c0",
          1554 => x"b9",
          1555 => x"ff",
          1556 => x"55",
          1557 => x"cc",
          1558 => x"c2",
          1559 => x"80",
          1560 => x"83",
          1561 => x"83",
          1562 => x"fc",
          1563 => x"51",
          1564 => x"33",
          1565 => x"d7",
          1566 => x"82",
          1567 => x"80",
          1568 => x"f2",
          1569 => x"ff",
          1570 => x"56",
          1571 => x"39",
          1572 => x"c4",
          1573 => x"d5",
          1574 => x"38",
          1575 => x"83",
          1576 => x"83",
          1577 => x"fb",
          1578 => x"08",
          1579 => x"83",
          1580 => x"83",
          1581 => x"fb",
          1582 => x"08",
          1583 => x"83",
          1584 => x"83",
          1585 => x"fa",
          1586 => x"08",
          1587 => x"83",
          1588 => x"83",
          1589 => x"fa",
          1590 => x"08",
          1591 => x"83",
          1592 => x"83",
          1593 => x"fa",
          1594 => x"08",
          1595 => x"83",
          1596 => x"83",
          1597 => x"f9",
          1598 => x"51",
          1599 => x"51",
          1600 => x"33",
          1601 => x"c4",
          1602 => x"33",
          1603 => x"10",
          1604 => x"08",
          1605 => x"df",
          1606 => x"ac",
          1607 => x"0d",
          1608 => x"c7",
          1609 => x"bc",
          1610 => x"0d",
          1611 => x"af",
          1612 => x"cc",
          1613 => x"0d",
          1614 => x"0b",
          1615 => x"f2",
          1616 => x"04",
          1617 => x"3d",
          1618 => x"80",
          1619 => x"88",
          1620 => x"ed",
          1621 => x"f3",
          1622 => x"76",
          1623 => x"c8",
          1624 => x"c0",
          1625 => x"17",
          1626 => x"08",
          1627 => x"ff",
          1628 => x"34",
          1629 => x"9f",
          1630 => x"85",
          1631 => x"b4",
          1632 => x"87",
          1633 => x"38",
          1634 => x"b9",
          1635 => x"e1",
          1636 => x"76",
          1637 => x"52",
          1638 => x"ff",
          1639 => x"84",
          1640 => x"83",
          1641 => x"80",
          1642 => x"0d",
          1643 => x"ad",
          1644 => x"57",
          1645 => x"91",
          1646 => x"75",
          1647 => x"70",
          1648 => x"84",
          1649 => x"08",
          1650 => x"08",
          1651 => x"81",
          1652 => x"99",
          1653 => x"57",
          1654 => x"54",
          1655 => x"0d",
          1656 => x"84",
          1657 => x"bd",
          1658 => x"d1",
          1659 => x"51",
          1660 => x"81",
          1661 => x"38",
          1662 => x"54",
          1663 => x"b6",
          1664 => x"76",
          1665 => x"5b",
          1666 => x"09",
          1667 => x"26",
          1668 => x"56",
          1669 => x"08",
          1670 => x"82",
          1671 => x"80",
          1672 => x"80",
          1673 => x"3f",
          1674 => x"38",
          1675 => x"b9",
          1676 => x"c8",
          1677 => x"08",
          1678 => x"77",
          1679 => x"83",
          1680 => x"3f",
          1681 => x"b2",
          1682 => x"aa",
          1683 => x"3d",
          1684 => x"5a",
          1685 => x"83",
          1686 => x"56",
          1687 => x"b0",
          1688 => x"cb",
          1689 => x"81",
          1690 => x"a0",
          1691 => x"93",
          1692 => x"eb",
          1693 => x"2b",
          1694 => x"2e",
          1695 => x"d1",
          1696 => x"2c",
          1697 => x"70",
          1698 => x"10",
          1699 => x"15",
          1700 => x"52",
          1701 => x"79",
          1702 => x"81",
          1703 => x"81",
          1704 => x"55",
          1705 => x"10",
          1706 => x"0b",
          1707 => x"77",
          1708 => x"15",
          1709 => x"75",
          1710 => x"c2",
          1711 => x"57",
          1712 => x"1b",
          1713 => x"d1",
          1714 => x"2c",
          1715 => x"83",
          1716 => x"5d",
          1717 => x"81",
          1718 => x"fe",
          1719 => x"38",
          1720 => x"0a",
          1721 => x"06",
          1722 => x"c0",
          1723 => x"51",
          1724 => x"33",
          1725 => x"83",
          1726 => x"42",
          1727 => x"76",
          1728 => x"39",
          1729 => x"38",
          1730 => x"39",
          1731 => x"84",
          1732 => x"34",
          1733 => x"55",
          1734 => x"10",
          1735 => x"08",
          1736 => x"0c",
          1737 => x"0b",
          1738 => x"d1",
          1739 => x"85",
          1740 => x"51",
          1741 => x"33",
          1742 => x"34",
          1743 => x"70",
          1744 => x"5b",
          1745 => x"38",
          1746 => x"58",
          1747 => x"70",
          1748 => x"fc",
          1749 => x"38",
          1750 => x"70",
          1751 => x"75",
          1752 => x"84",
          1753 => x"56",
          1754 => x"d5",
          1755 => x"95",
          1756 => x"51",
          1757 => x"08",
          1758 => x"84",
          1759 => x"84",
          1760 => x"55",
          1761 => x"ff",
          1762 => x"cd",
          1763 => x"08",
          1764 => x"10",
          1765 => x"57",
          1766 => x"56",
          1767 => x"51",
          1768 => x"08",
          1769 => x"08",
          1770 => x"52",
          1771 => x"d1",
          1772 => x"56",
          1773 => x"d5",
          1774 => x"fd",
          1775 => x"51",
          1776 => x"08",
          1777 => x"84",
          1778 => x"84",
          1779 => x"55",
          1780 => x"81",
          1781 => x"57",
          1782 => x"84",
          1783 => x"76",
          1784 => x"33",
          1785 => x"d1",
          1786 => x"d1",
          1787 => x"27",
          1788 => x"52",
          1789 => x"34",
          1790 => x"b2",
          1791 => x"81",
          1792 => x"57",
          1793 => x"f9",
          1794 => x"d1",
          1795 => x"f9",
          1796 => x"d1",
          1797 => x"2c",
          1798 => x"60",
          1799 => x"ac",
          1800 => x"3f",
          1801 => x"70",
          1802 => x"57",
          1803 => x"38",
          1804 => x"ff",
          1805 => x"29",
          1806 => x"84",
          1807 => x"7b",
          1808 => x"08",
          1809 => x"74",
          1810 => x"05",
          1811 => x"5d",
          1812 => x"38",
          1813 => x"18",
          1814 => x"52",
          1815 => x"75",
          1816 => x"05",
          1817 => x"5b",
          1818 => x"38",
          1819 => x"34",
          1820 => x"51",
          1821 => x"0a",
          1822 => x"2c",
          1823 => x"78",
          1824 => x"39",
          1825 => x"2e",
          1826 => x"52",
          1827 => x"d1",
          1828 => x"d1",
          1829 => x"dd",
          1830 => x"5f",
          1831 => x"52",
          1832 => x"d1",
          1833 => x"84",
          1834 => x"77",
          1835 => x"57",
          1836 => x"f3",
          1837 => x"e0",
          1838 => x"8b",
          1839 => x"06",
          1840 => x"53",
          1841 => x"b9",
          1842 => x"33",
          1843 => x"70",
          1844 => x"38",
          1845 => x"2e",
          1846 => x"77",
          1847 => x"84",
          1848 => x"88",
          1849 => x"3d",
          1850 => x"74",
          1851 => x"08",
          1852 => x"84",
          1853 => x"af",
          1854 => x"88",
          1855 => x"8c",
          1856 => x"8c",
          1857 => x"cc",
          1858 => x"f7",
          1859 => x"80",
          1860 => x"39",
          1861 => x"34",
          1862 => x"2e",
          1863 => x"88",
          1864 => x"ac",
          1865 => x"3f",
          1866 => x"ff",
          1867 => x"ff",
          1868 => x"7c",
          1869 => x"83",
          1870 => x"80",
          1871 => x"84",
          1872 => x"0c",
          1873 => x"33",
          1874 => x"80",
          1875 => x"33",
          1876 => x"34",
          1877 => x"34",
          1878 => x"ff",
          1879 => x"70",
          1880 => x"88",
          1881 => x"24",
          1882 => x"52",
          1883 => x"d1",
          1884 => x"2c",
          1885 => x"56",
          1886 => x"d5",
          1887 => x"f5",
          1888 => x"80",
          1889 => x"88",
          1890 => x"f3",
          1891 => x"88",
          1892 => x"80",
          1893 => x"98",
          1894 => x"55",
          1895 => x"a5",
          1896 => x"77",
          1897 => x"33",
          1898 => x"80",
          1899 => x"98",
          1900 => x"5b",
          1901 => x"16",
          1902 => x"d5",
          1903 => x"ab",
          1904 => x"81",
          1905 => x"d1",
          1906 => x"24",
          1907 => x"d1",
          1908 => x"58",
          1909 => x"d1",
          1910 => x"38",
          1911 => x"41",
          1912 => x"5b",
          1913 => x"80",
          1914 => x"98",
          1915 => x"58",
          1916 => x"55",
          1917 => x"ff",
          1918 => x"7a",
          1919 => x"60",
          1920 => x"84",
          1921 => x"8c",
          1922 => x"ff",
          1923 => x"ff",
          1924 => x"24",
          1925 => x"98",
          1926 => x"59",
          1927 => x"d5",
          1928 => x"ad",
          1929 => x"80",
          1930 => x"88",
          1931 => x"f1",
          1932 => x"88",
          1933 => x"80",
          1934 => x"98",
          1935 => x"41",
          1936 => x"dd",
          1937 => x"80",
          1938 => x"ad",
          1939 => x"d1",
          1940 => x"ff",
          1941 => x"51",
          1942 => x"33",
          1943 => x"80",
          1944 => x"08",
          1945 => x"84",
          1946 => x"a9",
          1947 => x"88",
          1948 => x"8c",
          1949 => x"8c",
          1950 => x"39",
          1951 => x"b9",
          1952 => x"b9",
          1953 => x"f3",
          1954 => x"c3",
          1955 => x"16",
          1956 => x"3f",
          1957 => x"0a",
          1958 => x"33",
          1959 => x"38",
          1960 => x"70",
          1961 => x"58",
          1962 => x"38",
          1963 => x"80",
          1964 => x"57",
          1965 => x"38",
          1966 => x"80",
          1967 => x"b8",
          1968 => x"80",
          1969 => x"e7",
          1970 => x"80",
          1971 => x"b4",
          1972 => x"ee",
          1973 => x"3f",
          1974 => x"58",
          1975 => x"ff",
          1976 => x"3f",
          1977 => x"34",
          1978 => x"81",
          1979 => x"ab",
          1980 => x"33",
          1981 => x"74",
          1982 => x"ac",
          1983 => x"3f",
          1984 => x"ff",
          1985 => x"52",
          1986 => x"d1",
          1987 => x"d1",
          1988 => x"c7",
          1989 => x"d1",
          1990 => x"34",
          1991 => x"0d",
          1992 => x"84",
          1993 => x"84",
          1994 => x"05",
          1995 => x"91",
          1996 => x"84",
          1997 => x"58",
          1998 => x"93",
          1999 => x"51",
          2000 => x"08",
          2001 => x"84",
          2002 => x"a5",
          2003 => x"05",
          2004 => x"81",
          2005 => x"ff",
          2006 => x"84",
          2007 => x"81",
          2008 => x"7b",
          2009 => x"70",
          2010 => x"84",
          2011 => x"74",
          2012 => x"ac",
          2013 => x"3f",
          2014 => x"ff",
          2015 => x"52",
          2016 => x"d1",
          2017 => x"d1",
          2018 => x"c7",
          2019 => x"83",
          2020 => x"fc",
          2021 => x"70",
          2022 => x"3f",
          2023 => x"f3",
          2024 => x"e0",
          2025 => x"80",
          2026 => x"52",
          2027 => x"f3",
          2028 => x"06",
          2029 => x"38",
          2030 => x"39",
          2031 => x"53",
          2032 => x"3f",
          2033 => x"82",
          2034 => x"51",
          2035 => x"d1",
          2036 => x"34",
          2037 => x"0d",
          2038 => x"c8",
          2039 => x"b9",
          2040 => x"c8",
          2041 => x"b4",
          2042 => x"82",
          2043 => x"5a",
          2044 => x"81",
          2045 => x"08",
          2046 => x"c8",
          2047 => x"08",
          2048 => x"08",
          2049 => x"77",
          2050 => x"b8",
          2051 => x"05",
          2052 => x"80",
          2053 => x"06",
          2054 => x"53",
          2055 => x"b9",
          2056 => x"33",
          2057 => x"70",
          2058 => x"81",
          2059 => x"93",
          2060 => x"ff",
          2061 => x"77",
          2062 => x"53",
          2063 => x"3f",
          2064 => x"81",
          2065 => x"80",
          2066 => x"34",
          2067 => x"f8",
          2068 => x"2b",
          2069 => x"81",
          2070 => x"d9",
          2071 => x"0c",
          2072 => x"83",
          2073 => x"41",
          2074 => x"9e",
          2075 => x"f7",
          2076 => x"c0",
          2077 => x"8a",
          2078 => x"39",
          2079 => x"33",
          2080 => x"5b",
          2081 => x"72",
          2082 => x"25",
          2083 => x"a8",
          2084 => x"a7",
          2085 => x"9f",
          2086 => x"75",
          2087 => x"f9",
          2088 => x"f8",
          2089 => x"2b",
          2090 => x"7a",
          2091 => x"27",
          2092 => x"56",
          2093 => x"0c",
          2094 => x"27",
          2095 => x"98",
          2096 => x"55",
          2097 => x"74",
          2098 => x"53",
          2099 => x"86",
          2100 => x"33",
          2101 => x"33",
          2102 => x"41",
          2103 => x"0b",
          2104 => x"06",
          2105 => x"06",
          2106 => x"ff",
          2107 => x"58",
          2108 => x"87",
          2109 => x"79",
          2110 => x"7c",
          2111 => x"06",
          2112 => x"14",
          2113 => x"74",
          2114 => x"74",
          2115 => x"59",
          2116 => x"2e",
          2117 => x"72",
          2118 => x"70",
          2119 => x"33",
          2120 => x"39",
          2121 => x"b0",
          2122 => x"81",
          2123 => x"81",
          2124 => x"74",
          2125 => x"5e",
          2126 => x"73",
          2127 => x"71",
          2128 => x"80",
          2129 => x"f8",
          2130 => x"34",
          2131 => x"71",
          2132 => x"71",
          2133 => x"76",
          2134 => x"39",
          2135 => x"33",
          2136 => x"11",
          2137 => x"11",
          2138 => x"5b",
          2139 => x"70",
          2140 => x"ff",
          2141 => x"ff",
          2142 => x"ff",
          2143 => x"5e",
          2144 => x"57",
          2145 => x"31",
          2146 => x"7d",
          2147 => x"71",
          2148 => x"62",
          2149 => x"5f",
          2150 => x"85",
          2151 => x"31",
          2152 => x"fd",
          2153 => x"fd",
          2154 => x"31",
          2155 => x"3d",
          2156 => x"8a",
          2157 => x"34",
          2158 => x"55",
          2159 => x"34",
          2160 => x"34",
          2161 => x"54",
          2162 => x"80",
          2163 => x"d8",
          2164 => x"54",
          2165 => x"f8",
          2166 => x"72",
          2167 => x"06",
          2168 => x"34",
          2169 => x"06",
          2170 => x"81",
          2171 => x"88",
          2172 => x"0b",
          2173 => x"b9",
          2174 => x"b7",
          2175 => x"f7",
          2176 => x"84",
          2177 => x"33",
          2178 => x"26",
          2179 => x"83",
          2180 => x"72",
          2181 => x"11",
          2182 => x"59",
          2183 => x"ff",
          2184 => x"58",
          2185 => x"83",
          2186 => x"83",
          2187 => x"76",
          2188 => x"ff",
          2189 => x"82",
          2190 => x"f8",
          2191 => x"83",
          2192 => x"5c",
          2193 => x"38",
          2194 => x"54",
          2195 => x"ac",
          2196 => x"55",
          2197 => x"34",
          2198 => x"70",
          2199 => x"84",
          2200 => x"9f",
          2201 => x"33",
          2202 => x"0b",
          2203 => x"81",
          2204 => x"9f",
          2205 => x"33",
          2206 => x"23",
          2207 => x"83",
          2208 => x"26",
          2209 => x"05",
          2210 => x"58",
          2211 => x"80",
          2212 => x"ff",
          2213 => x"29",
          2214 => x"27",
          2215 => x"e0",
          2216 => x"13",
          2217 => x"73",
          2218 => x"81",
          2219 => x"bc",
          2220 => x"29",
          2221 => x"26",
          2222 => x"c8",
          2223 => x"f8",
          2224 => x"83",
          2225 => x"5c",
          2226 => x"38",
          2227 => x"81",
          2228 => x"33",
          2229 => x"06",
          2230 => x"05",
          2231 => x"78",
          2232 => x"73",
          2233 => x"f4",
          2234 => x"31",
          2235 => x"16",
          2236 => x"34",
          2237 => x"8a",
          2238 => x"75",
          2239 => x"13",
          2240 => x"80",
          2241 => x"fe",
          2242 => x"59",
          2243 => x"84",
          2244 => x"fc",
          2245 => x"05",
          2246 => x"38",
          2247 => x"51",
          2248 => x"51",
          2249 => x"f8",
          2250 => x"0c",
          2251 => x"f8",
          2252 => x"81",
          2253 => x"e2",
          2254 => x"f8",
          2255 => x"86",
          2256 => x"70",
          2257 => x"72",
          2258 => x"f8",
          2259 => x"33",
          2260 => x"11",
          2261 => x"38",
          2262 => x"80",
          2263 => x"0d",
          2264 => x"31",
          2265 => x"54",
          2266 => x"34",
          2267 => x"3d",
          2268 => x"05",
          2269 => x"55",
          2270 => x"53",
          2271 => x"84",
          2272 => x"80",
          2273 => x"f8",
          2274 => x"56",
          2275 => x"81",
          2276 => x"fe",
          2277 => x"05",
          2278 => x"70",
          2279 => x"70",
          2280 => x"80",
          2281 => x"06",
          2282 => x"53",
          2283 => x"06",
          2284 => x"f4",
          2285 => x"83",
          2286 => x"81",
          2287 => x"f8",
          2288 => x"0c",
          2289 => x"33",
          2290 => x"f4",
          2291 => x"81",
          2292 => x"f8",
          2293 => x"83",
          2294 => x"c8",
          2295 => x"f4",
          2296 => x"70",
          2297 => x"83",
          2298 => x"83",
          2299 => x"f8",
          2300 => x"51",
          2301 => x"39",
          2302 => x"83",
          2303 => x"ff",
          2304 => x"f9",
          2305 => x"f4",
          2306 => x"33",
          2307 => x"f4",
          2308 => x"33",
          2309 => x"70",
          2310 => x"83",
          2311 => x"07",
          2312 => x"ba",
          2313 => x"06",
          2314 => x"f4",
          2315 => x"33",
          2316 => x"70",
          2317 => x"83",
          2318 => x"07",
          2319 => x"82",
          2320 => x"06",
          2321 => x"f2",
          2322 => x"06",
          2323 => x"34",
          2324 => x"bf",
          2325 => x"05",
          2326 => x"f7",
          2327 => x"be",
          2328 => x"78",
          2329 => x"24",
          2330 => x"38",
          2331 => x"84",
          2332 => x"34",
          2333 => x"f8",
          2334 => x"83",
          2335 => x"0b",
          2336 => x"b7",
          2337 => x"34",
          2338 => x"0b",
          2339 => x"b7",
          2340 => x"56",
          2341 => x"7c",
          2342 => x"ff",
          2343 => x"34",
          2344 => x"83",
          2345 => x"23",
          2346 => x"0d",
          2347 => x"81",
          2348 => x"83",
          2349 => x"f9",
          2350 => x"84",
          2351 => x"33",
          2352 => x"55",
          2353 => x"e3",
          2354 => x"0b",
          2355 => x"79",
          2356 => x"9c",
          2357 => x"f0",
          2358 => x"70",
          2359 => x"52",
          2360 => x"83",
          2361 => x"7d",
          2362 => x"b7",
          2363 => x"7b",
          2364 => x"f9",
          2365 => x"84",
          2366 => x"c0",
          2367 => x"a8",
          2368 => x"83",
          2369 => x"ff",
          2370 => x"52",
          2371 => x"3f",
          2372 => x"92",
          2373 => x"27",
          2374 => x"33",
          2375 => x"cf",
          2376 => x"5a",
          2377 => x"02",
          2378 => x"bc",
          2379 => x"f8",
          2380 => x"a0",
          2381 => x"51",
          2382 => x"83",
          2383 => x"52",
          2384 => x"2e",
          2385 => x"f9",
          2386 => x"75",
          2387 => x"2e",
          2388 => x"83",
          2389 => x"72",
          2390 => x"b7",
          2391 => x"14",
          2392 => x"f9",
          2393 => x"29",
          2394 => x"f8",
          2395 => x"73",
          2396 => x"f4",
          2397 => x"84",
          2398 => x"83",
          2399 => x"72",
          2400 => x"57",
          2401 => x"14",
          2402 => x"59",
          2403 => x"84",
          2404 => x"38",
          2405 => x"34",
          2406 => x"2e",
          2407 => x"76",
          2408 => x"84",
          2409 => x"75",
          2410 => x"80",
          2411 => x"06",
          2412 => x"f1",
          2413 => x"34",
          2414 => x"33",
          2415 => x"34",
          2416 => x"89",
          2417 => x"fd",
          2418 => x"06",
          2419 => x"38",
          2420 => x"81",
          2421 => x"83",
          2422 => x"74",
          2423 => x"75",
          2424 => x"0b",
          2425 => x"04",
          2426 => x"fd",
          2427 => x"81",
          2428 => x"83",
          2429 => x"34",
          2430 => x"83",
          2431 => x"55",
          2432 => x"73",
          2433 => x"a0",
          2434 => x"81",
          2435 => x"90",
          2436 => x"3f",
          2437 => x"80",
          2438 => x"57",
          2439 => x"75",
          2440 => x"2e",
          2441 => x"d1",
          2442 => x"78",
          2443 => x"bc",
          2444 => x"f9",
          2445 => x"5c",
          2446 => x"a0",
          2447 => x"83",
          2448 => x"72",
          2449 => x"78",
          2450 => x"f8",
          2451 => x"5a",
          2452 => x"b0",
          2453 => x"70",
          2454 => x"83",
          2455 => x"42",
          2456 => x"33",
          2457 => x"70",
          2458 => x"26",
          2459 => x"5a",
          2460 => x"75",
          2461 => x"b9",
          2462 => x"b7",
          2463 => x"81",
          2464 => x"38",
          2465 => x"80",
          2466 => x"bc",
          2467 => x"f9",
          2468 => x"40",
          2469 => x"a0",
          2470 => x"83",
          2471 => x"72",
          2472 => x"78",
          2473 => x"f8",
          2474 => x"83",
          2475 => x"1b",
          2476 => x"ff",
          2477 => x"f9",
          2478 => x"43",
          2479 => x"84",
          2480 => x"77",
          2481 => x"fe",
          2482 => x"80",
          2483 => x"0d",
          2484 => x"78",
          2485 => x"2e",
          2486 => x"0b",
          2487 => x"b9",
          2488 => x"9b",
          2489 => x"75",
          2490 => x"c8",
          2491 => x"b8",
          2492 => x"34",
          2493 => x"84",
          2494 => x"b9",
          2495 => x"9b",
          2496 => x"b8",
          2497 => x"f8",
          2498 => x"72",
          2499 => x"c4",
          2500 => x"34",
          2501 => x"33",
          2502 => x"12",
          2503 => x"fa",
          2504 => x"71",
          2505 => x"33",
          2506 => x"b7",
          2507 => x"f8",
          2508 => x"72",
          2509 => x"83",
          2510 => x"05",
          2511 => x"81",
          2512 => x"0b",
          2513 => x"84",
          2514 => x"70",
          2515 => x"73",
          2516 => x"05",
          2517 => x"72",
          2518 => x"06",
          2519 => x"5a",
          2520 => x"78",
          2521 => x"76",
          2522 => x"f8",
          2523 => x"84",
          2524 => x"c9",
          2525 => x"80",
          2526 => x"84",
          2527 => x"c8",
          2528 => x"f8",
          2529 => x"f9",
          2530 => x"f7",
          2531 => x"84",
          2532 => x"c8",
          2533 => x"ff",
          2534 => x"83",
          2535 => x"70",
          2536 => x"70",
          2537 => x"86",
          2538 => x"22",
          2539 => x"83",
          2540 => x"44",
          2541 => x"81",
          2542 => x"06",
          2543 => x"75",
          2544 => x"81",
          2545 => x"81",
          2546 => x"40",
          2547 => x"a0",
          2548 => x"83",
          2549 => x"72",
          2550 => x"a0",
          2551 => x"f8",
          2552 => x"5a",
          2553 => x"b0",
          2554 => x"70",
          2555 => x"83",
          2556 => x"43",
          2557 => x"33",
          2558 => x"1a",
          2559 => x"7b",
          2560 => x"33",
          2561 => x"58",
          2562 => x"f9",
          2563 => x"05",
          2564 => x"95",
          2565 => x"38",
          2566 => x"b8",
          2567 => x"ff",
          2568 => x"c8",
          2569 => x"05",
          2570 => x"f8",
          2571 => x"9f",
          2572 => x"9c",
          2573 => x"84",
          2574 => x"83",
          2575 => x"72",
          2576 => x"05",
          2577 => x"7b",
          2578 => x"83",
          2579 => x"59",
          2580 => x"38",
          2581 => x"81",
          2582 => x"72",
          2583 => x"e4",
          2584 => x"84",
          2585 => x"83",
          2586 => x"5e",
          2587 => x"fa",
          2588 => x"71",
          2589 => x"33",
          2590 => x"b7",
          2591 => x"f8",
          2592 => x"72",
          2593 => x"83",
          2594 => x"34",
          2595 => x"5b",
          2596 => x"84",
          2597 => x"38",
          2598 => x"34",
          2599 => x"59",
          2600 => x"f8",
          2601 => x"f8",
          2602 => x"81",
          2603 => x"72",
          2604 => x"5b",
          2605 => x"80",
          2606 => x"f8",
          2607 => x"71",
          2608 => x"0b",
          2609 => x"f8",
          2610 => x"83",
          2611 => x"1a",
          2612 => x"ff",
          2613 => x"f9",
          2614 => x"5a",
          2615 => x"98",
          2616 => x"81",
          2617 => x"fe",
          2618 => x"fe",
          2619 => x"0c",
          2620 => x"3d",
          2621 => x"59",
          2622 => x"83",
          2623 => x"58",
          2624 => x"0b",
          2625 => x"b9",
          2626 => x"f8",
          2627 => x"1b",
          2628 => x"84",
          2629 => x"5b",
          2630 => x"84",
          2631 => x"53",
          2632 => x"84",
          2633 => x"38",
          2634 => x"5a",
          2635 => x"83",
          2636 => x"22",
          2637 => x"cf",
          2638 => x"84",
          2639 => x"f8",
          2640 => x"f8",
          2641 => x"39",
          2642 => x"33",
          2643 => x"05",
          2644 => x"33",
          2645 => x"84",
          2646 => x"83",
          2647 => x"5a",
          2648 => x"18",
          2649 => x"29",
          2650 => x"60",
          2651 => x"b7",
          2652 => x"f8",
          2653 => x"72",
          2654 => x"83",
          2655 => x"34",
          2656 => x"58",
          2657 => x"b7",
          2658 => x"ff",
          2659 => x"80",
          2660 => x"bf",
          2661 => x"38",
          2662 => x"b4",
          2663 => x"3f",
          2664 => x"3d",
          2665 => x"f8",
          2666 => x"f8",
          2667 => x"76",
          2668 => x"83",
          2669 => x"83",
          2670 => x"83",
          2671 => x"ff",
          2672 => x"7a",
          2673 => x"9c",
          2674 => x"06",
          2675 => x"81",
          2676 => x"05",
          2677 => x"94",
          2678 => x"3f",
          2679 => x"b9",
          2680 => x"cc",
          2681 => x"24",
          2682 => x"ac",
          2683 => x"39",
          2684 => x"58",
          2685 => x"27",
          2686 => x"9c",
          2687 => x"b1",
          2688 => x"83",
          2689 => x"84",
          2690 => x"8f",
          2691 => x"b9",
          2692 => x"70",
          2693 => x"5e",
          2694 => x"e7",
          2695 => x"80",
          2696 => x"33",
          2697 => x"b7",
          2698 => x"27",
          2699 => x"34",
          2700 => x"f9",
          2701 => x"ff",
          2702 => x"a7",
          2703 => x"f8",
          2704 => x"f8",
          2705 => x"b7",
          2706 => x"76",
          2707 => x"75",
          2708 => x"84",
          2709 => x"8d",
          2710 => x"b9",
          2711 => x"70",
          2712 => x"42",
          2713 => x"cf",
          2714 => x"80",
          2715 => x"22",
          2716 => x"fc",
          2717 => x"f8",
          2718 => x"71",
          2719 => x"83",
          2720 => x"71",
          2721 => x"06",
          2722 => x"80",
          2723 => x"82",
          2724 => x"83",
          2725 => x"b8",
          2726 => x"e7",
          2727 => x"99",
          2728 => x"81",
          2729 => x"39",
          2730 => x"2e",
          2731 => x"83",
          2732 => x"b7",
          2733 => x"75",
          2734 => x"83",
          2735 => x"b8",
          2736 => x"c8",
          2737 => x"f8",
          2738 => x"33",
          2739 => x"25",
          2740 => x"f8",
          2741 => x"51",
          2742 => x"b8",
          2743 => x"8b",
          2744 => x"05",
          2745 => x"51",
          2746 => x"81",
          2747 => x"58",
          2748 => x"c9",
          2749 => x"38",
          2750 => x"26",
          2751 => x"81",
          2752 => x"97",
          2753 => x"77",
          2754 => x"33",
          2755 => x"b9",
          2756 => x"06",
          2757 => x"06",
          2758 => x"5c",
          2759 => x"5a",
          2760 => x"ff",
          2761 => x"27",
          2762 => x"f8",
          2763 => x"57",
          2764 => x"7a",
          2765 => x"af",
          2766 => x"80",
          2767 => x"33",
          2768 => x"7f",
          2769 => x"33",
          2770 => x"06",
          2771 => x"11",
          2772 => x"f6",
          2773 => x"70",
          2774 => x"33",
          2775 => x"81",
          2776 => x"ff",
          2777 => x"7c",
          2778 => x"33",
          2779 => x"ff",
          2780 => x"7c",
          2781 => x"57",
          2782 => x"b7",
          2783 => x"ee",
          2784 => x"f8",
          2785 => x"f6",
          2786 => x"26",
          2787 => x"7e",
          2788 => x"5e",
          2789 => x"5b",
          2790 => x"06",
          2791 => x"1d",
          2792 => x"f7",
          2793 => x"e0",
          2794 => x"1f",
          2795 => x"76",
          2796 => x"81",
          2797 => x"bc",
          2798 => x"29",
          2799 => x"27",
          2800 => x"5f",
          2801 => x"81",
          2802 => x"58",
          2803 => x"81",
          2804 => x"bb",
          2805 => x"5e",
          2806 => x"f6",
          2807 => x"75",
          2808 => x"84",
          2809 => x"f6",
          2810 => x"33",
          2811 => x"59",
          2812 => x"84",
          2813 => x"09",
          2814 => x"f9",
          2815 => x"f8",
          2816 => x"ff",
          2817 => x"33",
          2818 => x"7e",
          2819 => x"f5",
          2820 => x"27",
          2821 => x"10",
          2822 => x"86",
          2823 => x"5a",
          2824 => x"06",
          2825 => x"79",
          2826 => x"83",
          2827 => x"90",
          2828 => x"07",
          2829 => x"7a",
          2830 => x"05",
          2831 => x"58",
          2832 => x"b7",
          2833 => x"5f",
          2834 => x"06",
          2835 => x"64",
          2836 => x"26",
          2837 => x"7b",
          2838 => x"1d",
          2839 => x"38",
          2840 => x"18",
          2841 => x"34",
          2842 => x"81",
          2843 => x"38",
          2844 => x"78",
          2845 => x"57",
          2846 => x"39",
          2847 => x"58",
          2848 => x"70",
          2849 => x"f0",
          2850 => x"57",
          2851 => x"be",
          2852 => x"34",
          2853 => x"56",
          2854 => x"33",
          2855 => x"34",
          2856 => x"33",
          2857 => x"33",
          2858 => x"83",
          2859 => x"83",
          2860 => x"ff",
          2861 => x"f8",
          2862 => x"56",
          2863 => x"83",
          2864 => x"07",
          2865 => x"39",
          2866 => x"81",
          2867 => x"c3",
          2868 => x"06",
          2869 => x"34",
          2870 => x"f8",
          2871 => x"06",
          2872 => x"f4",
          2873 => x"f8",
          2874 => x"f4",
          2875 => x"75",
          2876 => x"83",
          2877 => x"e0",
          2878 => x"fe",
          2879 => x"cf",
          2880 => x"f8",
          2881 => x"f4",
          2882 => x"75",
          2883 => x"83",
          2884 => x"07",
          2885 => x"b3",
          2886 => x"06",
          2887 => x"34",
          2888 => x"81",
          2889 => x"f8",
          2890 => x"f4",
          2891 => x"f8",
          2892 => x"f4",
          2893 => x"f8",
          2894 => x"f4",
          2895 => x"f8",
          2896 => x"f4",
          2897 => x"56",
          2898 => x"39",
          2899 => x"b0",
          2900 => x"fd",
          2901 => x"34",
          2902 => x"ec",
          2903 => x"f8",
          2904 => x"f8",
          2905 => x"78",
          2906 => x"b8",
          2907 => x"84",
          2908 => x"c8",
          2909 => x"f8",
          2910 => x"81",
          2911 => x"cf",
          2912 => x"dc",
          2913 => x"fd",
          2914 => x"84",
          2915 => x"80",
          2916 => x"84",
          2917 => x"77",
          2918 => x"84",
          2919 => x"7a",
          2920 => x"fe",
          2921 => x"84",
          2922 => x"b8",
          2923 => x"f8",
          2924 => x"97",
          2925 => x"ff",
          2926 => x"39",
          2927 => x"52",
          2928 => x"39",
          2929 => x"8f",
          2930 => x"70",
          2931 => x"5f",
          2932 => x"51",
          2933 => x"75",
          2934 => x"f8",
          2935 => x"f8",
          2936 => x"2c",
          2937 => x"39",
          2938 => x"b7",
          2939 => x"75",
          2940 => x"f3",
          2941 => x"81",
          2942 => x"ee",
          2943 => x"b7",
          2944 => x"f8",
          2945 => x"a7",
          2946 => x"5f",
          2947 => x"ff",
          2948 => x"5b",
          2949 => x"81",
          2950 => x"ff",
          2951 => x"89",
          2952 => x"76",
          2953 => x"75",
          2954 => x"06",
          2955 => x"83",
          2956 => x"76",
          2957 => x"56",
          2958 => x"ff",
          2959 => x"80",
          2960 => x"77",
          2961 => x"71",
          2962 => x"86",
          2963 => x"80",
          2964 => x"06",
          2965 => x"5d",
          2966 => x"98",
          2967 => x"5e",
          2968 => x"81",
          2969 => x"58",
          2970 => x"81",
          2971 => x"bb",
          2972 => x"5d",
          2973 => x"e0",
          2974 => x"1e",
          2975 => x"76",
          2976 => x"81",
          2977 => x"bc",
          2978 => x"29",
          2979 => x"26",
          2980 => x"f8",
          2981 => x"1c",
          2982 => x"84",
          2983 => x"84",
          2984 => x"fd",
          2985 => x"b7",
          2986 => x"11",
          2987 => x"38",
          2988 => x"77",
          2989 => x"80",
          2990 => x"83",
          2991 => x"70",
          2992 => x"56",
          2993 => x"56",
          2994 => x"39",
          2995 => x"b7",
          2996 => x"75",
          2997 => x"ef",
          2998 => x"06",
          2999 => x"70",
          3000 => x"7a",
          3001 => x"09",
          3002 => x"39",
          3003 => x"34",
          3004 => x"83",
          3005 => x"7b",
          3006 => x"f2",
          3007 => x"7a",
          3008 => x"81",
          3009 => x"77",
          3010 => x"26",
          3011 => x"05",
          3012 => x"70",
          3013 => x"d4",
          3014 => x"56",
          3015 => x"39",
          3016 => x"ad",
          3017 => x"84",
          3018 => x"f1",
          3019 => x"34",
          3020 => x"33",
          3021 => x"34",
          3022 => x"a7",
          3023 => x"33",
          3024 => x"80",
          3025 => x"3f",
          3026 => x"3d",
          3027 => x"ab",
          3028 => x"85",
          3029 => x"bf",
          3030 => x"cc",
          3031 => x"ac",
          3032 => x"80",
          3033 => x"75",
          3034 => x"84",
          3035 => x"83",
          3036 => x"80",
          3037 => x"30",
          3038 => x"56",
          3039 => x"0c",
          3040 => x"09",
          3041 => x"83",
          3042 => x"07",
          3043 => x"c4",
          3044 => x"f9",
          3045 => x"29",
          3046 => x"f8",
          3047 => x"29",
          3048 => x"f7",
          3049 => x"81",
          3050 => x"73",
          3051 => x"87",
          3052 => x"88",
          3053 => x"86",
          3054 => x"f4",
          3055 => x"ff",
          3056 => x"cf",
          3057 => x"33",
          3058 => x"16",
          3059 => x"85",
          3060 => x"b4",
          3061 => x"75",
          3062 => x"2e",
          3063 => x"15",
          3064 => x"f6",
          3065 => x"ff",
          3066 => x"b3",
          3067 => x"2b",
          3068 => x"83",
          3069 => x"70",
          3070 => x"51",
          3071 => x"38",
          3072 => x"09",
          3073 => x"e4",
          3074 => x"80",
          3075 => x"a8",
          3076 => x"f7",
          3077 => x"5d",
          3078 => x"fc",
          3079 => x"8d",
          3080 => x"73",
          3081 => x"86",
          3082 => x"8b",
          3083 => x"73",
          3084 => x"54",
          3085 => x"f7",
          3086 => x"81",
          3087 => x"72",
          3088 => x"f7",
          3089 => x"84",
          3090 => x"e8",
          3091 => x"54",
          3092 => x"0b",
          3093 => x"9c",
          3094 => x"06",
          3095 => x"38",
          3096 => x"f7",
          3097 => x"9c",
          3098 => x"83",
          3099 => x"83",
          3100 => x"91",
          3101 => x"9c",
          3102 => x"dc",
          3103 => x"54",
          3104 => x"54",
          3105 => x"98",
          3106 => x"81",
          3107 => x"38",
          3108 => x"b7",
          3109 => x"54",
          3110 => x"53",
          3111 => x"81",
          3112 => x"34",
          3113 => x"58",
          3114 => x"83",
          3115 => x"77",
          3116 => x"7d",
          3117 => x"2e",
          3118 => x"59",
          3119 => x"54",
          3120 => x"2e",
          3121 => x"06",
          3122 => x"27",
          3123 => x"54",
          3124 => x"10",
          3125 => x"2b",
          3126 => x"33",
          3127 => x"9c",
          3128 => x"ea",
          3129 => x"a8",
          3130 => x"a0",
          3131 => x"ff",
          3132 => x"b7",
          3133 => x"83",
          3134 => x"70",
          3135 => x"7d",
          3136 => x"06",
          3137 => x"c6",
          3138 => x"83",
          3139 => x"78",
          3140 => x"70",
          3141 => x"27",
          3142 => x"72",
          3143 => x"c0",
          3144 => x"81",
          3145 => x"3f",
          3146 => x"0d",
          3147 => x"f9",
          3148 => x"38",
          3149 => x"5b",
          3150 => x"c9",
          3151 => x"34",
          3152 => x"ff",
          3153 => x"b1",
          3154 => x"81",
          3155 => x"90",
          3156 => x"8a",
          3157 => x"81",
          3158 => x"83",
          3159 => x"c0",
          3160 => x"27",
          3161 => x"08",
          3162 => x"06",
          3163 => x"f6",
          3164 => x"83",
          3165 => x"53",
          3166 => x"a2",
          3167 => x"83",
          3168 => x"70",
          3169 => x"33",
          3170 => x"fa",
          3171 => x"06",
          3172 => x"2e",
          3173 => x"81",
          3174 => x"ef",
          3175 => x"39",
          3176 => x"54",
          3177 => x"b7",
          3178 => x"80",
          3179 => x"76",
          3180 => x"be",
          3181 => x"53",
          3182 => x"83",
          3183 => x"f6",
          3184 => x"81",
          3185 => x"80",
          3186 => x"83",
          3187 => x"ff",
          3188 => x"38",
          3189 => x"84",
          3190 => x"56",
          3191 => x"38",
          3192 => x"ff",
          3193 => x"51",
          3194 => x"aa",
          3195 => x"14",
          3196 => x"de",
          3197 => x"34",
          3198 => x"39",
          3199 => x"3f",
          3200 => x"80",
          3201 => x"02",
          3202 => x"f3",
          3203 => x"85",
          3204 => x"fe",
          3205 => x"f0",
          3206 => x"08",
          3207 => x"90",
          3208 => x"52",
          3209 => x"72",
          3210 => x"c0",
          3211 => x"27",
          3212 => x"38",
          3213 => x"55",
          3214 => x"55",
          3215 => x"c0",
          3216 => x"53",
          3217 => x"c0",
          3218 => x"f6",
          3219 => x"9c",
          3220 => x"38",
          3221 => x"c0",
          3222 => x"83",
          3223 => x"70",
          3224 => x"2e",
          3225 => x"71",
          3226 => x"38",
          3227 => x"0d",
          3228 => x"88",
          3229 => x"02",
          3230 => x"80",
          3231 => x"2b",
          3232 => x"98",
          3233 => x"83",
          3234 => x"84",
          3235 => x"85",
          3236 => x"f3",
          3237 => x"83",
          3238 => x"34",
          3239 => x"56",
          3240 => x"86",
          3241 => x"9c",
          3242 => x"ce",
          3243 => x"08",
          3244 => x"70",
          3245 => x"87",
          3246 => x"73",
          3247 => x"db",
          3248 => x"ff",
          3249 => x"71",
          3250 => x"87",
          3251 => x"05",
          3252 => x"87",
          3253 => x"2e",
          3254 => x"98",
          3255 => x"87",
          3256 => x"87",
          3257 => x"26",
          3258 => x"16",
          3259 => x"80",
          3260 => x"06",
          3261 => x"70",
          3262 => x"80",
          3263 => x"52",
          3264 => x"70",
          3265 => x"05",
          3266 => x"76",
          3267 => x"04",
          3268 => x"3d",
          3269 => x"3d",
          3270 => x"33",
          3271 => x"08",
          3272 => x"06",
          3273 => x"55",
          3274 => x"2a",
          3275 => x"2a",
          3276 => x"15",
          3277 => x"c6",
          3278 => x"51",
          3279 => x"81",
          3280 => x"54",
          3281 => x"f3",
          3282 => x"83",
          3283 => x"34",
          3284 => x"56",
          3285 => x"86",
          3286 => x"9c",
          3287 => x"ce",
          3288 => x"08",
          3289 => x"70",
          3290 => x"87",
          3291 => x"73",
          3292 => x"db",
          3293 => x"ff",
          3294 => x"71",
          3295 => x"87",
          3296 => x"05",
          3297 => x"87",
          3298 => x"2e",
          3299 => x"98",
          3300 => x"87",
          3301 => x"87",
          3302 => x"26",
          3303 => x"16",
          3304 => x"80",
          3305 => x"52",
          3306 => x"81",
          3307 => x"38",
          3308 => x"88",
          3309 => x"fb",
          3310 => x"80",
          3311 => x"d4",
          3312 => x"34",
          3313 => x"87",
          3314 => x"08",
          3315 => x"c0",
          3316 => x"9c",
          3317 => x"81",
          3318 => x"52",
          3319 => x"81",
          3320 => x"a4",
          3321 => x"80",
          3322 => x"80",
          3323 => x"80",
          3324 => x"9c",
          3325 => x"51",
          3326 => x"33",
          3327 => x"73",
          3328 => x"2e",
          3329 => x"51",
          3330 => x"71",
          3331 => x"57",
          3332 => x"81",
          3333 => x"ff",
          3334 => x"51",
          3335 => x"04",
          3336 => x"7a",
          3337 => x"ff",
          3338 => x"33",
          3339 => x"83",
          3340 => x"12",
          3341 => x"07",
          3342 => x"59",
          3343 => x"81",
          3344 => x"83",
          3345 => x"2b",
          3346 => x"33",
          3347 => x"57",
          3348 => x"71",
          3349 => x"85",
          3350 => x"2b",
          3351 => x"54",
          3352 => x"81",
          3353 => x"84",
          3354 => x"33",
          3355 => x"70",
          3356 => x"77",
          3357 => x"84",
          3358 => x"86",
          3359 => x"84",
          3360 => x"34",
          3361 => x"08",
          3362 => x"88",
          3363 => x"88",
          3364 => x"34",
          3365 => x"04",
          3366 => x"8b",
          3367 => x"84",
          3368 => x"2b",
          3369 => x"51",
          3370 => x"72",
          3371 => x"70",
          3372 => x"71",
          3373 => x"5a",
          3374 => x"87",
          3375 => x"88",
          3376 => x"13",
          3377 => x"b8",
          3378 => x"71",
          3379 => x"70",
          3380 => x"72",
          3381 => x"b8",
          3382 => x"33",
          3383 => x"74",
          3384 => x"88",
          3385 => x"f8",
          3386 => x"52",
          3387 => x"77",
          3388 => x"84",
          3389 => x"81",
          3390 => x"2b",
          3391 => x"33",
          3392 => x"06",
          3393 => x"5a",
          3394 => x"81",
          3395 => x"17",
          3396 => x"8b",
          3397 => x"70",
          3398 => x"71",
          3399 => x"5a",
          3400 => x"e4",
          3401 => x"88",
          3402 => x"88",
          3403 => x"77",
          3404 => x"70",
          3405 => x"8b",
          3406 => x"82",
          3407 => x"2b",
          3408 => x"52",
          3409 => x"34",
          3410 => x"04",
          3411 => x"08",
          3412 => x"77",
          3413 => x"90",
          3414 => x"f4",
          3415 => x"0b",
          3416 => x"53",
          3417 => x"d3",
          3418 => x"76",
          3419 => x"84",
          3420 => x"34",
          3421 => x"b8",
          3422 => x"0b",
          3423 => x"84",
          3424 => x"80",
          3425 => x"88",
          3426 => x"17",
          3427 => x"b4",
          3428 => x"b8",
          3429 => x"82",
          3430 => x"fe",
          3431 => x"80",
          3432 => x"38",
          3433 => x"83",
          3434 => x"ff",
          3435 => x"11",
          3436 => x"07",
          3437 => x"ff",
          3438 => x"38",
          3439 => x"81",
          3440 => x"81",
          3441 => x"ff",
          3442 => x"5c",
          3443 => x"38",
          3444 => x"55",
          3445 => x"71",
          3446 => x"38",
          3447 => x"77",
          3448 => x"78",
          3449 => x"88",
          3450 => x"56",
          3451 => x"2e",
          3452 => x"73",
          3453 => x"80",
          3454 => x"82",
          3455 => x"78",
          3456 => x"88",
          3457 => x"74",
          3458 => x"b8",
          3459 => x"71",
          3460 => x"84",
          3461 => x"81",
          3462 => x"83",
          3463 => x"7e",
          3464 => x"5c",
          3465 => x"82",
          3466 => x"72",
          3467 => x"18",
          3468 => x"34",
          3469 => x"11",
          3470 => x"71",
          3471 => x"5c",
          3472 => x"85",
          3473 => x"16",
          3474 => x"12",
          3475 => x"2a",
          3476 => x"34",
          3477 => x"08",
          3478 => x"33",
          3479 => x"74",
          3480 => x"86",
          3481 => x"b9",
          3482 => x"84",
          3483 => x"2b",
          3484 => x"59",
          3485 => x"34",
          3486 => x"51",
          3487 => x"0d",
          3488 => x"71",
          3489 => x"05",
          3490 => x"88",
          3491 => x"59",
          3492 => x"76",
          3493 => x"70",
          3494 => x"71",
          3495 => x"05",
          3496 => x"88",
          3497 => x"5f",
          3498 => x"1a",
          3499 => x"b8",
          3500 => x"71",
          3501 => x"70",
          3502 => x"77",
          3503 => x"b8",
          3504 => x"39",
          3505 => x"08",
          3506 => x"77",
          3507 => x"c8",
          3508 => x"fb",
          3509 => x"b9",
          3510 => x"ff",
          3511 => x"80",
          3512 => x"80",
          3513 => x"fe",
          3514 => x"55",
          3515 => x"34",
          3516 => x"15",
          3517 => x"b9",
          3518 => x"81",
          3519 => x"08",
          3520 => x"80",
          3521 => x"70",
          3522 => x"88",
          3523 => x"b9",
          3524 => x"b9",
          3525 => x"76",
          3526 => x"34",
          3527 => x"38",
          3528 => x"67",
          3529 => x"08",
          3530 => x"aa",
          3531 => x"7f",
          3532 => x"84",
          3533 => x"83",
          3534 => x"06",
          3535 => x"7f",
          3536 => x"ff",
          3537 => x"33",
          3538 => x"70",
          3539 => x"70",
          3540 => x"2b",
          3541 => x"71",
          3542 => x"90",
          3543 => x"54",
          3544 => x"5f",
          3545 => x"82",
          3546 => x"2b",
          3547 => x"33",
          3548 => x"90",
          3549 => x"56",
          3550 => x"62",
          3551 => x"77",
          3552 => x"2e",
          3553 => x"62",
          3554 => x"61",
          3555 => x"70",
          3556 => x"71",
          3557 => x"81",
          3558 => x"2b",
          3559 => x"5b",
          3560 => x"76",
          3561 => x"71",
          3562 => x"11",
          3563 => x"8b",
          3564 => x"84",
          3565 => x"2b",
          3566 => x"52",
          3567 => x"77",
          3568 => x"84",
          3569 => x"33",
          3570 => x"83",
          3571 => x"87",
          3572 => x"88",
          3573 => x"41",
          3574 => x"16",
          3575 => x"33",
          3576 => x"81",
          3577 => x"5c",
          3578 => x"1a",
          3579 => x"82",
          3580 => x"2b",
          3581 => x"33",
          3582 => x"70",
          3583 => x"5a",
          3584 => x"1a",
          3585 => x"70",
          3586 => x"71",
          3587 => x"33",
          3588 => x"70",
          3589 => x"5a",
          3590 => x"83",
          3591 => x"1f",
          3592 => x"88",
          3593 => x"83",
          3594 => x"84",
          3595 => x"b9",
          3596 => x"05",
          3597 => x"44",
          3598 => x"7e",
          3599 => x"3d",
          3600 => x"b9",
          3601 => x"b4",
          3602 => x"84",
          3603 => x"84",
          3604 => x"81",
          3605 => x"08",
          3606 => x"85",
          3607 => x"60",
          3608 => x"34",
          3609 => x"22",
          3610 => x"83",
          3611 => x"5a",
          3612 => x"89",
          3613 => x"10",
          3614 => x"f8",
          3615 => x"81",
          3616 => x"08",
          3617 => x"2e",
          3618 => x"2e",
          3619 => x"3f",
          3620 => x"0c",
          3621 => x"b9",
          3622 => x"5e",
          3623 => x"33",
          3624 => x"06",
          3625 => x"40",
          3626 => x"61",
          3627 => x"2a",
          3628 => x"83",
          3629 => x"1f",
          3630 => x"2b",
          3631 => x"06",
          3632 => x"70",
          3633 => x"5b",
          3634 => x"81",
          3635 => x"34",
          3636 => x"7b",
          3637 => x"b9",
          3638 => x"88",
          3639 => x"75",
          3640 => x"54",
          3641 => x"06",
          3642 => x"82",
          3643 => x"2b",
          3644 => x"33",
          3645 => x"90",
          3646 => x"58",
          3647 => x"38",
          3648 => x"83",
          3649 => x"77",
          3650 => x"27",
          3651 => x"ff",
          3652 => x"80",
          3653 => x"80",
          3654 => x"fe",
          3655 => x"5a",
          3656 => x"34",
          3657 => x"1a",
          3658 => x"b9",
          3659 => x"81",
          3660 => x"08",
          3661 => x"80",
          3662 => x"70",
          3663 => x"64",
          3664 => x"34",
          3665 => x"10",
          3666 => x"42",
          3667 => x"61",
          3668 => x"7a",
          3669 => x"ff",
          3670 => x"38",
          3671 => x"bd",
          3672 => x"54",
          3673 => x"0d",
          3674 => x"12",
          3675 => x"07",
          3676 => x"33",
          3677 => x"7e",
          3678 => x"71",
          3679 => x"44",
          3680 => x"45",
          3681 => x"64",
          3682 => x"70",
          3683 => x"71",
          3684 => x"05",
          3685 => x"88",
          3686 => x"42",
          3687 => x"86",
          3688 => x"84",
          3689 => x"12",
          3690 => x"ff",
          3691 => x"5d",
          3692 => x"84",
          3693 => x"33",
          3694 => x"83",
          3695 => x"15",
          3696 => x"2a",
          3697 => x"54",
          3698 => x"84",
          3699 => x"81",
          3700 => x"2b",
          3701 => x"15",
          3702 => x"2a",
          3703 => x"55",
          3704 => x"34",
          3705 => x"11",
          3706 => x"07",
          3707 => x"42",
          3708 => x"51",
          3709 => x"08",
          3710 => x"06",
          3711 => x"f4",
          3712 => x"0b",
          3713 => x"53",
          3714 => x"c0",
          3715 => x"7f",
          3716 => x"84",
          3717 => x"34",
          3718 => x"b8",
          3719 => x"0b",
          3720 => x"84",
          3721 => x"80",
          3722 => x"88",
          3723 => x"1f",
          3724 => x"b4",
          3725 => x"b8",
          3726 => x"82",
          3727 => x"7e",
          3728 => x"c0",
          3729 => x"71",
          3730 => x"05",
          3731 => x"88",
          3732 => x"5e",
          3733 => x"34",
          3734 => x"b8",
          3735 => x"12",
          3736 => x"07",
          3737 => x"33",
          3738 => x"41",
          3739 => x"79",
          3740 => x"05",
          3741 => x"33",
          3742 => x"81",
          3743 => x"42",
          3744 => x"19",
          3745 => x"70",
          3746 => x"71",
          3747 => x"81",
          3748 => x"83",
          3749 => x"63",
          3750 => x"40",
          3751 => x"7b",
          3752 => x"70",
          3753 => x"8b",
          3754 => x"70",
          3755 => x"07",
          3756 => x"48",
          3757 => x"60",
          3758 => x"61",
          3759 => x"39",
          3760 => x"8b",
          3761 => x"84",
          3762 => x"2b",
          3763 => x"52",
          3764 => x"85",
          3765 => x"19",
          3766 => x"8b",
          3767 => x"86",
          3768 => x"2b",
          3769 => x"52",
          3770 => x"05",
          3771 => x"b9",
          3772 => x"33",
          3773 => x"06",
          3774 => x"77",
          3775 => x"b9",
          3776 => x"12",
          3777 => x"07",
          3778 => x"71",
          3779 => x"ff",
          3780 => x"56",
          3781 => x"55",
          3782 => x"34",
          3783 => x"33",
          3784 => x"83",
          3785 => x"12",
          3786 => x"ff",
          3787 => x"58",
          3788 => x"76",
          3789 => x"70",
          3790 => x"71",
          3791 => x"11",
          3792 => x"8b",
          3793 => x"84",
          3794 => x"2b",
          3795 => x"52",
          3796 => x"57",
          3797 => x"34",
          3798 => x"11",
          3799 => x"71",
          3800 => x"33",
          3801 => x"70",
          3802 => x"57",
          3803 => x"87",
          3804 => x"70",
          3805 => x"07",
          3806 => x"5a",
          3807 => x"81",
          3808 => x"1f",
          3809 => x"8b",
          3810 => x"73",
          3811 => x"07",
          3812 => x"5f",
          3813 => x"81",
          3814 => x"1f",
          3815 => x"2b",
          3816 => x"14",
          3817 => x"07",
          3818 => x"5f",
          3819 => x"75",
          3820 => x"70",
          3821 => x"71",
          3822 => x"70",
          3823 => x"05",
          3824 => x"84",
          3825 => x"65",
          3826 => x"5d",
          3827 => x"33",
          3828 => x"83",
          3829 => x"85",
          3830 => x"88",
          3831 => x"7a",
          3832 => x"05",
          3833 => x"84",
          3834 => x"2b",
          3835 => x"14",
          3836 => x"07",
          3837 => x"5c",
          3838 => x"34",
          3839 => x"b8",
          3840 => x"71",
          3841 => x"70",
          3842 => x"75",
          3843 => x"b8",
          3844 => x"33",
          3845 => x"74",
          3846 => x"88",
          3847 => x"f8",
          3848 => x"44",
          3849 => x"74",
          3850 => x"84",
          3851 => x"81",
          3852 => x"2b",
          3853 => x"33",
          3854 => x"06",
          3855 => x"46",
          3856 => x"81",
          3857 => x"5b",
          3858 => x"e5",
          3859 => x"84",
          3860 => x"62",
          3861 => x"51",
          3862 => x"88",
          3863 => x"b7",
          3864 => x"7a",
          3865 => x"58",
          3866 => x"77",
          3867 => x"89",
          3868 => x"3f",
          3869 => x"c8",
          3870 => x"80",
          3871 => x"b7",
          3872 => x"89",
          3873 => x"84",
          3874 => x"b9",
          3875 => x"52",
          3876 => x"3f",
          3877 => x"34",
          3878 => x"b8",
          3879 => x"0b",
          3880 => x"56",
          3881 => x"17",
          3882 => x"b4",
          3883 => x"70",
          3884 => x"58",
          3885 => x"73",
          3886 => x"70",
          3887 => x"05",
          3888 => x"34",
          3889 => x"77",
          3890 => x"39",
          3891 => x"51",
          3892 => x"84",
          3893 => x"b9",
          3894 => x"3d",
          3895 => x"53",
          3896 => x"d4",
          3897 => x"ff",
          3898 => x"b9",
          3899 => x"33",
          3900 => x"3d",
          3901 => x"60",
          3902 => x"5c",
          3903 => x"87",
          3904 => x"73",
          3905 => x"38",
          3906 => x"8c",
          3907 => x"d5",
          3908 => x"ff",
          3909 => x"87",
          3910 => x"38",
          3911 => x"80",
          3912 => x"38",
          3913 => x"c8",
          3914 => x"16",
          3915 => x"55",
          3916 => x"d5",
          3917 => x"02",
          3918 => x"57",
          3919 => x"38",
          3920 => x"81",
          3921 => x"73",
          3922 => x"0c",
          3923 => x"8e",
          3924 => x"06",
          3925 => x"c0",
          3926 => x"79",
          3927 => x"80",
          3928 => x"81",
          3929 => x"0c",
          3930 => x"81",
          3931 => x"56",
          3932 => x"39",
          3933 => x"9b",
          3934 => x"33",
          3935 => x"26",
          3936 => x"53",
          3937 => x"9b",
          3938 => x"0c",
          3939 => x"72",
          3940 => x"9a",
          3941 => x"0c",
          3942 => x"75",
          3943 => x"3d",
          3944 => x"0b",
          3945 => x"04",
          3946 => x"11",
          3947 => x"70",
          3948 => x"80",
          3949 => x"08",
          3950 => x"8c",
          3951 => x"0c",
          3952 => x"08",
          3953 => x"9b",
          3954 => x"ee",
          3955 => x"7c",
          3956 => x"5b",
          3957 => x"06",
          3958 => x"2e",
          3959 => x"81",
          3960 => x"b9",
          3961 => x"59",
          3962 => x"0d",
          3963 => x"b8",
          3964 => x"5a",
          3965 => x"c8",
          3966 => x"38",
          3967 => x"b4",
          3968 => x"a0",
          3969 => x"58",
          3970 => x"38",
          3971 => x"09",
          3972 => x"75",
          3973 => x"51",
          3974 => x"59",
          3975 => x"fb",
          3976 => x"2e",
          3977 => x"18",
          3978 => x"75",
          3979 => x"57",
          3980 => x"b6",
          3981 => x"19",
          3982 => x"0b",
          3983 => x"19",
          3984 => x"80",
          3985 => x"f2",
          3986 => x"0b",
          3987 => x"84",
          3988 => x"74",
          3989 => x"5b",
          3990 => x"2a",
          3991 => x"98",
          3992 => x"90",
          3993 => x"34",
          3994 => x"19",
          3995 => x"a6",
          3996 => x"84",
          3997 => x"05",
          3998 => x"7a",
          3999 => x"fa",
          4000 => x"53",
          4001 => x"d8",
          4002 => x"fd",
          4003 => x"0d",
          4004 => x"81",
          4005 => x"76",
          4006 => x"b9",
          4007 => x"77",
          4008 => x"cc",
          4009 => x"74",
          4010 => x"75",
          4011 => x"19",
          4012 => x"17",
          4013 => x"33",
          4014 => x"83",
          4015 => x"17",
          4016 => x"3f",
          4017 => x"38",
          4018 => x"0c",
          4019 => x"06",
          4020 => x"89",
          4021 => x"5d",
          4022 => x"38",
          4023 => x"56",
          4024 => x"84",
          4025 => x"17",
          4026 => x"3f",
          4027 => x"38",
          4028 => x"0c",
          4029 => x"06",
          4030 => x"7e",
          4031 => x"53",
          4032 => x"38",
          4033 => x"0c",
          4034 => x"a8",
          4035 => x"79",
          4036 => x"33",
          4037 => x"09",
          4038 => x"78",
          4039 => x"51",
          4040 => x"80",
          4041 => x"78",
          4042 => x"75",
          4043 => x"05",
          4044 => x"2b",
          4045 => x"8f",
          4046 => x"81",
          4047 => x"a8",
          4048 => x"79",
          4049 => x"33",
          4050 => x"09",
          4051 => x"78",
          4052 => x"51",
          4053 => x"80",
          4054 => x"78",
          4055 => x"75",
          4056 => x"b8",
          4057 => x"71",
          4058 => x"14",
          4059 => x"33",
          4060 => x"07",
          4061 => x"59",
          4062 => x"54",
          4063 => x"53",
          4064 => x"3f",
          4065 => x"2e",
          4066 => x"b9",
          4067 => x"08",
          4068 => x"08",
          4069 => x"fe",
          4070 => x"82",
          4071 => x"81",
          4072 => x"05",
          4073 => x"f6",
          4074 => x"81",
          4075 => x"70",
          4076 => x"81",
          4077 => x"09",
          4078 => x"c8",
          4079 => x"a8",
          4080 => x"08",
          4081 => x"7d",
          4082 => x"c8",
          4083 => x"b4",
          4084 => x"81",
          4085 => x"81",
          4086 => x"09",
          4087 => x"c8",
          4088 => x"a8",
          4089 => x"5b",
          4090 => x"c5",
          4091 => x"2e",
          4092 => x"54",
          4093 => x"53",
          4094 => x"f1",
          4095 => x"54",
          4096 => x"53",
          4097 => x"3f",
          4098 => x"2e",
          4099 => x"b9",
          4100 => x"08",
          4101 => x"08",
          4102 => x"fb",
          4103 => x"82",
          4104 => x"81",
          4105 => x"05",
          4106 => x"f4",
          4107 => x"81",
          4108 => x"05",
          4109 => x"f3",
          4110 => x"7a",
          4111 => x"3d",
          4112 => x"82",
          4113 => x"9c",
          4114 => x"55",
          4115 => x"24",
          4116 => x"8a",
          4117 => x"3d",
          4118 => x"08",
          4119 => x"58",
          4120 => x"83",
          4121 => x"2e",
          4122 => x"54",
          4123 => x"33",
          4124 => x"08",
          4125 => x"5a",
          4126 => x"ff",
          4127 => x"79",
          4128 => x"5e",
          4129 => x"5a",
          4130 => x"1a",
          4131 => x"3d",
          4132 => x"06",
          4133 => x"1a",
          4134 => x"08",
          4135 => x"38",
          4136 => x"7c",
          4137 => x"81",
          4138 => x"19",
          4139 => x"c8",
          4140 => x"81",
          4141 => x"79",
          4142 => x"fc",
          4143 => x"33",
          4144 => x"f0",
          4145 => x"7d",
          4146 => x"b9",
          4147 => x"ba",
          4148 => x"bb",
          4149 => x"fe",
          4150 => x"89",
          4151 => x"08",
          4152 => x"38",
          4153 => x"56",
          4154 => x"82",
          4155 => x"19",
          4156 => x"3f",
          4157 => x"38",
          4158 => x"0c",
          4159 => x"83",
          4160 => x"77",
          4161 => x"7c",
          4162 => x"9f",
          4163 => x"07",
          4164 => x"83",
          4165 => x"08",
          4166 => x"56",
          4167 => x"81",
          4168 => x"81",
          4169 => x"81",
          4170 => x"09",
          4171 => x"c8",
          4172 => x"70",
          4173 => x"84",
          4174 => x"74",
          4175 => x"55",
          4176 => x"54",
          4177 => x"51",
          4178 => x"80",
          4179 => x"75",
          4180 => x"7d",
          4181 => x"84",
          4182 => x"88",
          4183 => x"8f",
          4184 => x"81",
          4185 => x"81",
          4186 => x"81",
          4187 => x"81",
          4188 => x"09",
          4189 => x"c8",
          4190 => x"70",
          4191 => x"84",
          4192 => x"7e",
          4193 => x"33",
          4194 => x"fb",
          4195 => x"7c",
          4196 => x"3f",
          4197 => x"76",
          4198 => x"33",
          4199 => x"84",
          4200 => x"06",
          4201 => x"83",
          4202 => x"1b",
          4203 => x"c8",
          4204 => x"27",
          4205 => x"74",
          4206 => x"38",
          4207 => x"81",
          4208 => x"5c",
          4209 => x"b8",
          4210 => x"57",
          4211 => x"c8",
          4212 => x"c5",
          4213 => x"34",
          4214 => x"31",
          4215 => x"5d",
          4216 => x"87",
          4217 => x"2e",
          4218 => x"54",
          4219 => x"33",
          4220 => x"e7",
          4221 => x"52",
          4222 => x"7e",
          4223 => x"83",
          4224 => x"ff",
          4225 => x"34",
          4226 => x"34",
          4227 => x"39",
          4228 => x"7a",
          4229 => x"98",
          4230 => x"06",
          4231 => x"7d",
          4232 => x"1d",
          4233 => x"1d",
          4234 => x"1d",
          4235 => x"7c",
          4236 => x"81",
          4237 => x"80",
          4238 => x"08",
          4239 => x"70",
          4240 => x"38",
          4241 => x"56",
          4242 => x"26",
          4243 => x"82",
          4244 => x"f5",
          4245 => x"81",
          4246 => x"08",
          4247 => x"08",
          4248 => x"25",
          4249 => x"73",
          4250 => x"81",
          4251 => x"84",
          4252 => x"81",
          4253 => x"08",
          4254 => x"f0",
          4255 => x"c8",
          4256 => x"08",
          4257 => x"ce",
          4258 => x"08",
          4259 => x"39",
          4260 => x"26",
          4261 => x"51",
          4262 => x"c8",
          4263 => x"b9",
          4264 => x"07",
          4265 => x"c8",
          4266 => x"ff",
          4267 => x"2e",
          4268 => x"74",
          4269 => x"08",
          4270 => x"57",
          4271 => x"8e",
          4272 => x"f5",
          4273 => x"b9",
          4274 => x"08",
          4275 => x"80",
          4276 => x"90",
          4277 => x"94",
          4278 => x"86",
          4279 => x"19",
          4280 => x"34",
          4281 => x"8c",
          4282 => x"c8",
          4283 => x"c8",
          4284 => x"2e",
          4285 => x"78",
          4286 => x"08",
          4287 => x"08",
          4288 => x"04",
          4289 => x"38",
          4290 => x"0d",
          4291 => x"73",
          4292 => x"73",
          4293 => x"73",
          4294 => x"74",
          4295 => x"82",
          4296 => x"53",
          4297 => x"72",
          4298 => x"98",
          4299 => x"18",
          4300 => x"94",
          4301 => x"0c",
          4302 => x"9c",
          4303 => x"c8",
          4304 => x"84",
          4305 => x"ac",
          4306 => x"ac",
          4307 => x"57",
          4308 => x"17",
          4309 => x"56",
          4310 => x"8a",
          4311 => x"08",
          4312 => x"ff",
          4313 => x"cd",
          4314 => x"b9",
          4315 => x"0b",
          4316 => x"38",
          4317 => x"08",
          4318 => x"31",
          4319 => x"aa",
          4320 => x"8a",
          4321 => x"70",
          4322 => x"5a",
          4323 => x"38",
          4324 => x"08",
          4325 => x"38",
          4326 => x"38",
          4327 => x"75",
          4328 => x"22",
          4329 => x"38",
          4330 => x"0c",
          4331 => x"80",
          4332 => x"3d",
          4333 => x"19",
          4334 => x"5c",
          4335 => x"eb",
          4336 => x"82",
          4337 => x"27",
          4338 => x"08",
          4339 => x"84",
          4340 => x"60",
          4341 => x"08",
          4342 => x"b9",
          4343 => x"c8",
          4344 => x"56",
          4345 => x"91",
          4346 => x"ff",
          4347 => x"08",
          4348 => x"ea",
          4349 => x"05",
          4350 => x"8d",
          4351 => x"b0",
          4352 => x"1a",
          4353 => x"57",
          4354 => x"34",
          4355 => x"56",
          4356 => x"81",
          4357 => x"77",
          4358 => x"3f",
          4359 => x"81",
          4360 => x"0c",
          4361 => x"3d",
          4362 => x"53",
          4363 => x"52",
          4364 => x"08",
          4365 => x"83",
          4366 => x"08",
          4367 => x"fe",
          4368 => x"82",
          4369 => x"81",
          4370 => x"05",
          4371 => x"e3",
          4372 => x"22",
          4373 => x"74",
          4374 => x"7c",
          4375 => x"08",
          4376 => x"7d",
          4377 => x"76",
          4378 => x"19",
          4379 => x"84",
          4380 => x"ee",
          4381 => x"7c",
          4382 => x"1e",
          4383 => x"82",
          4384 => x"80",
          4385 => x"d1",
          4386 => x"74",
          4387 => x"38",
          4388 => x"81",
          4389 => x"b9",
          4390 => x"5a",
          4391 => x"5b",
          4392 => x"70",
          4393 => x"81",
          4394 => x"81",
          4395 => x"34",
          4396 => x"ae",
          4397 => x"80",
          4398 => x"74",
          4399 => x"56",
          4400 => x"60",
          4401 => x"80",
          4402 => x"b9",
          4403 => x"81",
          4404 => x"fe",
          4405 => x"94",
          4406 => x"08",
          4407 => x"e1",
          4408 => x"08",
          4409 => x"38",
          4410 => x"b4",
          4411 => x"b9",
          4412 => x"08",
          4413 => x"41",
          4414 => x"a8",
          4415 => x"1a",
          4416 => x"33",
          4417 => x"90",
          4418 => x"81",
          4419 => x"5b",
          4420 => x"33",
          4421 => x"08",
          4422 => x"76",
          4423 => x"74",
          4424 => x"60",
          4425 => x"c1",
          4426 => x"0c",
          4427 => x"0d",
          4428 => x"18",
          4429 => x"06",
          4430 => x"33",
          4431 => x"58",
          4432 => x"33",
          4433 => x"05",
          4434 => x"e5",
          4435 => x"33",
          4436 => x"44",
          4437 => x"79",
          4438 => x"10",
          4439 => x"23",
          4440 => x"77",
          4441 => x"2a",
          4442 => x"90",
          4443 => x"38",
          4444 => x"23",
          4445 => x"41",
          4446 => x"2e",
          4447 => x"39",
          4448 => x"74",
          4449 => x"78",
          4450 => x"05",
          4451 => x"56",
          4452 => x"fd",
          4453 => x"7a",
          4454 => x"04",
          4455 => x"5c",
          4456 => x"84",
          4457 => x"08",
          4458 => x"5d",
          4459 => x"5e",
          4460 => x"1b",
          4461 => x"1b",
          4462 => x"09",
          4463 => x"75",
          4464 => x"51",
          4465 => x"80",
          4466 => x"75",
          4467 => x"b2",
          4468 => x"59",
          4469 => x"19",
          4470 => x"57",
          4471 => x"e5",
          4472 => x"81",
          4473 => x"38",
          4474 => x"81",
          4475 => x"56",
          4476 => x"81",
          4477 => x"5a",
          4478 => x"06",
          4479 => x"38",
          4480 => x"1c",
          4481 => x"8b",
          4482 => x"81",
          4483 => x"5a",
          4484 => x"58",
          4485 => x"38",
          4486 => x"5d",
          4487 => x"7b",
          4488 => x"08",
          4489 => x"fe",
          4490 => x"93",
          4491 => x"08",
          4492 => x"dc",
          4493 => x"08",
          4494 => x"38",
          4495 => x"b4",
          4496 => x"b9",
          4497 => x"08",
          4498 => x"5a",
          4499 => x"dd",
          4500 => x"1c",
          4501 => x"33",
          4502 => x"c5",
          4503 => x"1c",
          4504 => x"55",
          4505 => x"81",
          4506 => x"8d",
          4507 => x"90",
          4508 => x"5e",
          4509 => x"ff",
          4510 => x"f4",
          4511 => x"84",
          4512 => x"38",
          4513 => x"c2",
          4514 => x"1d",
          4515 => x"57",
          4516 => x"38",
          4517 => x"1b",
          4518 => x"40",
          4519 => x"bf",
          4520 => x"81",
          4521 => x"33",
          4522 => x"71",
          4523 => x"80",
          4524 => x"26",
          4525 => x"8a",
          4526 => x"61",
          4527 => x"5b",
          4528 => x"b9",
          4529 => x"de",
          4530 => x"78",
          4531 => x"86",
          4532 => x"2e",
          4533 => x"79",
          4534 => x"7f",
          4535 => x"ff",
          4536 => x"0b",
          4537 => x"04",
          4538 => x"38",
          4539 => x"3d",
          4540 => x"33",
          4541 => x"86",
          4542 => x"1d",
          4543 => x"80",
          4544 => x"17",
          4545 => x"38",
          4546 => x"60",
          4547 => x"05",
          4548 => x"34",
          4549 => x"80",
          4550 => x"56",
          4551 => x"c0",
          4552 => x"3d",
          4553 => x"59",
          4554 => x"70",
          4555 => x"05",
          4556 => x"38",
          4557 => x"79",
          4558 => x"38",
          4559 => x"75",
          4560 => x"2a",
          4561 => x"2a",
          4562 => x"80",
          4563 => x"32",
          4564 => x"d7",
          4565 => x"87",
          4566 => x"58",
          4567 => x"75",
          4568 => x"76",
          4569 => x"2a",
          4570 => x"1f",
          4571 => x"58",
          4572 => x"33",
          4573 => x"16",
          4574 => x"75",
          4575 => x"2e",
          4576 => x"56",
          4577 => x"98",
          4578 => x"71",
          4579 => x"87",
          4580 => x"f8",
          4581 => x"38",
          4582 => x"fe",
          4583 => x"2e",
          4584 => x"56",
          4585 => x"81",
          4586 => x"05",
          4587 => x"84",
          4588 => x"75",
          4589 => x"7e",
          4590 => x"1d",
          4591 => x"c8",
          4592 => x"ed",
          4593 => x"84",
          4594 => x"b9",
          4595 => x"1e",
          4596 => x"76",
          4597 => x"40",
          4598 => x"a3",
          4599 => x"52",
          4600 => x"84",
          4601 => x"ff",
          4602 => x"76",
          4603 => x"70",
          4604 => x"81",
          4605 => x"78",
          4606 => x"c9",
          4607 => x"86",
          4608 => x"83",
          4609 => x"b9",
          4610 => x"87",
          4611 => x"75",
          4612 => x"40",
          4613 => x"57",
          4614 => x"83",
          4615 => x"82",
          4616 => x"52",
          4617 => x"84",
          4618 => x"ff",
          4619 => x"75",
          4620 => x"9c",
          4621 => x"81",
          4622 => x"f4",
          4623 => x"58",
          4624 => x"33",
          4625 => x"15",
          4626 => x"ab",
          4627 => x"8c",
          4628 => x"77",
          4629 => x"3d",
          4630 => x"25",
          4631 => x"b9",
          4632 => x"ec",
          4633 => x"84",
          4634 => x"38",
          4635 => x"08",
          4636 => x"d3",
          4637 => x"2e",
          4638 => x"b9",
          4639 => x"08",
          4640 => x"19",
          4641 => x"41",
          4642 => x"b9",
          4643 => x"85",
          4644 => x"58",
          4645 => x"c8",
          4646 => x"ef",
          4647 => x"58",
          4648 => x"80",
          4649 => x"33",
          4650 => x"ff",
          4651 => x"74",
          4652 => x"98",
          4653 => x"08",
          4654 => x"5b",
          4655 => x"c9",
          4656 => x"52",
          4657 => x"84",
          4658 => x"ff",
          4659 => x"75",
          4660 => x"08",
          4661 => x"5f",
          4662 => x"0b",
          4663 => x"75",
          4664 => x"7c",
          4665 => x"58",
          4666 => x"38",
          4667 => x"5b",
          4668 => x"7b",
          4669 => x"57",
          4670 => x"34",
          4671 => x"81",
          4672 => x"76",
          4673 => x"78",
          4674 => x"80",
          4675 => x"81",
          4676 => x"51",
          4677 => x"58",
          4678 => x"7f",
          4679 => x"fb",
          4680 => x"53",
          4681 => x"52",
          4682 => x"b9",
          4683 => x"c8",
          4684 => x"a8",
          4685 => x"57",
          4686 => x"c9",
          4687 => x"2e",
          4688 => x"54",
          4689 => x"53",
          4690 => x"d1",
          4691 => x"9c",
          4692 => x"74",
          4693 => x"ba",
          4694 => x"57",
          4695 => x"d7",
          4696 => x"d4",
          4697 => x"61",
          4698 => x"3f",
          4699 => x"81",
          4700 => x"83",
          4701 => x"08",
          4702 => x"8a",
          4703 => x"2e",
          4704 => x"fc",
          4705 => x"7f",
          4706 => x"39",
          4707 => x"70",
          4708 => x"38",
          4709 => x"08",
          4710 => x"81",
          4711 => x"c1",
          4712 => x"19",
          4713 => x"33",
          4714 => x"f3",
          4715 => x"5e",
          4716 => x"1c",
          4717 => x"1c",
          4718 => x"70",
          4719 => x"57",
          4720 => x"bc",
          4721 => x"81",
          4722 => x"38",
          4723 => x"ff",
          4724 => x"82",
          4725 => x"70",
          4726 => x"38",
          4727 => x"7a",
          4728 => x"05",
          4729 => x"70",
          4730 => x"08",
          4731 => x"53",
          4732 => x"2e",
          4733 => x"30",
          4734 => x"54",
          4735 => x"2e",
          4736 => x"59",
          4737 => x"81",
          4738 => x"76",
          4739 => x"05",
          4740 => x"1d",
          4741 => x"f3",
          4742 => x"57",
          4743 => x"82",
          4744 => x"33",
          4745 => x"1e",
          4746 => x"33",
          4747 => x"11",
          4748 => x"90",
          4749 => x"33",
          4750 => x"71",
          4751 => x"96",
          4752 => x"41",
          4753 => x"86",
          4754 => x"33",
          4755 => x"84",
          4756 => x"e5",
          4757 => x"11",
          4758 => x"83",
          4759 => x"51",
          4760 => x"08",
          4761 => x"75",
          4762 => x"b3",
          4763 => x"34",
          4764 => x"58",
          4765 => x"78",
          4766 => x"54",
          4767 => x"74",
          4768 => x"25",
          4769 => x"75",
          4770 => x"78",
          4771 => x"56",
          4772 => x"33",
          4773 => x"88",
          4774 => x"54",
          4775 => x"54",
          4776 => x"08",
          4777 => x"27",
          4778 => x"81",
          4779 => x"a0",
          4780 => x"53",
          4781 => x"81",
          4782 => x"13",
          4783 => x"ff",
          4784 => x"2a",
          4785 => x"80",
          4786 => x"5f",
          4787 => x"63",
          4788 => x"65",
          4789 => x"2e",
          4790 => x"2e",
          4791 => x"d9",
          4792 => x"73",
          4793 => x"55",
          4794 => x"42",
          4795 => x"70",
          4796 => x"73",
          4797 => x"ff",
          4798 => x"74",
          4799 => x"80",
          4800 => x"ff",
          4801 => x"9f",
          4802 => x"5b",
          4803 => x"80",
          4804 => x"ff",
          4805 => x"83",
          4806 => x"56",
          4807 => x"38",
          4808 => x"70",
          4809 => x"56",
          4810 => x"5b",
          4811 => x"26",
          4812 => x"74",
          4813 => x"81",
          4814 => x"80",
          4815 => x"81",
          4816 => x"80",
          4817 => x"72",
          4818 => x"46",
          4819 => x"af",
          4820 => x"70",
          4821 => x"54",
          4822 => x"0c",
          4823 => x"42",
          4824 => x"b4",
          4825 => x"8d",
          4826 => x"ff",
          4827 => x"86",
          4828 => x"3d",
          4829 => x"81",
          4830 => x"fe",
          4831 => x"ab",
          4832 => x"8d",
          4833 => x"c8",
          4834 => x"80",
          4835 => x"73",
          4836 => x"2e",
          4837 => x"70",
          4838 => x"dd",
          4839 => x"70",
          4840 => x"7d",
          4841 => x"27",
          4842 => x"f8",
          4843 => x"76",
          4844 => x"76",
          4845 => x"70",
          4846 => x"52",
          4847 => x"2e",
          4848 => x"57",
          4849 => x"56",
          4850 => x"c7",
          4851 => x"ff",
          4852 => x"a0",
          4853 => x"ff",
          4854 => x"38",
          4855 => x"fe",
          4856 => x"2e",
          4857 => x"54",
          4858 => x"38",
          4859 => x"ae",
          4860 => x"0b",
          4861 => x"81",
          4862 => x"f4",
          4863 => x"16",
          4864 => x"5d",
          4865 => x"a0",
          4866 => x"70",
          4867 => x"75",
          4868 => x"bb",
          4869 => x"38",
          4870 => x"70",
          4871 => x"51",
          4872 => x"e0",
          4873 => x"75",
          4874 => x"5a",
          4875 => x"88",
          4876 => x"06",
          4877 => x"70",
          4878 => x"ff",
          4879 => x"81",
          4880 => x"2e",
          4881 => x"77",
          4882 => x"06",
          4883 => x"79",
          4884 => x"38",
          4885 => x"85",
          4886 => x"2a",
          4887 => x"38",
          4888 => x"34",
          4889 => x"c8",
          4890 => x"b9",
          4891 => x"84",
          4892 => x"06",
          4893 => x"06",
          4894 => x"74",
          4895 => x"98",
          4896 => x"42",
          4897 => x"ce",
          4898 => x"70",
          4899 => x"2e",
          4900 => x"38",
          4901 => x"82",
          4902 => x"81",
          4903 => x"73",
          4904 => x"38",
          4905 => x"80",
          4906 => x"76",
          4907 => x"75",
          4908 => x"53",
          4909 => x"07",
          4910 => x"e3",
          4911 => x"1d",
          4912 => x"fe",
          4913 => x"58",
          4914 => x"70",
          4915 => x"80",
          4916 => x"83",
          4917 => x"33",
          4918 => x"07",
          4919 => x"83",
          4920 => x"0c",
          4921 => x"39",
          4922 => x"f0",
          4923 => x"38",
          4924 => x"17",
          4925 => x"2b",
          4926 => x"5e",
          4927 => x"95",
          4928 => x"39",
          4929 => x"2e",
          4930 => x"39",
          4931 => x"0b",
          4932 => x"04",
          4933 => x"ff",
          4934 => x"59",
          4935 => x"83",
          4936 => x"fc",
          4937 => x"b5",
          4938 => x"84",
          4939 => x"70",
          4940 => x"80",
          4941 => x"83",
          4942 => x"81",
          4943 => x"2e",
          4944 => x"83",
          4945 => x"56",
          4946 => x"38",
          4947 => x"70",
          4948 => x"59",
          4949 => x"59",
          4950 => x"54",
          4951 => x"07",
          4952 => x"9f",
          4953 => x"7d",
          4954 => x"17",
          4955 => x"5f",
          4956 => x"79",
          4957 => x"fa",
          4958 => x"83",
          4959 => x"5a",
          4960 => x"80",
          4961 => x"05",
          4962 => x"1b",
          4963 => x"80",
          4964 => x"90",
          4965 => x"5a",
          4966 => x"05",
          4967 => x"34",
          4968 => x"5b",
          4969 => x"9c",
          4970 => x"58",
          4971 => x"06",
          4972 => x"82",
          4973 => x"38",
          4974 => x"3d",
          4975 => x"02",
          4976 => x"42",
          4977 => x"70",
          4978 => x"d7",
          4979 => x"70",
          4980 => x"85",
          4981 => x"2e",
          4982 => x"56",
          4983 => x"10",
          4984 => x"58",
          4985 => x"96",
          4986 => x"06",
          4987 => x"9b",
          4988 => x"b0",
          4989 => x"06",
          4990 => x"2e",
          4991 => x"16",
          4992 => x"18",
          4993 => x"ff",
          4994 => x"81",
          4995 => x"83",
          4996 => x"2e",
          4997 => x"41",
          4998 => x"5b",
          4999 => x"18",
          5000 => x"7a",
          5001 => x"33",
          5002 => x"b9",
          5003 => x"55",
          5004 => x"56",
          5005 => x"84",
          5006 => x"56",
          5007 => x"2e",
          5008 => x"38",
          5009 => x"85",
          5010 => x"83",
          5011 => x"83",
          5012 => x"c3",
          5013 => x"59",
          5014 => x"83",
          5015 => x"ce",
          5016 => x"5a",
          5017 => x"11",
          5018 => x"71",
          5019 => x"72",
          5020 => x"56",
          5021 => x"a0",
          5022 => x"18",
          5023 => x"70",
          5024 => x"58",
          5025 => x"81",
          5026 => x"19",
          5027 => x"23",
          5028 => x"38",
          5029 => x"bb",
          5030 => x"18",
          5031 => x"74",
          5032 => x"5e",
          5033 => x"80",
          5034 => x"71",
          5035 => x"38",
          5036 => x"12",
          5037 => x"07",
          5038 => x"2b",
          5039 => x"58",
          5040 => x"80",
          5041 => x"5d",
          5042 => x"ce",
          5043 => x"5a",
          5044 => x"52",
          5045 => x"3f",
          5046 => x"c8",
          5047 => x"b9",
          5048 => x"26",
          5049 => x"f5",
          5050 => x"f5",
          5051 => x"16",
          5052 => x"0c",
          5053 => x"1d",
          5054 => x"2e",
          5055 => x"8d",
          5056 => x"7d",
          5057 => x"7c",
          5058 => x"70",
          5059 => x"5a",
          5060 => x"58",
          5061 => x"ff",
          5062 => x"18",
          5063 => x"7c",
          5064 => x"34",
          5065 => x"7c",
          5066 => x"23",
          5067 => x"80",
          5068 => x"84",
          5069 => x"8b",
          5070 => x"0d",
          5071 => x"ff",
          5072 => x"91",
          5073 => x"d0",
          5074 => x"fe",
          5075 => x"5f",
          5076 => x"7a",
          5077 => x"81",
          5078 => x"58",
          5079 => x"16",
          5080 => x"9f",
          5081 => x"e0",
          5082 => x"75",
          5083 => x"77",
          5084 => x"ff",
          5085 => x"70",
          5086 => x"58",
          5087 => x"81",
          5088 => x"25",
          5089 => x"39",
          5090 => x"82",
          5091 => x"fe",
          5092 => x"7a",
          5093 => x"2e",
          5094 => x"75",
          5095 => x"25",
          5096 => x"ad",
          5097 => x"38",
          5098 => x"83",
          5099 => x"80",
          5100 => x"84",
          5101 => x"88",
          5102 => x"72",
          5103 => x"71",
          5104 => x"77",
          5105 => x"19",
          5106 => x"ff",
          5107 => x"70",
          5108 => x"9b",
          5109 => x"84",
          5110 => x"42",
          5111 => x"2e",
          5112 => x"34",
          5113 => x"80",
          5114 => x"54",
          5115 => x"33",
          5116 => x"c8",
          5117 => x"81",
          5118 => x"75",
          5119 => x"71",
          5120 => x"7b",
          5121 => x"a8",
          5122 => x"58",
          5123 => x"75",
          5124 => x"25",
          5125 => x"38",
          5126 => x"58",
          5127 => x"84",
          5128 => x"78",
          5129 => x"58",
          5130 => x"80",
          5131 => x"1a",
          5132 => x"38",
          5133 => x"18",
          5134 => x"70",
          5135 => x"05",
          5136 => x"5b",
          5137 => x"c5",
          5138 => x"0b",
          5139 => x"5d",
          5140 => x"7e",
          5141 => x"31",
          5142 => x"80",
          5143 => x"e1",
          5144 => x"58",
          5145 => x"c8",
          5146 => x"75",
          5147 => x"81",
          5148 => x"58",
          5149 => x"c8",
          5150 => x"80",
          5151 => x"58",
          5152 => x"70",
          5153 => x"ff",
          5154 => x"2e",
          5155 => x"38",
          5156 => x"fc",
          5157 => x"5a",
          5158 => x"71",
          5159 => x"40",
          5160 => x"80",
          5161 => x"5a",
          5162 => x"fd",
          5163 => x"e8",
          5164 => x"55",
          5165 => x"d5",
          5166 => x"17",
          5167 => x"33",
          5168 => x"82",
          5169 => x"17",
          5170 => x"d2",
          5171 => x"85",
          5172 => x"18",
          5173 => x"18",
          5174 => x"18",
          5175 => x"75",
          5176 => x"f8",
          5177 => x"82",
          5178 => x"2b",
          5179 => x"88",
          5180 => x"59",
          5181 => x"85",
          5182 => x"cd",
          5183 => x"82",
          5184 => x"2b",
          5185 => x"88",
          5186 => x"40",
          5187 => x"85",
          5188 => x"9d",
          5189 => x"82",
          5190 => x"2b",
          5191 => x"88",
          5192 => x"0c",
          5193 => x"82",
          5194 => x"2b",
          5195 => x"88",
          5196 => x"05",
          5197 => x"40",
          5198 => x"84",
          5199 => x"84",
          5200 => x"84",
          5201 => x"0b",
          5202 => x"83",
          5203 => x"0c",
          5204 => x"17",
          5205 => x"18",
          5206 => x"84",
          5207 => x"06",
          5208 => x"83",
          5209 => x"08",
          5210 => x"8b",
          5211 => x"2e",
          5212 => x"5a",
          5213 => x"2e",
          5214 => x"18",
          5215 => x"ab",
          5216 => x"18",
          5217 => x"8d",
          5218 => x"22",
          5219 => x"17",
          5220 => x"90",
          5221 => x"33",
          5222 => x"71",
          5223 => x"2b",
          5224 => x"d8",
          5225 => x"e8",
          5226 => x"80",
          5227 => x"57",
          5228 => x"5a",
          5229 => x"75",
          5230 => x"05",
          5231 => x"ff",
          5232 => x"3d",
          5233 => x"70",
          5234 => x"76",
          5235 => x"38",
          5236 => x"9f",
          5237 => x"e2",
          5238 => x"80",
          5239 => x"80",
          5240 => x"10",
          5241 => x"55",
          5242 => x"34",
          5243 => x"80",
          5244 => x"7c",
          5245 => x"53",
          5246 => x"ef",
          5247 => x"73",
          5248 => x"04",
          5249 => x"3d",
          5250 => x"81",
          5251 => x"26",
          5252 => x"06",
          5253 => x"80",
          5254 => x"b8",
          5255 => x"5a",
          5256 => x"70",
          5257 => x"59",
          5258 => x"e0",
          5259 => x"ff",
          5260 => x"38",
          5261 => x"54",
          5262 => x"74",
          5263 => x"76",
          5264 => x"30",
          5265 => x"5c",
          5266 => x"81",
          5267 => x"25",
          5268 => x"39",
          5269 => x"60",
          5270 => x"0d",
          5271 => x"33",
          5272 => x"a6",
          5273 => x"3d",
          5274 => x"52",
          5275 => x"08",
          5276 => x"8f",
          5277 => x"84",
          5278 => x"7e",
          5279 => x"5a",
          5280 => x"57",
          5281 => x"ba",
          5282 => x"2e",
          5283 => x"c1",
          5284 => x"77",
          5285 => x"77",
          5286 => x"2e",
          5287 => x"9a",
          5288 => x"70",
          5289 => x"83",
          5290 => x"17",
          5291 => x"0b",
          5292 => x"17",
          5293 => x"34",
          5294 => x"17",
          5295 => x"33",
          5296 => x"66",
          5297 => x"0b",
          5298 => x"34",
          5299 => x"81",
          5300 => x"80",
          5301 => x"7c",
          5302 => x"27",
          5303 => x"83",
          5304 => x"fe",
          5305 => x"70",
          5306 => x"fe",
          5307 => x"57",
          5308 => x"38",
          5309 => x"2a",
          5310 => x"38",
          5311 => x"80",
          5312 => x"79",
          5313 => x"06",
          5314 => x"80",
          5315 => x"a0",
          5316 => x"9b",
          5317 => x"2b",
          5318 => x"5a",
          5319 => x"88",
          5320 => x"82",
          5321 => x"2b",
          5322 => x"88",
          5323 => x"8c",
          5324 => x"41",
          5325 => x"84",
          5326 => x"0b",
          5327 => x"0c",
          5328 => x"80",
          5329 => x"84",
          5330 => x"1a",
          5331 => x"58",
          5332 => x"56",
          5333 => x"81",
          5334 => x"2e",
          5335 => x"ff",
          5336 => x"58",
          5337 => x"38",
          5338 => x"2e",
          5339 => x"c0",
          5340 => x"06",
          5341 => x"81",
          5342 => x"38",
          5343 => x"39",
          5344 => x"39",
          5345 => x"39",
          5346 => x"c8",
          5347 => x"fb",
          5348 => x"7b",
          5349 => x"16",
          5350 => x"71",
          5351 => x"5c",
          5352 => x"27",
          5353 => x"ff",
          5354 => x"5d",
          5355 => x"a7",
          5356 => x"fc",
          5357 => x"2e",
          5358 => x"76",
          5359 => x"c8",
          5360 => x"fe",
          5361 => x"75",
          5362 => x"94",
          5363 => x"55",
          5364 => x"7d",
          5365 => x"80",
          5366 => x"17",
          5367 => x"94",
          5368 => x"2b",
          5369 => x"0b",
          5370 => x"34",
          5371 => x"0b",
          5372 => x"8b",
          5373 => x"0b",
          5374 => x"34",
          5375 => x"81",
          5376 => x"80",
          5377 => x"b4",
          5378 => x"16",
          5379 => x"06",
          5380 => x"16",
          5381 => x"ba",
          5382 => x"85",
          5383 => x"17",
          5384 => x"18",
          5385 => x"38",
          5386 => x"54",
          5387 => x"53",
          5388 => x"81",
          5389 => x"09",
          5390 => x"c8",
          5391 => x"a8",
          5392 => x"5c",
          5393 => x"92",
          5394 => x"2e",
          5395 => x"54",
          5396 => x"53",
          5397 => x"a3",
          5398 => x"74",
          5399 => x"39",
          5400 => x"38",
          5401 => x"2e",
          5402 => x"12",
          5403 => x"7d",
          5404 => x"78",
          5405 => x"5c",
          5406 => x"89",
          5407 => x"f7",
          5408 => x"56",
          5409 => x"0c",
          5410 => x"57",
          5411 => x"7f",
          5412 => x"0d",
          5413 => x"5a",
          5414 => x"2e",
          5415 => x"2e",
          5416 => x"2e",
          5417 => x"22",
          5418 => x"38",
          5419 => x"82",
          5420 => x"82",
          5421 => x"57",
          5422 => x"38",
          5423 => x"31",
          5424 => x"38",
          5425 => x"59",
          5426 => x"e3",
          5427 => x"89",
          5428 => x"83",
          5429 => x"75",
          5430 => x"83",
          5431 => x"59",
          5432 => x"08",
          5433 => x"83",
          5434 => x"29",
          5435 => x"80",
          5436 => x"89",
          5437 => x"81",
          5438 => x"85",
          5439 => x"76",
          5440 => x"ff",
          5441 => x"83",
          5442 => x"59",
          5443 => x"08",
          5444 => x"38",
          5445 => x"1b",
          5446 => x"57",
          5447 => x"ff",
          5448 => x"2b",
          5449 => x"7f",
          5450 => x"70",
          5451 => x"fe",
          5452 => x"c8",
          5453 => x"b9",
          5454 => x"5c",
          5455 => x"75",
          5456 => x"59",
          5457 => x"58",
          5458 => x"b6",
          5459 => x"5d",
          5460 => x"06",
          5461 => x"b8",
          5462 => x"9e",
          5463 => x"2e",
          5464 => x"b4",
          5465 => x"94",
          5466 => x"7f",
          5467 => x"80",
          5468 => x"05",
          5469 => x"34",
          5470 => x"d1",
          5471 => x"77",
          5472 => x"56",
          5473 => x"54",
          5474 => x"53",
          5475 => x"c9",
          5476 => x"7f",
          5477 => x"84",
          5478 => x"19",
          5479 => x"c8",
          5480 => x"27",
          5481 => x"74",
          5482 => x"38",
          5483 => x"08",
          5484 => x"51",
          5485 => x"bb",
          5486 => x"08",
          5487 => x"52",
          5488 => x"b9",
          5489 => x"16",
          5490 => x"b9",
          5491 => x"b8",
          5492 => x"b2",
          5493 => x"0b",
          5494 => x"04",
          5495 => x"84",
          5496 => x"f0",
          5497 => x"40",
          5498 => x"79",
          5499 => x"75",
          5500 => x"74",
          5501 => x"84",
          5502 => x"85",
          5503 => x"55",
          5504 => x"55",
          5505 => x"70",
          5506 => x"56",
          5507 => x"1a",
          5508 => x"27",
          5509 => x"2e",
          5510 => x"5f",
          5511 => x"22",
          5512 => x"56",
          5513 => x"88",
          5514 => x"b1",
          5515 => x"74",
          5516 => x"1b",
          5517 => x"88",
          5518 => x"9c",
          5519 => x"1a",
          5520 => x"05",
          5521 => x"38",
          5522 => x"18",
          5523 => x"85",
          5524 => x"59",
          5525 => x"77",
          5526 => x"76",
          5527 => x"7c",
          5528 => x"a1",
          5529 => x"38",
          5530 => x"57",
          5531 => x"0b",
          5532 => x"58",
          5533 => x"77",
          5534 => x"56",
          5535 => x"1a",
          5536 => x"31",
          5537 => x"94",
          5538 => x"0c",
          5539 => x"5b",
          5540 => x"75",
          5541 => x"90",
          5542 => x"5b",
          5543 => x"84",
          5544 => x"74",
          5545 => x"04",
          5546 => x"38",
          5547 => x"1b",
          5548 => x"84",
          5549 => x"27",
          5550 => x"16",
          5551 => x"83",
          5552 => x"7f",
          5553 => x"81",
          5554 => x"16",
          5555 => x"b9",
          5556 => x"57",
          5557 => x"83",
          5558 => x"ff",
          5559 => x"59",
          5560 => x"76",
          5561 => x"81",
          5562 => x"ef",
          5563 => x"34",
          5564 => x"08",
          5565 => x"33",
          5566 => x"5c",
          5567 => x"81",
          5568 => x"08",
          5569 => x"17",
          5570 => x"55",
          5571 => x"38",
          5572 => x"09",
          5573 => x"b4",
          5574 => x"7f",
          5575 => x"a9",
          5576 => x"1a",
          5577 => x"93",
          5578 => x"b9",
          5579 => x"1b",
          5580 => x"0c",
          5581 => x"52",
          5582 => x"b9",
          5583 => x"fb",
          5584 => x"ab",
          5585 => x"cc",
          5586 => x"b9",
          5587 => x"81",
          5588 => x"70",
          5589 => x"97",
          5590 => x"b8",
          5591 => x"34",
          5592 => x"58",
          5593 => x"38",
          5594 => x"09",
          5595 => x"b4",
          5596 => x"76",
          5597 => x"f9",
          5598 => x"16",
          5599 => x"b9",
          5600 => x"f2",
          5601 => x"ec",
          5602 => x"b8",
          5603 => x"57",
          5604 => x"08",
          5605 => x"83",
          5606 => x"08",
          5607 => x"fe",
          5608 => x"82",
          5609 => x"81",
          5610 => x"05",
          5611 => x"ff",
          5612 => x"0c",
          5613 => x"39",
          5614 => x"84",
          5615 => x"82",
          5616 => x"b9",
          5617 => x"3d",
          5618 => x"2e",
          5619 => x"2e",
          5620 => x"2e",
          5621 => x"22",
          5622 => x"38",
          5623 => x"81",
          5624 => x"2a",
          5625 => x"81",
          5626 => x"57",
          5627 => x"83",
          5628 => x"81",
          5629 => x"17",
          5630 => x"b9",
          5631 => x"59",
          5632 => x"81",
          5633 => x"33",
          5634 => x"34",
          5635 => x"ff",
          5636 => x"18",
          5637 => x"18",
          5638 => x"5c",
          5639 => x"38",
          5640 => x"74",
          5641 => x"74",
          5642 => x"74",
          5643 => x"80",
          5644 => x"a1",
          5645 => x"99",
          5646 => x"80",
          5647 => x"0b",
          5648 => x"94",
          5649 => x"33",
          5650 => x"19",
          5651 => x"3d",
          5652 => x"53",
          5653 => x"52",
          5654 => x"84",
          5655 => x"b9",
          5656 => x"08",
          5657 => x"08",
          5658 => x"fe",
          5659 => x"82",
          5660 => x"81",
          5661 => x"05",
          5662 => x"ff",
          5663 => x"39",
          5664 => x"34",
          5665 => x"34",
          5666 => x"74",
          5667 => x"74",
          5668 => x"74",
          5669 => x"80",
          5670 => x"a1",
          5671 => x"99",
          5672 => x"80",
          5673 => x"0b",
          5674 => x"c4",
          5675 => x"33",
          5676 => x"19",
          5677 => x"51",
          5678 => x"08",
          5679 => x"74",
          5680 => x"f9",
          5681 => x"fe",
          5682 => x"b9",
          5683 => x"80",
          5684 => x"80",
          5685 => x"80",
          5686 => x"16",
          5687 => x"38",
          5688 => x"84",
          5689 => x"c8",
          5690 => x"33",
          5691 => x"c8",
          5692 => x"73",
          5693 => x"3d",
          5694 => x"75",
          5695 => x"05",
          5696 => x"71",
          5697 => x"71",
          5698 => x"33",
          5699 => x"84",
          5700 => x"c8",
          5701 => x"84",
          5702 => x"78",
          5703 => x"53",
          5704 => x"82",
          5705 => x"59",
          5706 => x"80",
          5707 => x"08",
          5708 => x"58",
          5709 => x"ff",
          5710 => x"26",
          5711 => x"06",
          5712 => x"99",
          5713 => x"ff",
          5714 => x"2a",
          5715 => x"06",
          5716 => x"76",
          5717 => x"2a",
          5718 => x"2e",
          5719 => x"58",
          5720 => x"51",
          5721 => x"38",
          5722 => x"ea",
          5723 => x"05",
          5724 => x"84",
          5725 => x"08",
          5726 => x"c8",
          5727 => x"68",
          5728 => x"94",
          5729 => x"b9",
          5730 => x"d7",
          5731 => x"80",
          5732 => x"05",
          5733 => x"59",
          5734 => x"9b",
          5735 => x"2b",
          5736 => x"58",
          5737 => x"19",
          5738 => x"3d",
          5739 => x"2e",
          5740 => x"0b",
          5741 => x"04",
          5742 => x"98",
          5743 => x"98",
          5744 => x"7e",
          5745 => x"c8",
          5746 => x"3d",
          5747 => x"3d",
          5748 => x"53",
          5749 => x"80",
          5750 => x"b9",
          5751 => x"83",
          5752 => x"7f",
          5753 => x"0c",
          5754 => x"79",
          5755 => x"3d",
          5756 => x"51",
          5757 => x"08",
          5758 => x"38",
          5759 => x"b4",
          5760 => x"b9",
          5761 => x"7d",
          5762 => x"b8",
          5763 => x"8b",
          5764 => x"2e",
          5765 => x"b4",
          5766 => x"df",
          5767 => x"33",
          5768 => x"5d",
          5769 => x"82",
          5770 => x"80",
          5771 => x"84",
          5772 => x"08",
          5773 => x"ff",
          5774 => x"59",
          5775 => x"df",
          5776 => x"33",
          5777 => x"42",
          5778 => x"81",
          5779 => x"84",
          5780 => x"a4",
          5781 => x"84",
          5782 => x"38",
          5783 => x"81",
          5784 => x"05",
          5785 => x"78",
          5786 => x"80",
          5787 => x"17",
          5788 => x"7c",
          5789 => x"26",
          5790 => x"38",
          5791 => x"80",
          5792 => x"19",
          5793 => x"34",
          5794 => x"3d",
          5795 => x"80",
          5796 => x"38",
          5797 => x"0b",
          5798 => x"83",
          5799 => x"43",
          5800 => x"8d",
          5801 => x"57",
          5802 => x"5b",
          5803 => x"76",
          5804 => x"7e",
          5805 => x"81",
          5806 => x"ba",
          5807 => x"ff",
          5808 => x"91",
          5809 => x"c8",
          5810 => x"16",
          5811 => x"71",
          5812 => x"5e",
          5813 => x"17",
          5814 => x"07",
          5815 => x"5d",
          5816 => x"3f",
          5817 => x"c8",
          5818 => x"b1",
          5819 => x"b8",
          5820 => x"5e",
          5821 => x"b9",
          5822 => x"c8",
          5823 => x"a8",
          5824 => x"5a",
          5825 => x"83",
          5826 => x"2e",
          5827 => x"54",
          5828 => x"53",
          5829 => x"88",
          5830 => x"ff",
          5831 => x"58",
          5832 => x"a4",
          5833 => x"05",
          5834 => x"5e",
          5835 => x"fd",
          5836 => x"3d",
          5837 => x"33",
          5838 => x"60",
          5839 => x"08",
          5840 => x"7c",
          5841 => x"26",
          5842 => x"80",
          5843 => x"80",
          5844 => x"7b",
          5845 => x"2e",
          5846 => x"2e",
          5847 => x"2e",
          5848 => x"22",
          5849 => x"38",
          5850 => x"81",
          5851 => x"81",
          5852 => x"76",
          5853 => x"54",
          5854 => x"38",
          5855 => x"52",
          5856 => x"38",
          5857 => x"9c",
          5858 => x"77",
          5859 => x"8c",
          5860 => x"81",
          5861 => x"94",
          5862 => x"08",
          5863 => x"98",
          5864 => x"76",
          5865 => x"17",
          5866 => x"81",
          5867 => x"81",
          5868 => x"99",
          5869 => x"84",
          5870 => x"38",
          5871 => x"27",
          5872 => x"14",
          5873 => x"16",
          5874 => x"16",
          5875 => x"0c",
          5876 => x"70",
          5877 => x"fe",
          5878 => x"57",
          5879 => x"06",
          5880 => x"94",
          5881 => x"38",
          5882 => x"80",
          5883 => x"73",
          5884 => x"8c",
          5885 => x"38",
          5886 => x"b9",
          5887 => x"0b",
          5888 => x"73",
          5889 => x"16",
          5890 => x"fe",
          5891 => x"94",
          5892 => x"83",
          5893 => x"38",
          5894 => x"05",
          5895 => x"f6",
          5896 => x"b0",
          5897 => x"5a",
          5898 => x"38",
          5899 => x"73",
          5900 => x"84",
          5901 => x"81",
          5902 => x"84",
          5903 => x"fc",
          5904 => x"fc",
          5905 => x"97",
          5906 => x"84",
          5907 => x"84",
          5908 => x"38",
          5909 => x"73",
          5910 => x"0b",
          5911 => x"c8",
          5912 => x"0d",
          5913 => x"a2",
          5914 => x"52",
          5915 => x"3f",
          5916 => x"c8",
          5917 => x"0c",
          5918 => x"8c",
          5919 => x"52",
          5920 => x"b9",
          5921 => x"80",
          5922 => x"2b",
          5923 => x"86",
          5924 => x"5b",
          5925 => x"9c",
          5926 => x"33",
          5927 => x"5d",
          5928 => x"b3",
          5929 => x"86",
          5930 => x"75",
          5931 => x"c8",
          5932 => x"74",
          5933 => x"0c",
          5934 => x"0c",
          5935 => x"18",
          5936 => x"07",
          5937 => x"ff",
          5938 => x"89",
          5939 => x"08",
          5940 => x"33",
          5941 => x"13",
          5942 => x"76",
          5943 => x"73",
          5944 => x"b9",
          5945 => x"13",
          5946 => x"b9",
          5947 => x"38",
          5948 => x"f8",
          5949 => x"56",
          5950 => x"54",
          5951 => x"53",
          5952 => x"22",
          5953 => x"2e",
          5954 => x"75",
          5955 => x"2e",
          5956 => x"ff",
          5957 => x"53",
          5958 => x"38",
          5959 => x"52",
          5960 => x"52",
          5961 => x"b9",
          5962 => x"72",
          5963 => x"06",
          5964 => x"0c",
          5965 => x"75",
          5966 => x"52",
          5967 => x"b9",
          5968 => x"72",
          5969 => x"06",
          5970 => x"74",
          5971 => x"c8",
          5972 => x"0d",
          5973 => x"e8",
          5974 => x"53",
          5975 => x"54",
          5976 => x"66",
          5977 => x"97",
          5978 => x"b9",
          5979 => x"80",
          5980 => x"0c",
          5981 => x"51",
          5982 => x"08",
          5983 => x"02",
          5984 => x"55",
          5985 => x"80",
          5986 => x"ff",
          5987 => x"0c",
          5988 => x"b9",
          5989 => x"3d",
          5990 => x"95",
          5991 => x"c0",
          5992 => x"84",
          5993 => x"0c",
          5994 => x"94",
          5995 => x"75",
          5996 => x"84",
          5997 => x"84",
          5998 => x"78",
          5999 => x"18",
          6000 => x"59",
          6001 => x"71",
          6002 => x"2e",
          6003 => x"5f",
          6004 => x"75",
          6005 => x"51",
          6006 => x"08",
          6007 => x"5e",
          6008 => x"57",
          6009 => x"7d",
          6010 => x"b8",
          6011 => x"71",
          6012 => x"14",
          6013 => x"33",
          6014 => x"07",
          6015 => x"60",
          6016 => x"05",
          6017 => x"58",
          6018 => x"7a",
          6019 => x"17",
          6020 => x"34",
          6021 => x"0d",
          6022 => x"b8",
          6023 => x"5d",
          6024 => x"b9",
          6025 => x"c8",
          6026 => x"a8",
          6027 => x"5f",
          6028 => x"bd",
          6029 => x"2e",
          6030 => x"54",
          6031 => x"53",
          6032 => x"fb",
          6033 => x"82",
          6034 => x"52",
          6035 => x"b9",
          6036 => x"84",
          6037 => x"38",
          6038 => x"b9",
          6039 => x"81",
          6040 => x"17",
          6041 => x"0c",
          6042 => x"81",
          6043 => x"c8",
          6044 => x"33",
          6045 => x"30",
          6046 => x"ff",
          6047 => x"5f",
          6048 => x"8f",
          6049 => x"60",
          6050 => x"18",
          6051 => x"77",
          6052 => x"60",
          6053 => x"7b",
          6054 => x"38",
          6055 => x"38",
          6056 => x"38",
          6057 => x"59",
          6058 => x"54",
          6059 => x"17",
          6060 => x"17",
          6061 => x"58",
          6062 => x"38",
          6063 => x"08",
          6064 => x"88",
          6065 => x"74",
          6066 => x"26",
          6067 => x"18",
          6068 => x"77",
          6069 => x"34",
          6070 => x"18",
          6071 => x"0c",
          6072 => x"78",
          6073 => x"51",
          6074 => x"08",
          6075 => x"80",
          6076 => x"2e",
          6077 => x"ff",
          6078 => x"52",
          6079 => x"b9",
          6080 => x"08",
          6081 => x"58",
          6082 => x"15",
          6083 => x"07",
          6084 => x"77",
          6085 => x"81",
          6086 => x"84",
          6087 => x"fe",
          6088 => x"fe",
          6089 => x"59",
          6090 => x"0c",
          6091 => x"76",
          6092 => x"c8",
          6093 => x"b9",
          6094 => x"75",
          6095 => x"c8",
          6096 => x"38",
          6097 => x"78",
          6098 => x"b9",
          6099 => x"b9",
          6100 => x"96",
          6101 => x"53",
          6102 => x"3f",
          6103 => x"c8",
          6104 => x"51",
          6105 => x"08",
          6106 => x"80",
          6107 => x"2e",
          6108 => x"ff",
          6109 => x"52",
          6110 => x"b9",
          6111 => x"08",
          6112 => x"58",
          6113 => x"94",
          6114 => x"54",
          6115 => x"79",
          6116 => x"56",
          6117 => x"81",
          6118 => x"18",
          6119 => x"56",
          6120 => x"59",
          6121 => x"08",
          6122 => x"39",
          6123 => x"fd",
          6124 => x"c0",
          6125 => x"3d",
          6126 => x"05",
          6127 => x"3f",
          6128 => x"c8",
          6129 => x"b9",
          6130 => x"4b",
          6131 => x"52",
          6132 => x"c8",
          6133 => x"38",
          6134 => x"2a",
          6135 => x"cd",
          6136 => x"24",
          6137 => x"70",
          6138 => x"ff",
          6139 => x"11",
          6140 => x"07",
          6141 => x"7c",
          6142 => x"2a",
          6143 => x"ed",
          6144 => x"2e",
          6145 => x"84",
          6146 => x"52",
          6147 => x"c8",
          6148 => x"e5",
          6149 => x"51",
          6150 => x"08",
          6151 => x"87",
          6152 => x"0d",
          6153 => x"71",
          6154 => x"07",
          6155 => x"b9",
          6156 => x"b9",
          6157 => x"6f",
          6158 => x"ff",
          6159 => x"51",
          6160 => x"08",
          6161 => x"be",
          6162 => x"25",
          6163 => x"74",
          6164 => x"58",
          6165 => x"17",
          6166 => x"56",
          6167 => x"f5",
          6168 => x"b9",
          6169 => x"17",
          6170 => x"b4",
          6171 => x"83",
          6172 => x"2e",
          6173 => x"54",
          6174 => x"33",
          6175 => x"c8",
          6176 => x"81",
          6177 => x"77",
          6178 => x"78",
          6179 => x"19",
          6180 => x"52",
          6181 => x"b9",
          6182 => x"80",
          6183 => x"09",
          6184 => x"fe",
          6185 => x"53",
          6186 => x"f2",
          6187 => x"08",
          6188 => x"38",
          6189 => x"b4",
          6190 => x"b9",
          6191 => x"08",
          6192 => x"55",
          6193 => x"de",
          6194 => x"18",
          6195 => x"33",
          6196 => x"fe",
          6197 => x"80",
          6198 => x"f6",
          6199 => x"84",
          6200 => x"38",
          6201 => x"e6",
          6202 => x"80",
          6203 => x"51",
          6204 => x"08",
          6205 => x"94",
          6206 => x"27",
          6207 => x"0c",
          6208 => x"84",
          6209 => x"ff",
          6210 => x"79",
          6211 => x"08",
          6212 => x"90",
          6213 => x"3d",
          6214 => x"ff",
          6215 => x"56",
          6216 => x"38",
          6217 => x"0d",
          6218 => x"70",
          6219 => x"b9",
          6220 => x"8b",
          6221 => x"9f",
          6222 => x"84",
          6223 => x"80",
          6224 => x"06",
          6225 => x"38",
          6226 => x"52",
          6227 => x"c8",
          6228 => x"08",
          6229 => x"08",
          6230 => x"c8",
          6231 => x"81",
          6232 => x"83",
          6233 => x"e2",
          6234 => x"05",
          6235 => x"8d",
          6236 => x"b0",
          6237 => x"18",
          6238 => x"57",
          6239 => x"34",
          6240 => x"58",
          6241 => x"81",
          6242 => x"78",
          6243 => x"c9",
          6244 => x"38",
          6245 => x"ff",
          6246 => x"53",
          6247 => x"52",
          6248 => x"84",
          6249 => x"c8",
          6250 => x"a8",
          6251 => x"08",
          6252 => x"5b",
          6253 => x"e1",
          6254 => x"18",
          6255 => x"33",
          6256 => x"39",
          6257 => x"81",
          6258 => x"18",
          6259 => x"7c",
          6260 => x"c8",
          6261 => x"2e",
          6262 => x"81",
          6263 => x"08",
          6264 => x"74",
          6265 => x"84",
          6266 => x"17",
          6267 => x"5c",
          6268 => x"18",
          6269 => x"07",
          6270 => x"78",
          6271 => x"b9",
          6272 => x"17",
          6273 => x"57",
          6274 => x"06",
          6275 => x"56",
          6276 => x"34",
          6277 => x"57",
          6278 => x"90",
          6279 => x"75",
          6280 => x"1a",
          6281 => x"80",
          6282 => x"7c",
          6283 => x"80",
          6284 => x"7a",
          6285 => x"74",
          6286 => x"a0",
          6287 => x"58",
          6288 => x"77",
          6289 => x"56",
          6290 => x"80",
          6291 => x"ff",
          6292 => x"f2",
          6293 => x"80",
          6294 => x"83",
          6295 => x"0b",
          6296 => x"96",
          6297 => x"b9",
          6298 => x"84",
          6299 => x"b9",
          6300 => x"98",
          6301 => x"34",
          6302 => x"34",
          6303 => x"34",
          6304 => x"d9",
          6305 => x"34",
          6306 => x"7d",
          6307 => x"c8",
          6308 => x"9f",
          6309 => x"74",
          6310 => x"57",
          6311 => x"39",
          6312 => x"17",
          6313 => x"cd",
          6314 => x"d8",
          6315 => x"a1",
          6316 => x"18",
          6317 => x"18",
          6318 => x"34",
          6319 => x"7d",
          6320 => x"c8",
          6321 => x"0d",
          6322 => x"5b",
          6323 => x"70",
          6324 => x"56",
          6325 => x"74",
          6326 => x"38",
          6327 => x"52",
          6328 => x"84",
          6329 => x"08",
          6330 => x"c8",
          6331 => x"3d",
          6332 => x"70",
          6333 => x"b9",
          6334 => x"dc",
          6335 => x"a0",
          6336 => x"a0",
          6337 => x"58",
          6338 => x"77",
          6339 => x"55",
          6340 => x"78",
          6341 => x"05",
          6342 => x"34",
          6343 => x"3d",
          6344 => x"3f",
          6345 => x"c8",
          6346 => x"08",
          6347 => x"b9",
          6348 => x"33",
          6349 => x"57",
          6350 => x"17",
          6351 => x"59",
          6352 => x"7f",
          6353 => x"5d",
          6354 => x"05",
          6355 => x"33",
          6356 => x"99",
          6357 => x"ff",
          6358 => x"77",
          6359 => x"81",
          6360 => x"9f",
          6361 => x"81",
          6362 => x"78",
          6363 => x"9f",
          6364 => x"80",
          6365 => x"5e",
          6366 => x"7c",
          6367 => x"7b",
          6368 => x"0c",
          6369 => x"52",
          6370 => x"84",
          6371 => x"08",
          6372 => x"aa",
          6373 => x"ac",
          6374 => x"84",
          6375 => x"08",
          6376 => x"8d",
          6377 => x"58",
          6378 => x"33",
          6379 => x"1a",
          6380 => x"05",
          6381 => x"70",
          6382 => x"89",
          6383 => x"19",
          6384 => x"34",
          6385 => x"06",
          6386 => x"38",
          6387 => x"38",
          6388 => x"71",
          6389 => x"5c",
          6390 => x"fe",
          6391 => x"56",
          6392 => x"17",
          6393 => x"05",
          6394 => x"38",
          6395 => x"76",
          6396 => x"7e",
          6397 => x"b8",
          6398 => x"e3",
          6399 => x"2e",
          6400 => x"b4",
          6401 => x"18",
          6402 => x"15",
          6403 => x"06",
          6404 => x"06",
          6405 => x"7b",
          6406 => x"34",
          6407 => x"81",
          6408 => x"7d",
          6409 => x"56",
          6410 => x"81",
          6411 => x"3d",
          6412 => x"74",
          6413 => x"51",
          6414 => x"08",
          6415 => x"38",
          6416 => x"80",
          6417 => x"38",
          6418 => x"7a",
          6419 => x"81",
          6420 => x"16",
          6421 => x"b9",
          6422 => x"57",
          6423 => x"55",
          6424 => x"e5",
          6425 => x"90",
          6426 => x"52",
          6427 => x"b9",
          6428 => x"80",
          6429 => x"84",
          6430 => x"f9",
          6431 => x"3f",
          6432 => x"0c",
          6433 => x"b9",
          6434 => x"18",
          6435 => x"71",
          6436 => x"5c",
          6437 => x"84",
          6438 => x"08",
          6439 => x"b9",
          6440 => x"54",
          6441 => x"16",
          6442 => x"58",
          6443 => x"81",
          6444 => x"08",
          6445 => x"17",
          6446 => x"55",
          6447 => x"38",
          6448 => x"09",
          6449 => x"b4",
          6450 => x"7b",
          6451 => x"c9",
          6452 => x"54",
          6453 => x"53",
          6454 => x"b1",
          6455 => x"fc",
          6456 => x"18",
          6457 => x"31",
          6458 => x"a0",
          6459 => x"17",
          6460 => x"06",
          6461 => x"08",
          6462 => x"81",
          6463 => x"79",
          6464 => x"02",
          6465 => x"80",
          6466 => x"96",
          6467 => x"ff",
          6468 => x"56",
          6469 => x"38",
          6470 => x"0d",
          6471 => x"d0",
          6472 => x"b9",
          6473 => x"e0",
          6474 => x"a0",
          6475 => x"74",
          6476 => x"33",
          6477 => x"56",
          6478 => x"55",
          6479 => x"fe",
          6480 => x"84",
          6481 => x"ec",
          6482 => x"3d",
          6483 => x"a1",
          6484 => x"84",
          6485 => x"74",
          6486 => x"04",
          6487 => x"05",
          6488 => x"c8",
          6489 => x"38",
          6490 => x"06",
          6491 => x"84",
          6492 => x"2b",
          6493 => x"34",
          6494 => x"34",
          6495 => x"34",
          6496 => x"34",
          6497 => x"78",
          6498 => x"c8",
          6499 => x"0d",
          6500 => x"5b",
          6501 => x"9b",
          6502 => x"b9",
          6503 => x"70",
          6504 => x"51",
          6505 => x"81",
          6506 => x"a4",
          6507 => x"25",
          6508 => x"38",
          6509 => x"80",
          6510 => x"08",
          6511 => x"77",
          6512 => x"7a",
          6513 => x"06",
          6514 => x"b8",
          6515 => x"dc",
          6516 => x"2e",
          6517 => x"b4",
          6518 => x"7c",
          6519 => x"74",
          6520 => x"74",
          6521 => x"18",
          6522 => x"33",
          6523 => x"81",
          6524 => x"75",
          6525 => x"5e",
          6526 => x"0c",
          6527 => x"40",
          6528 => x"fe",
          6529 => x"57",
          6530 => x"8d",
          6531 => x"fe",
          6532 => x"fe",
          6533 => x"53",
          6534 => x"52",
          6535 => x"84",
          6536 => x"06",
          6537 => x"83",
          6538 => x"08",
          6539 => x"74",
          6540 => x"82",
          6541 => x"81",
          6542 => x"16",
          6543 => x"52",
          6544 => x"3f",
          6545 => x"16",
          6546 => x"d2",
          6547 => x"fe",
          6548 => x"74",
          6549 => x"c8",
          6550 => x"e1",
          6551 => x"c8",
          6552 => x"81",
          6553 => x"33",
          6554 => x"27",
          6555 => x"80",
          6556 => x"38",
          6557 => x"57",
          6558 => x"e1",
          6559 => x"3d",
          6560 => x"05",
          6561 => x"3f",
          6562 => x"c8",
          6563 => x"8b",
          6564 => x"05",
          6565 => x"38",
          6566 => x"81",
          6567 => x"78",
          6568 => x"3d",
          6569 => x"18",
          6570 => x"7c",
          6571 => x"ff",
          6572 => x"b5",
          6573 => x"dc",
          6574 => x"ff",
          6575 => x"38",
          6576 => x"33",
          6577 => x"78",
          6578 => x"78",
          6579 => x"33",
          6580 => x"74",
          6581 => x"09",
          6582 => x"06",
          6583 => x"77",
          6584 => x"81",
          6585 => x"38",
          6586 => x"81",
          6587 => x"7b",
          6588 => x"a3",
          6589 => x"06",
          6590 => x"fe",
          6591 => x"56",
          6592 => x"80",
          6593 => x"79",
          6594 => x"2e",
          6595 => x"5a",
          6596 => x"80",
          6597 => x"ef",
          6598 => x"84",
          6599 => x"74",
          6600 => x"3d",
          6601 => x"9e",
          6602 => x"ff",
          6603 => x"86",
          6604 => x"3d",
          6605 => x"fe",
          6606 => x"f4",
          6607 => x"84",
          6608 => x"80",
          6609 => x"59",
          6610 => x"33",
          6611 => x"15",
          6612 => x"0b",
          6613 => x"ec",
          6614 => x"56",
          6615 => x"8a",
          6616 => x"b9",
          6617 => x"fe",
          6618 => x"fe",
          6619 => x"52",
          6620 => x"c8",
          6621 => x"2e",
          6622 => x"b9",
          6623 => x"16",
          6624 => x"77",
          6625 => x"74",
          6626 => x"38",
          6627 => x"81",
          6628 => x"84",
          6629 => x"ff",
          6630 => x"78",
          6631 => x"08",
          6632 => x"e5",
          6633 => x"80",
          6634 => x"2e",
          6635 => x"81",
          6636 => x"fe",
          6637 => x"57",
          6638 => x"86",
          6639 => x"bf",
          6640 => x"a0",
          6641 => x"05",
          6642 => x"38",
          6643 => x"8b",
          6644 => x"81",
          6645 => x"58",
          6646 => x"fd",
          6647 => x"33",
          6648 => x"15",
          6649 => x"6b",
          6650 => x"0b",
          6651 => x"bc",
          6652 => x"ce",
          6653 => x"54",
          6654 => x"18",
          6655 => x"b9",
          6656 => x"80",
          6657 => x"19",
          6658 => x"31",
          6659 => x"38",
          6660 => x"b1",
          6661 => x"e8",
          6662 => x"fe",
          6663 => x"57",
          6664 => x"b6",
          6665 => x"59",
          6666 => x"a1",
          6667 => x"19",
          6668 => x"33",
          6669 => x"39",
          6670 => x"05",
          6671 => x"89",
          6672 => x"08",
          6673 => x"33",
          6674 => x"15",
          6675 => x"78",
          6676 => x"5f",
          6677 => x"56",
          6678 => x"81",
          6679 => x"38",
          6680 => x"06",
          6681 => x"38",
          6682 => x"70",
          6683 => x"87",
          6684 => x"30",
          6685 => x"c8",
          6686 => x"53",
          6687 => x"38",
          6688 => x"82",
          6689 => x"74",
          6690 => x"81",
          6691 => x"75",
          6692 => x"c8",
          6693 => x"b9",
          6694 => x"84",
          6695 => x"19",
          6696 => x"78",
          6697 => x"56",
          6698 => x"90",
          6699 => x"c8",
          6700 => x"33",
          6701 => x"c8",
          6702 => x"38",
          6703 => x"39",
          6704 => x"7d",
          6705 => x"81",
          6706 => x"38",
          6707 => x"dd",
          6708 => x"84",
          6709 => x"81",
          6710 => x"d7",
          6711 => x"7b",
          6712 => x"18",
          6713 => x"33",
          6714 => x"34",
          6715 => x"08",
          6716 => x"38",
          6717 => x"15",
          6718 => x"34",
          6719 => x"ff",
          6720 => x"be",
          6721 => x"54",
          6722 => x"a1",
          6723 => x"0d",
          6724 => x"88",
          6725 => x"5f",
          6726 => x"5b",
          6727 => x"79",
          6728 => x"26",
          6729 => x"38",
          6730 => x"92",
          6731 => x"76",
          6732 => x"84",
          6733 => x"74",
          6734 => x"75",
          6735 => x"b9",
          6736 => x"52",
          6737 => x"b9",
          6738 => x"06",
          6739 => x"38",
          6740 => x"57",
          6741 => x"05",
          6742 => x"b0",
          6743 => x"38",
          6744 => x"38",
          6745 => x"38",
          6746 => x"ff",
          6747 => x"80",
          6748 => x"80",
          6749 => x"7f",
          6750 => x"89",
          6751 => x"89",
          6752 => x"80",
          6753 => x"80",
          6754 => x"74",
          6755 => x"df",
          6756 => x"79",
          6757 => x"84",
          6758 => x"83",
          6759 => x"33",
          6760 => x"57",
          6761 => x"06",
          6762 => x"05",
          6763 => x"80",
          6764 => x"83",
          6765 => x"2b",
          6766 => x"70",
          6767 => x"07",
          6768 => x"12",
          6769 => x"07",
          6770 => x"2b",
          6771 => x"0c",
          6772 => x"44",
          6773 => x"4b",
          6774 => x"27",
          6775 => x"80",
          6776 => x"70",
          6777 => x"83",
          6778 => x"82",
          6779 => x"66",
          6780 => x"4a",
          6781 => x"8a",
          6782 => x"2a",
          6783 => x"56",
          6784 => x"77",
          6785 => x"77",
          6786 => x"58",
          6787 => x"27",
          6788 => x"81",
          6789 => x"84",
          6790 => x"f5",
          6791 => x"c8",
          6792 => x"71",
          6793 => x"43",
          6794 => x"5c",
          6795 => x"05",
          6796 => x"72",
          6797 => x"2e",
          6798 => x"90",
          6799 => x"74",
          6800 => x"31",
          6801 => x"52",
          6802 => x"c8",
          6803 => x"38",
          6804 => x"dd",
          6805 => x"c8",
          6806 => x"f9",
          6807 => x"26",
          6808 => x"39",
          6809 => x"9f",
          6810 => x"81",
          6811 => x"b9",
          6812 => x"d4",
          6813 => x"81",
          6814 => x"26",
          6815 => x"06",
          6816 => x"81",
          6817 => x"5f",
          6818 => x"70",
          6819 => x"05",
          6820 => x"57",
          6821 => x"70",
          6822 => x"18",
          6823 => x"18",
          6824 => x"30",
          6825 => x"2e",
          6826 => x"be",
          6827 => x"72",
          6828 => x"4a",
          6829 => x"1c",
          6830 => x"ff",
          6831 => x"9f",
          6832 => x"51",
          6833 => x"b9",
          6834 => x"2a",
          6835 => x"56",
          6836 => x"8e",
          6837 => x"74",
          6838 => x"56",
          6839 => x"ba",
          6840 => x"f9",
          6841 => x"57",
          6842 => x"6e",
          6843 => x"39",
          6844 => x"9d",
          6845 => x"81",
          6846 => x"57",
          6847 => x"0d",
          6848 => x"62",
          6849 => x"60",
          6850 => x"8e",
          6851 => x"61",
          6852 => x"58",
          6853 => x"8b",
          6854 => x"76",
          6855 => x"81",
          6856 => x"ef",
          6857 => x"34",
          6858 => x"8d",
          6859 => x"4b",
          6860 => x"2a",
          6861 => x"61",
          6862 => x"30",
          6863 => x"78",
          6864 => x"92",
          6865 => x"ff",
          6866 => x"ff",
          6867 => x"74",
          6868 => x"34",
          6869 => x"98",
          6870 => x"ff",
          6871 => x"05",
          6872 => x"88",
          6873 => x"7e",
          6874 => x"34",
          6875 => x"84",
          6876 => x"62",
          6877 => x"a7",
          6878 => x"a1",
          6879 => x"aa",
          6880 => x"55",
          6881 => x"2a",
          6882 => x"80",
          6883 => x"05",
          6884 => x"90",
          6885 => x"58",
          6886 => x"ff",
          6887 => x"fe",
          6888 => x"83",
          6889 => x"81",
          6890 => x"fe",
          6891 => x"c8",
          6892 => x"62",
          6893 => x"57",
          6894 => x"34",
          6895 => x"75",
          6896 => x"38",
          6897 => x"2e",
          6898 => x"76",
          6899 => x"70",
          6900 => x"59",
          6901 => x"76",
          6902 => x"57",
          6903 => x"76",
          6904 => x"79",
          6905 => x"c8",
          6906 => x"57",
          6907 => x"34",
          6908 => x"1b",
          6909 => x"38",
          6910 => x"ff",
          6911 => x"83",
          6912 => x"26",
          6913 => x"53",
          6914 => x"3f",
          6915 => x"74",
          6916 => x"db",
          6917 => x"38",
          6918 => x"8a",
          6919 => x"38",
          6920 => x"83",
          6921 => x"38",
          6922 => x"70",
          6923 => x"78",
          6924 => x"aa",
          6925 => x"78",
          6926 => x"81",
          6927 => x"05",
          6928 => x"43",
          6929 => x"fc",
          6930 => x"34",
          6931 => x"07",
          6932 => x"b9",
          6933 => x"61",
          6934 => x"c7",
          6935 => x"34",
          6936 => x"05",
          6937 => x"62",
          6938 => x"05",
          6939 => x"83",
          6940 => x"7e",
          6941 => x"78",
          6942 => x"f1",
          6943 => x"f7",
          6944 => x"51",
          6945 => x"b9",
          6946 => x"c8",
          6947 => x"0d",
          6948 => x"f9",
          6949 => x"5c",
          6950 => x"91",
          6951 => x"22",
          6952 => x"74",
          6953 => x"56",
          6954 => x"57",
          6955 => x"75",
          6956 => x"fc",
          6957 => x"10",
          6958 => x"5e",
          6959 => x"c8",
          6960 => x"fd",
          6961 => x"38",
          6962 => x"c8",
          6963 => x"38",
          6964 => x"5b",
          6965 => x"c8",
          6966 => x"2e",
          6967 => x"39",
          6968 => x"2a",
          6969 => x"90",
          6970 => x"75",
          6971 => x"34",
          6972 => x"05",
          6973 => x"a1",
          6974 => x"61",
          6975 => x"05",
          6976 => x"a5",
          6977 => x"61",
          6978 => x"75",
          6979 => x"05",
          6980 => x"61",
          6981 => x"34",
          6982 => x"b1",
          6983 => x"80",
          6984 => x"80",
          6985 => x"05",
          6986 => x"e5",
          6987 => x"05",
          6988 => x"34",
          6989 => x"cd",
          6990 => x"76",
          6991 => x"55",
          6992 => x"54",
          6993 => x"be",
          6994 => x"08",
          6995 => x"05",
          6996 => x"76",
          6997 => x"52",
          6998 => x"c3",
          6999 => x"9f",
          7000 => x"f8",
          7001 => x"81",
          7002 => x"05",
          7003 => x"84",
          7004 => x"ff",
          7005 => x"05",
          7006 => x"61",
          7007 => x"34",
          7008 => x"39",
          7009 => x"79",
          7010 => x"61",
          7011 => x"57",
          7012 => x"60",
          7013 => x"5e",
          7014 => x"81",
          7015 => x"81",
          7016 => x"80",
          7017 => x"f2",
          7018 => x"61",
          7019 => x"83",
          7020 => x"7a",
          7021 => x"2a",
          7022 => x"7a",
          7023 => x"05",
          7024 => x"83",
          7025 => x"05",
          7026 => x"76",
          7027 => x"83",
          7028 => x"ff",
          7029 => x"53",
          7030 => x"3f",
          7031 => x"79",
          7032 => x"57",
          7033 => x"7e",
          7034 => x"05",
          7035 => x"38",
          7036 => x"54",
          7037 => x"9a",
          7038 => x"06",
          7039 => x"8d",
          7040 => x"05",
          7041 => x"2e",
          7042 => x"80",
          7043 => x"76",
          7044 => x"3d",
          7045 => x"84",
          7046 => x"8a",
          7047 => x"56",
          7048 => x"08",
          7049 => x"75",
          7050 => x"8e",
          7051 => x"88",
          7052 => x"3d",
          7053 => x"52",
          7054 => x"74",
          7055 => x"9f",
          7056 => x"1c",
          7057 => x"39",
          7058 => x"ff",
          7059 => x"ff",
          7060 => x"cc",
          7061 => x"05",
          7062 => x"38",
          7063 => x"2e",
          7064 => x"24",
          7065 => x"05",
          7066 => x"55",
          7067 => x"18",
          7068 => x"55",
          7069 => x"ff",
          7070 => x"52",
          7071 => x"84",
          7072 => x"2e",
          7073 => x"0c",
          7074 => x"b0",
          7075 => x"76",
          7076 => x"7b",
          7077 => x"2a",
          7078 => x"a5",
          7079 => x"3f",
          7080 => x"0c",
          7081 => x"75",
          7082 => x"53",
          7083 => x"38",
          7084 => x"84",
          7085 => x"83",
          7086 => x"b5",
          7087 => x"80",
          7088 => x"51",
          7089 => x"70",
          7090 => x"80",
          7091 => x"e7",
          7092 => x"39",
          7093 => x"84",
          7094 => x"04",
          7095 => x"02",
          7096 => x"80",
          7097 => x"70",
          7098 => x"3d",
          7099 => x"81",
          7100 => x"e9",
          7101 => x"70",
          7102 => x"3d",
          7103 => x"70",
          7104 => x"70",
          7105 => x"56",
          7106 => x"38",
          7107 => x"71",
          7108 => x"07",
          7109 => x"71",
          7110 => x"88",
          7111 => x"14",
          7112 => x"71",
          7113 => x"82",
          7114 => x"80",
          7115 => x"52",
          7116 => x"70",
          7117 => x"04",
          7118 => x"71",
          7119 => x"83",
          7120 => x"c7",
          7121 => x"57",
          7122 => x"16",
          7123 => x"f1",
          7124 => x"06",
          7125 => x"83",
          7126 => x"d0",
          7127 => x"51",
          7128 => x"ff",
          7129 => x"70",
          7130 => x"b9",
          7131 => x"71",
          7132 => x"52",
          7133 => x"10",
          7134 => x"ef",
          7135 => x"ff",
          7136 => x"ff",
          7137 => x"00",
          7138 => x"00",
          7139 => x"00",
          7140 => x"00",
          7141 => x"00",
          7142 => x"00",
          7143 => x"00",
          7144 => x"00",
          7145 => x"00",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"64",
          7374 => x"64",
          7375 => x"66",
          7376 => x"66",
          7377 => x"66",
          7378 => x"6d",
          7379 => x"6d",
          7380 => x"6d",
          7381 => x"6d",
          7382 => x"6d",
          7383 => x"6d",
          7384 => x"68",
          7385 => x"68",
          7386 => x"00",
          7387 => x"72",
          7388 => x"72",
          7389 => x"69",
          7390 => x"74",
          7391 => x"63",
          7392 => x"74",
          7393 => x"6d",
          7394 => x"6b",
          7395 => x"65",
          7396 => x"6f",
          7397 => x"72",
          7398 => x"6d",
          7399 => x"6e",
          7400 => x"2e",
          7401 => x"6d",
          7402 => x"6e",
          7403 => x"00",
          7404 => x"66",
          7405 => x"20",
          7406 => x"00",
          7407 => x"20",
          7408 => x"65",
          7409 => x"6f",
          7410 => x"72",
          7411 => x"61",
          7412 => x"2e",
          7413 => x"61",
          7414 => x"65",
          7415 => x"6f",
          7416 => x"65",
          7417 => x"73",
          7418 => x"6e",
          7419 => x"73",
          7420 => x"20",
          7421 => x"62",
          7422 => x"44",
          7423 => x"6d",
          7424 => x"69",
          7425 => x"00",
          7426 => x"73",
          7427 => x"70",
          7428 => x"64",
          7429 => x"20",
          7430 => x"69",
          7431 => x"00",
          7432 => x"20",
          7433 => x"20",
          7434 => x"00",
          7435 => x"73",
          7436 => x"64",
          7437 => x"6c",
          7438 => x"6e",
          7439 => x"4e",
          7440 => x"66",
          7441 => x"4e",
          7442 => x"66",
          7443 => x"44",
          7444 => x"20",
          7445 => x"49",
          7446 => x"20",
          7447 => x"44",
          7448 => x"6f",
          7449 => x"65",
          7450 => x"0a",
          7451 => x"65",
          7452 => x"20",
          7453 => x"65",
          7454 => x"00",
          7455 => x"00",
          7456 => x"58",
          7457 => x"25",
          7458 => x"20",
          7459 => x"20",
          7460 => x"00",
          7461 => x"20",
          7462 => x"7a",
          7463 => x"73",
          7464 => x"34",
          7465 => x"76",
          7466 => x"20",
          7467 => x"76",
          7468 => x"25",
          7469 => x"0a",
          7470 => x"20",
          7471 => x"20",
          7472 => x"20",
          7473 => x"20",
          7474 => x"30",
          7475 => x"20",
          7476 => x"41",
          7477 => x"20",
          7478 => x"20",
          7479 => x"30",
          7480 => x"5a",
          7481 => x"72",
          7482 => x"6e",
          7483 => x"55",
          7484 => x"20",
          7485 => x"70",
          7486 => x"31",
          7487 => x"65",
          7488 => x"55",
          7489 => x"20",
          7490 => x"70",
          7491 => x"30",
          7492 => x"65",
          7493 => x"49",
          7494 => x"20",
          7495 => x"70",
          7496 => x"4c",
          7497 => x"65",
          7498 => x"50",
          7499 => x"72",
          7500 => x"54",
          7501 => x"74",
          7502 => x"53",
          7503 => x"75",
          7504 => x"2e",
          7505 => x"6c",
          7506 => x"65",
          7507 => x"61",
          7508 => x"2e",
          7509 => x"7a",
          7510 => x"68",
          7511 => x"65",
          7512 => x"69",
          7513 => x"20",
          7514 => x"20",
          7515 => x"73",
          7516 => x"6d",
          7517 => x"2e",
          7518 => x"25",
          7519 => x"30",
          7520 => x"63",
          7521 => x"00",
          7522 => x"62",
          7523 => x"25",
          7524 => x"00",
          7525 => x"20",
          7526 => x"6e",
          7527 => x"52",
          7528 => x"6e",
          7529 => x"63",
          7530 => x"2e",
          7531 => x"69",
          7532 => x"20",
          7533 => x"20",
          7534 => x"43",
          7535 => x"75",
          7536 => x"64",
          7537 => x"0a",
          7538 => x"75",
          7539 => x"64",
          7540 => x"6c",
          7541 => x"25",
          7542 => x"38",
          7543 => x"25",
          7544 => x"34",
          7545 => x"61",
          7546 => x"00",
          7547 => x"78",
          7548 => x"3e",
          7549 => x"30",
          7550 => x"43",
          7551 => x"2e",
          7552 => x"58",
          7553 => x"43",
          7554 => x"2e",
          7555 => x"44",
          7556 => x"6f",
          7557 => x"70",
          7558 => x"25",
          7559 => x"73",
          7560 => x"72",
          7561 => x"73",
          7562 => x"6e",
          7563 => x"63",
          7564 => x"6d",
          7565 => x"3f",
          7566 => x"64",
          7567 => x"25",
          7568 => x"25",
          7569 => x"43",
          7570 => x"61",
          7571 => x"3a",
          7572 => x"73",
          7573 => x"65",
          7574 => x"41",
          7575 => x"73",
          7576 => x"43",
          7577 => x"74",
          7578 => x"20",
          7579 => x"20",
          7580 => x"00",
          7581 => x"43",
          7582 => x"72",
          7583 => x"20",
          7584 => x"20",
          7585 => x"00",
          7586 => x"53",
          7587 => x"61",
          7588 => x"65",
          7589 => x"20",
          7590 => x"00",
          7591 => x"3a",
          7592 => x"5a",
          7593 => x"20",
          7594 => x"20",
          7595 => x"20",
          7596 => x"00",
          7597 => x"53",
          7598 => x"6c",
          7599 => x"71",
          7600 => x"20",
          7601 => x"34",
          7602 => x"20",
          7603 => x"62",
          7604 => x"41",
          7605 => x"20",
          7606 => x"64",
          7607 => x"7a",
          7608 => x"53",
          7609 => x"6f",
          7610 => x"20",
          7611 => x"20",
          7612 => x"34",
          7613 => x"20",
          7614 => x"20",
          7615 => x"20",
          7616 => x"4c",
          7617 => x"57",
          7618 => x"20",
          7619 => x"42",
          7620 => x"00",
          7621 => x"49",
          7622 => x"4c",
          7623 => x"65",
          7624 => x"29",
          7625 => x"54",
          7626 => x"20",
          7627 => x"73",
          7628 => x"29",
          7629 => x"53",
          7630 => x"20",
          7631 => x"65",
          7632 => x"29",
          7633 => x"52",
          7634 => x"20",
          7635 => x"25",
          7636 => x"20",
          7637 => x"20",
          7638 => x"30",
          7639 => x"29",
          7640 => x"49",
          7641 => x"4d",
          7642 => x"25",
          7643 => x"20",
          7644 => x"4d",
          7645 => x"30",
          7646 => x"29",
          7647 => x"57",
          7648 => x"20",
          7649 => x"25",
          7650 => x"20",
          7651 => x"6f",
          7652 => x"67",
          7653 => x"6f",
          7654 => x"00",
          7655 => x"6c",
          7656 => x"75",
          7657 => x"00",
          7658 => x"00",
          7659 => x"00",
          7660 => x"01",
          7661 => x"00",
          7662 => x"00",
          7663 => x"01",
          7664 => x"00",
          7665 => x"00",
          7666 => x"01",
          7667 => x"00",
          7668 => x"00",
          7669 => x"01",
          7670 => x"00",
          7671 => x"00",
          7672 => x"01",
          7673 => x"00",
          7674 => x"00",
          7675 => x"04",
          7676 => x"00",
          7677 => x"00",
          7678 => x"04",
          7679 => x"00",
          7680 => x"00",
          7681 => x"04",
          7682 => x"00",
          7683 => x"00",
          7684 => x"04",
          7685 => x"00",
          7686 => x"00",
          7687 => x"03",
          7688 => x"00",
          7689 => x"00",
          7690 => x"03",
          7691 => x"1b",
          7692 => x"1b",
          7693 => x"1b",
          7694 => x"1b",
          7695 => x"1b",
          7696 => x"1b",
          7697 => x"0e",
          7698 => x"0b",
          7699 => x"06",
          7700 => x"04",
          7701 => x"02",
          7702 => x"43",
          7703 => x"70",
          7704 => x"74",
          7705 => x"72",
          7706 => x"20",
          7707 => x"6e",
          7708 => x"6f",
          7709 => x"00",
          7710 => x"25",
          7711 => x"73",
          7712 => x"65",
          7713 => x"73",
          7714 => x"68",
          7715 => x"66",
          7716 => x"45",
          7717 => x"3e",
          7718 => x"1b",
          7719 => x"1b",
          7720 => x"1b",
          7721 => x"1b",
          7722 => x"1b",
          7723 => x"1b",
          7724 => x"1b",
          7725 => x"1b",
          7726 => x"1b",
          7727 => x"1b",
          7728 => x"1b",
          7729 => x"1b",
          7730 => x"1b",
          7731 => x"1b",
          7732 => x"1b",
          7733 => x"1b",
          7734 => x"00",
          7735 => x"00",
          7736 => x"2c",
          7737 => x"64",
          7738 => x"25",
          7739 => x"44",
          7740 => x"25",
          7741 => x"2c",
          7742 => x"25",
          7743 => x"3a",
          7744 => x"2c",
          7745 => x"64",
          7746 => x"52",
          7747 => x"75",
          7748 => x"55",
          7749 => x"25",
          7750 => x"44",
          7751 => x"25",
          7752 => x"48",
          7753 => x"00",
          7754 => x"65",
          7755 => x"6e",
          7756 => x"53",
          7757 => x"3e",
          7758 => x"2b",
          7759 => x"46",
          7760 => x"32",
          7761 => x"53",
          7762 => x"4e",
          7763 => x"20",
          7764 => x"20",
          7765 => x"41",
          7766 => x"41",
          7767 => x"00",
          7768 => x"00",
          7769 => x"01",
          7770 => x"14",
          7771 => x"80",
          7772 => x"45",
          7773 => x"90",
          7774 => x"59",
          7775 => x"41",
          7776 => x"a8",
          7777 => x"b0",
          7778 => x"b8",
          7779 => x"c0",
          7780 => x"c8",
          7781 => x"d0",
          7782 => x"d8",
          7783 => x"e0",
          7784 => x"e8",
          7785 => x"f0",
          7786 => x"f8",
          7787 => x"2b",
          7788 => x"5c",
          7789 => x"7f",
          7790 => x"00",
          7791 => x"00",
          7792 => x"00",
          7793 => x"00",
          7794 => x"00",
          7795 => x"00",
          7796 => x"00",
          7797 => x"00",
          7798 => x"00",
          7799 => x"00",
          7800 => x"00",
          7801 => x"20",
          7802 => x"00",
          7803 => x"00",
          7804 => x"00",
          7805 => x"00",
          7806 => x"25",
          7807 => x"25",
          7808 => x"25",
          7809 => x"25",
          7810 => x"25",
          7811 => x"25",
          7812 => x"25",
          7813 => x"25",
          7814 => x"25",
          7815 => x"25",
          7816 => x"25",
          7817 => x"25",
          7818 => x"03",
          7819 => x"00",
          7820 => x"03",
          7821 => x"03",
          7822 => x"22",
          7823 => x"00",
          7824 => x"00",
          7825 => x"25",
          7826 => x"00",
          7827 => x"00",
          7828 => x"01",
          7829 => x"01",
          7830 => x"01",
          7831 => x"01",
          7832 => x"01",
          7833 => x"01",
          7834 => x"01",
          7835 => x"01",
          7836 => x"01",
          7837 => x"01",
          7838 => x"01",
          7839 => x"01",
          7840 => x"01",
          7841 => x"01",
          7842 => x"01",
          7843 => x"01",
          7844 => x"01",
          7845 => x"01",
          7846 => x"01",
          7847 => x"01",
          7848 => x"01",
          7849 => x"01",
          7850 => x"01",
          7851 => x"01",
          7852 => x"00",
          7853 => x"01",
          7854 => x"02",
          7855 => x"02",
          7856 => x"02",
          7857 => x"01",
          7858 => x"01",
          7859 => x"02",
          7860 => x"02",
          7861 => x"01",
          7862 => x"02",
          7863 => x"01",
          7864 => x"02",
          7865 => x"02",
          7866 => x"02",
          7867 => x"02",
          7868 => x"02",
          7869 => x"01",
          7870 => x"02",
          7871 => x"01",
          7872 => x"02",
          7873 => x"02",
          7874 => x"00",
          7875 => x"03",
          7876 => x"03",
          7877 => x"03",
          7878 => x"03",
          7879 => x"03",
          7880 => x"01",
          7881 => x"03",
          7882 => x"03",
          7883 => x"03",
          7884 => x"07",
          7885 => x"01",
          7886 => x"00",
          7887 => x"05",
          7888 => x"1d",
          7889 => x"01",
          7890 => x"06",
          7891 => x"06",
          7892 => x"06",
          7893 => x"1f",
          7894 => x"1f",
          7895 => x"1f",
          7896 => x"1f",
          7897 => x"1f",
          7898 => x"1f",
          7899 => x"1f",
          7900 => x"1f",
          7901 => x"1f",
          7902 => x"1f",
          7903 => x"06",
          7904 => x"00",
          7905 => x"1f",
          7906 => x"21",
          7907 => x"21",
          7908 => x"04",
          7909 => x"01",
          7910 => x"01",
          7911 => x"03",
          7912 => x"00",
          7913 => x"00",
          7914 => x"00",
          7915 => x"00",
          7916 => x"00",
          7917 => x"00",
          7918 => x"00",
          7919 => x"00",
          7920 => x"00",
          7921 => x"00",
          7922 => x"00",
          7923 => x"00",
          7924 => x"00",
          7925 => x"00",
          7926 => x"00",
          7927 => x"00",
          7928 => x"00",
          7929 => x"00",
          7930 => x"00",
          7931 => x"00",
          7932 => x"00",
          7933 => x"00",
          7934 => x"00",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"00",
          7963 => x"00",
          7964 => x"00",
          7965 => x"00",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"01",
          7974 => x"00",
          7975 => x"00",
          7976 => x"05",
          7977 => x"00",
          7978 => x"01",
          7979 => x"01",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"00",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"01",
          7993 => x"01",
          7994 => x"02",
          7995 => x"1b",
          7996 => x"79",
          7997 => x"71",
          7998 => x"69",
          7999 => x"61",
          8000 => x"31",
          8001 => x"5c",
          8002 => x"f6",
          8003 => x"08",
          8004 => x"80",
          8005 => x"1b",
          8006 => x"59",
          8007 => x"51",
          8008 => x"49",
          8009 => x"41",
          8010 => x"31",
          8011 => x"5c",
          8012 => x"f6",
          8013 => x"08",
          8014 => x"80",
          8015 => x"1b",
          8016 => x"59",
          8017 => x"51",
          8018 => x"49",
          8019 => x"41",
          8020 => x"21",
          8021 => x"7c",
          8022 => x"f7",
          8023 => x"fb",
          8024 => x"85",
          8025 => x"1b",
          8026 => x"19",
          8027 => x"11",
          8028 => x"09",
          8029 => x"01",
          8030 => x"f0",
          8031 => x"f0",
          8032 => x"f0",
          8033 => x"f0",
          8034 => x"80",
          8035 => x"bf",
          8036 => x"35",
          8037 => x"7c",
          8038 => x"3d",
          8039 => x"46",
          8040 => x"3f",
          8041 => x"d3",
          8042 => x"c6",
          8043 => x"f0",
          8044 => x"80",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"ce",
          9082 => x"fc",
          9083 => x"c4",
          9084 => x"eb",
          9085 => x"64",
          9086 => x"2f",
          9087 => x"24",
          9088 => x"51",
          9089 => x"04",
          9090 => x"0c",
          9091 => x"14",
          9092 => x"59",
          9093 => x"84",
          9094 => x"8c",
          9095 => x"94",
          9096 => x"80",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
        others => X"00"
    );

    shared variable RAM4 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"80",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"09",
             9 => x"83",
            10 => x"00",
            11 => x"00",
            12 => x"73",
            13 => x"83",
            14 => x"ff",
            15 => x"00",
            16 => x"73",
            17 => x"06",
            18 => x"00",
            19 => x"00",
            20 => x"53",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"72",
            26 => x"06",
            27 => x"00",
            28 => x"53",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"04",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"0b",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"2a",
            49 => x"05",
            50 => x"00",
            51 => x"00",
            52 => x"83",
            53 => x"2b",
            54 => x"51",
            55 => x"00",
            56 => x"70",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"70",
            61 => x"06",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"51",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"06",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"09",
            77 => x"2a",
            78 => x"00",
            79 => x"00",
            80 => x"bd",
            81 => x"08",
            82 => x"00",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"88",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"88",
            91 => x"00",
            92 => x"0a",
            93 => x"06",
            94 => x"06",
            95 => x"00",
            96 => x"0a",
            97 => x"71",
            98 => x"05",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"52",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"51",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"8c",
           134 => x"04",
           135 => x"0b",
           136 => x"8c",
           137 => x"04",
           138 => x"0b",
           139 => x"8d",
           140 => x"04",
           141 => x"0b",
           142 => x"8d",
           143 => x"04",
           144 => x"0b",
           145 => x"8e",
           146 => x"04",
           147 => x"0b",
           148 => x"8e",
           149 => x"04",
           150 => x"0b",
           151 => x"8f",
           152 => x"04",
           153 => x"0b",
           154 => x"8f",
           155 => x"04",
           156 => x"0b",
           157 => x"90",
           158 => x"04",
           159 => x"0b",
           160 => x"90",
           161 => x"04",
           162 => x"0b",
           163 => x"91",
           164 => x"04",
           165 => x"0b",
           166 => x"91",
           167 => x"04",
           168 => x"0b",
           169 => x"92",
           170 => x"04",
           171 => x"0b",
           172 => x"92",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"d4",
           193 => x"d4",
           194 => x"b9",
           195 => x"d4",
           196 => x"b9",
           197 => x"d4",
           198 => x"b9",
           199 => x"d4",
           200 => x"b9",
           201 => x"d4",
           202 => x"b9",
           203 => x"d4",
           204 => x"b9",
           205 => x"d4",
           206 => x"b9",
           207 => x"d4",
           208 => x"b9",
           209 => x"d4",
           210 => x"b9",
           211 => x"d4",
           212 => x"b9",
           213 => x"d4",
           214 => x"b9",
           215 => x"d4",
           216 => x"b9",
           217 => x"b9",
           218 => x"84",
           219 => x"84",
           220 => x"04",
           221 => x"2d",
           222 => x"90",
           223 => x"db",
           224 => x"80",
           225 => x"c9",
           226 => x"c0",
           227 => x"82",
           228 => x"80",
           229 => x"0c",
           230 => x"08",
           231 => x"d4",
           232 => x"d4",
           233 => x"b9",
           234 => x"b9",
           235 => x"84",
           236 => x"84",
           237 => x"04",
           238 => x"2d",
           239 => x"90",
           240 => x"be",
           241 => x"80",
           242 => x"f3",
           243 => x"c0",
           244 => x"82",
           245 => x"80",
           246 => x"0c",
           247 => x"08",
           248 => x"d4",
           249 => x"d4",
           250 => x"b9",
           251 => x"b9",
           252 => x"84",
           253 => x"84",
           254 => x"04",
           255 => x"2d",
           256 => x"90",
           257 => x"88",
           258 => x"80",
           259 => x"e5",
           260 => x"c0",
           261 => x"82",
           262 => x"80",
           263 => x"0c",
           264 => x"08",
           265 => x"d4",
           266 => x"d4",
           267 => x"b9",
           268 => x"b9",
           269 => x"84",
           270 => x"84",
           271 => x"04",
           272 => x"2d",
           273 => x"90",
           274 => x"ff",
           275 => x"80",
           276 => x"a4",
           277 => x"c0",
           278 => x"83",
           279 => x"80",
           280 => x"0c",
           281 => x"08",
           282 => x"d4",
           283 => x"d4",
           284 => x"b9",
           285 => x"b9",
           286 => x"84",
           287 => x"84",
           288 => x"04",
           289 => x"2d",
           290 => x"90",
           291 => x"fa",
           292 => x"80",
           293 => x"d7",
           294 => x"c0",
           295 => x"b1",
           296 => x"c0",
           297 => x"81",
           298 => x"80",
           299 => x"0c",
           300 => x"08",
           301 => x"d4",
           302 => x"d4",
           303 => x"b9",
           304 => x"b9",
           305 => x"3c",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"ff",
           311 => x"83",
           312 => x"fc",
           313 => x"80",
           314 => x"06",
           315 => x"0a",
           316 => x"51",
           317 => x"b4",
           318 => x"05",
           319 => x"04",
           320 => x"00",
           321 => x"84",
           322 => x"84",
           323 => x"86",
           324 => x"7a",
           325 => x"06",
           326 => x"57",
           327 => x"06",
           328 => x"8a",
           329 => x"2a",
           330 => x"25",
           331 => x"75",
           332 => x"08",
           333 => x"ae",
           334 => x"81",
           335 => x"32",
           336 => x"51",
           337 => x"38",
           338 => x"b9",
           339 => x"0b",
           340 => x"04",
           341 => x"84",
           342 => x"0a",
           343 => x"52",
           344 => x"73",
           345 => x"0d",
           346 => x"05",
           347 => x"85",
           348 => x"63",
           349 => x"1f",
           350 => x"81",
           351 => x"54",
           352 => x"d2",
           353 => x"80",
           354 => x"54",
           355 => x"d0",
           356 => x"38",
           357 => x"25",
           358 => x"80",
           359 => x"81",
           360 => x"2e",
           361 => x"7b",
           362 => x"1d",
           363 => x"91",
           364 => x"78",
           365 => x"98",
           366 => x"80",
           367 => x"2c",
           368 => x"24",
           369 => x"72",
           370 => x"58",
           371 => x"76",
           372 => x"81",
           373 => x"33",
           374 => x"9e",
           375 => x"3f",
           376 => x"ff",
           377 => x"06",
           378 => x"74",
           379 => x"17",
           380 => x"72",
           381 => x"73",
           382 => x"80",
           383 => x"76",
           384 => x"58",
           385 => x"39",
           386 => x"5a",
           387 => x"83",
           388 => x"84",
           389 => x"93",
           390 => x"ff",
           391 => x"05",
           392 => x"84",
           393 => x"7e",
           394 => x"75",
           395 => x"08",
           396 => x"7d",
           397 => x"b2",
           398 => x"38",
           399 => x"80",
           400 => x"86",
           401 => x"80",
           402 => x"29",
           403 => x"2e",
           404 => x"fc",
           405 => x"58",
           406 => x"55",
           407 => x"2c",
           408 => x"73",
           409 => x"f7",
           410 => x"41",
           411 => x"80",
           412 => x"90",
           413 => x"06",
           414 => x"96",
           415 => x"73",
           416 => x"06",
           417 => x"2a",
           418 => x"7e",
           419 => x"7a",
           420 => x"2e",
           421 => x"29",
           422 => x"5a",
           423 => x"7c",
           424 => x"78",
           425 => x"05",
           426 => x"80",
           427 => x"72",
           428 => x"80",
           429 => x"98",
           430 => x"9d",
           431 => x"3f",
           432 => x"ff",
           433 => x"55",
           434 => x"2a",
           435 => x"2e",
           436 => x"84",
           437 => x"ca",
           438 => x"38",
           439 => x"7c",
           440 => x"87",
           441 => x"09",
           442 => x"5b",
           443 => x"78",
           444 => x"05",
           445 => x"75",
           446 => x"51",
           447 => x"07",
           448 => x"5b",
           449 => x"7a",
           450 => x"90",
           451 => x"83",
           452 => x"5a",
           453 => x"77",
           454 => x"70",
           455 => x"80",
           456 => x"2c",
           457 => x"7a",
           458 => x"7a",
           459 => x"80",
           460 => x"2c",
           461 => x"b3",
           462 => x"3f",
           463 => x"ff",
           464 => x"2e",
           465 => x"81",
           466 => x"e2",
           467 => x"06",
           468 => x"fe",
           469 => x"05",
           470 => x"39",
           471 => x"07",
           472 => x"80",
           473 => x"80",
           474 => x"5d",
           475 => x"fb",
           476 => x"70",
           477 => x"82",
           478 => x"5b",
           479 => x"7a",
           480 => x"f8",
           481 => x"07",
           482 => x"f7",
           483 => x"84",
           484 => x"58",
           485 => x"51",
           486 => x"83",
           487 => x"2b",
           488 => x"87",
           489 => x"58",
           490 => x"39",
           491 => x"81",
           492 => x"cf",
           493 => x"b9",
           494 => x"71",
           495 => x"7a",
           496 => x"76",
           497 => x"78",
           498 => x"05",
           499 => x"74",
           500 => x"51",
           501 => x"b0",
           502 => x"09",
           503 => x"76",
           504 => x"81",
           505 => x"38",
           506 => x"71",
           507 => x"83",
           508 => x"fa",
           509 => x"ad",
           510 => x"54",
           511 => x"ad",
           512 => x"82",
           513 => x"80",
           514 => x"78",
           515 => x"5a",
           516 => x"51",
           517 => x"a0",
           518 => x"78",
           519 => x"b9",
           520 => x"71",
           521 => x"39",
           522 => x"ff",
           523 => x"39",
           524 => x"53",
           525 => x"84",
           526 => x"55",
           527 => x"11",
           528 => x"81",
           529 => x"56",
           530 => x"d5",
           531 => x"53",
           532 => x"ac",
           533 => x"53",
           534 => x"2e",
           535 => x"05",
           536 => x"38",
           537 => x"84",
           538 => x"08",
           539 => x"74",
           540 => x"83",
           541 => x"b9",
           542 => x"3d",
           543 => x"85",
           544 => x"70",
           545 => x"56",
           546 => x"38",
           547 => x"72",
           548 => x"76",
           549 => x"3d",
           550 => x"33",
           551 => x"52",
           552 => x"2d",
           553 => x"38",
           554 => x"54",
           555 => x"3d",
           556 => x"51",
           557 => x"3d",
           558 => x"81",
           559 => x"56",
           560 => x"82",
           561 => x"ac",
           562 => x"16",
           563 => x"76",
           564 => x"0c",
           565 => x"16",
           566 => x"0c",
           567 => x"81",
           568 => x"73",
           569 => x"e3",
           570 => x"16",
           571 => x"0d",
           572 => x"06",
           573 => x"56",
           574 => x"86",
           575 => x"72",
           576 => x"2e",
           577 => x"53",
           578 => x"81",
           579 => x"05",
           580 => x"54",
           581 => x"0d",
           582 => x"85",
           583 => x"8c",
           584 => x"c8",
           585 => x"94",
           586 => x"c8",
           587 => x"25",
           588 => x"90",
           589 => x"ff",
           590 => x"72",
           591 => x"b9",
           592 => x"a0",
           593 => x"54",
           594 => x"71",
           595 => x"53",
           596 => x"52",
           597 => x"70",
           598 => x"f0",
           599 => x"3d",
           600 => x"71",
           601 => x"2e",
           602 => x"70",
           603 => x"05",
           604 => x"34",
           605 => x"84",
           606 => x"70",
           607 => x"70",
           608 => x"13",
           609 => x"11",
           610 => x"13",
           611 => x"34",
           612 => x"39",
           613 => x"71",
           614 => x"f7",
           615 => x"b9",
           616 => x"fd",
           617 => x"54",
           618 => x"70",
           619 => x"f0",
           620 => x"3d",
           621 => x"71",
           622 => x"2e",
           623 => x"33",
           624 => x"11",
           625 => x"c8",
           626 => x"0d",
           627 => x"80",
           628 => x"81",
           629 => x"2e",
           630 => x"54",
           631 => x"53",
           632 => x"b9",
           633 => x"80",
           634 => x"51",
           635 => x"33",
           636 => x"38",
           637 => x"86",
           638 => x"0c",
           639 => x"77",
           640 => x"3f",
           641 => x"08",
           642 => x"3f",
           643 => x"c8",
           644 => x"c8",
           645 => x"53",
           646 => x"fe",
           647 => x"73",
           648 => x"04",
           649 => x"54",
           650 => x"38",
           651 => x"70",
           652 => x"71",
           653 => x"ff",
           654 => x"84",
           655 => x"fd",
           656 => x"53",
           657 => x"72",
           658 => x"11",
           659 => x"c8",
           660 => x"0d",
           661 => x"80",
           662 => x"3f",
           663 => x"53",
           664 => x"80",
           665 => x"31",
           666 => x"cb",
           667 => x"c3",
           668 => x"72",
           669 => x"55",
           670 => x"72",
           671 => x"77",
           672 => x"2c",
           673 => x"71",
           674 => x"55",
           675 => x"10",
           676 => x"0c",
           677 => x"76",
           678 => x"70",
           679 => x"90",
           680 => x"fe",
           681 => x"83",
           682 => x"70",
           683 => x"25",
           684 => x"2a",
           685 => x"06",
           686 => x"71",
           687 => x"81",
           688 => x"74",
           689 => x"c8",
           690 => x"56",
           691 => x"56",
           692 => x"86",
           693 => x"77",
           694 => x"94",
           695 => x"74",
           696 => x"85",
           697 => x"7a",
           698 => x"8b",
           699 => x"b9",
           700 => x"80",
           701 => x"3f",
           702 => x"73",
           703 => x"80",
           704 => x"12",
           705 => x"71",
           706 => x"74",
           707 => x"9f",
           708 => x"72",
           709 => x"06",
           710 => x"1c",
           711 => x"53",
           712 => x"0c",
           713 => x"78",
           714 => x"2c",
           715 => x"73",
           716 => x"75",
           717 => x"fc",
           718 => x"32",
           719 => x"3d",
           720 => x"5b",
           721 => x"70",
           722 => x"09",
           723 => x"78",
           724 => x"2e",
           725 => x"38",
           726 => x"14",
           727 => x"db",
           728 => x"27",
           729 => x"89",
           730 => x"55",
           731 => x"51",
           732 => x"13",
           733 => x"73",
           734 => x"81",
           735 => x"16",
           736 => x"56",
           737 => x"80",
           738 => x"7a",
           739 => x"0c",
           740 => x"70",
           741 => x"73",
           742 => x"38",
           743 => x"55",
           744 => x"90",
           745 => x"81",
           746 => x"14",
           747 => x"27",
           748 => x"0c",
           749 => x"15",
           750 => x"80",
           751 => x"b9",
           752 => x"3d",
           753 => x"7b",
           754 => x"59",
           755 => x"38",
           756 => x"55",
           757 => x"ad",
           758 => x"81",
           759 => x"77",
           760 => x"80",
           761 => x"80",
           762 => x"70",
           763 => x"70",
           764 => x"27",
           765 => x"06",
           766 => x"38",
           767 => x"76",
           768 => x"70",
           769 => x"ff",
           770 => x"75",
           771 => x"75",
           772 => x"04",
           773 => x"33",
           774 => x"81",
           775 => x"78",
           776 => x"e2",
           777 => x"f8",
           778 => x"27",
           779 => x"88",
           780 => x"75",
           781 => x"04",
           782 => x"70",
           783 => x"39",
           784 => x"3d",
           785 => x"b9",
           786 => x"c8",
           787 => x"71",
           788 => x"83",
           789 => x"83",
           790 => x"3d",
           791 => x"b3",
           792 => x"c4",
           793 => x"04",
           794 => x"83",
           795 => x"ef",
           796 => x"cf",
           797 => x"0d",
           798 => x"3f",
           799 => x"51",
           800 => x"83",
           801 => x"3d",
           802 => x"db",
           803 => x"8c",
           804 => x"04",
           805 => x"83",
           806 => x"ee",
           807 => x"d0",
           808 => x"0d",
           809 => x"3f",
           810 => x"51",
           811 => x"83",
           812 => x"3d",
           813 => x"83",
           814 => x"a8",
           815 => x"04",
           816 => x"83",
           817 => x"ed",
           818 => x"3d",
           819 => x"05",
           820 => x"70",
           821 => x"59",
           822 => x"38",
           823 => x"ff",
           824 => x"e2",
           825 => x"70",
           826 => x"b9",
           827 => x"80",
           828 => x"af",
           829 => x"80",
           830 => x"06",
           831 => x"aa",
           832 => x"74",
           833 => x"52",
           834 => x"3f",
           835 => x"f4",
           836 => x"df",
           837 => x"96",
           838 => x"87",
           839 => x"08",
           840 => x"80",
           841 => x"ce",
           842 => x"b9",
           843 => x"74",
           844 => x"75",
           845 => x"52",
           846 => x"c8",
           847 => x"84",
           848 => x"53",
           849 => x"f8",
           850 => x"7c",
           851 => x"59",
           852 => x"51",
           853 => x"8b",
           854 => x"81",
           855 => x"0c",
           856 => x"d5",
           857 => x"b9",
           858 => x"2d",
           859 => x"0c",
           860 => x"7f",
           861 => x"05",
           862 => x"5c",
           863 => x"83",
           864 => x"51",
           865 => x"dd",
           866 => x"b2",
           867 => x"7c",
           868 => x"53",
           869 => x"33",
           870 => x"3f",
           871 => x"54",
           872 => x"26",
           873 => x"b8",
           874 => x"c0",
           875 => x"80",
           876 => x"55",
           877 => x"81",
           878 => x"06",
           879 => x"80",
           880 => x"d5",
           881 => x"3f",
           882 => x"38",
           883 => x"78",
           884 => x"9d",
           885 => x"2b",
           886 => x"2e",
           887 => x"c3",
           888 => x"fe",
           889 => x"0c",
           890 => x"51",
           891 => x"ac",
           892 => x"3f",
           893 => x"da",
           894 => x"3f",
           895 => x"54",
           896 => x"27",
           897 => x"7a",
           898 => x"d2",
           899 => x"84",
           900 => x"ea",
           901 => x"fe",
           902 => x"d0",
           903 => x"53",
           904 => x"79",
           905 => x"72",
           906 => x"83",
           907 => x"14",
           908 => x"51",
           909 => x"38",
           910 => x"52",
           911 => x"56",
           912 => x"84",
           913 => x"88",
           914 => x"a0",
           915 => x"06",
           916 => x"39",
           917 => x"c8",
           918 => x"a0",
           919 => x"30",
           920 => x"51",
           921 => x"80",
           922 => x"94",
           923 => x"70",
           924 => x"72",
           925 => x"73",
           926 => x"57",
           927 => x"38",
           928 => x"c8",
           929 => x"0d",
           930 => x"d7",
           931 => x"d3",
           932 => x"9c",
           933 => x"06",
           934 => x"82",
           935 => x"82",
           936 => x"06",
           937 => x"84",
           938 => x"81",
           939 => x"06",
           940 => x"86",
           941 => x"80",
           942 => x"06",
           943 => x"2a",
           944 => x"ef",
           945 => x"9c",
           946 => x"a5",
           947 => x"d7",
           948 => x"9b",
           949 => x"8d",
           950 => x"88",
           951 => x"c6",
           952 => x"3f",
           953 => x"80",
           954 => x"70",
           955 => x"ff",
           956 => x"bd",
           957 => x"3f",
           958 => x"2a",
           959 => x"2e",
           960 => x"51",
           961 => x"9b",
           962 => x"72",
           963 => x"71",
           964 => x"39",
           965 => x"bc",
           966 => x"ed",
           967 => x"51",
           968 => x"ff",
           969 => x"83",
           970 => x"51",
           971 => x"81",
           972 => x"e6",
           973 => x"b5",
           974 => x"3f",
           975 => x"2a",
           976 => x"2e",
           977 => x"3d",
           978 => x"84",
           979 => x"51",
           980 => x"08",
           981 => x"78",
           982 => x"b4",
           983 => x"83",
           984 => x"48",
           985 => x"eb",
           986 => x"33",
           987 => x"80",
           988 => x"83",
           989 => x"7d",
           990 => x"5a",
           991 => x"79",
           992 => x"06",
           993 => x"5a",
           994 => x"7b",
           995 => x"83",
           996 => x"e7",
           997 => x"b9",
           998 => x"52",
           999 => x"08",
          1000 => x"81",
          1001 => x"81",
          1002 => x"c4",
          1003 => x"2e",
          1004 => x"51",
          1005 => x"5e",
          1006 => x"c9",
          1007 => x"3d",
          1008 => x"84",
          1009 => x"5c",
          1010 => x"b9",
          1011 => x"b9",
          1012 => x"81",
          1013 => x"2e",
          1014 => x"e2",
          1015 => x"7b",
          1016 => x"7c",
          1017 => x"58",
          1018 => x"55",
          1019 => x"80",
          1020 => x"84",
          1021 => x"09",
          1022 => x"51",
          1023 => x"26",
          1024 => x"59",
          1025 => x"70",
          1026 => x"95",
          1027 => x"07",
          1028 => x"2e",
          1029 => x"e1",
          1030 => x"3f",
          1031 => x"7e",
          1032 => x"ee",
          1033 => x"59",
          1034 => x"d5",
          1035 => x"88",
          1036 => x"c5",
          1037 => x"bc",
          1038 => x"52",
          1039 => x"b9",
          1040 => x"b9",
          1041 => x"0b",
          1042 => x"06",
          1043 => x"06",
          1044 => x"d8",
          1045 => x"0b",
          1046 => x"a8",
          1047 => x"d4",
          1048 => x"b7",
          1049 => x"85",
          1050 => x"fd",
          1051 => x"d4",
          1052 => x"83",
          1053 => x"3f",
          1054 => x"51",
          1055 => x"08",
          1056 => x"38",
          1057 => x"fb",
          1058 => x"db",
          1059 => x"fe",
          1060 => x"55",
          1061 => x"d6",
          1062 => x"fd",
          1063 => x"ff",
          1064 => x"81",
          1065 => x"ef",
          1066 => x"39",
          1067 => x"80",
          1068 => x"de",
          1069 => x"39",
          1070 => x"80",
          1071 => x"c8",
          1072 => x"52",
          1073 => x"68",
          1074 => x"80",
          1075 => x"08",
          1076 => x"3f",
          1077 => x"11",
          1078 => x"3f",
          1079 => x"ff",
          1080 => x"d0",
          1081 => x"3d",
          1082 => x"51",
          1083 => x"80",
          1084 => x"f0",
          1085 => x"92",
          1086 => x"38",
          1087 => x"83",
          1088 => x"d5",
          1089 => x"51",
          1090 => x"59",
          1091 => x"9f",
          1092 => x"70",
          1093 => x"f4",
          1094 => x"ca",
          1095 => x"f8",
          1096 => x"53",
          1097 => x"84",
          1098 => x"59",
          1099 => x"b8",
          1100 => x"08",
          1101 => x"b3",
          1102 => x"ae",
          1103 => x"87",
          1104 => x"59",
          1105 => x"53",
          1106 => x"84",
          1107 => x"38",
          1108 => x"80",
          1109 => x"c8",
          1110 => x"3d",
          1111 => x"51",
          1112 => x"80",
          1113 => x"51",
          1114 => x"78",
          1115 => x"33",
          1116 => x"2e",
          1117 => x"33",
          1118 => x"ce",
          1119 => x"19",
          1120 => x"3d",
          1121 => x"51",
          1122 => x"80",
          1123 => x"fc",
          1124 => x"de",
          1125 => x"f7",
          1126 => x"53",
          1127 => x"84",
          1128 => x"38",
          1129 => x"68",
          1130 => x"65",
          1131 => x"7c",
          1132 => x"b8",
          1133 => x"05",
          1134 => x"08",
          1135 => x"fe",
          1136 => x"e7",
          1137 => x"38",
          1138 => x"fc",
          1139 => x"08",
          1140 => x"fb",
          1141 => x"ae",
          1142 => x"84",
          1143 => x"39",
          1144 => x"79",
          1145 => x"fe",
          1146 => x"e7",
          1147 => x"2e",
          1148 => x"db",
          1149 => x"49",
          1150 => x"80",
          1151 => x"c8",
          1152 => x"b8",
          1153 => x"05",
          1154 => x"08",
          1155 => x"fe",
          1156 => x"e6",
          1157 => x"2e",
          1158 => x"11",
          1159 => x"3f",
          1160 => x"b9",
          1161 => x"cb",
          1162 => x"7a",
          1163 => x"70",
          1164 => x"f5",
          1165 => x"cf",
          1166 => x"87",
          1167 => x"3d",
          1168 => x"3f",
          1169 => x"78",
          1170 => x"08",
          1171 => x"c8",
          1172 => x"39",
          1173 => x"80",
          1174 => x"c8",
          1175 => x"5a",
          1176 => x"f2",
          1177 => x"11",
          1178 => x"3f",
          1179 => x"f2",
          1180 => x"8a",
          1181 => x"3d",
          1182 => x"51",
          1183 => x"80",
          1184 => x"7a",
          1185 => x"90",
          1186 => x"2a",
          1187 => x"2e",
          1188 => x"88",
          1189 => x"3f",
          1190 => x"52",
          1191 => x"a4",
          1192 => x"64",
          1193 => x"45",
          1194 => x"80",
          1195 => x"c8",
          1196 => x"64",
          1197 => x"b8",
          1198 => x"05",
          1199 => x"08",
          1200 => x"02",
          1201 => x"05",
          1202 => x"f0",
          1203 => x"e2",
          1204 => x"f2",
          1205 => x"05",
          1206 => x"7d",
          1207 => x"ff",
          1208 => x"b9",
          1209 => x"39",
          1210 => x"80",
          1211 => x"c8",
          1212 => x"5c",
          1213 => x"68",
          1214 => x"3d",
          1215 => x"51",
          1216 => x"80",
          1217 => x"0c",
          1218 => x"f7",
          1219 => x"06",
          1220 => x"90",
          1221 => x"7c",
          1222 => x"7b",
          1223 => x"8c",
          1224 => x"3f",
          1225 => x"11",
          1226 => x"3f",
          1227 => x"38",
          1228 => x"79",
          1229 => x"f7",
          1230 => x"7b",
          1231 => x"90",
          1232 => x"cd",
          1233 => x"83",
          1234 => x"83",
          1235 => x"59",
          1236 => x"d3",
          1237 => x"83",
          1238 => x"a5",
          1239 => x"8b",
          1240 => x"3f",
          1241 => x"59",
          1242 => x"98",
          1243 => x"cf",
          1244 => x"83",
          1245 => x"83",
          1246 => x"9b",
          1247 => x"ee",
          1248 => x"80",
          1249 => x"49",
          1250 => x"5d",
          1251 => x"a8",
          1252 => x"b4",
          1253 => x"39",
          1254 => x"fb",
          1255 => x"84",
          1256 => x"70",
          1257 => x"74",
          1258 => x"08",
          1259 => x"84",
          1260 => x"74",
          1261 => x"87",
          1262 => x"87",
          1263 => x"3f",
          1264 => x"08",
          1265 => x"51",
          1266 => x"08",
          1267 => x"87",
          1268 => x"0b",
          1269 => x"f2",
          1270 => x"84",
          1271 => x"d5",
          1272 => x"0c",
          1273 => x"56",
          1274 => x"97",
          1275 => x"83",
          1276 => x"c4",
          1277 => x"52",
          1278 => x"54",
          1279 => x"52",
          1280 => x"8d",
          1281 => x"e3",
          1282 => x"c3",
          1283 => x"d3",
          1284 => x"3f",
          1285 => x"08",
          1286 => x"73",
          1287 => x"81",
          1288 => x"09",
          1289 => x"33",
          1290 => x"70",
          1291 => x"06",
          1292 => x"74",
          1293 => x"80",
          1294 => x"54",
          1295 => x"54",
          1296 => x"2e",
          1297 => x"80",
          1298 => x"a0",
          1299 => x"54",
          1300 => x"25",
          1301 => x"2e",
          1302 => x"54",
          1303 => x"84",
          1304 => x"70",
          1305 => x"ff",
          1306 => x"33",
          1307 => x"70",
          1308 => x"39",
          1309 => x"72",
          1310 => x"38",
          1311 => x"72",
          1312 => x"c8",
          1313 => x"fc",
          1314 => x"84",
          1315 => x"74",
          1316 => x"04",
          1317 => x"ff",
          1318 => x"26",
          1319 => x"05",
          1320 => x"8a",
          1321 => x"70",
          1322 => x"33",
          1323 => x"f2",
          1324 => x"74",
          1325 => x"22",
          1326 => x"80",
          1327 => x"52",
          1328 => x"81",
          1329 => x"22",
          1330 => x"33",
          1331 => x"33",
          1332 => x"33",
          1333 => x"33",
          1334 => x"33",
          1335 => x"c0",
          1336 => x"a0",
          1337 => x"0c",
          1338 => x"86",
          1339 => x"5b",
          1340 => x"0c",
          1341 => x"7b",
          1342 => x"7b",
          1343 => x"08",
          1344 => x"98",
          1345 => x"87",
          1346 => x"1c",
          1347 => x"7b",
          1348 => x"08",
          1349 => x"98",
          1350 => x"80",
          1351 => x"59",
          1352 => x"1b",
          1353 => x"1b",
          1354 => x"1b",
          1355 => x"52",
          1356 => x"3f",
          1357 => x"02",
          1358 => x"a8",
          1359 => x"84",
          1360 => x"2c",
          1361 => x"06",
          1362 => x"71",
          1363 => x"04",
          1364 => x"b9",
          1365 => x"51",
          1366 => x"df",
          1367 => x"84",
          1368 => x"2c",
          1369 => x"c7",
          1370 => x"52",
          1371 => x"e7",
          1372 => x"2b",
          1373 => x"2e",
          1374 => x"54",
          1375 => x"84",
          1376 => x"fc",
          1377 => x"f2",
          1378 => x"55",
          1379 => x"87",
          1380 => x"70",
          1381 => x"2e",
          1382 => x"06",
          1383 => x"32",
          1384 => x"38",
          1385 => x"cf",
          1386 => x"c0",
          1387 => x"38",
          1388 => x"0c",
          1389 => x"0d",
          1390 => x"51",
          1391 => x"81",
          1392 => x"71",
          1393 => x"2e",
          1394 => x"70",
          1395 => x"52",
          1396 => x"0d",
          1397 => x"9f",
          1398 => x"80",
          1399 => x"0d",
          1400 => x"52",
          1401 => x"81",
          1402 => x"ff",
          1403 => x"80",
          1404 => x"70",
          1405 => x"52",
          1406 => x"2a",
          1407 => x"38",
          1408 => x"80",
          1409 => x"06",
          1410 => x"06",
          1411 => x"80",
          1412 => x"52",
          1413 => x"55",
          1414 => x"b9",
          1415 => x"91",
          1416 => x"98",
          1417 => x"72",
          1418 => x"81",
          1419 => x"38",
          1420 => x"2a",
          1421 => x"ce",
          1422 => x"c0",
          1423 => x"06",
          1424 => x"38",
          1425 => x"84",
          1426 => x"f2",
          1427 => x"83",
          1428 => x"08",
          1429 => x"9c",
          1430 => x"9e",
          1431 => x"c0",
          1432 => x"87",
          1433 => x"0c",
          1434 => x"a4",
          1435 => x"f2",
          1436 => x"83",
          1437 => x"08",
          1438 => x"c4",
          1439 => x"9e",
          1440 => x"23",
          1441 => x"bc",
          1442 => x"f2",
          1443 => x"83",
          1444 => x"c8",
          1445 => x"08",
          1446 => x"52",
          1447 => x"c9",
          1448 => x"08",
          1449 => x"52",
          1450 => x"71",
          1451 => x"c0",
          1452 => x"06",
          1453 => x"38",
          1454 => x"80",
          1455 => x"88",
          1456 => x"80",
          1457 => x"f2",
          1458 => x"90",
          1459 => x"52",
          1460 => x"52",
          1461 => x"87",
          1462 => x"80",
          1463 => x"83",
          1464 => x"34",
          1465 => x"70",
          1466 => x"70",
          1467 => x"83",
          1468 => x"9e",
          1469 => x"51",
          1470 => x"81",
          1471 => x"0b",
          1472 => x"80",
          1473 => x"2e",
          1474 => x"d1",
          1475 => x"08",
          1476 => x"52",
          1477 => x"71",
          1478 => x"c0",
          1479 => x"51",
          1480 => x"81",
          1481 => x"c0",
          1482 => x"8a",
          1483 => x"34",
          1484 => x"70",
          1485 => x"80",
          1486 => x"f2",
          1487 => x"83",
          1488 => x"71",
          1489 => x"c0",
          1490 => x"52",
          1491 => x"52",
          1492 => x"9e",
          1493 => x"f2",
          1494 => x"52",
          1495 => x"d9",
          1496 => x"f2",
          1497 => x"83",
          1498 => x"f2",
          1499 => x"83",
          1500 => x"38",
          1501 => x"9d",
          1502 => x"84",
          1503 => x"73",
          1504 => x"56",
          1505 => x"33",
          1506 => x"d5",
          1507 => x"f2",
          1508 => x"83",
          1509 => x"38",
          1510 => x"88",
          1511 => x"82",
          1512 => x"73",
          1513 => x"c2",
          1514 => x"83",
          1515 => x"83",
          1516 => x"51",
          1517 => x"08",
          1518 => x"90",
          1519 => x"3f",
          1520 => x"bc",
          1521 => x"bc",
          1522 => x"51",
          1523 => x"bd",
          1524 => x"54",
          1525 => x"e4",
          1526 => x"cf",
          1527 => x"ca",
          1528 => x"0d",
          1529 => x"84",
          1530 => x"84",
          1531 => x"76",
          1532 => x"08",
          1533 => x"98",
          1534 => x"c0",
          1535 => x"51",
          1536 => x"bd",
          1537 => x"54",
          1538 => x"bc",
          1539 => x"ca",
          1540 => x"38",
          1541 => x"c0",
          1542 => x"bb",
          1543 => x"d9",
          1544 => x"f2",
          1545 => x"ff",
          1546 => x"52",
          1547 => x"3f",
          1548 => x"83",
          1549 => x"51",
          1550 => x"08",
          1551 => x"c8",
          1552 => x"84",
          1553 => x"84",
          1554 => x"51",
          1555 => x"33",
          1556 => x"fe",
          1557 => x"bf",
          1558 => x"73",
          1559 => x"39",
          1560 => x"3f",
          1561 => x"2e",
          1562 => x"84",
          1563 => x"d0",
          1564 => x"38",
          1565 => x"bf",
          1566 => x"73",
          1567 => x"83",
          1568 => x"51",
          1569 => x"33",
          1570 => x"d2",
          1571 => x"dc",
          1572 => x"f2",
          1573 => x"ee",
          1574 => x"52",
          1575 => x"3f",
          1576 => x"2e",
          1577 => x"94",
          1578 => x"52",
          1579 => x"3f",
          1580 => x"2e",
          1581 => x"8c",
          1582 => x"52",
          1583 => x"3f",
          1584 => x"2e",
          1585 => x"84",
          1586 => x"52",
          1587 => x"3f",
          1588 => x"2e",
          1589 => x"9c",
          1590 => x"52",
          1591 => x"3f",
          1592 => x"2e",
          1593 => x"a4",
          1594 => x"52",
          1595 => x"3f",
          1596 => x"2e",
          1597 => x"90",
          1598 => x"98",
          1599 => x"ca",
          1600 => x"38",
          1601 => x"05",
          1602 => x"71",
          1603 => x"71",
          1604 => x"af",
          1605 => x"de",
          1606 => x"3d",
          1607 => x"af",
          1608 => x"de",
          1609 => x"3d",
          1610 => x"af",
          1611 => x"de",
          1612 => x"3d",
          1613 => x"80",
          1614 => x"83",
          1615 => x"0c",
          1616 => x"ad",
          1617 => x"58",
          1618 => x"82",
          1619 => x"80",
          1620 => x"83",
          1621 => x"52",
          1622 => x"b9",
          1623 => x"51",
          1624 => x"81",
          1625 => x"c8",
          1626 => x"08",
          1627 => x"74",
          1628 => x"07",
          1629 => x"2e",
          1630 => x"f3",
          1631 => x"82",
          1632 => x"8f",
          1633 => x"84",
          1634 => x"83",
          1635 => x"78",
          1636 => x"76",
          1637 => x"51",
          1638 => x"56",
          1639 => x"52",
          1640 => x"3f",
          1641 => x"3d",
          1642 => x"08",
          1643 => x"33",
          1644 => x"81",
          1645 => x"56",
          1646 => x"05",
          1647 => x"3f",
          1648 => x"73",
          1649 => x"c8",
          1650 => x"73",
          1651 => x"2e",
          1652 => x"06",
          1653 => x"80",
          1654 => x"3d",
          1655 => x"ff",
          1656 => x"c7",
          1657 => x"2e",
          1658 => x"76",
          1659 => x"08",
          1660 => x"c9",
          1661 => x"57",
          1662 => x"ff",
          1663 => x"76",
          1664 => x"70",
          1665 => x"2e",
          1666 => x"75",
          1667 => x"59",
          1668 => x"c8",
          1669 => x"56",
          1670 => x"08",
          1671 => x"53",
          1672 => x"fd",
          1673 => x"ba",
          1674 => x"84",
          1675 => x"b9",
          1676 => x"c8",
          1677 => x"80",
          1678 => x"16",
          1679 => x"88",
          1680 => x"ff",
          1681 => x"0c",
          1682 => x"b5",
          1683 => x"08",
          1684 => x"34",
          1685 => x"08",
          1686 => x"f3",
          1687 => x"82",
          1688 => x"38",
          1689 => x"90",
          1690 => x"38",
          1691 => x"51",
          1692 => x"98",
          1693 => x"ff",
          1694 => x"84",
          1695 => x"98",
          1696 => x"2b",
          1697 => x"70",
          1698 => x"08",
          1699 => x"46",
          1700 => x"74",
          1701 => x"27",
          1702 => x"29",
          1703 => x"57",
          1704 => x"75",
          1705 => x"80",
          1706 => x"57",
          1707 => x"d0",
          1708 => x"78",
          1709 => x"2e",
          1710 => x"81",
          1711 => x"81",
          1712 => x"84",
          1713 => x"97",
          1714 => x"2b",
          1715 => x"5f",
          1716 => x"2e",
          1717 => x"34",
          1718 => x"ba",
          1719 => x"80",
          1720 => x"ff",
          1721 => x"80",
          1722 => x"2b",
          1723 => x"16",
          1724 => x"38",
          1725 => x"33",
          1726 => x"38",
          1727 => x"f2",
          1728 => x"ab",
          1729 => x"b2",
          1730 => x"76",
          1731 => x"80",
          1732 => x"62",
          1733 => x"74",
          1734 => x"76",
          1735 => x"7f",
          1736 => x"80",
          1737 => x"84",
          1738 => x"fd",
          1739 => x"88",
          1740 => x"8c",
          1741 => x"8c",
          1742 => x"33",
          1743 => x"33",
          1744 => x"d6",
          1745 => x"15",
          1746 => x"16",
          1747 => x"3f",
          1748 => x"da",
          1749 => x"05",
          1750 => x"38",
          1751 => x"34",
          1752 => x"33",
          1753 => x"84",
          1754 => x"b5",
          1755 => x"a0",
          1756 => x"ac",
          1757 => x"3f",
          1758 => x"7a",
          1759 => x"06",
          1760 => x"a5",
          1761 => x"fb",
          1762 => x"ac",
          1763 => x"10",
          1764 => x"08",
          1765 => x"08",
          1766 => x"75",
          1767 => x"c8",
          1768 => x"c8",
          1769 => x"75",
          1770 => x"84",
          1771 => x"56",
          1772 => x"84",
          1773 => x"b3",
          1774 => x"a0",
          1775 => x"ac",
          1776 => x"3f",
          1777 => x"74",
          1778 => x"06",
          1779 => x"70",
          1780 => x"5b",
          1781 => x"38",
          1782 => x"57",
          1783 => x"70",
          1784 => x"84",
          1785 => x"84",
          1786 => x"78",
          1787 => x"08",
          1788 => x"8c",
          1789 => x"ff",
          1790 => x"70",
          1791 => x"5a",
          1792 => x"38",
          1793 => x"84",
          1794 => x"2e",
          1795 => x"84",
          1796 => x"98",
          1797 => x"5a",
          1798 => x"d5",
          1799 => x"ae",
          1800 => x"2b",
          1801 => x"5a",
          1802 => x"86",
          1803 => x"51",
          1804 => x"0a",
          1805 => x"2c",
          1806 => x"74",
          1807 => x"ac",
          1808 => x"3f",
          1809 => x"0a",
          1810 => x"33",
          1811 => x"b9",
          1812 => x"81",
          1813 => x"08",
          1814 => x"3f",
          1815 => x"0a",
          1816 => x"33",
          1817 => x"e6",
          1818 => x"78",
          1819 => x"33",
          1820 => x"80",
          1821 => x"98",
          1822 => x"55",
          1823 => x"b6",
          1824 => x"80",
          1825 => x"08",
          1826 => x"84",
          1827 => x"84",
          1828 => x"55",
          1829 => x"05",
          1830 => x"08",
          1831 => x"84",
          1832 => x"3f",
          1833 => x"58",
          1834 => x"33",
          1835 => x"83",
          1836 => x"f2",
          1837 => x"74",
          1838 => x"fc",
          1839 => x"70",
          1840 => x"84",
          1841 => x"b8",
          1842 => x"05",
          1843 => x"ad",
          1844 => x"80",
          1845 => x"58",
          1846 => x"0b",
          1847 => x"d1",
          1848 => x"b4",
          1849 => x"55",
          1850 => x"ac",
          1851 => x"3f",
          1852 => x"ff",
          1853 => x"52",
          1854 => x"d1",
          1855 => x"d1",
          1856 => x"74",
          1857 => x"9f",
          1858 => x"34",
          1859 => x"be",
          1860 => x"1d",
          1861 => x"80",
          1862 => x"52",
          1863 => x"d5",
          1864 => x"a6",
          1865 => x"51",
          1866 => x"33",
          1867 => x"34",
          1868 => x"38",
          1869 => x"3f",
          1870 => x"0b",
          1871 => x"c8",
          1872 => x"8c",
          1873 => x"7a",
          1874 => x"88",
          1875 => x"88",
          1876 => x"8c",
          1877 => x"51",
          1878 => x"33",
          1879 => x"d1",
          1880 => x"76",
          1881 => x"08",
          1882 => x"84",
          1883 => x"98",
          1884 => x"59",
          1885 => x"84",
          1886 => x"ac",
          1887 => x"81",
          1888 => x"d1",
          1889 => x"24",
          1890 => x"52",
          1891 => x"81",
          1892 => x"70",
          1893 => x"51",
          1894 => x"f3",
          1895 => x"33",
          1896 => x"76",
          1897 => x"81",
          1898 => x"70",
          1899 => x"57",
          1900 => x"7b",
          1901 => x"84",
          1902 => x"ff",
          1903 => x"29",
          1904 => x"84",
          1905 => x"76",
          1906 => x"84",
          1907 => x"58",
          1908 => x"84",
          1909 => x"ae",
          1910 => x"57",
          1911 => x"16",
          1912 => x"81",
          1913 => x"70",
          1914 => x"57",
          1915 => x"18",
          1916 => x"81",
          1917 => x"33",
          1918 => x"76",
          1919 => x"75",
          1920 => x"d1",
          1921 => x"81",
          1922 => x"81",
          1923 => x"76",
          1924 => x"70",
          1925 => x"57",
          1926 => x"84",
          1927 => x"aa",
          1928 => x"81",
          1929 => x"d1",
          1930 => x"25",
          1931 => x"52",
          1932 => x"81",
          1933 => x"70",
          1934 => x"57",
          1935 => x"f0",
          1936 => x"75",
          1937 => x"ff",
          1938 => x"84",
          1939 => x"81",
          1940 => x"7b",
          1941 => x"88",
          1942 => x"74",
          1943 => x"ac",
          1944 => x"3f",
          1945 => x"ff",
          1946 => x"52",
          1947 => x"d1",
          1948 => x"d1",
          1949 => x"c7",
          1950 => x"84",
          1951 => x"84",
          1952 => x"83",
          1953 => x"80",
          1954 => x"7b",
          1955 => x"ce",
          1956 => x"80",
          1957 => x"88",
          1958 => x"da",
          1959 => x"2b",
          1960 => x"5d",
          1961 => x"8e",
          1962 => x"08",
          1963 => x"e0",
          1964 => x"bb",
          1965 => x"75",
          1966 => x"f3",
          1967 => x"74",
          1968 => x"81",
          1969 => x"51",
          1970 => x"f3",
          1971 => x"5f",
          1972 => x"e9",
          1973 => x"18",
          1974 => x"38",
          1975 => x"e8",
          1976 => x"88",
          1977 => x"06",
          1978 => x"ff",
          1979 => x"88",
          1980 => x"5d",
          1981 => x"d5",
          1982 => x"f6",
          1983 => x"51",
          1984 => x"08",
          1985 => x"84",
          1986 => x"84",
          1987 => x"55",
          1988 => x"84",
          1989 => x"88",
          1990 => x"3d",
          1991 => x"3f",
          1992 => x"34",
          1993 => x"81",
          1994 => x"aa",
          1995 => x"06",
          1996 => x"33",
          1997 => x"f1",
          1998 => x"88",
          1999 => x"ac",
          2000 => x"3f",
          2001 => x"ff",
          2002 => x"ff",
          2003 => x"76",
          2004 => x"51",
          2005 => x"08",
          2006 => x"08",
          2007 => x"52",
          2008 => x"1d",
          2009 => x"33",
          2010 => x"58",
          2011 => x"d5",
          2012 => x"86",
          2013 => x"51",
          2014 => x"08",
          2015 => x"84",
          2016 => x"84",
          2017 => x"55",
          2018 => x"3f",
          2019 => x"87",
          2020 => x"19",
          2021 => x"d1",
          2022 => x"83",
          2023 => x"f2",
          2024 => x"74",
          2025 => x"7b",
          2026 => x"83",
          2027 => x"ff",
          2028 => x"f2",
          2029 => x"b1",
          2030 => x"76",
          2031 => x"c0",
          2032 => x"51",
          2033 => x"08",
          2034 => x"84",
          2035 => x"88",
          2036 => x"3d",
          2037 => x"b9",
          2038 => x"84",
          2039 => x"b9",
          2040 => x"f3",
          2041 => x"51",
          2042 => x"08",
          2043 => x"09",
          2044 => x"c8",
          2045 => x"b9",
          2046 => x"c8",
          2047 => x"c8",
          2048 => x"80",
          2049 => x"f3",
          2050 => x"e0",
          2051 => x"74",
          2052 => x"fc",
          2053 => x"70",
          2054 => x"84",
          2055 => x"b8",
          2056 => x"05",
          2057 => x"38",
          2058 => x"57",
          2059 => x"75",
          2060 => x"38",
          2061 => x"76",
          2062 => x"f2",
          2063 => x"70",
          2064 => x"27",
          2065 => x"b8",
          2066 => x"d3",
          2067 => x"82",
          2068 => x"05",
          2069 => x"80",
          2070 => x"75",
          2071 => x"10",
          2072 => x"40",
          2073 => x"ff",
          2074 => x"fe",
          2075 => x"f1",
          2076 => x"9f",
          2077 => x"e4",
          2078 => x"05",
          2079 => x"33",
          2080 => x"38",
          2081 => x"73",
          2082 => x"82",
          2083 => x"86",
          2084 => x"56",
          2085 => x"38",
          2086 => x"f8",
          2087 => x"83",
          2088 => x"90",
          2089 => x"07",
          2090 => x"77",
          2091 => x"05",
          2092 => x"55",
          2093 => x"78",
          2094 => x"84",
          2095 => x"55",
          2096 => x"74",
          2097 => x"13",
          2098 => x"04",
          2099 => x"f8",
          2100 => x"f9",
          2101 => x"5b",
          2102 => x"80",
          2103 => x"ff",
          2104 => x"ff",
          2105 => x"ff",
          2106 => x"5d",
          2107 => x"26",
          2108 => x"56",
          2109 => x"06",
          2110 => x"ff",
          2111 => x"29",
          2112 => x"74",
          2113 => x"33",
          2114 => x"1b",
          2115 => x"80",
          2116 => x"53",
          2117 => x"73",
          2118 => x"f4",
          2119 => x"e8",
          2120 => x"a7",
          2121 => x"70",
          2122 => x"70",
          2123 => x"70",
          2124 => x"56",
          2125 => x"38",
          2126 => x"06",
          2127 => x"79",
          2128 => x"83",
          2129 => x"f9",
          2130 => x"2b",
          2131 => x"07",
          2132 => x"5b",
          2133 => x"be",
          2134 => x"f8",
          2135 => x"10",
          2136 => x"29",
          2137 => x"57",
          2138 => x"80",
          2139 => x"81",
          2140 => x"81",
          2141 => x"83",
          2142 => x"05",
          2143 => x"5e",
          2144 => x"7a",
          2145 => x"53",
          2146 => x"06",
          2147 => x"06",
          2148 => x"58",
          2149 => x"26",
          2150 => x"73",
          2151 => x"79",
          2152 => x"7b",
          2153 => x"78",
          2154 => x"fb",
          2155 => x"ff",
          2156 => x"73",
          2157 => x"9c",
          2158 => x"75",
          2159 => x"76",
          2160 => x"94",
          2161 => x"ff",
          2162 => x"fa",
          2163 => x"08",
          2164 => x"81",
          2165 => x"55",
          2166 => x"ff",
          2167 => x"75",
          2168 => x"77",
          2169 => x"a0",
          2170 => x"06",
          2171 => x"d0",
          2172 => x"84",
          2173 => x"84",
          2174 => x"04",
          2175 => x"02",
          2176 => x"bb",
          2177 => x"79",
          2178 => x"33",
          2179 => x"33",
          2180 => x"80",
          2181 => x"57",
          2182 => x"ff",
          2183 => x"57",
          2184 => x"38",
          2185 => x"74",
          2186 => x"33",
          2187 => x"81",
          2188 => x"26",
          2189 => x"83",
          2190 => x"70",
          2191 => x"33",
          2192 => x"89",
          2193 => x"29",
          2194 => x"26",
          2195 => x"54",
          2196 => x"16",
          2197 => x"75",
          2198 => x"54",
          2199 => x"73",
          2200 => x"f4",
          2201 => x"a0",
          2202 => x"70",
          2203 => x"9f",
          2204 => x"ba",
          2205 => x"f6",
          2206 => x"77",
          2207 => x"73",
          2208 => x"81",
          2209 => x"29",
          2210 => x"a0",
          2211 => x"81",
          2212 => x"71",
          2213 => x"79",
          2214 => x"54",
          2215 => x"c4",
          2216 => x"34",
          2217 => x"70",
          2218 => x"b7",
          2219 => x"71",
          2220 => x"75",
          2221 => x"b9",
          2222 => x"83",
          2223 => x"70",
          2224 => x"33",
          2225 => x"f9",
          2226 => x"78",
          2227 => x"f8",
          2228 => x"81",
          2229 => x"81",
          2230 => x"29",
          2231 => x"54",
          2232 => x"f8",
          2233 => x"76",
          2234 => x"e0",
          2235 => x"57",
          2236 => x"fe",
          2237 => x"34",
          2238 => x"ff",
          2239 => x"39",
          2240 => x"56",
          2241 => x"33",
          2242 => x"34",
          2243 => x"39",
          2244 => x"9f",
          2245 => x"9b",
          2246 => x"05",
          2247 => x"33",
          2248 => x"83",
          2249 => x"c8",
          2250 => x"83",
          2251 => x"70",
          2252 => x"2e",
          2253 => x"f8",
          2254 => x"0c",
          2255 => x"33",
          2256 => x"2c",
          2257 => x"83",
          2258 => x"f8",
          2259 => x"ff",
          2260 => x"83",
          2261 => x"34",
          2262 => x"3d",
          2263 => x"73",
          2264 => x"06",
          2265 => x"f9",
          2266 => x"86",
          2267 => x"72",
          2268 => x"55",
          2269 => x"70",
          2270 => x"0b",
          2271 => x"04",
          2272 => x"f8",
          2273 => x"05",
          2274 => x"38",
          2275 => x"34",
          2276 => x"8f",
          2277 => x"38",
          2278 => x"51",
          2279 => x"70",
          2280 => x"f0",
          2281 => x"52",
          2282 => x"81",
          2283 => x"f8",
          2284 => x"0c",
          2285 => x"33",
          2286 => x"83",
          2287 => x"c8",
          2288 => x"f4",
          2289 => x"f8",
          2290 => x"33",
          2291 => x"83",
          2292 => x"0b",
          2293 => x"b9",
          2294 => x"f8",
          2295 => x"51",
          2296 => x"39",
          2297 => x"70",
          2298 => x"83",
          2299 => x"07",
          2300 => x"93",
          2301 => x"06",
          2302 => x"34",
          2303 => x"81",
          2304 => x"f8",
          2305 => x"f4",
          2306 => x"f8",
          2307 => x"f4",
          2308 => x"51",
          2309 => x"39",
          2310 => x"b0",
          2311 => x"fe",
          2312 => x"ef",
          2313 => x"f8",
          2314 => x"f4",
          2315 => x"51",
          2316 => x"39",
          2317 => x"a0",
          2318 => x"fe",
          2319 => x"8f",
          2320 => x"fd",
          2321 => x"fa",
          2322 => x"f4",
          2323 => x"02",
          2324 => x"c3",
          2325 => x"f8",
          2326 => x"b7",
          2327 => x"59",
          2328 => x"82",
          2329 => x"82",
          2330 => x"0b",
          2331 => x"f8",
          2332 => x"83",
          2333 => x"78",
          2334 => x"80",
          2335 => x"84",
          2336 => x"f8",
          2337 => x"82",
          2338 => x"84",
          2339 => x"33",
          2340 => x"54",
          2341 => x"51",
          2342 => x"be",
          2343 => x"7a",
          2344 => x"f6",
          2345 => x"3d",
          2346 => x"34",
          2347 => x"0b",
          2348 => x"f8",
          2349 => x"23",
          2350 => x"ca",
          2351 => x"79",
          2352 => x"83",
          2353 => x"80",
          2354 => x"79",
          2355 => x"b9",
          2356 => x"e3",
          2357 => x"1a",
          2358 => x"33",
          2359 => x"38",
          2360 => x"3f",
          2361 => x"84",
          2362 => x"34",
          2363 => x"f8",
          2364 => x"0b",
          2365 => x"b7",
          2366 => x"34",
          2367 => x"0b",
          2368 => x"51",
          2369 => x"08",
          2370 => x"f0",
          2371 => x"ff",
          2372 => x"08",
          2373 => x"19",
          2374 => x"ff",
          2375 => x"06",
          2376 => x"7a",
          2377 => x"b7",
          2378 => x"f8",
          2379 => x"a7",
          2380 => x"53",
          2381 => x"70",
          2382 => x"33",
          2383 => x"81",
          2384 => x"81",
          2385 => x"38",
          2386 => x"88",
          2387 => x"33",
          2388 => x"33",
          2389 => x"84",
          2390 => x"80",
          2391 => x"f8",
          2392 => x"71",
          2393 => x"83",
          2394 => x"33",
          2395 => x"f8",
          2396 => x"34",
          2397 => x"06",
          2398 => x"33",
          2399 => x"55",
          2400 => x"9a",
          2401 => x"06",
          2402 => x"38",
          2403 => x"ea",
          2404 => x"f9",
          2405 => x"80",
          2406 => x"57",
          2407 => x"0b",
          2408 => x"04",
          2409 => x"24",
          2410 => x"81",
          2411 => x"51",
          2412 => x"f9",
          2413 => x"15",
          2414 => x"74",
          2415 => x"fe",
          2416 => x"51",
          2417 => x"ff",
          2418 => x"91",
          2419 => x"3f",
          2420 => x"54",
          2421 => x"39",
          2422 => x"39",
          2423 => x"80",
          2424 => x"0d",
          2425 => x"06",
          2426 => x"70",
          2427 => x"73",
          2428 => x"f9",
          2429 => x"3f",
          2430 => x"06",
          2431 => x"38",
          2432 => x"fe",
          2433 => x"34",
          2434 => x"fe",
          2435 => x"d8",
          2436 => x"02",
          2437 => x"08",
          2438 => x"38",
          2439 => x"8a",
          2440 => x"82",
          2441 => x"38",
          2442 => x"b7",
          2443 => x"f8",
          2444 => x"5e",
          2445 => x"a7",
          2446 => x"33",
          2447 => x"22",
          2448 => x"40",
          2449 => x"f8",
          2450 => x"40",
          2451 => x"a7",
          2452 => x"33",
          2453 => x"22",
          2454 => x"11",
          2455 => x"f4",
          2456 => x"1d",
          2457 => x"61",
          2458 => x"33",
          2459 => x"56",
          2460 => x"84",
          2461 => x"78",
          2462 => x"25",
          2463 => x"b3",
          2464 => x"38",
          2465 => x"b7",
          2466 => x"f8",
          2467 => x"40",
          2468 => x"a7",
          2469 => x"33",
          2470 => x"22",
          2471 => x"56",
          2472 => x"f8",
          2473 => x"57",
          2474 => x"80",
          2475 => x"81",
          2476 => x"f8",
          2477 => x"42",
          2478 => x"60",
          2479 => x"58",
          2480 => x"27",
          2481 => x"34",
          2482 => x"3d",
          2483 => x"38",
          2484 => x"8d",
          2485 => x"80",
          2486 => x"84",
          2487 => x"78",
          2488 => x"56",
          2489 => x"b8",
          2490 => x"84",
          2491 => x"18",
          2492 => x"0b",
          2493 => x"84",
          2494 => x"78",
          2495 => x"84",
          2496 => x"83",
          2497 => x"72",
          2498 => x"b7",
          2499 => x"1d",
          2500 => x"f9",
          2501 => x"29",
          2502 => x"f8",
          2503 => x"76",
          2504 => x"f4",
          2505 => x"84",
          2506 => x"83",
          2507 => x"72",
          2508 => x"59",
          2509 => x"9a",
          2510 => x"39",
          2511 => x"80",
          2512 => x"39",
          2513 => x"33",
          2514 => x"33",
          2515 => x"80",
          2516 => x"5d",
          2517 => x"ff",
          2518 => x"59",
          2519 => x"38",
          2520 => x"57",
          2521 => x"83",
          2522 => x"0b",
          2523 => x"b8",
          2524 => x"34",
          2525 => x"0b",
          2526 => x"b9",
          2527 => x"f8",
          2528 => x"f8",
          2529 => x"f8",
          2530 => x"0b",
          2531 => x"b9",
          2532 => x"80",
          2533 => x"38",
          2534 => x"33",
          2535 => x"33",
          2536 => x"11",
          2537 => x"f6",
          2538 => x"70",
          2539 => x"33",
          2540 => x"7d",
          2541 => x"ff",
          2542 => x"38",
          2543 => x"7b",
          2544 => x"78",
          2545 => x"5f",
          2546 => x"a7",
          2547 => x"33",
          2548 => x"22",
          2549 => x"40",
          2550 => x"83",
          2551 => x"05",
          2552 => x"a7",
          2553 => x"33",
          2554 => x"22",
          2555 => x"11",
          2556 => x"f4",
          2557 => x"81",
          2558 => x"7c",
          2559 => x"bd",
          2560 => x"19",
          2561 => x"f8",
          2562 => x"ff",
          2563 => x"2e",
          2564 => x"d7",
          2565 => x"84",
          2566 => x"38",
          2567 => x"84",
          2568 => x"d0",
          2569 => x"83",
          2570 => x"e7",
          2571 => x"0c",
          2572 => x"33",
          2573 => x"06",
          2574 => x"06",
          2575 => x"80",
          2576 => x"72",
          2577 => x"06",
          2578 => x"5c",
          2579 => x"ef",
          2580 => x"7a",
          2581 => x"72",
          2582 => x"b7",
          2583 => x"34",
          2584 => x"33",
          2585 => x"12",
          2586 => x"f8",
          2587 => x"76",
          2588 => x"f4",
          2589 => x"84",
          2590 => x"83",
          2591 => x"72",
          2592 => x"59",
          2593 => x"18",
          2594 => x"06",
          2595 => x"38",
          2596 => x"fb",
          2597 => x"f9",
          2598 => x"5d",
          2599 => x"83",
          2600 => x"83",
          2601 => x"72",
          2602 => x"72",
          2603 => x"5b",
          2604 => x"a0",
          2605 => x"83",
          2606 => x"72",
          2607 => x"a0",
          2608 => x"f8",
          2609 => x"5e",
          2610 => x"80",
          2611 => x"81",
          2612 => x"f8",
          2613 => x"44",
          2614 => x"84",
          2615 => x"70",
          2616 => x"27",
          2617 => x"34",
          2618 => x"c4",
          2619 => x"9c",
          2620 => x"33",
          2621 => x"34",
          2622 => x"06",
          2623 => x"81",
          2624 => x"84",
          2625 => x"83",
          2626 => x"c4",
          2627 => x"33",
          2628 => x"33",
          2629 => x"39",
          2630 => x"11",
          2631 => x"3f",
          2632 => x"f0",
          2633 => x"57",
          2634 => x"10",
          2635 => x"05",
          2636 => x"fb",
          2637 => x"5c",
          2638 => x"83",
          2639 => x"83",
          2640 => x"e5",
          2641 => x"f8",
          2642 => x"29",
          2643 => x"19",
          2644 => x"34",
          2645 => x"33",
          2646 => x"12",
          2647 => x"fa",
          2648 => x"71",
          2649 => x"33",
          2650 => x"84",
          2651 => x"83",
          2652 => x"72",
          2653 => x"5a",
          2654 => x"1e",
          2655 => x"5c",
          2656 => x"84",
          2657 => x"38",
          2658 => x"34",
          2659 => x"b7",
          2660 => x"bd",
          2661 => x"f3",
          2662 => x"e4",
          2663 => x"9c",
          2664 => x"83",
          2665 => x"83",
          2666 => x"57",
          2667 => x"39",
          2668 => x"34",
          2669 => x"34",
          2670 => x"34",
          2671 => x"5b",
          2672 => x"b9",
          2673 => x"81",
          2674 => x"33",
          2675 => x"81",
          2676 => x"52",
          2677 => x"f8",
          2678 => x"84",
          2679 => x"f7",
          2680 => x"a0",
          2681 => x"f7",
          2682 => x"c0",
          2683 => x"5b",
          2684 => x"7b",
          2685 => x"b9",
          2686 => x"75",
          2687 => x"10",
          2688 => x"04",
          2689 => x"2e",
          2690 => x"84",
          2691 => x"09",
          2692 => x"59",
          2693 => x"fd",
          2694 => x"75",
          2695 => x"9d",
          2696 => x"84",
          2697 => x"7b",
          2698 => x"f9",
          2699 => x"f8",
          2700 => x"81",
          2701 => x"fd",
          2702 => x"f8",
          2703 => x"83",
          2704 => x"84",
          2705 => x"76",
          2706 => x"56",
          2707 => x"39",
          2708 => x"2e",
          2709 => x"84",
          2710 => x"09",
          2711 => x"59",
          2712 => x"fc",
          2713 => x"7a",
          2714 => x"9c",
          2715 => x"06",
          2716 => x"83",
          2717 => x"72",
          2718 => x"11",
          2719 => x"58",
          2720 => x"ff",
          2721 => x"fe",
          2722 => x"84",
          2723 => x"0b",
          2724 => x"84",
          2725 => x"fb",
          2726 => x"77",
          2727 => x"38",
          2728 => x"d0",
          2729 => x"80",
          2730 => x"33",
          2731 => x"84",
          2732 => x"56",
          2733 => x"76",
          2734 => x"84",
          2735 => x"8c",
          2736 => x"f8",
          2737 => x"bb",
          2738 => x"60",
          2739 => x"f8",
          2740 => x"90",
          2741 => x"84",
          2742 => x"27",
          2743 => x"9c",
          2744 => x"f0",
          2745 => x"70",
          2746 => x"58",
          2747 => x"b8",
          2748 => x"8d",
          2749 => x"83",
          2750 => x"76",
          2751 => x"fa",
          2752 => x"81",
          2753 => x"9f",
          2754 => x"84",
          2755 => x"ff",
          2756 => x"ff",
          2757 => x"59",
          2758 => x"77",
          2759 => x"81",
          2760 => x"7f",
          2761 => x"f8",
          2762 => x"11",
          2763 => x"38",
          2764 => x"f9",
          2765 => x"7e",
          2766 => x"9d",
          2767 => x"7a",
          2768 => x"f8",
          2769 => x"ff",
          2770 => x"29",
          2771 => x"f8",
          2772 => x"05",
          2773 => x"ce",
          2774 => x"60",
          2775 => x"ff",
          2776 => x"80",
          2777 => x"bb",
          2778 => x"38",
          2779 => x"23",
          2780 => x"41",
          2781 => x"84",
          2782 => x"8d",
          2783 => x"f8",
          2784 => x"f8",
          2785 => x"76",
          2786 => x"05",
          2787 => x"5c",
          2788 => x"80",
          2789 => x"ff",
          2790 => x"29",
          2791 => x"27",
          2792 => x"57",
          2793 => x"c4",
          2794 => x"34",
          2795 => x"70",
          2796 => x"b7",
          2797 => x"71",
          2798 => x"60",
          2799 => x"33",
          2800 => x"70",
          2801 => x"05",
          2802 => x"34",
          2803 => x"b7",
          2804 => x"40",
          2805 => x"38",
          2806 => x"56",
          2807 => x"52",
          2808 => x"3f",
          2809 => x"bc",
          2810 => x"5d",
          2811 => x"38",
          2812 => x"2e",
          2813 => x"f8",
          2814 => x"83",
          2815 => x"76",
          2816 => x"bb",
          2817 => x"38",
          2818 => x"26",
          2819 => x"7d",
          2820 => x"7a",
          2821 => x"05",
          2822 => x"5d",
          2823 => x"83",
          2824 => x"38",
          2825 => x"38",
          2826 => x"71",
          2827 => x"71",
          2828 => x"77",
          2829 => x"84",
          2830 => x"05",
          2831 => x"84",
          2832 => x"41",
          2833 => x"ff",
          2834 => x"29",
          2835 => x"77",
          2836 => x"70",
          2837 => x"76",
          2838 => x"e0",
          2839 => x"9a",
          2840 => x"19",
          2841 => x"34",
          2842 => x"c0",
          2843 => x"79",
          2844 => x"17",
          2845 => x"a8",
          2846 => x"5d",
          2847 => x"33",
          2848 => x"80",
          2849 => x"5d",
          2850 => x"06",
          2851 => x"f4",
          2852 => x"59",
          2853 => x"17",
          2854 => x"7c",
          2855 => x"bc",
          2856 => x"bb",
          2857 => x"39",
          2858 => x"75",
          2859 => x"81",
          2860 => x"83",
          2861 => x"07",
          2862 => x"39",
          2863 => x"83",
          2864 => x"d4",
          2865 => x"06",
          2866 => x"34",
          2867 => x"9f",
          2868 => x"f4",
          2869 => x"83",
          2870 => x"ff",
          2871 => x"f8",
          2872 => x"83",
          2873 => x"f8",
          2874 => x"56",
          2875 => x"39",
          2876 => x"80",
          2877 => x"34",
          2878 => x"81",
          2879 => x"83",
          2880 => x"f8",
          2881 => x"56",
          2882 => x"39",
          2883 => x"86",
          2884 => x"fe",
          2885 => x"fc",
          2886 => x"f4",
          2887 => x"33",
          2888 => x"83",
          2889 => x"f8",
          2890 => x"83",
          2891 => x"f8",
          2892 => x"83",
          2893 => x"f8",
          2894 => x"83",
          2895 => x"f8",
          2896 => x"07",
          2897 => x"cc",
          2898 => x"06",
          2899 => x"34",
          2900 => x"f9",
          2901 => x"3f",
          2902 => x"83",
          2903 => x"83",
          2904 => x"59",
          2905 => x"84",
          2906 => x"0b",
          2907 => x"b9",
          2908 => x"83",
          2909 => x"70",
          2910 => x"e7",
          2911 => x"3d",
          2912 => x"f8",
          2913 => x"38",
          2914 => x"0c",
          2915 => x"0b",
          2916 => x"04",
          2917 => x"39",
          2918 => x"5c",
          2919 => x"83",
          2920 => x"22",
          2921 => x"84",
          2922 => x"83",
          2923 => x"d1",
          2924 => x"81",
          2925 => x"d8",
          2926 => x"80",
          2927 => x"98",
          2928 => x"ef",
          2929 => x"05",
          2930 => x"58",
          2931 => x"81",
          2932 => x"40",
          2933 => x"83",
          2934 => x"f8",
          2935 => x"9f",
          2936 => x"e2",
          2937 => x"84",
          2938 => x"56",
          2939 => x"57",
          2940 => x"70",
          2941 => x"26",
          2942 => x"84",
          2943 => x"83",
          2944 => x"86",
          2945 => x"22",
          2946 => x"83",
          2947 => x"5d",
          2948 => x"2e",
          2949 => x"06",
          2950 => x"84",
          2951 => x"76",
          2952 => x"56",
          2953 => x"ff",
          2954 => x"24",
          2955 => x"56",
          2956 => x"16",
          2957 => x"81",
          2958 => x"57",
          2959 => x"75",
          2960 => x"06",
          2961 => x"58",
          2962 => x"b0",
          2963 => x"ff",
          2964 => x"42",
          2965 => x"84",
          2966 => x"33",
          2967 => x"70",
          2968 => x"05",
          2969 => x"34",
          2970 => x"b7",
          2971 => x"41",
          2972 => x"38",
          2973 => x"c4",
          2974 => x"34",
          2975 => x"70",
          2976 => x"b7",
          2977 => x"71",
          2978 => x"78",
          2979 => x"83",
          2980 => x"c4",
          2981 => x"33",
          2982 => x"22",
          2983 => x"5d",
          2984 => x"84",
          2985 => x"ff",
          2986 => x"83",
          2987 => x"23",
          2988 => x"5a",
          2989 => x"76",
          2990 => x"33",
          2991 => x"59",
          2992 => x"80",
          2993 => x"88",
          2994 => x"84",
          2995 => x"56",
          2996 => x"57",
          2997 => x"81",
          2998 => x"33",
          2999 => x"33",
          3000 => x"2e",
          3001 => x"a1",
          3002 => x"f8",
          3003 => x"75",
          3004 => x"7c",
          3005 => x"34",
          3006 => x"77",
          3007 => x"70",
          3008 => x"33",
          3009 => x"7a",
          3010 => x"81",
          3011 => x"77",
          3012 => x"27",
          3013 => x"31",
          3014 => x"a8",
          3015 => x"fc",
          3016 => x"fc",
          3017 => x"23",
          3018 => x"f8",
          3019 => x"18",
          3020 => x"77",
          3021 => x"e9",
          3022 => x"05",
          3023 => x"72",
          3024 => x"9c",
          3025 => x"85",
          3026 => x"d7",
          3027 => x"0c",
          3028 => x"02",
          3029 => x"f7",
          3030 => x"f7",
          3031 => x"74",
          3032 => x"56",
          3033 => x"78",
          3034 => x"04",
          3035 => x"73",
          3036 => x"70",
          3037 => x"2a",
          3038 => x"a8",
          3039 => x"2e",
          3040 => x"7b",
          3041 => x"76",
          3042 => x"85",
          3043 => x"f8",
          3044 => x"71",
          3045 => x"83",
          3046 => x"79",
          3047 => x"83",
          3048 => x"74",
          3049 => x"54",
          3050 => x"0b",
          3051 => x"98",
          3052 => x"38",
          3053 => x"83",
          3054 => x"81",
          3055 => x"27",
          3056 => x"14",
          3057 => x"f2",
          3058 => x"2e",
          3059 => x"86",
          3060 => x"34",
          3061 => x"ff",
          3062 => x"86",
          3063 => x"83",
          3064 => x"81",
          3065 => x"ff",
          3066 => x"98",
          3067 => x"75",
          3068 => x"06",
          3069 => x"06",
          3070 => x"e7",
          3071 => x"73",
          3072 => x"85",
          3073 => x"34",
          3074 => x"f7",
          3075 => x"83",
          3076 => x"5d",
          3077 => x"f6",
          3078 => x"2e",
          3079 => x"54",
          3080 => x"f7",
          3081 => x"2e",
          3082 => x"54",
          3083 => x"06",
          3084 => x"83",
          3085 => x"2e",
          3086 => x"53",
          3087 => x"83",
          3088 => x"27",
          3089 => x"87",
          3090 => x"54",
          3091 => x"81",
          3092 => x"f7",
          3093 => x"ff",
          3094 => x"f6",
          3095 => x"83",
          3096 => x"72",
          3097 => x"10",
          3098 => x"04",
          3099 => x"2e",
          3100 => x"98",
          3101 => x"fc",
          3102 => x"33",
          3103 => x"74",
          3104 => x"c0",
          3105 => x"73",
          3106 => x"94",
          3107 => x"84",
          3108 => x"f0",
          3109 => x"08",
          3110 => x"72",
          3111 => x"76",
          3112 => x"80",
          3113 => x"57",
          3114 => x"79",
          3115 => x"38",
          3116 => x"81",
          3117 => x"06",
          3118 => x"54",
          3119 => x"80",
          3120 => x"ff",
          3121 => x"72",
          3122 => x"58",
          3123 => x"10",
          3124 => x"83",
          3125 => x"70",
          3126 => x"98",
          3127 => x"fd",
          3128 => x"ff",
          3129 => x"ff",
          3130 => x"78",
          3131 => x"84",
          3132 => x"2e",
          3133 => x"30",
          3134 => x"56",
          3135 => x"81",
          3136 => x"f9",
          3137 => x"10",
          3138 => x"54",
          3139 => x"13",
          3140 => x"73",
          3141 => x"53",
          3142 => x"b7",
          3143 => x"78",
          3144 => x"d4",
          3145 => x"3d",
          3146 => x"54",
          3147 => x"92",
          3148 => x"05",
          3149 => x"fa",
          3150 => x"15",
          3151 => x"34",
          3152 => x"fa",
          3153 => x"72",
          3154 => x"f7",
          3155 => x"fc",
          3156 => x"73",
          3157 => x"38",
          3158 => x"87",
          3159 => x"73",
          3160 => x"9c",
          3161 => x"ff",
          3162 => x"83",
          3163 => x"72",
          3164 => x"06",
          3165 => x"f7",
          3166 => x"33",
          3167 => x"33",
          3168 => x"a3",
          3169 => x"56",
          3170 => x"81",
          3171 => x"81",
          3172 => x"09",
          3173 => x"39",
          3174 => x"98",
          3175 => x"57",
          3176 => x"84",
          3177 => x"39",
          3178 => x"54",
          3179 => x"b7",
          3180 => x"81",
          3181 => x"f7",
          3182 => x"0c",
          3183 => x"70",
          3184 => x"54",
          3185 => x"74",
          3186 => x"06",
          3187 => x"83",
          3188 => x"34",
          3189 => x"06",
          3190 => x"83",
          3191 => x"34",
          3192 => x"83",
          3193 => x"f6",
          3194 => x"84",
          3195 => x"fe",
          3196 => x"cc",
          3197 => x"bb",
          3198 => x"ac",
          3199 => x"0d",
          3200 => x"57",
          3201 => x"83",
          3202 => x"34",
          3203 => x"56",
          3204 => x"86",
          3205 => x"9c",
          3206 => x"ce",
          3207 => x"08",
          3208 => x"70",
          3209 => x"87",
          3210 => x"73",
          3211 => x"db",
          3212 => x"ff",
          3213 => x"71",
          3214 => x"87",
          3215 => x"05",
          3216 => x"87",
          3217 => x"2e",
          3218 => x"98",
          3219 => x"87",
          3220 => x"87",
          3221 => x"26",
          3222 => x"16",
          3223 => x"80",
          3224 => x"52",
          3225 => x"8a",
          3226 => x"3d",
          3227 => x"0c",
          3228 => x"79",
          3229 => x"52",
          3230 => x"88",
          3231 => x"75",
          3232 => x"71",
          3233 => x"70",
          3234 => x"75",
          3235 => x"83",
          3236 => x"34",
          3237 => x"71",
          3238 => x"55",
          3239 => x"0b",
          3240 => x"98",
          3241 => x"80",
          3242 => x"9c",
          3243 => x"51",
          3244 => x"33",
          3245 => x"74",
          3246 => x"2e",
          3247 => x"51",
          3248 => x"38",
          3249 => x"38",
          3250 => x"90",
          3251 => x"52",
          3252 => x"72",
          3253 => x"c0",
          3254 => x"27",
          3255 => x"38",
          3256 => x"75",
          3257 => x"ff",
          3258 => x"75",
          3259 => x"ff",
          3260 => x"51",
          3261 => x"38",
          3262 => x"55",
          3263 => x"71",
          3264 => x"81",
          3265 => x"38",
          3266 => x"0d",
          3267 => x"88",
          3268 => x"fa",
          3269 => x"05",
          3270 => x"d4",
          3271 => x"80",
          3272 => x"55",
          3273 => x"90",
          3274 => x"90",
          3275 => x"86",
          3276 => x"80",
          3277 => x"55",
          3278 => x"70",
          3279 => x"05",
          3280 => x"83",
          3281 => x"34",
          3282 => x"75",
          3283 => x"55",
          3284 => x"0b",
          3285 => x"98",
          3286 => x"80",
          3287 => x"9c",
          3288 => x"51",
          3289 => x"33",
          3290 => x"74",
          3291 => x"2e",
          3292 => x"51",
          3293 => x"38",
          3294 => x"38",
          3295 => x"90",
          3296 => x"52",
          3297 => x"72",
          3298 => x"c0",
          3299 => x"27",
          3300 => x"38",
          3301 => x"75",
          3302 => x"ff",
          3303 => x"75",
          3304 => x"06",
          3305 => x"70",
          3306 => x"83",
          3307 => x"0c",
          3308 => x"39",
          3309 => x"51",
          3310 => x"f3",
          3311 => x"16",
          3312 => x"34",
          3313 => x"d4",
          3314 => x"87",
          3315 => x"98",
          3316 => x"38",
          3317 => x"08",
          3318 => x"71",
          3319 => x"98",
          3320 => x"27",
          3321 => x"2e",
          3322 => x"08",
          3323 => x"98",
          3324 => x"08",
          3325 => x"15",
          3326 => x"52",
          3327 => x"ff",
          3328 => x"08",
          3329 => x"52",
          3330 => x"06",
          3331 => x"72",
          3332 => x"38",
          3333 => x"cc",
          3334 => x"0d",
          3335 => x"08",
          3336 => x"ff",
          3337 => x"70",
          3338 => x"71",
          3339 => x"81",
          3340 => x"2b",
          3341 => x"57",
          3342 => x"24",
          3343 => x"33",
          3344 => x"83",
          3345 => x"12",
          3346 => x"07",
          3347 => x"80",
          3348 => x"33",
          3349 => x"83",
          3350 => x"52",
          3351 => x"73",
          3352 => x"34",
          3353 => x"12",
          3354 => x"07",
          3355 => x"51",
          3356 => x"34",
          3357 => x"0b",
          3358 => x"34",
          3359 => x"14",
          3360 => x"b8",
          3361 => x"71",
          3362 => x"70",
          3363 => x"72",
          3364 => x"0d",
          3365 => x"71",
          3366 => x"11",
          3367 => x"88",
          3368 => x"54",
          3369 => x"34",
          3370 => x"08",
          3371 => x"33",
          3372 => x"56",
          3373 => x"33",
          3374 => x"70",
          3375 => x"86",
          3376 => x"b9",
          3377 => x"33",
          3378 => x"06",
          3379 => x"76",
          3380 => x"b9",
          3381 => x"12",
          3382 => x"07",
          3383 => x"71",
          3384 => x"ff",
          3385 => x"54",
          3386 => x"52",
          3387 => x"34",
          3388 => x"33",
          3389 => x"83",
          3390 => x"12",
          3391 => x"ff",
          3392 => x"55",
          3393 => x"70",
          3394 => x"70",
          3395 => x"71",
          3396 => x"05",
          3397 => x"2b",
          3398 => x"52",
          3399 => x"fc",
          3400 => x"71",
          3401 => x"70",
          3402 => x"34",
          3403 => x"08",
          3404 => x"71",
          3405 => x"05",
          3406 => x"88",
          3407 => x"5c",
          3408 => x"15",
          3409 => x"0d",
          3410 => x"b8",
          3411 => x"38",
          3412 => x"fb",
          3413 => x"ff",
          3414 => x"80",
          3415 => x"80",
          3416 => x"fe",
          3417 => x"55",
          3418 => x"34",
          3419 => x"15",
          3420 => x"b9",
          3421 => x"81",
          3422 => x"08",
          3423 => x"80",
          3424 => x"70",
          3425 => x"88",
          3426 => x"b9",
          3427 => x"b9",
          3428 => x"76",
          3429 => x"34",
          3430 => x"52",
          3431 => x"8e",
          3432 => x"70",
          3433 => x"83",
          3434 => x"84",
          3435 => x"2b",
          3436 => x"81",
          3437 => x"cc",
          3438 => x"33",
          3439 => x"70",
          3440 => x"83",
          3441 => x"53",
          3442 => x"8a",
          3443 => x"73",
          3444 => x"33",
          3445 => x"c1",
          3446 => x"38",
          3447 => x"2b",
          3448 => x"71",
          3449 => x"06",
          3450 => x"79",
          3451 => x"74",
          3452 => x"78",
          3453 => x"2e",
          3454 => x"2b",
          3455 => x"70",
          3456 => x"76",
          3457 => x"b9",
          3458 => x"53",
          3459 => x"34",
          3460 => x"33",
          3461 => x"70",
          3462 => x"05",
          3463 => x"2a",
          3464 => x"75",
          3465 => x"53",
          3466 => x"08",
          3467 => x"15",
          3468 => x"86",
          3469 => x"2b",
          3470 => x"5c",
          3471 => x"72",
          3472 => x"70",
          3473 => x"87",
          3474 => x"88",
          3475 => x"15",
          3476 => x"b8",
          3477 => x"12",
          3478 => x"07",
          3479 => x"75",
          3480 => x"84",
          3481 => x"05",
          3482 => x"88",
          3483 => x"57",
          3484 => x"15",
          3485 => x"05",
          3486 => x"3d",
          3487 => x"33",
          3488 => x"79",
          3489 => x"71",
          3490 => x"5b",
          3491 => x"34",
          3492 => x"08",
          3493 => x"33",
          3494 => x"74",
          3495 => x"71",
          3496 => x"5d",
          3497 => x"86",
          3498 => x"b9",
          3499 => x"33",
          3500 => x"06",
          3501 => x"75",
          3502 => x"b9",
          3503 => x"f1",
          3504 => x"b8",
          3505 => x"38",
          3506 => x"b9",
          3507 => x"51",
          3508 => x"84",
          3509 => x"84",
          3510 => x"a0",
          3511 => x"80",
          3512 => x"51",
          3513 => x"08",
          3514 => x"16",
          3515 => x"84",
          3516 => x"84",
          3517 => x"34",
          3518 => x"b8",
          3519 => x"fe",
          3520 => x"06",
          3521 => x"74",
          3522 => x"84",
          3523 => x"84",
          3524 => x"55",
          3525 => x"15",
          3526 => x"dd",
          3527 => x"65",
          3528 => x"b8",
          3529 => x"84",
          3530 => x"38",
          3531 => x"54",
          3532 => x"05",
          3533 => x"ff",
          3534 => x"06",
          3535 => x"ff",
          3536 => x"70",
          3537 => x"07",
          3538 => x"06",
          3539 => x"83",
          3540 => x"33",
          3541 => x"70",
          3542 => x"53",
          3543 => x"5e",
          3544 => x"38",
          3545 => x"88",
          3546 => x"70",
          3547 => x"71",
          3548 => x"56",
          3549 => x"7a",
          3550 => x"58",
          3551 => x"80",
          3552 => x"77",
          3553 => x"59",
          3554 => x"1e",
          3555 => x"2b",
          3556 => x"33",
          3557 => x"90",
          3558 => x"57",
          3559 => x"38",
          3560 => x"33",
          3561 => x"7a",
          3562 => x"71",
          3563 => x"05",
          3564 => x"88",
          3565 => x"48",
          3566 => x"56",
          3567 => x"34",
          3568 => x"11",
          3569 => x"71",
          3570 => x"33",
          3571 => x"70",
          3572 => x"57",
          3573 => x"87",
          3574 => x"70",
          3575 => x"07",
          3576 => x"5a",
          3577 => x"81",
          3578 => x"1f",
          3579 => x"8b",
          3580 => x"73",
          3581 => x"07",
          3582 => x"5f",
          3583 => x"81",
          3584 => x"1f",
          3585 => x"2b",
          3586 => x"14",
          3587 => x"07",
          3588 => x"5f",
          3589 => x"75",
          3590 => x"70",
          3591 => x"71",
          3592 => x"70",
          3593 => x"05",
          3594 => x"84",
          3595 => x"65",
          3596 => x"5d",
          3597 => x"38",
          3598 => x"95",
          3599 => x"84",
          3600 => x"b9",
          3601 => x"52",
          3602 => x"3f",
          3603 => x"34",
          3604 => x"b8",
          3605 => x"0b",
          3606 => x"5c",
          3607 => x"1d",
          3608 => x"b4",
          3609 => x"70",
          3610 => x"5c",
          3611 => x"77",
          3612 => x"70",
          3613 => x"05",
          3614 => x"34",
          3615 => x"b8",
          3616 => x"80",
          3617 => x"80",
          3618 => x"9b",
          3619 => x"c8",
          3620 => x"84",
          3621 => x"11",
          3622 => x"12",
          3623 => x"ff",
          3624 => x"5e",
          3625 => x"34",
          3626 => x"88",
          3627 => x"7b",
          3628 => x"70",
          3629 => x"88",
          3630 => x"f8",
          3631 => x"06",
          3632 => x"5e",
          3633 => x"76",
          3634 => x"05",
          3635 => x"63",
          3636 => x"84",
          3637 => x"ed",
          3638 => x"7b",
          3639 => x"42",
          3640 => x"ff",
          3641 => x"06",
          3642 => x"88",
          3643 => x"70",
          3644 => x"71",
          3645 => x"58",
          3646 => x"f7",
          3647 => x"fa",
          3648 => x"38",
          3649 => x"7b",
          3650 => x"84",
          3651 => x"a0",
          3652 => x"80",
          3653 => x"51",
          3654 => x"08",
          3655 => x"1b",
          3656 => x"84",
          3657 => x"84",
          3658 => x"34",
          3659 => x"b8",
          3660 => x"fe",
          3661 => x"06",
          3662 => x"74",
          3663 => x"05",
          3664 => x"10",
          3665 => x"05",
          3666 => x"81",
          3667 => x"80",
          3668 => x"ff",
          3669 => x"c0",
          3670 => x"82",
          3671 => x"7f",
          3672 => x"3d",
          3673 => x"83",
          3674 => x"2b",
          3675 => x"12",
          3676 => x"07",
          3677 => x"33",
          3678 => x"43",
          3679 => x"5c",
          3680 => x"7a",
          3681 => x"08",
          3682 => x"33",
          3683 => x"74",
          3684 => x"71",
          3685 => x"41",
          3686 => x"64",
          3687 => x"34",
          3688 => x"81",
          3689 => x"ff",
          3690 => x"5a",
          3691 => x"34",
          3692 => x"11",
          3693 => x"71",
          3694 => x"81",
          3695 => x"88",
          3696 => x"45",
          3697 => x"34",
          3698 => x"33",
          3699 => x"83",
          3700 => x"83",
          3701 => x"88",
          3702 => x"55",
          3703 => x"18",
          3704 => x"82",
          3705 => x"2b",
          3706 => x"2b",
          3707 => x"05",
          3708 => x"b8",
          3709 => x"ff",
          3710 => x"ff",
          3711 => x"80",
          3712 => x"80",
          3713 => x"fe",
          3714 => x"56",
          3715 => x"34",
          3716 => x"16",
          3717 => x"b9",
          3718 => x"81",
          3719 => x"08",
          3720 => x"80",
          3721 => x"70",
          3722 => x"88",
          3723 => x"b9",
          3724 => x"b9",
          3725 => x"7f",
          3726 => x"34",
          3727 => x"fc",
          3728 => x"33",
          3729 => x"79",
          3730 => x"71",
          3731 => x"48",
          3732 => x"05",
          3733 => x"b9",
          3734 => x"85",
          3735 => x"2b",
          3736 => x"15",
          3737 => x"2a",
          3738 => x"40",
          3739 => x"87",
          3740 => x"70",
          3741 => x"07",
          3742 => x"59",
          3743 => x"81",
          3744 => x"1f",
          3745 => x"2b",
          3746 => x"33",
          3747 => x"70",
          3748 => x"05",
          3749 => x"5d",
          3750 => x"34",
          3751 => x"08",
          3752 => x"71",
          3753 => x"05",
          3754 => x"2b",
          3755 => x"2a",
          3756 => x"5b",
          3757 => x"34",
          3758 => x"b3",
          3759 => x"71",
          3760 => x"05",
          3761 => x"88",
          3762 => x"5a",
          3763 => x"79",
          3764 => x"70",
          3765 => x"71",
          3766 => x"05",
          3767 => x"88",
          3768 => x"5e",
          3769 => x"86",
          3770 => x"84",
          3771 => x"12",
          3772 => x"ff",
          3773 => x"55",
          3774 => x"84",
          3775 => x"81",
          3776 => x"2b",
          3777 => x"33",
          3778 => x"8f",
          3779 => x"2a",
          3780 => x"5e",
          3781 => x"17",
          3782 => x"70",
          3783 => x"71",
          3784 => x"81",
          3785 => x"ff",
          3786 => x"5e",
          3787 => x"34",
          3788 => x"08",
          3789 => x"33",
          3790 => x"74",
          3791 => x"71",
          3792 => x"05",
          3793 => x"88",
          3794 => x"49",
          3795 => x"57",
          3796 => x"1d",
          3797 => x"84",
          3798 => x"2b",
          3799 => x"14",
          3800 => x"07",
          3801 => x"40",
          3802 => x"7b",
          3803 => x"16",
          3804 => x"2b",
          3805 => x"2a",
          3806 => x"79",
          3807 => x"70",
          3808 => x"71",
          3809 => x"05",
          3810 => x"2b",
          3811 => x"5d",
          3812 => x"75",
          3813 => x"70",
          3814 => x"8b",
          3815 => x"82",
          3816 => x"2b",
          3817 => x"5d",
          3818 => x"34",
          3819 => x"08",
          3820 => x"33",
          3821 => x"56",
          3822 => x"7e",
          3823 => x"3f",
          3824 => x"61",
          3825 => x"06",
          3826 => x"19",
          3827 => x"71",
          3828 => x"33",
          3829 => x"70",
          3830 => x"55",
          3831 => x"85",
          3832 => x"1e",
          3833 => x"8b",
          3834 => x"86",
          3835 => x"2b",
          3836 => x"48",
          3837 => x"05",
          3838 => x"b9",
          3839 => x"33",
          3840 => x"06",
          3841 => x"78",
          3842 => x"b9",
          3843 => x"12",
          3844 => x"07",
          3845 => x"71",
          3846 => x"ff",
          3847 => x"5d",
          3848 => x"40",
          3849 => x"34",
          3850 => x"33",
          3851 => x"83",
          3852 => x"12",
          3853 => x"ff",
          3854 => x"58",
          3855 => x"78",
          3856 => x"06",
          3857 => x"54",
          3858 => x"5f",
          3859 => x"38",
          3860 => x"08",
          3861 => x"df",
          3862 => x"ef",
          3863 => x"0d",
          3864 => x"58",
          3865 => x"54",
          3866 => x"0c",
          3867 => x"d3",
          3868 => x"b9",
          3869 => x"53",
          3870 => x"fe",
          3871 => x"0c",
          3872 => x"0b",
          3873 => x"84",
          3874 => x"76",
          3875 => x"df",
          3876 => x"75",
          3877 => x"b9",
          3878 => x"81",
          3879 => x"08",
          3880 => x"87",
          3881 => x"b9",
          3882 => x"07",
          3883 => x"2a",
          3884 => x"34",
          3885 => x"22",
          3886 => x"08",
          3887 => x"15",
          3888 => x"54",
          3889 => x"cc",
          3890 => x"33",
          3891 => x"38",
          3892 => x"84",
          3893 => x"fe",
          3894 => x"83",
          3895 => x"51",
          3896 => x"81",
          3897 => x"84",
          3898 => x"12",
          3899 => x"84",
          3900 => x"7e",
          3901 => x"5a",
          3902 => x"26",
          3903 => x"54",
          3904 => x"bd",
          3905 => x"98",
          3906 => x"51",
          3907 => x"81",
          3908 => x"38",
          3909 => x"e2",
          3910 => x"fc",
          3911 => x"83",
          3912 => x"b9",
          3913 => x"80",
          3914 => x"5a",
          3915 => x"38",
          3916 => x"60",
          3917 => x"5c",
          3918 => x"87",
          3919 => x"73",
          3920 => x"38",
          3921 => x"8c",
          3922 => x"d7",
          3923 => x"ff",
          3924 => x"87",
          3925 => x"38",
          3926 => x"80",
          3927 => x"38",
          3928 => x"c8",
          3929 => x"16",
          3930 => x"55",
          3931 => x"d5",
          3932 => x"05",
          3933 => x"05",
          3934 => x"73",
          3935 => x"33",
          3936 => x"73",
          3937 => x"8c",
          3938 => x"38",
          3939 => x"2e",
          3940 => x"c8",
          3941 => x"0a",
          3942 => x"86",
          3943 => x"80",
          3944 => x"0d",
          3945 => x"8c",
          3946 => x"08",
          3947 => x"70",
          3948 => x"8c",
          3949 => x"98",
          3950 => x"72",
          3951 => x"71",
          3952 => x"ff",
          3953 => x"73",
          3954 => x"0d",
          3955 => x"71",
          3956 => x"81",
          3957 => x"83",
          3958 => x"52",
          3959 => x"84",
          3960 => x"81",
          3961 => x"3d",
          3962 => x"53",
          3963 => x"52",
          3964 => x"b9",
          3965 => x"d9",
          3966 => x"34",
          3967 => x"31",
          3968 => x"5c",
          3969 => x"9b",
          3970 => x"2e",
          3971 => x"54",
          3972 => x"33",
          3973 => x"57",
          3974 => x"fe",
          3975 => x"81",
          3976 => x"b8",
          3977 => x"80",
          3978 => x"17",
          3979 => x"84",
          3980 => x"b7",
          3981 => x"d2",
          3982 => x"ba",
          3983 => x"34",
          3984 => x"80",
          3985 => x"c1",
          3986 => x"0b",
          3987 => x"55",
          3988 => x"2a",
          3989 => x"90",
          3990 => x"74",
          3991 => x"34",
          3992 => x"19",
          3993 => x"a5",
          3994 => x"84",
          3995 => x"74",
          3996 => x"81",
          3997 => x"54",
          3998 => x"51",
          3999 => x"80",
          4000 => x"fb",
          4001 => x"2e",
          4002 => x"3d",
          4003 => x"56",
          4004 => x"08",
          4005 => x"84",
          4006 => x"ff",
          4007 => x"81",
          4008 => x"38",
          4009 => x"38",
          4010 => x"a8",
          4011 => x"b4",
          4012 => x"17",
          4013 => x"06",
          4014 => x"b8",
          4015 => x"e3",
          4016 => x"85",
          4017 => x"18",
          4018 => x"ff",
          4019 => x"70",
          4020 => x"5d",
          4021 => x"b5",
          4022 => x"5c",
          4023 => x"06",
          4024 => x"b8",
          4025 => x"93",
          4026 => x"85",
          4027 => x"18",
          4028 => x"ff",
          4029 => x"2b",
          4030 => x"2a",
          4031 => x"ae",
          4032 => x"c8",
          4033 => x"2a",
          4034 => x"08",
          4035 => x"18",
          4036 => x"2e",
          4037 => x"54",
          4038 => x"33",
          4039 => x"08",
          4040 => x"5a",
          4041 => x"38",
          4042 => x"b8",
          4043 => x"88",
          4044 => x"5b",
          4045 => x"09",
          4046 => x"2a",
          4047 => x"08",
          4048 => x"18",
          4049 => x"2e",
          4050 => x"54",
          4051 => x"33",
          4052 => x"08",
          4053 => x"5a",
          4054 => x"38",
          4055 => x"05",
          4056 => x"33",
          4057 => x"81",
          4058 => x"75",
          4059 => x"06",
          4060 => x"5e",
          4061 => x"81",
          4062 => x"70",
          4063 => x"e2",
          4064 => x"7b",
          4065 => x"84",
          4066 => x"17",
          4067 => x"c8",
          4068 => x"27",
          4069 => x"74",
          4070 => x"38",
          4071 => x"08",
          4072 => x"51",
          4073 => x"39",
          4074 => x"17",
          4075 => x"f6",
          4076 => x"2e",
          4077 => x"b9",
          4078 => x"08",
          4079 => x"18",
          4080 => x"5e",
          4081 => x"b9",
          4082 => x"54",
          4083 => x"53",
          4084 => x"3f",
          4085 => x"2e",
          4086 => x"b9",
          4087 => x"08",
          4088 => x"08",
          4089 => x"fd",
          4090 => x"82",
          4091 => x"81",
          4092 => x"05",
          4093 => x"f4",
          4094 => x"81",
          4095 => x"70",
          4096 => x"da",
          4097 => x"7d",
          4098 => x"84",
          4099 => x"17",
          4100 => x"c8",
          4101 => x"27",
          4102 => x"74",
          4103 => x"38",
          4104 => x"08",
          4105 => x"51",
          4106 => x"39",
          4107 => x"08",
          4108 => x"51",
          4109 => x"5b",
          4110 => x"f2",
          4111 => x"59",
          4112 => x"75",
          4113 => x"33",
          4114 => x"78",
          4115 => x"82",
          4116 => x"90",
          4117 => x"1a",
          4118 => x"08",
          4119 => x"38",
          4120 => x"7c",
          4121 => x"81",
          4122 => x"19",
          4123 => x"c8",
          4124 => x"81",
          4125 => x"79",
          4126 => x"06",
          4127 => x"58",
          4128 => x"2a",
          4129 => x"83",
          4130 => x"90",
          4131 => x"81",
          4132 => x"a8",
          4133 => x"1a",
          4134 => x"e1",
          4135 => x"7c",
          4136 => x"38",
          4137 => x"81",
          4138 => x"b9",
          4139 => x"58",
          4140 => x"58",
          4141 => x"83",
          4142 => x"11",
          4143 => x"7e",
          4144 => x"5c",
          4145 => x"75",
          4146 => x"79",
          4147 => x"7a",
          4148 => x"34",
          4149 => x"70",
          4150 => x"1b",
          4151 => x"b7",
          4152 => x"5e",
          4153 => x"06",
          4154 => x"b8",
          4155 => x"83",
          4156 => x"85",
          4157 => x"1a",
          4158 => x"79",
          4159 => x"1b",
          4160 => x"55",
          4161 => x"2b",
          4162 => x"71",
          4163 => x"0b",
          4164 => x"1a",
          4165 => x"08",
          4166 => x"38",
          4167 => x"53",
          4168 => x"3f",
          4169 => x"2e",
          4170 => x"b9",
          4171 => x"08",
          4172 => x"08",
          4173 => x"5c",
          4174 => x"33",
          4175 => x"81",
          4176 => x"33",
          4177 => x"08",
          4178 => x"58",
          4179 => x"38",
          4180 => x"7b",
          4181 => x"7a",
          4182 => x"71",
          4183 => x"34",
          4184 => x"39",
          4185 => x"53",
          4186 => x"3f",
          4187 => x"2e",
          4188 => x"b9",
          4189 => x"08",
          4190 => x"08",
          4191 => x"5e",
          4192 => x"19",
          4193 => x"06",
          4194 => x"53",
          4195 => x"c2",
          4196 => x"54",
          4197 => x"1a",
          4198 => x"5c",
          4199 => x"81",
          4200 => x"08",
          4201 => x"a8",
          4202 => x"b9",
          4203 => x"7e",
          4204 => x"55",
          4205 => x"e3",
          4206 => x"52",
          4207 => x"7c",
          4208 => x"53",
          4209 => x"52",
          4210 => x"b9",
          4211 => x"fb",
          4212 => x"1a",
          4213 => x"08",
          4214 => x"08",
          4215 => x"fb",
          4216 => x"82",
          4217 => x"81",
          4218 => x"19",
          4219 => x"fa",
          4220 => x"76",
          4221 => x"3f",
          4222 => x"10",
          4223 => x"ff",
          4224 => x"1f",
          4225 => x"1f",
          4226 => x"88",
          4227 => x"06",
          4228 => x"70",
          4229 => x"0a",
          4230 => x"7d",
          4231 => x"b9",
          4232 => x"ba",
          4233 => x"bb",
          4234 => x"0d",
          4235 => x"7a",
          4236 => x"76",
          4237 => x"1a",
          4238 => x"08",
          4239 => x"d7",
          4240 => x"76",
          4241 => x"76",
          4242 => x"26",
          4243 => x"f0",
          4244 => x"2e",
          4245 => x"c8",
          4246 => x"c8",
          4247 => x"80",
          4248 => x"55",
          4249 => x"09",
          4250 => x"74",
          4251 => x"04",
          4252 => x"c8",
          4253 => x"51",
          4254 => x"b9",
          4255 => x"c8",
          4256 => x"2e",
          4257 => x"c8",
          4258 => x"dd",
          4259 => x"76",
          4260 => x"79",
          4261 => x"b9",
          4262 => x"84",
          4263 => x"72",
          4264 => x"b9",
          4265 => x"73",
          4266 => x"80",
          4267 => x"81",
          4268 => x"1a",
          4269 => x"57",
          4270 => x"fe",
          4271 => x"51",
          4272 => x"84",
          4273 => x"c8",
          4274 => x"7a",
          4275 => x"75",
          4276 => x"05",
          4277 => x"26",
          4278 => x"84",
          4279 => x"1a",
          4280 => x"0c",
          4281 => x"b9",
          4282 => x"b9",
          4283 => x"80",
          4284 => x"52",
          4285 => x"c8",
          4286 => x"c8",
          4287 => x"0d",
          4288 => x"b9",
          4289 => x"3d",
          4290 => x"58",
          4291 => x"38",
          4292 => x"38",
          4293 => x"55",
          4294 => x"75",
          4295 => x"2a",
          4296 => x"56",
          4297 => x"08",
          4298 => x"98",
          4299 => x"2e",
          4300 => x"19",
          4301 => x"05",
          4302 => x"b9",
          4303 => x"0b",
          4304 => x"04",
          4305 => x"ff",
          4306 => x"2b",
          4307 => x"9c",
          4308 => x"54",
          4309 => x"38",
          4310 => x"19",
          4311 => x"0c",
          4312 => x"ec",
          4313 => x"84",
          4314 => x"81",
          4315 => x"9e",
          4316 => x"c8",
          4317 => x"76",
          4318 => x"ff",
          4319 => x"0c",
          4320 => x"7f",
          4321 => x"5c",
          4322 => x"86",
          4323 => x"17",
          4324 => x"b2",
          4325 => x"9d",
          4326 => x"58",
          4327 => x"1a",
          4328 => x"f5",
          4329 => x"18",
          4330 => x"0c",
          4331 => x"8f",
          4332 => x"8a",
          4333 => x"06",
          4334 => x"51",
          4335 => x"5d",
          4336 => x"08",
          4337 => x"c8",
          4338 => x"08",
          4339 => x"38",
          4340 => x"17",
          4341 => x"84",
          4342 => x"b9",
          4343 => x"82",
          4344 => x"ff",
          4345 => x"08",
          4346 => x"c8",
          4347 => x"80",
          4348 => x"fe",
          4349 => x"27",
          4350 => x"29",
          4351 => x"b4",
          4352 => x"78",
          4353 => x"58",
          4354 => x"74",
          4355 => x"27",
          4356 => x"53",
          4357 => x"b2",
          4358 => x"38",
          4359 => x"18",
          4360 => x"8f",
          4361 => x"08",
          4362 => x"33",
          4363 => x"c8",
          4364 => x"08",
          4365 => x"1a",
          4366 => x"27",
          4367 => x"7b",
          4368 => x"38",
          4369 => x"08",
          4370 => x"51",
          4371 => x"19",
          4372 => x"55",
          4373 => x"38",
          4374 => x"1a",
          4375 => x"75",
          4376 => x"22",
          4377 => x"98",
          4378 => x"0b",
          4379 => x"04",
          4380 => x"84",
          4381 => x"98",
          4382 => x"2e",
          4383 => x"5a",
          4384 => x"82",
          4385 => x"55",
          4386 => x"94",
          4387 => x"52",
          4388 => x"84",
          4389 => x"ff",
          4390 => x"76",
          4391 => x"08",
          4392 => x"82",
          4393 => x"70",
          4394 => x"1d",
          4395 => x"78",
          4396 => x"71",
          4397 => x"55",
          4398 => x"43",
          4399 => x"75",
          4400 => x"5d",
          4401 => x"84",
          4402 => x"08",
          4403 => x"75",
          4404 => x"0c",
          4405 => x"19",
          4406 => x"51",
          4407 => x"c8",
          4408 => x"ef",
          4409 => x"34",
          4410 => x"84",
          4411 => x"1a",
          4412 => x"33",
          4413 => x"fe",
          4414 => x"a0",
          4415 => x"19",
          4416 => x"fe",
          4417 => x"06",
          4418 => x"06",
          4419 => x"18",
          4420 => x"1f",
          4421 => x"5e",
          4422 => x"55",
          4423 => x"75",
          4424 => x"38",
          4425 => x"1d",
          4426 => x"3d",
          4427 => x"8d",
          4428 => x"81",
          4429 => x"19",
          4430 => x"07",
          4431 => x"77",
          4432 => x"f3",
          4433 => x"83",
          4434 => x"11",
          4435 => x"52",
          4436 => x"38",
          4437 => x"79",
          4438 => x"62",
          4439 => x"8c",
          4440 => x"86",
          4441 => x"2e",
          4442 => x"dd",
          4443 => x"63",
          4444 => x"5e",
          4445 => x"ff",
          4446 => x"c0",
          4447 => x"57",
          4448 => x"05",
          4449 => x"7f",
          4450 => x"59",
          4451 => x"2e",
          4452 => x"0c",
          4453 => x"0d",
          4454 => x"5c",
          4455 => x"3f",
          4456 => x"c8",
          4457 => x"40",
          4458 => x"1b",
          4459 => x"b4",
          4460 => x"83",
          4461 => x"2e",
          4462 => x"54",
          4463 => x"33",
          4464 => x"08",
          4465 => x"57",
          4466 => x"81",
          4467 => x"58",
          4468 => x"8b",
          4469 => x"06",
          4470 => x"81",
          4471 => x"2a",
          4472 => x"ef",
          4473 => x"2e",
          4474 => x"7d",
          4475 => x"75",
          4476 => x"05",
          4477 => x"ff",
          4478 => x"e4",
          4479 => x"ab",
          4480 => x"38",
          4481 => x"70",
          4482 => x"05",
          4483 => x"5a",
          4484 => x"dc",
          4485 => x"ff",
          4486 => x"52",
          4487 => x"c8",
          4488 => x"2e",
          4489 => x"0c",
          4490 => x"1b",
          4491 => x"51",
          4492 => x"c8",
          4493 => x"a4",
          4494 => x"34",
          4495 => x"84",
          4496 => x"1c",
          4497 => x"33",
          4498 => x"fd",
          4499 => x"a0",
          4500 => x"1b",
          4501 => x"fd",
          4502 => x"ab",
          4503 => x"42",
          4504 => x"2a",
          4505 => x"38",
          4506 => x"70",
          4507 => x"59",
          4508 => x"81",
          4509 => x"51",
          4510 => x"5a",
          4511 => x"d9",
          4512 => x"fe",
          4513 => x"ac",
          4514 => x"33",
          4515 => x"c7",
          4516 => x"9a",
          4517 => x"42",
          4518 => x"70",
          4519 => x"55",
          4520 => x"18",
          4521 => x"33",
          4522 => x"75",
          4523 => x"fe",
          4524 => x"a1",
          4525 => x"10",
          4526 => x"1b",
          4527 => x"84",
          4528 => x"fe",
          4529 => x"8c",
          4530 => x"70",
          4531 => x"80",
          4532 => x"38",
          4533 => x"41",
          4534 => x"81",
          4535 => x"84",
          4536 => x"0d",
          4537 => x"bc",
          4538 => x"ea",
          4539 => x"13",
          4540 => x"5e",
          4541 => x"8c",
          4542 => x"74",
          4543 => x"10",
          4544 => x"f4",
          4545 => x"8c",
          4546 => x"81",
          4547 => x"59",
          4548 => x"02",
          4549 => x"58",
          4550 => x"80",
          4551 => x"94",
          4552 => x"58",
          4553 => x"77",
          4554 => x"81",
          4555 => x"ef",
          4556 => x"7a",
          4557 => x"b8",
          4558 => x"58",
          4559 => x"81",
          4560 => x"90",
          4561 => x"60",
          4562 => x"a1",
          4563 => x"25",
          4564 => x"38",
          4565 => x"57",
          4566 => x"b9",
          4567 => x"74",
          4568 => x"84",
          4569 => x"77",
          4570 => x"7a",
          4571 => x"79",
          4572 => x"81",
          4573 => x"38",
          4574 => x"a0",
          4575 => x"16",
          4576 => x"38",
          4577 => x"19",
          4578 => x"34",
          4579 => x"51",
          4580 => x"8b",
          4581 => x"27",
          4582 => x"e4",
          4583 => x"08",
          4584 => x"09",
          4585 => x"db",
          4586 => x"02",
          4587 => x"58",
          4588 => x"5b",
          4589 => x"8c",
          4590 => x"b9",
          4591 => x"51",
          4592 => x"56",
          4593 => x"84",
          4594 => x"98",
          4595 => x"08",
          4596 => x"33",
          4597 => x"82",
          4598 => x"18",
          4599 => x"3f",
          4600 => x"38",
          4601 => x"0c",
          4602 => x"08",
          4603 => x"2e",
          4604 => x"25",
          4605 => x"81",
          4606 => x"2e",
          4607 => x"ee",
          4608 => x"84",
          4609 => x"38",
          4610 => x"38",
          4611 => x"1b",
          4612 => x"08",
          4613 => x"38",
          4614 => x"84",
          4615 => x"1c",
          4616 => x"3f",
          4617 => x"38",
          4618 => x"0c",
          4619 => x"0b",
          4620 => x"70",
          4621 => x"74",
          4622 => x"7b",
          4623 => x"57",
          4624 => x"ff",
          4625 => x"08",
          4626 => x"7c",
          4627 => x"34",
          4628 => x"98",
          4629 => x"80",
          4630 => x"fe",
          4631 => x"51",
          4632 => x"56",
          4633 => x"c7",
          4634 => x"18",
          4635 => x"51",
          4636 => x"77",
          4637 => x"84",
          4638 => x"18",
          4639 => x"a0",
          4640 => x"33",
          4641 => x"84",
          4642 => x"7f",
          4643 => x"53",
          4644 => x"b9",
          4645 => x"fe",
          4646 => x"56",
          4647 => x"81",
          4648 => x"5a",
          4649 => x"06",
          4650 => x"38",
          4651 => x"41",
          4652 => x"1c",
          4653 => x"33",
          4654 => x"82",
          4655 => x"1c",
          4656 => x"3f",
          4657 => x"38",
          4658 => x"0c",
          4659 => x"1c",
          4660 => x"06",
          4661 => x"8f",
          4662 => x"34",
          4663 => x"34",
          4664 => x"5a",
          4665 => x"8b",
          4666 => x"1b",
          4667 => x"33",
          4668 => x"05",
          4669 => x"75",
          4670 => x"57",
          4671 => x"38",
          4672 => x"38",
          4673 => x"76",
          4674 => x"34",
          4675 => x"7d",
          4676 => x"08",
          4677 => x"38",
          4678 => x"38",
          4679 => x"08",
          4680 => x"33",
          4681 => x"84",
          4682 => x"b9",
          4683 => x"08",
          4684 => x"08",
          4685 => x"fb",
          4686 => x"82",
          4687 => x"81",
          4688 => x"05",
          4689 => x"cf",
          4690 => x"76",
          4691 => x"56",
          4692 => x"fa",
          4693 => x"57",
          4694 => x"fa",
          4695 => x"fe",
          4696 => x"53",
          4697 => x"92",
          4698 => x"09",
          4699 => x"08",
          4700 => x"1d",
          4701 => x"27",
          4702 => x"82",
          4703 => x"56",
          4704 => x"58",
          4705 => x"87",
          4706 => x"81",
          4707 => x"fe",
          4708 => x"1c",
          4709 => x"52",
          4710 => x"fc",
          4711 => x"a0",
          4712 => x"18",
          4713 => x"39",
          4714 => x"40",
          4715 => x"98",
          4716 => x"ac",
          4717 => x"80",
          4718 => x"22",
          4719 => x"2e",
          4720 => x"22",
          4721 => x"95",
          4722 => x"ff",
          4723 => x"26",
          4724 => x"11",
          4725 => x"d4",
          4726 => x"30",
          4727 => x"94",
          4728 => x"80",
          4729 => x"1c",
          4730 => x"56",
          4731 => x"85",
          4732 => x"70",
          4733 => x"5b",
          4734 => x"80",
          4735 => x"05",
          4736 => x"70",
          4737 => x"8a",
          4738 => x"88",
          4739 => x"96",
          4740 => x"81",
          4741 => x"81",
          4742 => x"0b",
          4743 => x"11",
          4744 => x"89",
          4745 => x"13",
          4746 => x"9c",
          4747 => x"71",
          4748 => x"14",
          4749 => x"33",
          4750 => x"33",
          4751 => x"5f",
          4752 => x"77",
          4753 => x"16",
          4754 => x"7b",
          4755 => x"81",
          4756 => x"96",
          4757 => x"57",
          4758 => x"07",
          4759 => x"c8",
          4760 => x"ff",
          4761 => x"81",
          4762 => x"7a",
          4763 => x"05",
          4764 => x"5b",
          4765 => x"57",
          4766 => x"39",
          4767 => x"80",
          4768 => x"57",
          4769 => x"81",
          4770 => x"08",
          4771 => x"1f",
          4772 => x"fe",
          4773 => x"59",
          4774 => x"5a",
          4775 => x"1c",
          4776 => x"76",
          4777 => x"72",
          4778 => x"38",
          4779 => x"55",
          4780 => x"34",
          4781 => x"89",
          4782 => x"79",
          4783 => x"83",
          4784 => x"70",
          4785 => x"5d",
          4786 => x"0d",
          4787 => x"80",
          4788 => x"af",
          4789 => x"dc",
          4790 => x"81",
          4791 => x"0c",
          4792 => x"42",
          4793 => x"73",
          4794 => x"61",
          4795 => x"53",
          4796 => x"73",
          4797 => x"ff",
          4798 => x"56",
          4799 => x"83",
          4800 => x"30",
          4801 => x"57",
          4802 => x"74",
          4803 => x"80",
          4804 => x"0b",
          4805 => x"06",
          4806 => x"ab",
          4807 => x"16",
          4808 => x"54",
          4809 => x"06",
          4810 => x"fe",
          4811 => x"5d",
          4812 => x"70",
          4813 => x"73",
          4814 => x"39",
          4815 => x"70",
          4816 => x"55",
          4817 => x"70",
          4818 => x"72",
          4819 => x"32",
          4820 => x"51",
          4821 => x"1d",
          4822 => x"41",
          4823 => x"38",
          4824 => x"81",
          4825 => x"83",
          4826 => x"38",
          4827 => x"93",
          4828 => x"70",
          4829 => x"2e",
          4830 => x"0b",
          4831 => x"de",
          4832 => x"b9",
          4833 => x"73",
          4834 => x"25",
          4835 => x"80",
          4836 => x"62",
          4837 => x"2e",
          4838 => x"30",
          4839 => x"59",
          4840 => x"75",
          4841 => x"84",
          4842 => x"38",
          4843 => x"38",
          4844 => x"22",
          4845 => x"2a",
          4846 => x"ae",
          4847 => x"17",
          4848 => x"19",
          4849 => x"fe",
          4850 => x"ff",
          4851 => x"7a",
          4852 => x"ff",
          4853 => x"f1",
          4854 => x"19",
          4855 => x"ae",
          4856 => x"05",
          4857 => x"8f",
          4858 => x"7c",
          4859 => x"8b",
          4860 => x"70",
          4861 => x"72",
          4862 => x"78",
          4863 => x"54",
          4864 => x"74",
          4865 => x"32",
          4866 => x"54",
          4867 => x"83",
          4868 => x"83",
          4869 => x"30",
          4870 => x"07",
          4871 => x"83",
          4872 => x"38",
          4873 => x"07",
          4874 => x"56",
          4875 => x"fc",
          4876 => x"15",
          4877 => x"74",
          4878 => x"76",
          4879 => x"88",
          4880 => x"58",
          4881 => x"83",
          4882 => x"38",
          4883 => x"9d",
          4884 => x"2e",
          4885 => x"82",
          4886 => x"85",
          4887 => x"1d",
          4888 => x"b9",
          4889 => x"84",
          4890 => x"38",
          4891 => x"81",
          4892 => x"81",
          4893 => x"38",
          4894 => x"82",
          4895 => x"73",
          4896 => x"f9",
          4897 => x"11",
          4898 => x"a0",
          4899 => x"85",
          4900 => x"39",
          4901 => x"09",
          4902 => x"54",
          4903 => x"a0",
          4904 => x"23",
          4905 => x"54",
          4906 => x"73",
          4907 => x"13",
          4908 => x"a0",
          4909 => x"51",
          4910 => x"ab",
          4911 => x"08",
          4912 => x"06",
          4913 => x"33",
          4914 => x"74",
          4915 => x"08",
          4916 => x"11",
          4917 => x"2b",
          4918 => x"7d",
          4919 => x"1d",
          4920 => x"b7",
          4921 => x"fe",
          4922 => x"88",
          4923 => x"76",
          4924 => x"82",
          4925 => x"59",
          4926 => x"fd",
          4927 => x"98",
          4928 => x"88",
          4929 => x"d6",
          4930 => x"80",
          4931 => x"0d",
          4932 => x"81",
          4933 => x"1d",
          4934 => x"79",
          4935 => x"5a",
          4936 => x"83",
          4937 => x"3f",
          4938 => x"06",
          4939 => x"78",
          4940 => x"06",
          4941 => x"74",
          4942 => x"80",
          4943 => x"0b",
          4944 => x"06",
          4945 => x"e0",
          4946 => x"19",
          4947 => x"54",
          4948 => x"06",
          4949 => x"15",
          4950 => x"82",
          4951 => x"ff",
          4952 => x"38",
          4953 => x"e0",
          4954 => x"56",
          4955 => x"74",
          4956 => x"55",
          4957 => x"39",
          4958 => x"06",
          4959 => x"38",
          4960 => x"a0",
          4961 => x"81",
          4962 => x"33",
          4963 => x"71",
          4964 => x"0c",
          4965 => x"a0",
          4966 => x"74",
          4967 => x"5a",
          4968 => x"ff",
          4969 => x"33",
          4970 => x"81",
          4971 => x"74",
          4972 => x"f2",
          4973 => x"93",
          4974 => x"69",
          4975 => x"42",
          4976 => x"08",
          4977 => x"85",
          4978 => x"33",
          4979 => x"2e",
          4980 => x"ba",
          4981 => x"33",
          4982 => x"75",
          4983 => x"08",
          4984 => x"85",
          4985 => x"fe",
          4986 => x"2e",
          4987 => x"bb",
          4988 => x"ff",
          4989 => x"80",
          4990 => x"75",
          4991 => x"81",
          4992 => x"51",
          4993 => x"08",
          4994 => x"56",
          4995 => x"80",
          4996 => x"06",
          4997 => x"80",
          4998 => x"b4",
          4999 => x"54",
          5000 => x"18",
          5001 => x"84",
          5002 => x"ff",
          5003 => x"84",
          5004 => x"33",
          5005 => x"07",
          5006 => x"d5",
          5007 => x"8b",
          5008 => x"61",
          5009 => x"2e",
          5010 => x"26",
          5011 => x"80",
          5012 => x"5e",
          5013 => x"06",
          5014 => x"80",
          5015 => x"57",
          5016 => x"83",
          5017 => x"2b",
          5018 => x"70",
          5019 => x"07",
          5020 => x"75",
          5021 => x"82",
          5022 => x"11",
          5023 => x"8d",
          5024 => x"78",
          5025 => x"c5",
          5026 => x"18",
          5027 => x"c4",
          5028 => x"87",
          5029 => x"c9",
          5030 => x"40",
          5031 => x"06",
          5032 => x"38",
          5033 => x"33",
          5034 => x"a4",
          5035 => x"82",
          5036 => x"2b",
          5037 => x"88",
          5038 => x"5a",
          5039 => x"33",
          5040 => x"07",
          5041 => x"81",
          5042 => x"05",
          5043 => x"78",
          5044 => x"fd",
          5045 => x"b9",
          5046 => x"84",
          5047 => x"f5",
          5048 => x"ff",
          5049 => x"9f",
          5050 => x"82",
          5051 => x"19",
          5052 => x"7b",
          5053 => x"83",
          5054 => x"5c",
          5055 => x"38",
          5056 => x"55",
          5057 => x"19",
          5058 => x"56",
          5059 => x"8d",
          5060 => x"38",
          5061 => x"90",
          5062 => x"34",
          5063 => x"77",
          5064 => x"5d",
          5065 => x"18",
          5066 => x"0c",
          5067 => x"77",
          5068 => x"04",
          5069 => x"3d",
          5070 => x"81",
          5071 => x"26",
          5072 => x"06",
          5073 => x"87",
          5074 => x"b8",
          5075 => x"5b",
          5076 => x"70",
          5077 => x"5a",
          5078 => x"e0",
          5079 => x"ff",
          5080 => x"38",
          5081 => x"55",
          5082 => x"75",
          5083 => x"77",
          5084 => x"30",
          5085 => x"5d",
          5086 => x"38",
          5087 => x"7c",
          5088 => x"a9",
          5089 => x"77",
          5090 => x"7d",
          5091 => x"39",
          5092 => x"e9",
          5093 => x"59",
          5094 => x"80",
          5095 => x"83",
          5096 => x"a6",
          5097 => x"59",
          5098 => x"7a",
          5099 => x"33",
          5100 => x"71",
          5101 => x"70",
          5102 => x"33",
          5103 => x"40",
          5104 => x"ff",
          5105 => x"25",
          5106 => x"33",
          5107 => x"31",
          5108 => x"05",
          5109 => x"5b",
          5110 => x"80",
          5111 => x"18",
          5112 => x"55",
          5113 => x"81",
          5114 => x"17",
          5115 => x"b9",
          5116 => x"55",
          5117 => x"58",
          5118 => x"33",
          5119 => x"58",
          5120 => x"06",
          5121 => x"57",
          5122 => x"38",
          5123 => x"80",
          5124 => x"bc",
          5125 => x"82",
          5126 => x"0b",
          5127 => x"7b",
          5128 => x"81",
          5129 => x"77",
          5130 => x"84",
          5131 => x"d1",
          5132 => x"ee",
          5133 => x"7b",
          5134 => x"81",
          5135 => x"1b",
          5136 => x"80",
          5137 => x"85",
          5138 => x"40",
          5139 => x"33",
          5140 => x"71",
          5141 => x"77",
          5142 => x"2e",
          5143 => x"8d",
          5144 => x"b9",
          5145 => x"58",
          5146 => x"0b",
          5147 => x"5d",
          5148 => x"b9",
          5149 => x"0b",
          5150 => x"5a",
          5151 => x"7a",
          5152 => x"31",
          5153 => x"80",
          5154 => x"e1",
          5155 => x"e4",
          5156 => x"05",
          5157 => x"33",
          5158 => x"42",
          5159 => x"75",
          5160 => x"57",
          5161 => x"58",
          5162 => x"80",
          5163 => x"57",
          5164 => x"f9",
          5165 => x"b4",
          5166 => x"17",
          5167 => x"06",
          5168 => x"b8",
          5169 => x"b0",
          5170 => x"2e",
          5171 => x"b4",
          5172 => x"84",
          5173 => x"b6",
          5174 => x"5e",
          5175 => x"06",
          5176 => x"33",
          5177 => x"88",
          5178 => x"07",
          5179 => x"41",
          5180 => x"8b",
          5181 => x"f8",
          5182 => x"33",
          5183 => x"88",
          5184 => x"07",
          5185 => x"44",
          5186 => x"8a",
          5187 => x"f8",
          5188 => x"33",
          5189 => x"88",
          5190 => x"07",
          5191 => x"1e",
          5192 => x"33",
          5193 => x"88",
          5194 => x"07",
          5195 => x"90",
          5196 => x"45",
          5197 => x"34",
          5198 => x"7c",
          5199 => x"23",
          5200 => x"80",
          5201 => x"7b",
          5202 => x"7f",
          5203 => x"b4",
          5204 => x"81",
          5205 => x"3f",
          5206 => x"81",
          5207 => x"08",
          5208 => x"18",
          5209 => x"27",
          5210 => x"82",
          5211 => x"08",
          5212 => x"80",
          5213 => x"8a",
          5214 => x"fc",
          5215 => x"e2",
          5216 => x"5a",
          5217 => x"17",
          5218 => x"e4",
          5219 => x"71",
          5220 => x"14",
          5221 => x"33",
          5222 => x"82",
          5223 => x"f5",
          5224 => x"f9",
          5225 => x"75",
          5226 => x"77",
          5227 => x"75",
          5228 => x"39",
          5229 => x"08",
          5230 => x"51",
          5231 => x"f0",
          5232 => x"64",
          5233 => x"ff",
          5234 => x"e9",
          5235 => x"70",
          5236 => x"80",
          5237 => x"2e",
          5238 => x"54",
          5239 => x"10",
          5240 => x"55",
          5241 => x"74",
          5242 => x"38",
          5243 => x"0c",
          5244 => x"80",
          5245 => x"51",
          5246 => x"54",
          5247 => x"0d",
          5248 => x"92",
          5249 => x"70",
          5250 => x"89",
          5251 => x"ff",
          5252 => x"2e",
          5253 => x"e5",
          5254 => x"59",
          5255 => x"78",
          5256 => x"12",
          5257 => x"38",
          5258 => x"54",
          5259 => x"89",
          5260 => x"57",
          5261 => x"54",
          5262 => x"38",
          5263 => x"70",
          5264 => x"07",
          5265 => x"38",
          5266 => x"7b",
          5267 => x"98",
          5268 => x"79",
          5269 => x"3d",
          5270 => x"05",
          5271 => x"2e",
          5272 => x"9d",
          5273 => x"05",
          5274 => x"c8",
          5275 => x"2e",
          5276 => x"75",
          5277 => x"04",
          5278 => x"52",
          5279 => x"08",
          5280 => x"81",
          5281 => x"80",
          5282 => x"83",
          5283 => x"38",
          5284 => x"38",
          5285 => x"80",
          5286 => x"33",
          5287 => x"61",
          5288 => x"7d",
          5289 => x"8e",
          5290 => x"a1",
          5291 => x"91",
          5292 => x"17",
          5293 => x"9a",
          5294 => x"7d",
          5295 => x"38",
          5296 => x"80",
          5297 => x"1c",
          5298 => x"55",
          5299 => x"2e",
          5300 => x"7d",
          5301 => x"7c",
          5302 => x"26",
          5303 => x"0c",
          5304 => x"33",
          5305 => x"25",
          5306 => x"5e",
          5307 => x"82",
          5308 => x"84",
          5309 => x"91",
          5310 => x"7d",
          5311 => x"5a",
          5312 => x"81",
          5313 => x"77",
          5314 => x"08",
          5315 => x"67",
          5316 => x"88",
          5317 => x"57",
          5318 => x"7a",
          5319 => x"33",
          5320 => x"88",
          5321 => x"07",
          5322 => x"60",
          5323 => x"52",
          5324 => x"22",
          5325 => x"80",
          5326 => x"1a",
          5327 => x"74",
          5328 => x"2e",
          5329 => x"8a",
          5330 => x"5b",
          5331 => x"25",
          5332 => x"38",
          5333 => x"80",
          5334 => x"51",
          5335 => x"08",
          5336 => x"83",
          5337 => x"ff",
          5338 => x"56",
          5339 => x"91",
          5340 => x"2a",
          5341 => x"b8",
          5342 => x"ed",
          5343 => x"e5",
          5344 => x"dd",
          5345 => x"b9",
          5346 => x"76",
          5347 => x"76",
          5348 => x"95",
          5349 => x"2b",
          5350 => x"5e",
          5351 => x"7b",
          5352 => x"51",
          5353 => x"08",
          5354 => x"81",
          5355 => x"2e",
          5356 => x"ff",
          5357 => x"52",
          5358 => x"b9",
          5359 => x"08",
          5360 => x"5b",
          5361 => x"16",
          5362 => x"07",
          5363 => x"7a",
          5364 => x"39",
          5365 => x"95",
          5366 => x"33",
          5367 => x"90",
          5368 => x"80",
          5369 => x"17",
          5370 => x"cc",
          5371 => x"0b",
          5372 => x"80",
          5373 => x"17",
          5374 => x"09",
          5375 => x"39",
          5376 => x"5d",
          5377 => x"83",
          5378 => x"81",
          5379 => x"b8",
          5380 => x"a3",
          5381 => x"2e",
          5382 => x"b4",
          5383 => x"90",
          5384 => x"bc",
          5385 => x"81",
          5386 => x"70",
          5387 => x"a4",
          5388 => x"2e",
          5389 => x"b9",
          5390 => x"08",
          5391 => x"08",
          5392 => x"ff",
          5393 => x"82",
          5394 => x"81",
          5395 => x"05",
          5396 => x"ff",
          5397 => x"39",
          5398 => x"af",
          5399 => x"a2",
          5400 => x"80",
          5401 => x"9c",
          5402 => x"77",
          5403 => x"22",
          5404 => x"56",
          5405 => x"75",
          5406 => x"56",
          5407 => x"76",
          5408 => x"79",
          5409 => x"08",
          5410 => x"81",
          5411 => x"3d",
          5412 => x"5d",
          5413 => x"80",
          5414 => x"80",
          5415 => x"80",
          5416 => x"1b",
          5417 => x"b7",
          5418 => x"76",
          5419 => x"74",
          5420 => x"06",
          5421 => x"ed",
          5422 => x"71",
          5423 => x"ef",
          5424 => x"60",
          5425 => x"81",
          5426 => x"76",
          5427 => x"75",
          5428 => x"81",
          5429 => x"2e",
          5430 => x"60",
          5431 => x"1a",
          5432 => x"27",
          5433 => x"78",
          5434 => x"74",
          5435 => x"7c",
          5436 => x"83",
          5437 => x"27",
          5438 => x"54",
          5439 => x"51",
          5440 => x"08",
          5441 => x"57",
          5442 => x"19",
          5443 => x"9e",
          5444 => x"b8",
          5445 => x"05",
          5446 => x"34",
          5447 => x"89",
          5448 => x"19",
          5449 => x"1a",
          5450 => x"7b",
          5451 => x"b9",
          5452 => x"84",
          5453 => x"74",
          5454 => x"57",
          5455 => x"31",
          5456 => x"7b",
          5457 => x"2e",
          5458 => x"71",
          5459 => x"81",
          5460 => x"53",
          5461 => x"ff",
          5462 => x"80",
          5463 => x"75",
          5464 => x"60",
          5465 => x"79",
          5466 => x"77",
          5467 => x"81",
          5468 => x"59",
          5469 => x"fe",
          5470 => x"33",
          5471 => x"16",
          5472 => x"81",
          5473 => x"70",
          5474 => x"9e",
          5475 => x"08",
          5476 => x"38",
          5477 => x"b4",
          5478 => x"b9",
          5479 => x"08",
          5480 => x"55",
          5481 => x"d4",
          5482 => x"1a",
          5483 => x"33",
          5484 => x"fe",
          5485 => x"1a",
          5486 => x"08",
          5487 => x"84",
          5488 => x"81",
          5489 => x"84",
          5490 => x"fb",
          5491 => x"fb",
          5492 => x"81",
          5493 => x"0d",
          5494 => x"0b",
          5495 => x"04",
          5496 => x"40",
          5497 => x"57",
          5498 => x"56",
          5499 => x"55",
          5500 => x"22",
          5501 => x"2e",
          5502 => x"76",
          5503 => x"33",
          5504 => x"33",
          5505 => x"87",
          5506 => x"94",
          5507 => x"77",
          5508 => x"80",
          5509 => x"06",
          5510 => x"11",
          5511 => x"5a",
          5512 => x"38",
          5513 => x"84",
          5514 => x"38",
          5515 => x"98",
          5516 => x"74",
          5517 => x"08",
          5518 => x"98",
          5519 => x"fe",
          5520 => x"f0",
          5521 => x"b0",
          5522 => x"2e",
          5523 => x"2a",
          5524 => x"38",
          5525 => x"38",
          5526 => x"53",
          5527 => x"9b",
          5528 => x"a1",
          5529 => x"56",
          5530 => x"80",
          5531 => x"57",
          5532 => x"33",
          5533 => x"16",
          5534 => x"83",
          5535 => x"79",
          5536 => x"1e",
          5537 => x"1f",
          5538 => x"5e",
          5539 => x"56",
          5540 => x"38",
          5541 => x"07",
          5542 => x"75",
          5543 => x"04",
          5544 => x"0d",
          5545 => x"c8",
          5546 => x"9c",
          5547 => x"06",
          5548 => x"79",
          5549 => x"b4",
          5550 => x"0b",
          5551 => x"7f",
          5552 => x"38",
          5553 => x"81",
          5554 => x"84",
          5555 => x"ff",
          5556 => x"7b",
          5557 => x"83",
          5558 => x"7e",
          5559 => x"38",
          5560 => x"70",
          5561 => x"75",
          5562 => x"19",
          5563 => x"16",
          5564 => x"17",
          5565 => x"81",
          5566 => x"09",
          5567 => x"c8",
          5568 => x"a8",
          5569 => x"5d",
          5570 => x"f0",
          5571 => x"2e",
          5572 => x"54",
          5573 => x"53",
          5574 => x"98",
          5575 => x"94",
          5576 => x"26",
          5577 => x"81",
          5578 => x"94",
          5579 => x"1c",
          5580 => x"08",
          5581 => x"84",
          5582 => x"08",
          5583 => x"fd",
          5584 => x"ab",
          5585 => x"84",
          5586 => x"39",
          5587 => x"16",
          5588 => x"ff",
          5589 => x"81",
          5590 => x"17",
          5591 => x"31",
          5592 => x"89",
          5593 => x"2e",
          5594 => x"54",
          5595 => x"53",
          5596 => x"96",
          5597 => x"81",
          5598 => x"84",
          5599 => x"f9",
          5600 => x"f9",
          5601 => x"53",
          5602 => x"52",
          5603 => x"c8",
          5604 => x"08",
          5605 => x"17",
          5606 => x"27",
          5607 => x"77",
          5608 => x"38",
          5609 => x"08",
          5610 => x"51",
          5611 => x"12",
          5612 => x"f4",
          5613 => x"0b",
          5614 => x"04",
          5615 => x"84",
          5616 => x"f5",
          5617 => x"80",
          5618 => x"80",
          5619 => x"80",
          5620 => x"19",
          5621 => x"b5",
          5622 => x"79",
          5623 => x"86",
          5624 => x"2e",
          5625 => x"5a",
          5626 => x"38",
          5627 => x"38",
          5628 => x"81",
          5629 => x"84",
          5630 => x"ff",
          5631 => x"75",
          5632 => x"11",
          5633 => x"18",
          5634 => x"83",
          5635 => x"9a",
          5636 => x"9b",
          5637 => x"19",
          5638 => x"c1",
          5639 => x"34",
          5640 => x"34",
          5641 => x"34",
          5642 => x"34",
          5643 => x"34",
          5644 => x"0b",
          5645 => x"34",
          5646 => x"81",
          5647 => x"96",
          5648 => x"19",
          5649 => x"90",
          5650 => x"8d",
          5651 => x"08",
          5652 => x"33",
          5653 => x"56",
          5654 => x"84",
          5655 => x"17",
          5656 => x"c8",
          5657 => x"27",
          5658 => x"74",
          5659 => x"38",
          5660 => x"08",
          5661 => x"51",
          5662 => x"e8",
          5663 => x"18",
          5664 => x"18",
          5665 => x"34",
          5666 => x"34",
          5667 => x"34",
          5668 => x"34",
          5669 => x"34",
          5670 => x"0b",
          5671 => x"34",
          5672 => x"81",
          5673 => x"94",
          5674 => x"19",
          5675 => x"90",
          5676 => x"33",
          5677 => x"c8",
          5678 => x"38",
          5679 => x"39",
          5680 => x"fb",
          5681 => x"84",
          5682 => x"74",
          5683 => x"72",
          5684 => x"71",
          5685 => x"84",
          5686 => x"96",
          5687 => x"75",
          5688 => x"b9",
          5689 => x"13",
          5690 => x"b9",
          5691 => x"38",
          5692 => x"f6",
          5693 => x"5b",
          5694 => x"81",
          5695 => x"52",
          5696 => x"38",
          5697 => x"a4",
          5698 => x"70",
          5699 => x"b9",
          5700 => x"0b",
          5701 => x"04",
          5702 => x"06",
          5703 => x"38",
          5704 => x"05",
          5705 => x"38",
          5706 => x"79",
          5707 => x"05",
          5708 => x"33",
          5709 => x"99",
          5710 => x"ff",
          5711 => x"70",
          5712 => x"81",
          5713 => x"9f",
          5714 => x"81",
          5715 => x"74",
          5716 => x"9f",
          5717 => x"80",
          5718 => x"5b",
          5719 => x"7a",
          5720 => x"f7",
          5721 => x"39",
          5722 => x"cc",
          5723 => x"3f",
          5724 => x"c8",
          5725 => x"b9",
          5726 => x"5c",
          5727 => x"c5",
          5728 => x"84",
          5729 => x"80",
          5730 => x"5a",
          5731 => x"b2",
          5732 => x"57",
          5733 => x"63",
          5734 => x"88",
          5735 => x"57",
          5736 => x"98",
          5737 => x"98",
          5738 => x"84",
          5739 => x"85",
          5740 => x"0d",
          5741 => x"71",
          5742 => x"07",
          5743 => x"7a",
          5744 => x"b9",
          5745 => x"9e",
          5746 => x"e6",
          5747 => x"80",
          5748 => x"52",
          5749 => x"84",
          5750 => x"08",
          5751 => x"0c",
          5752 => x"3d",
          5753 => x"58",
          5754 => x"d8",
          5755 => x"7a",
          5756 => x"c8",
          5757 => x"92",
          5758 => x"56",
          5759 => x"84",
          5760 => x"5d",
          5761 => x"53",
          5762 => x"ff",
          5763 => x"80",
          5764 => x"76",
          5765 => x"80",
          5766 => x"12",
          5767 => x"33",
          5768 => x"2e",
          5769 => x"0c",
          5770 => x"3f",
          5771 => x"c8",
          5772 => x"51",
          5773 => x"08",
          5774 => x"80",
          5775 => x"12",
          5776 => x"33",
          5777 => x"2e",
          5778 => x"38",
          5779 => x"ff",
          5780 => x"59",
          5781 => x"b4",
          5782 => x"78",
          5783 => x"b8",
          5784 => x"3f",
          5785 => x"79",
          5786 => x"81",
          5787 => x"57",
          5788 => x"78",
          5789 => x"9c",
          5790 => x"18",
          5791 => x"ff",
          5792 => x"75",
          5793 => x"e6",
          5794 => x"34",
          5795 => x"bd",
          5796 => x"80",
          5797 => x"10",
          5798 => x"33",
          5799 => x"2e",
          5800 => x"33",
          5801 => x"1a",
          5802 => x"57",
          5803 => x"5f",
          5804 => x"34",
          5805 => x"38",
          5806 => x"76",
          5807 => x"38",
          5808 => x"b9",
          5809 => x"95",
          5810 => x"2b",
          5811 => x"56",
          5812 => x"94",
          5813 => x"2b",
          5814 => x"5a",
          5815 => x"ce",
          5816 => x"b9",
          5817 => x"ff",
          5818 => x"53",
          5819 => x"52",
          5820 => x"84",
          5821 => x"b9",
          5822 => x"08",
          5823 => x"08",
          5824 => x"fc",
          5825 => x"82",
          5826 => x"81",
          5827 => x"05",
          5828 => x"ff",
          5829 => x"39",
          5830 => x"5c",
          5831 => x"d1",
          5832 => x"b8",
          5833 => x"59",
          5834 => x"06",
          5835 => x"e5",
          5836 => x"79",
          5837 => x"77",
          5838 => x"3d",
          5839 => x"33",
          5840 => x"78",
          5841 => x"59",
          5842 => x"0c",
          5843 => x"0d",
          5844 => x"80",
          5845 => x"80",
          5846 => x"80",
          5847 => x"16",
          5848 => x"a0",
          5849 => x"75",
          5850 => x"72",
          5851 => x"76",
          5852 => x"08",
          5853 => x"cc",
          5854 => x"2b",
          5855 => x"f7",
          5856 => x"bb",
          5857 => x"15",
          5858 => x"bb",
          5859 => x"26",
          5860 => x"70",
          5861 => x"17",
          5862 => x"82",
          5863 => x"38",
          5864 => x"94",
          5865 => x"2a",
          5866 => x"2e",
          5867 => x"ff",
          5868 => x"54",
          5869 => x"a3",
          5870 => x"74",
          5871 => x"9c",
          5872 => x"98",
          5873 => x"91",
          5874 => x"c8",
          5875 => x"33",
          5876 => x"73",
          5877 => x"55",
          5878 => x"81",
          5879 => x"0c",
          5880 => x"90",
          5881 => x"33",
          5882 => x"34",
          5883 => x"2e",
          5884 => x"85",
          5885 => x"84",
          5886 => x"80",
          5887 => x"54",
          5888 => x"98",
          5889 => x"38",
          5890 => x"57",
          5891 => x"76",
          5892 => x"a9",
          5893 => x"fe",
          5894 => x"80",
          5895 => x"29",
          5896 => x"11",
          5897 => x"df",
          5898 => x"39",
          5899 => x"3f",
          5900 => x"39",
          5901 => x"3f",
          5902 => x"72",
          5903 => x"56",
          5904 => x"ff",
          5905 => x"54",
          5906 => x"38",
          5907 => x"ed",
          5908 => x"0c",
          5909 => x"82",
          5910 => x"b9",
          5911 => x"3d",
          5912 => x"2e",
          5913 => x"05",
          5914 => x"9b",
          5915 => x"b9",
          5916 => x"76",
          5917 => x"0c",
          5918 => x"7d",
          5919 => x"84",
          5920 => x"08",
          5921 => x"98",
          5922 => x"38",
          5923 => x"06",
          5924 => x"38",
          5925 => x"12",
          5926 => x"33",
          5927 => x"2e",
          5928 => x"58",
          5929 => x"52",
          5930 => x"b9",
          5931 => x"38",
          5932 => x"76",
          5933 => x"76",
          5934 => x"94",
          5935 => x"2b",
          5936 => x"5a",
          5937 => x"55",
          5938 => x"74",
          5939 => x"72",
          5940 => x"86",
          5941 => x"71",
          5942 => x"57",
          5943 => x"84",
          5944 => x"81",
          5945 => x"84",
          5946 => x"dc",
          5947 => x"39",
          5948 => x"89",
          5949 => x"08",
          5950 => x"33",
          5951 => x"14",
          5952 => x"78",
          5953 => x"59",
          5954 => x"80",
          5955 => x"51",
          5956 => x"08",
          5957 => x"b5",
          5958 => x"76",
          5959 => x"72",
          5960 => x"84",
          5961 => x"70",
          5962 => x"08",
          5963 => x"c8",
          5964 => x"53",
          5965 => x"72",
          5966 => x"84",
          5967 => x"70",
          5968 => x"08",
          5969 => x"52",
          5970 => x"b9",
          5971 => x"3d",
          5972 => x"fd",
          5973 => x"06",
          5974 => x"08",
          5975 => x"0d",
          5976 => x"53",
          5977 => x"84",
          5978 => x"08",
          5979 => x"c8",
          5980 => x"75",
          5981 => x"c8",
          5982 => x"38",
          5983 => x"2b",
          5984 => x"76",
          5985 => x"51",
          5986 => x"c8",
          5987 => x"84",
          5988 => x"ed",
          5989 => x"53",
          5990 => x"51",
          5991 => x"5a",
          5992 => x"75",
          5993 => x"11",
          5994 => x"75",
          5995 => x"79",
          5996 => x"04",
          5997 => x"5b",
          5998 => x"a8",
          5999 => x"5d",
          6000 => x"1d",
          6001 => x"76",
          6002 => x"78",
          6003 => x"54",
          6004 => x"33",
          6005 => x"c8",
          6006 => x"81",
          6007 => x"5b",
          6008 => x"5e",
          6009 => x"17",
          6010 => x"33",
          6011 => x"81",
          6012 => x"75",
          6013 => x"06",
          6014 => x"05",
          6015 => x"ff",
          6016 => x"53",
          6017 => x"38",
          6018 => x"84",
          6019 => x"18",
          6020 => x"3d",
          6021 => x"53",
          6022 => x"52",
          6023 => x"84",
          6024 => x"b9",
          6025 => x"08",
          6026 => x"08",
          6027 => x"fe",
          6028 => x"82",
          6029 => x"81",
          6030 => x"05",
          6031 => x"fe",
          6032 => x"39",
          6033 => x"75",
          6034 => x"84",
          6035 => x"38",
          6036 => x"f7",
          6037 => x"84",
          6038 => x"05",
          6039 => x"9c",
          6040 => x"7f",
          6041 => x"33",
          6042 => x"fe",
          6043 => x"11",
          6044 => x"70",
          6045 => x"83",
          6046 => x"59",
          6047 => x"fe",
          6048 => x"81",
          6049 => x"94",
          6050 => x"58",
          6051 => x"82",
          6052 => x"0d",
          6053 => x"9f",
          6054 => x"97",
          6055 => x"8f",
          6056 => x"59",
          6057 => x"80",
          6058 => x"91",
          6059 => x"90",
          6060 => x"55",
          6061 => x"c4",
          6062 => x"18",
          6063 => x"38",
          6064 => x"81",
          6065 => x"74",
          6066 => x"88",
          6067 => x"0c",
          6068 => x"18",
          6069 => x"91",
          6070 => x"c8",
          6071 => x"78",
          6072 => x"76",
          6073 => x"c8",
          6074 => x"2e",
          6075 => x"81",
          6076 => x"08",
          6077 => x"73",
          6078 => x"84",
          6079 => x"16",
          6080 => x"55",
          6081 => x"81",
          6082 => x"81",
          6083 => x"54",
          6084 => x"39",
          6085 => x"3f",
          6086 => x"73",
          6087 => x"56",
          6088 => x"33",
          6089 => x"18",
          6090 => x"52",
          6091 => x"b9",
          6092 => x"84",
          6093 => x"38",
          6094 => x"b9",
          6095 => x"a1",
          6096 => x"08",
          6097 => x"84",
          6098 => x"84",
          6099 => x"81",
          6100 => x"ff",
          6101 => x"c7",
          6102 => x"b9",
          6103 => x"76",
          6104 => x"c8",
          6105 => x"2e",
          6106 => x"81",
          6107 => x"08",
          6108 => x"73",
          6109 => x"84",
          6110 => x"16",
          6111 => x"55",
          6112 => x"15",
          6113 => x"07",
          6114 => x"77",
          6115 => x"74",
          6116 => x"39",
          6117 => x"90",
          6118 => x"82",
          6119 => x"33",
          6120 => x"c8",
          6121 => x"fa",
          6122 => x"54",
          6123 => x"56",
          6124 => x"db",
          6125 => x"9c",
          6126 => x"fb",
          6127 => x"b9",
          6128 => x"84",
          6129 => x"7d",
          6130 => x"70",
          6131 => x"b9",
          6132 => x"de",
          6133 => x"85",
          6134 => x"77",
          6135 => x"7b",
          6136 => x"33",
          6137 => x"7b",
          6138 => x"9b",
          6139 => x"2b",
          6140 => x"58",
          6141 => x"84",
          6142 => x"80",
          6143 => x"7b",
          6144 => x"41",
          6145 => x"70",
          6146 => x"b9",
          6147 => x"fe",
          6148 => x"74",
          6149 => x"c8",
          6150 => x"38",
          6151 => x"3d",
          6152 => x"33",
          6153 => x"7d",
          6154 => x"84",
          6155 => x"84",
          6156 => x"08",
          6157 => x"74",
          6158 => x"78",
          6159 => x"c8",
          6160 => x"2e",
          6161 => x"80",
          6162 => x"38",
          6163 => x"08",
          6164 => x"9c",
          6165 => x"82",
          6166 => x"fe",
          6167 => x"84",
          6168 => x"b8",
          6169 => x"5a",
          6170 => x"38",
          6171 => x"7a",
          6172 => x"81",
          6173 => x"17",
          6174 => x"b9",
          6175 => x"56",
          6176 => x"56",
          6177 => x"e5",
          6178 => x"90",
          6179 => x"80",
          6180 => x"84",
          6181 => x"08",
          6182 => x"2e",
          6183 => x"56",
          6184 => x"08",
          6185 => x"fe",
          6186 => x"c8",
          6187 => x"a6",
          6188 => x"34",
          6189 => x"84",
          6190 => x"18",
          6191 => x"33",
          6192 => x"fe",
          6193 => x"a0",
          6194 => x"17",
          6195 => x"58",
          6196 => x"27",
          6197 => x"fe",
          6198 => x"5a",
          6199 => x"cb",
          6200 => x"fd",
          6201 => x"2e",
          6202 => x"76",
          6203 => x"c8",
          6204 => x"11",
          6205 => x"7b",
          6206 => x"18",
          6207 => x"7b",
          6208 => x"26",
          6209 => x"39",
          6210 => x"c8",
          6211 => x"fd",
          6212 => x"9f",
          6213 => x"51",
          6214 => x"08",
          6215 => x"8a",
          6216 => x"3d",
          6217 => x"3d",
          6218 => x"84",
          6219 => x"08",
          6220 => x"0c",
          6221 => x"08",
          6222 => x"02",
          6223 => x"81",
          6224 => x"b9",
          6225 => x"70",
          6226 => x"b9",
          6227 => x"c8",
          6228 => x"c8",
          6229 => x"b9",
          6230 => x"75",
          6231 => x"08",
          6232 => x"80",
          6233 => x"fe",
          6234 => x"27",
          6235 => x"29",
          6236 => x"b4",
          6237 => x"79",
          6238 => x"58",
          6239 => x"74",
          6240 => x"27",
          6241 => x"53",
          6242 => x"ee",
          6243 => x"df",
          6244 => x"56",
          6245 => x"08",
          6246 => x"33",
          6247 => x"56",
          6248 => x"b9",
          6249 => x"08",
          6250 => x"18",
          6251 => x"33",
          6252 => x"fe",
          6253 => x"a0",
          6254 => x"17",
          6255 => x"ca",
          6256 => x"55",
          6257 => x"9c",
          6258 => x"52",
          6259 => x"b9",
          6260 => x"80",
          6261 => x"08",
          6262 => x"c8",
          6263 => x"53",
          6264 => x"3f",
          6265 => x"9c",
          6266 => x"5a",
          6267 => x"81",
          6268 => x"81",
          6269 => x"55",
          6270 => x"84",
          6271 => x"8a",
          6272 => x"06",
          6273 => x"81",
          6274 => x"1f",
          6275 => x"57",
          6276 => x"7d",
          6277 => x"58",
          6278 => x"59",
          6279 => x"cf",
          6280 => x"34",
          6281 => x"7d",
          6282 => x"77",
          6283 => x"5b",
          6284 => x"55",
          6285 => x"59",
          6286 => x"57",
          6287 => x"33",
          6288 => x"16",
          6289 => x"0b",
          6290 => x"83",
          6291 => x"80",
          6292 => x"7a",
          6293 => x"74",
          6294 => x"81",
          6295 => x"92",
          6296 => x"84",
          6297 => x"56",
          6298 => x"84",
          6299 => x"0b",
          6300 => x"17",
          6301 => x"18",
          6302 => x"18",
          6303 => x"80",
          6304 => x"16",
          6305 => x"34",
          6306 => x"b9",
          6307 => x"0c",
          6308 => x"55",
          6309 => x"2a",
          6310 => x"fd",
          6311 => x"cc",
          6312 => x"80",
          6313 => x"80",
          6314 => x"fe",
          6315 => x"94",
          6316 => x"95",
          6317 => x"16",
          6318 => x"34",
          6319 => x"b9",
          6320 => x"3d",
          6321 => x"59",
          6322 => x"79",
          6323 => x"26",
          6324 => x"38",
          6325 => x"af",
          6326 => x"05",
          6327 => x"3f",
          6328 => x"c8",
          6329 => x"b9",
          6330 => x"a6",
          6331 => x"3d",
          6332 => x"84",
          6333 => x"08",
          6334 => x"81",
          6335 => x"38",
          6336 => x"58",
          6337 => x"33",
          6338 => x"15",
          6339 => x"b0",
          6340 => x"81",
          6341 => x"59",
          6342 => x"b3",
          6343 => x"d5",
          6344 => x"b9",
          6345 => x"3d",
          6346 => x"84",
          6347 => x"76",
          6348 => x"57",
          6349 => x"82",
          6350 => x"5d",
          6351 => x"80",
          6352 => x"72",
          6353 => x"81",
          6354 => x"5b",
          6355 => x"77",
          6356 => x"81",
          6357 => x"58",
          6358 => x"70",
          6359 => x"70",
          6360 => x"09",
          6361 => x"38",
          6362 => x"07",
          6363 => x"7a",
          6364 => x"1e",
          6365 => x"38",
          6366 => x"39",
          6367 => x"7f",
          6368 => x"05",
          6369 => x"3f",
          6370 => x"c8",
          6371 => x"6c",
          6372 => x"fe",
          6373 => x"3f",
          6374 => x"c8",
          6375 => x"0b",
          6376 => x"05",
          6377 => x"57",
          6378 => x"ff",
          6379 => x"cb",
          6380 => x"33",
          6381 => x"7e",
          6382 => x"8b",
          6383 => x"1e",
          6384 => x"81",
          6385 => x"c5",
          6386 => x"bd",
          6387 => x"33",
          6388 => x"58",
          6389 => x"38",
          6390 => x"5e",
          6391 => x"8a",
          6392 => x"08",
          6393 => x"b5",
          6394 => x"08",
          6395 => x"5f",
          6396 => x"53",
          6397 => x"fe",
          6398 => x"80",
          6399 => x"77",
          6400 => x"d8",
          6401 => x"81",
          6402 => x"81",
          6403 => x"ff",
          6404 => x"34",
          6405 => x"18",
          6406 => x"09",
          6407 => x"5e",
          6408 => x"2a",
          6409 => x"57",
          6410 => x"aa",
          6411 => x"56",
          6412 => x"78",
          6413 => x"c8",
          6414 => x"f5",
          6415 => x"57",
          6416 => x"b4",
          6417 => x"7e",
          6418 => x"38",
          6419 => x"81",
          6420 => x"84",
          6421 => x"ff",
          6422 => x"77",
          6423 => x"5a",
          6424 => x"34",
          6425 => x"80",
          6426 => x"84",
          6427 => x"08",
          6428 => x"74",
          6429 => x"74",
          6430 => x"9d",
          6431 => x"c8",
          6432 => x"84",
          6433 => x"95",
          6434 => x"2b",
          6435 => x"56",
          6436 => x"08",
          6437 => x"c8",
          6438 => x"84",
          6439 => x"81",
          6440 => x"81",
          6441 => x"81",
          6442 => x"09",
          6443 => x"c8",
          6444 => x"a8",
          6445 => x"59",
          6446 => x"a0",
          6447 => x"2e",
          6448 => x"54",
          6449 => x"53",
          6450 => x"e1",
          6451 => x"81",
          6452 => x"70",
          6453 => x"e1",
          6454 => x"08",
          6455 => x"83",
          6456 => x"08",
          6457 => x"74",
          6458 => x"82",
          6459 => x"81",
          6460 => x"17",
          6461 => x"52",
          6462 => x"3f",
          6463 => x"0d",
          6464 => x"05",
          6465 => x"53",
          6466 => x"51",
          6467 => x"08",
          6468 => x"8a",
          6469 => x"3d",
          6470 => x"3d",
          6471 => x"84",
          6472 => x"08",
          6473 => x"81",
          6474 => x"38",
          6475 => x"12",
          6476 => x"51",
          6477 => x"78",
          6478 => x"51",
          6479 => x"08",
          6480 => x"04",
          6481 => x"96",
          6482 => x"ff",
          6483 => x"55",
          6484 => x"38",
          6485 => x"0d",
          6486 => x"d0",
          6487 => x"b9",
          6488 => x"e0",
          6489 => x"a0",
          6490 => x"60",
          6491 => x"90",
          6492 => x"17",
          6493 => x"17",
          6494 => x"17",
          6495 => x"17",
          6496 => x"34",
          6497 => x"b9",
          6498 => x"3d",
          6499 => x"5d",
          6500 => x"52",
          6501 => x"84",
          6502 => x"30",
          6503 => x"25",
          6504 => x"38",
          6505 => x"81",
          6506 => x"80",
          6507 => x"8c",
          6508 => x"78",
          6509 => x"11",
          6510 => x"08",
          6511 => x"33",
          6512 => x"81",
          6513 => x"53",
          6514 => x"fe",
          6515 => x"80",
          6516 => x"76",
          6517 => x"38",
          6518 => x"56",
          6519 => x"56",
          6520 => x"75",
          6521 => x"12",
          6522 => x"07",
          6523 => x"2b",
          6524 => x"5d",
          6525 => x"c8",
          6526 => x"80",
          6527 => x"55",
          6528 => x"08",
          6529 => x"81",
          6530 => x"06",
          6531 => x"57",
          6532 => x"08",
          6533 => x"33",
          6534 => x"59",
          6535 => x"81",
          6536 => x"08",
          6537 => x"17",
          6538 => x"55",
          6539 => x"38",
          6540 => x"09",
          6541 => x"b4",
          6542 => x"7a",
          6543 => x"e2",
          6544 => x"b8",
          6545 => x"da",
          6546 => x"2e",
          6547 => x"52",
          6548 => x"b9",
          6549 => x"fe",
          6550 => x"b9",
          6551 => x"18",
          6552 => x"75",
          6553 => x"78",
          6554 => x"58",
          6555 => x"f2",
          6556 => x"5c",
          6557 => x"fc",
          6558 => x"e1",
          6559 => x"b4",
          6560 => x"eb",
          6561 => x"b9",
          6562 => x"5d",
          6563 => x"81",
          6564 => x"f4",
          6565 => x"70",
          6566 => x"9f",
          6567 => x"90",
          6568 => x"81",
          6569 => x"75",
          6570 => x"81",
          6571 => x"83",
          6572 => x"9f",
          6573 => x"ff",
          6574 => x"e0",
          6575 => x"d8",
          6576 => x"58",
          6577 => x"56",
          6578 => x"70",
          6579 => x"58",
          6580 => x"2e",
          6581 => x"ff",
          6582 => x"ff",
          6583 => x"26",
          6584 => x"8f",
          6585 => x"70",
          6586 => x"76",
          6587 => x"1a",
          6588 => x"ff",
          6589 => x"26",
          6590 => x"86",
          6591 => x"79",
          6592 => x"56",
          6593 => x"a0",
          6594 => x"1a",
          6595 => x"47",
          6596 => x"fe",
          6597 => x"55",
          6598 => x"38",
          6599 => x"a1",
          6600 => x"51",
          6601 => x"83",
          6602 => x"38",
          6603 => x"a1",
          6604 => x"56",
          6605 => x"fe",
          6606 => x"55",
          6607 => x"79",
          6608 => x"7e",
          6609 => x"58",
          6610 => x"ff",
          6611 => x"81",
          6612 => x"d9",
          6613 => x"74",
          6614 => x"fe",
          6615 => x"84",
          6616 => x"06",
          6617 => x"2e",
          6618 => x"76",
          6619 => x"b9",
          6620 => x"75",
          6621 => x"84",
          6622 => x"98",
          6623 => x"08",
          6624 => x"55",
          6625 => x"d7",
          6626 => x"52",
          6627 => x"3f",
          6628 => x"38",
          6629 => x"0c",
          6630 => x"17",
          6631 => x"81",
          6632 => x"70",
          6633 => x"80",
          6634 => x"79",
          6635 => x"51",
          6636 => x"08",
          6637 => x"ff",
          6638 => x"fd",
          6639 => x"38",
          6640 => x"81",
          6641 => x"f4",
          6642 => x"34",
          6643 => x"70",
          6644 => x"05",
          6645 => x"2e",
          6646 => x"58",
          6647 => x"ff",
          6648 => x"39",
          6649 => x"81",
          6650 => x"d7",
          6651 => x"fd",
          6652 => x"81",
          6653 => x"81",
          6654 => x"84",
          6655 => x"06",
          6656 => x"83",
          6657 => x"08",
          6658 => x"8a",
          6659 => x"2e",
          6660 => x"fd",
          6661 => x"51",
          6662 => x"08",
          6663 => x"fd",
          6664 => x"58",
          6665 => x"fe",
          6666 => x"a0",
          6667 => x"18",
          6668 => x"a9",
          6669 => x"88",
          6670 => x"57",
          6671 => x"76",
          6672 => x"74",
          6673 => x"86",
          6674 => x"78",
          6675 => x"73",
          6676 => x"33",
          6677 => x"2e",
          6678 => x"9c",
          6679 => x"81",
          6680 => x"8c",
          6681 => x"2b",
          6682 => x"fd",
          6683 => x"70",
          6684 => x"b9",
          6685 => x"42",
          6686 => x"88",
          6687 => x"38",
          6688 => x"59",
          6689 => x"3f",
          6690 => x"08",
          6691 => x"b9",
          6692 => x"84",
          6693 => x"38",
          6694 => x"81",
          6695 => x"74",
          6696 => x"87",
          6697 => x"0c",
          6698 => x"b9",
          6699 => x"15",
          6700 => x"b9",
          6701 => x"ad",
          6702 => x"a7",
          6703 => x"7a",
          6704 => x"38",
          6705 => x"e6",
          6706 => x"fe",
          6707 => x"56",
          6708 => x"77",
          6709 => x"74",
          6710 => x"55",
          6711 => x"88",
          6712 => x"17",
          6713 => x"18",
          6714 => x"16",
          6715 => x"e9",
          6716 => x"84",
          6717 => x"16",
          6718 => x"54",
          6719 => x"fe",
          6720 => x"81",
          6721 => x"ff",
          6722 => x"3d",
          6723 => x"02",
          6724 => x"42",
          6725 => x"5f",
          6726 => x"38",
          6727 => x"9f",
          6728 => x"9b",
          6729 => x"85",
          6730 => x"80",
          6731 => x"10",
          6732 => x"5a",
          6733 => x"34",
          6734 => x"84",
          6735 => x"81",
          6736 => x"84",
          6737 => x"81",
          6738 => x"ab",
          6739 => x"8a",
          6740 => x"fc",
          6741 => x"d0",
          6742 => x"98",
          6743 => x"90",
          6744 => x"88",
          6745 => x"83",
          6746 => x"84",
          6747 => x"81",
          6748 => x"1f",
          6749 => x"7e",
          6750 => x"70",
          6751 => x"60",
          6752 => x"70",
          6753 => x"57",
          6754 => x"84",
          6755 => x"52",
          6756 => x"57",
          6757 => x"60",
          6758 => x"05",
          6759 => x"8e",
          6760 => x"81",
          6761 => x"61",
          6762 => x"62",
          6763 => x"18",
          6764 => x"90",
          6765 => x"33",
          6766 => x"71",
          6767 => x"82",
          6768 => x"2b",
          6769 => x"88",
          6770 => x"3d",
          6771 => x"0c",
          6772 => x"5a",
          6773 => x"79",
          6774 => x"81",
          6775 => x"2a",
          6776 => x"2e",
          6777 => x"64",
          6778 => x"47",
          6779 => x"30",
          6780 => x"2e",
          6781 => x"8c",
          6782 => x"22",
          6783 => x"74",
          6784 => x"56",
          6785 => x"57",
          6786 => x"75",
          6787 => x"fd",
          6788 => x"10",
          6789 => x"9f",
          6790 => x"b9",
          6791 => x"05",
          6792 => x"4c",
          6793 => x"81",
          6794 => x"68",
          6795 => x"06",
          6796 => x"83",
          6797 => x"77",
          6798 => x"57",
          6799 => x"7c",
          6800 => x"31",
          6801 => x"b9",
          6802 => x"f6",
          6803 => x"82",
          6804 => x"b9",
          6805 => x"89",
          6806 => x"c0",
          6807 => x"a3",
          6808 => x"0c",
          6809 => x"04",
          6810 => x"84",
          6811 => x"b9",
          6812 => x"70",
          6813 => x"89",
          6814 => x"ff",
          6815 => x"2e",
          6816 => x"b8",
          6817 => x"7a",
          6818 => x"81",
          6819 => x"59",
          6820 => x"17",
          6821 => x"9f",
          6822 => x"e0",
          6823 => x"76",
          6824 => x"78",
          6825 => x"ff",
          6826 => x"70",
          6827 => x"4a",
          6828 => x"81",
          6829 => x"25",
          6830 => x"39",
          6831 => x"79",
          6832 => x"84",
          6833 => x"83",
          6834 => x"40",
          6835 => x"55",
          6836 => x"38",
          6837 => x"81",
          6838 => x"ff",
          6839 => x"56",
          6840 => x"93",
          6841 => x"82",
          6842 => x"8b",
          6843 => x"26",
          6844 => x"5b",
          6845 => x"8e",
          6846 => x"3d",
          6847 => x"55",
          6848 => x"f5",
          6849 => x"5b",
          6850 => x"80",
          6851 => x"05",
          6852 => x"38",
          6853 => x"55",
          6854 => x"70",
          6855 => x"74",
          6856 => x"65",
          6857 => x"61",
          6858 => x"06",
          6859 => x"88",
          6860 => x"81",
          6861 => x"70",
          6862 => x"34",
          6863 => x"61",
          6864 => x"ff",
          6865 => x"ff",
          6866 => x"34",
          6867 => x"05",
          6868 => x"61",
          6869 => x"34",
          6870 => x"9b",
          6871 => x"7e",
          6872 => x"34",
          6873 => x"05",
          6874 => x"0c",
          6875 => x"34",
          6876 => x"61",
          6877 => x"34",
          6878 => x"61",
          6879 => x"06",
          6880 => x"88",
          6881 => x"ff",
          6882 => x"a6",
          6883 => x"e5",
          6884 => x"05",
          6885 => x"34",
          6886 => x"83",
          6887 => x"60",
          6888 => x"34",
          6889 => x"51",
          6890 => x"b9",
          6891 => x"5c",
          6892 => x"61",
          6893 => x"58",
          6894 => x"63",
          6895 => x"c0",
          6896 => x"81",
          6897 => x"34",
          6898 => x"64",
          6899 => x"2a",
          6900 => x"34",
          6901 => x"7c",
          6902 => x"38",
          6903 => x"52",
          6904 => x"b9",
          6905 => x"61",
          6906 => x"58",
          6907 => x"78",
          6908 => x"c9",
          6909 => x"2e",
          6910 => x"2e",
          6911 => x"66",
          6912 => x"7a",
          6913 => x"d2",
          6914 => x"38",
          6915 => x"75",
          6916 => x"93",
          6917 => x"26",
          6918 => x"83",
          6919 => x"61",
          6920 => x"b3",
          6921 => x"75",
          6922 => x"59",
          6923 => x"ff",
          6924 => x"47",
          6925 => x"34",
          6926 => x"83",
          6927 => x"6c",
          6928 => x"51",
          6929 => x"05",
          6930 => x"bf",
          6931 => x"84",
          6932 => x"7e",
          6933 => x"83",
          6934 => x"05",
          6935 => x"c9",
          6936 => x"34",
          6937 => x"cb",
          6938 => x"61",
          6939 => x"5f",
          6940 => x"54",
          6941 => x"c2",
          6942 => x"08",
          6943 => x"79",
          6944 => x"84",
          6945 => x"b9",
          6946 => x"3d",
          6947 => x"55",
          6948 => x"45",
          6949 => x"78",
          6950 => x"fc",
          6951 => x"38",
          6952 => x"fc",
          6953 => x"57",
          6954 => x"76",
          6955 => x"51",
          6956 => x"08",
          6957 => x"2a",
          6958 => x"b9",
          6959 => x"47",
          6960 => x"cb",
          6961 => x"b9",
          6962 => x"e6",
          6963 => x"2a",
          6964 => x"f8",
          6965 => x"80",
          6966 => x"ab",
          6967 => x"88",
          6968 => x"75",
          6969 => x"34",
          6970 => x"05",
          6971 => x"c3",
          6972 => x"34",
          6973 => x"cc",
          6974 => x"a4",
          6975 => x"61",
          6976 => x"78",
          6977 => x"56",
          6978 => x"ac",
          6979 => x"80",
          6980 => x"05",
          6981 => x"61",
          6982 => x"34",
          6983 => x"61",
          6984 => x"c2",
          6985 => x"83",
          6986 => x"81",
          6987 => x"58",
          6988 => x"f9",
          6989 => x"33",
          6990 => x"15",
          6991 => x"81",
          6992 => x"fe",
          6993 => x"c8",
          6994 => x"61",
          6995 => x"34",
          6996 => x"60",
          6997 => x"fc",
          6998 => x"0c",
          6999 => x"04",
          7000 => x"70",
          7001 => x"81",
          7002 => x"61",
          7003 => x"34",
          7004 => x"87",
          7005 => x"ff",
          7006 => x"05",
          7007 => x"b1",
          7008 => x"52",
          7009 => x"80",
          7010 => x"05",
          7011 => x"38",
          7012 => x"05",
          7013 => x"70",
          7014 => x"70",
          7015 => x"34",
          7016 => x"80",
          7017 => x"c1",
          7018 => x"61",
          7019 => x"5b",
          7020 => x"88",
          7021 => x"34",
          7022 => x"ea",
          7023 => x"61",
          7024 => x"ec",
          7025 => x"34",
          7026 => x"61",
          7027 => x"34",
          7028 => x"1f",
          7029 => x"b2",
          7030 => x"52",
          7031 => x"61",
          7032 => x"0d",
          7033 => x"ff",
          7034 => x"b8",
          7035 => x"05",
          7036 => x"ff",
          7037 => x"81",
          7038 => x"74",
          7039 => x"81",
          7040 => x"8a",
          7041 => x"38",
          7042 => x"38",
          7043 => x"8e",
          7044 => x"02",
          7045 => x"77",
          7046 => x"08",
          7047 => x"17",
          7048 => x"77",
          7049 => x"24",
          7050 => x"19",
          7051 => x"8b",
          7052 => x"17",
          7053 => x"3f",
          7054 => x"07",
          7055 => x"81",
          7056 => x"d3",
          7057 => x"3f",
          7058 => x"80",
          7059 => x"80",
          7060 => x"81",
          7061 => x"f4",
          7062 => x"8a",
          7063 => x"76",
          7064 => x"8c",
          7065 => x"16",
          7066 => x"84",
          7067 => x"7c",
          7068 => x"3d",
          7069 => x"05",
          7070 => x"3f",
          7071 => x"7a",
          7072 => x"c8",
          7073 => x"ff",
          7074 => x"52",
          7075 => x"74",
          7076 => x"9f",
          7077 => x"ff",
          7078 => x"eb",
          7079 => x"c8",
          7080 => x"0d",
          7081 => x"52",
          7082 => x"90",
          7083 => x"71",
          7084 => x"04",
          7085 => x"83",
          7086 => x"73",
          7087 => x"22",
          7088 => x"12",
          7089 => x"71",
          7090 => x"83",
          7091 => x"e1",
          7092 => x"06",
          7093 => x"0d",
          7094 => x"22",
          7095 => x"51",
          7096 => x"38",
          7097 => x"84",
          7098 => x"09",
          7099 => x"26",
          7100 => x"05",
          7101 => x"84",
          7102 => x"51",
          7103 => x"38",
          7104 => x"8c",
          7105 => x"d9",
          7106 => x"75",
          7107 => x"26",
          7108 => x"38",
          7109 => x"71",
          7110 => x"70",
          7111 => x"38",
          7112 => x"70",
          7113 => x"70",
          7114 => x"55",
          7115 => x"51",
          7116 => x"0d",
          7117 => x"39",
          7118 => x"10",
          7119 => x"04",
          7120 => x"06",
          7121 => x"b0",
          7122 => x"51",
          7123 => x"ff",
          7124 => x"70",
          7125 => x"39",
          7126 => x"57",
          7127 => x"ff",
          7128 => x"16",
          7129 => x"ff",
          7130 => x"76",
          7131 => x"58",
          7132 => x"31",
          7133 => x"fe",
          7134 => x"ff",
          7135 => x"ff",
          7136 => x"8b",
          7137 => x"75",
          7138 => x"5f",
          7139 => x"49",
          7140 => x"33",
          7141 => x"1d",
          7142 => x"07",
          7143 => x"f1",
          7144 => x"db",
          7145 => x"c5",
          7146 => x"bf",
          7147 => x"59",
          7148 => x"59",
          7149 => x"59",
          7150 => x"59",
          7151 => x"59",
          7152 => x"59",
          7153 => x"59",
          7154 => x"59",
          7155 => x"59",
          7156 => x"59",
          7157 => x"59",
          7158 => x"59",
          7159 => x"59",
          7160 => x"59",
          7161 => x"59",
          7162 => x"59",
          7163 => x"59",
          7164 => x"59",
          7165 => x"59",
          7166 => x"59",
          7167 => x"59",
          7168 => x"59",
          7169 => x"59",
          7170 => x"59",
          7171 => x"59",
          7172 => x"59",
          7173 => x"59",
          7174 => x"59",
          7175 => x"59",
          7176 => x"07",
          7177 => x"59",
          7178 => x"a8",
          7179 => x"2c",
          7180 => x"59",
          7181 => x"59",
          7182 => x"59",
          7183 => x"59",
          7184 => x"59",
          7185 => x"59",
          7186 => x"59",
          7187 => x"59",
          7188 => x"59",
          7189 => x"59",
          7190 => x"59",
          7191 => x"59",
          7192 => x"59",
          7193 => x"59",
          7194 => x"59",
          7195 => x"59",
          7196 => x"59",
          7197 => x"59",
          7198 => x"59",
          7199 => x"59",
          7200 => x"59",
          7201 => x"59",
          7202 => x"59",
          7203 => x"59",
          7204 => x"59",
          7205 => x"59",
          7206 => x"ab",
          7207 => x"59",
          7208 => x"59",
          7209 => x"59",
          7210 => x"59",
          7211 => x"63",
          7212 => x"59",
          7213 => x"59",
          7214 => x"47",
          7215 => x"22",
          7216 => x"46",
          7217 => x"5e",
          7218 => x"97",
          7219 => x"01",
          7220 => x"21",
          7221 => x"9b",
          7222 => x"cb",
          7223 => x"12",
          7224 => x"de",
          7225 => x"0b",
          7226 => x"de",
          7227 => x"12",
          7228 => x"74",
          7229 => x"7c",
          7230 => x"ba",
          7231 => x"3c",
          7232 => x"55",
          7233 => x"62",
          7234 => x"62",
          7235 => x"62",
          7236 => x"3b",
          7237 => x"62",
          7238 => x"62",
          7239 => x"62",
          7240 => x"62",
          7241 => x"62",
          7242 => x"62",
          7243 => x"62",
          7244 => x"62",
          7245 => x"62",
          7246 => x"62",
          7247 => x"62",
          7248 => x"68",
          7249 => x"42",
          7250 => x"30",
          7251 => x"85",
          7252 => x"85",
          7253 => x"8a",
          7254 => x"94",
          7255 => x"e9",
          7256 => x"c8",
          7257 => x"6c",
          7258 => x"77",
          7259 => x"a0",
          7260 => x"5c",
          7261 => x"02",
          7262 => x"dc",
          7263 => x"89",
          7264 => x"89",
          7265 => x"89",
          7266 => x"a5",
          7267 => x"6a",
          7268 => x"89",
          7269 => x"89",
          7270 => x"89",
          7271 => x"89",
          7272 => x"89",
          7273 => x"89",
          7274 => x"89",
          7275 => x"89",
          7276 => x"89",
          7277 => x"27",
          7278 => x"89",
          7279 => x"ca",
          7280 => x"7b",
          7281 => x"89",
          7282 => x"89",
          7283 => x"89",
          7284 => x"ac",
          7285 => x"21",
          7286 => x"21",
          7287 => x"21",
          7288 => x"21",
          7289 => x"21",
          7290 => x"21",
          7291 => x"21",
          7292 => x"21",
          7293 => x"21",
          7294 => x"21",
          7295 => x"21",
          7296 => x"21",
          7297 => x"21",
          7298 => x"21",
          7299 => x"be",
          7300 => x"f3",
          7301 => x"ce",
          7302 => x"7e",
          7303 => x"21",
          7304 => x"4e",
          7305 => x"2a",
          7306 => x"89",
          7307 => x"67",
          7308 => x"21",
          7309 => x"7b",
          7310 => x"d7",
          7311 => x"d7",
          7312 => x"d7",
          7313 => x"d7",
          7314 => x"d7",
          7315 => x"d7",
          7316 => x"f9",
          7317 => x"d7",
          7318 => x"d7",
          7319 => x"d7",
          7320 => x"d7",
          7321 => x"50",
          7322 => x"67",
          7323 => x"39",
          7324 => x"d2",
          7325 => x"bb",
          7326 => x"a5",
          7327 => x"8e",
          7328 => x"01",
          7329 => x"fd",
          7330 => x"fd",
          7331 => x"fd",
          7332 => x"fd",
          7333 => x"fd",
          7334 => x"fd",
          7335 => x"0d",
          7336 => x"fd",
          7337 => x"fd",
          7338 => x"fd",
          7339 => x"fd",
          7340 => x"fd",
          7341 => x"fd",
          7342 => x"fd",
          7343 => x"fd",
          7344 => x"fd",
          7345 => x"fd",
          7346 => x"fd",
          7347 => x"fd",
          7348 => x"fd",
          7349 => x"fd",
          7350 => x"fd",
          7351 => x"fd",
          7352 => x"fd",
          7353 => x"fd",
          7354 => x"fd",
          7355 => x"fd",
          7356 => x"17",
          7357 => x"fd",
          7358 => x"fd",
          7359 => x"fd",
          7360 => x"fd",
          7361 => x"fd",
          7362 => x"e1",
          7363 => x"b8",
          7364 => x"fd",
          7365 => x"fd",
          7366 => x"ff",
          7367 => x"fd",
          7368 => x"0f",
          7369 => x"fd",
          7370 => x"fd",
          7371 => x"fd",
          7372 => x"17",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"00",
          7383 => x"00",
          7384 => x"00",
          7385 => x"6c",
          7386 => x"00",
          7387 => x"00",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"00",
          7392 => x"00",
          7393 => x"00",
          7394 => x"00",
          7395 => x"6e",
          7396 => x"6f",
          7397 => x"61",
          7398 => x"69",
          7399 => x"74",
          7400 => x"20",
          7401 => x"65",
          7402 => x"2e",
          7403 => x"75",
          7404 => x"74",
          7405 => x"2e",
          7406 => x"65",
          7407 => x"6b",
          7408 => x"65",
          7409 => x"65",
          7410 => x"63",
          7411 => x"64",
          7412 => x"6d",
          7413 => x"74",
          7414 => x"63",
          7415 => x"6c",
          7416 => x"79",
          7417 => x"75",
          7418 => x"69",
          7419 => x"6b",
          7420 => x"61",
          7421 => x"00",
          7422 => x"75",
          7423 => x"20",
          7424 => x"2e",
          7425 => x"69",
          7426 => x"20",
          7427 => x"65",
          7428 => x"65",
          7429 => x"20",
          7430 => x"2e",
          7431 => x"65",
          7432 => x"79",
          7433 => x"2e",
          7434 => x"65",
          7435 => x"65",
          7436 => x"61",
          7437 => x"65",
          7438 => x"00",
          7439 => x"20",
          7440 => x"00",
          7441 => x"20",
          7442 => x"00",
          7443 => x"74",
          7444 => x"00",
          7445 => x"6c",
          7446 => x"00",
          7447 => x"72",
          7448 => x"63",
          7449 => x"00",
          7450 => x"74",
          7451 => x"74",
          7452 => x"74",
          7453 => x"0a",
          7454 => x"64",
          7455 => x"6c",
          7456 => x"00",
          7457 => x"00",
          7458 => x"00",
          7459 => x"58",
          7460 => x"20",
          7461 => x"00",
          7462 => x"25",
          7463 => x"30",
          7464 => x"00",
          7465 => x"00",
          7466 => x"65",
          7467 => x"20",
          7468 => x"2a",
          7469 => x"00",
          7470 => x"65",
          7471 => x"73",
          7472 => x"20",
          7473 => x"25",
          7474 => x"00",
          7475 => x"20",
          7476 => x"20",
          7477 => x"20",
          7478 => x"25",
          7479 => x"00",
          7480 => x"65",
          7481 => x"61",
          7482 => x"00",
          7483 => x"58",
          7484 => x"75",
          7485 => x"54",
          7486 => x"74",
          7487 => x"00",
          7488 => x"58",
          7489 => x"75",
          7490 => x"54",
          7491 => x"74",
          7492 => x"00",
          7493 => x"52",
          7494 => x"75",
          7495 => x"54",
          7496 => x"74",
          7497 => x"00",
          7498 => x"65",
          7499 => x"00",
          7500 => x"6e",
          7501 => x"00",
          7502 => x"20",
          7503 => x"72",
          7504 => x"62",
          7505 => x"6d",
          7506 => x"00",
          7507 => x"63",
          7508 => x"00",
          7509 => x"2e",
          7510 => x"6c",
          7511 => x"6e",
          7512 => x"65",
          7513 => x"64",
          7514 => x"61",
          7515 => x"20",
          7516 => x"79",
          7517 => x"00",
          7518 => x"00",
          7519 => x"20",
          7520 => x"2e",
          7521 => x"00",
          7522 => x"5c",
          7523 => x"73",
          7524 => x"64",
          7525 => x"69",
          7526 => x"00",
          7527 => x"69",
          7528 => x"69",
          7529 => x"2e",
          7530 => x"6c",
          7531 => x"65",
          7532 => x"78",
          7533 => x"00",
          7534 => x"74",
          7535 => x"6f",
          7536 => x"2e",
          7537 => x"63",
          7538 => x"6f",
          7539 => x"38",
          7540 => x"00",
          7541 => x"30",
          7542 => x"00",
          7543 => x"30",
          7544 => x"70",
          7545 => x"2e",
          7546 => x"6c",
          7547 => x"2d",
          7548 => x"25",
          7549 => x"00",
          7550 => x"2e",
          7551 => x"6c",
          7552 => x"00",
          7553 => x"67",
          7554 => x"00",
          7555 => x"6d",
          7556 => x"6d",
          7557 => x"00",
          7558 => x"25",
          7559 => x"6f",
          7560 => x"75",
          7561 => x"61",
          7562 => x"6f",
          7563 => x"6d",
          7564 => x"00",
          7565 => x"25",
          7566 => x"3a",
          7567 => x"64",
          7568 => x"20",
          7569 => x"72",
          7570 => x"00",
          7571 => x"65",
          7572 => x"6d",
          7573 => x"00",
          7574 => x"65",
          7575 => x"20",
          7576 => x"65",
          7577 => x"72",
          7578 => x"73",
          7579 => x"0a",
          7580 => x"20",
          7581 => x"6f",
          7582 => x"74",
          7583 => x"73",
          7584 => x"0a",
          7585 => x"20",
          7586 => x"74",
          7587 => x"72",
          7588 => x"20",
          7589 => x"0a",
          7590 => x"63",
          7591 => x"20",
          7592 => x"20",
          7593 => x"20",
          7594 => x"20",
          7595 => x"0a",
          7596 => x"20",
          7597 => x"43",
          7598 => x"65",
          7599 => x"20",
          7600 => x"30",
          7601 => x"00",
          7602 => x"68",
          7603 => x"52",
          7604 => x"6b",
          7605 => x"25",
          7606 => x"48",
          7607 => x"20",
          7608 => x"6c",
          7609 => x"71",
          7610 => x"20",
          7611 => x"30",
          7612 => x"00",
          7613 => x"00",
          7614 => x"00",
          7615 => x"54",
          7616 => x"20",
          7617 => x"00",
          7618 => x"48",
          7619 => x"53",
          7620 => x"20",
          7621 => x"52",
          7622 => x"6e",
          7623 => x"64",
          7624 => x"20",
          7625 => x"20",
          7626 => x"72",
          7627 => x"64",
          7628 => x"20",
          7629 => x"20",
          7630 => x"63",
          7631 => x"64",
          7632 => x"20",
          7633 => x"20",
          7634 => x"3a",
          7635 => x"00",
          7636 => x"4d",
          7637 => x"25",
          7638 => x"58",
          7639 => x"20",
          7640 => x"41",
          7641 => x"3a",
          7642 => x"00",
          7643 => x"41",
          7644 => x"25",
          7645 => x"58",
          7646 => x"20",
          7647 => x"4d",
          7648 => x"3a",
          7649 => x"00",
          7650 => x"53",
          7651 => x"69",
          7652 => x"6e",
          7653 => x"6d",
          7654 => x"6c",
          7655 => x"69",
          7656 => x"78",
          7657 => x"00",
          7658 => x"00",
          7659 => x"a8",
          7660 => x"03",
          7661 => x"00",
          7662 => x"a0",
          7663 => x"05",
          7664 => x"00",
          7665 => x"98",
          7666 => x"07",
          7667 => x"00",
          7668 => x"90",
          7669 => x"08",
          7670 => x"00",
          7671 => x"88",
          7672 => x"09",
          7673 => x"00",
          7674 => x"80",
          7675 => x"0d",
          7676 => x"00",
          7677 => x"78",
          7678 => x"0e",
          7679 => x"00",
          7680 => x"70",
          7681 => x"0f",
          7682 => x"00",
          7683 => x"68",
          7684 => x"11",
          7685 => x"00",
          7686 => x"60",
          7687 => x"13",
          7688 => x"00",
          7689 => x"58",
          7690 => x"15",
          7691 => x"00",
          7692 => x"00",
          7693 => x"7e",
          7694 => x"00",
          7695 => x"7e",
          7696 => x"00",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"6f",
          7703 => x"61",
          7704 => x"6f",
          7705 => x"2c",
          7706 => x"69",
          7707 => x"74",
          7708 => x"74",
          7709 => x"00",
          7710 => x"25",
          7711 => x"6c",
          7712 => x"65",
          7713 => x"20",
          7714 => x"20",
          7715 => x"20",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"00",
          7721 => x"00",
          7722 => x"00",
          7723 => x"00",
          7724 => x"00",
          7725 => x"00",
          7726 => x"00",
          7727 => x"00",
          7728 => x"00",
          7729 => x"00",
          7730 => x"00",
          7731 => x"00",
          7732 => x"00",
          7733 => x"7e",
          7734 => x"7e",
          7735 => x"64",
          7736 => x"25",
          7737 => x"3a",
          7738 => x"00",
          7739 => x"2d",
          7740 => x"64",
          7741 => x"00",
          7742 => x"64",
          7743 => x"78",
          7744 => x"25",
          7745 => x"00",
          7746 => x"43",
          7747 => x"00",
          7748 => x"20",
          7749 => x"00",
          7750 => x"20",
          7751 => x"00",
          7752 => x"20",
          7753 => x"74",
          7754 => x"69",
          7755 => x"00",
          7756 => x"3c",
          7757 => x"00",
          7758 => x"00",
          7759 => x"33",
          7760 => x"4d",
          7761 => x"00",
          7762 => x"20",
          7763 => x"20",
          7764 => x"4e",
          7765 => x"46",
          7766 => x"00",
          7767 => x"00",
          7768 => x"00",
          7769 => x"12",
          7770 => x"00",
          7771 => x"80",
          7772 => x"8f",
          7773 => x"55",
          7774 => x"9f",
          7775 => x"a7",
          7776 => x"af",
          7777 => x"b7",
          7778 => x"bf",
          7779 => x"c7",
          7780 => x"cf",
          7781 => x"d7",
          7782 => x"df",
          7783 => x"e7",
          7784 => x"ef",
          7785 => x"f7",
          7786 => x"ff",
          7787 => x"2f",
          7788 => x"7c",
          7789 => x"04",
          7790 => x"00",
          7791 => x"02",
          7792 => x"20",
          7793 => x"fc",
          7794 => x"e0",
          7795 => x"eb",
          7796 => x"ec",
          7797 => x"e6",
          7798 => x"f2",
          7799 => x"d6",
          7800 => x"a5",
          7801 => x"ed",
          7802 => x"d1",
          7803 => x"10",
          7804 => x"a1",
          7805 => x"92",
          7806 => x"61",
          7807 => x"63",
          7808 => x"5c",
          7809 => x"34",
          7810 => x"3c",
          7811 => x"54",
          7812 => x"50",
          7813 => x"64",
          7814 => x"52",
          7815 => x"18",
          7816 => x"8c",
          7817 => x"df",
          7818 => x"c3",
          7819 => x"98",
          7820 => x"c6",
          7821 => x"b1",
          7822 => x"21",
          7823 => x"19",
          7824 => x"b2",
          7825 => x"1a",
          7826 => x"07",
          7827 => x"00",
          7828 => x"39",
          7829 => x"79",
          7830 => x"43",
          7831 => x"84",
          7832 => x"87",
          7833 => x"8b",
          7834 => x"90",
          7835 => x"94",
          7836 => x"98",
          7837 => x"9c",
          7838 => x"a0",
          7839 => x"a4",
          7840 => x"a7",
          7841 => x"ac",
          7842 => x"af",
          7843 => x"b3",
          7844 => x"b8",
          7845 => x"bc",
          7846 => x"c0",
          7847 => x"c4",
          7848 => x"c8",
          7849 => x"ca",
          7850 => x"01",
          7851 => x"f3",
          7852 => x"f4",
          7853 => x"12",
          7854 => x"3b",
          7855 => x"3f",
          7856 => x"46",
          7857 => x"81",
          7858 => x"8a",
          7859 => x"90",
          7860 => x"5f",
          7861 => x"94",
          7862 => x"67",
          7863 => x"62",
          7864 => x"9c",
          7865 => x"73",
          7866 => x"77",
          7867 => x"7b",
          7868 => x"7f",
          7869 => x"a9",
          7870 => x"87",
          7871 => x"b2",
          7872 => x"8f",
          7873 => x"7b",
          7874 => x"ff",
          7875 => x"88",
          7876 => x"11",
          7877 => x"a3",
          7878 => x"03",
          7879 => x"d8",
          7880 => x"f9",
          7881 => x"f6",
          7882 => x"fa",
          7883 => x"50",
          7884 => x"8a",
          7885 => x"cf",
          7886 => x"44",
          7887 => x"00",
          7888 => x"00",
          7889 => x"00",
          7890 => x"20",
          7891 => x"40",
          7892 => x"59",
          7893 => x"5d",
          7894 => x"08",
          7895 => x"bb",
          7896 => x"cb",
          7897 => x"f9",
          7898 => x"fb",
          7899 => x"08",
          7900 => x"04",
          7901 => x"bc",
          7902 => x"d0",
          7903 => x"e5",
          7904 => x"01",
          7905 => x"32",
          7906 => x"01",
          7907 => x"30",
          7908 => x"67",
          7909 => x"80",
          7910 => x"41",
          7911 => x"00",
          7912 => x"00",
          7913 => x"00",
          7914 => x"00",
          7915 => x"00",
          7916 => x"00",
          7917 => x"00",
          7918 => x"00",
          7919 => x"00",
          7920 => x"00",
          7921 => x"00",
          7922 => x"00",
          7923 => x"00",
          7924 => x"00",
          7925 => x"00",
          7926 => x"00",
          7927 => x"00",
          7928 => x"00",
          7929 => x"00",
          7930 => x"00",
          7931 => x"00",
          7932 => x"00",
          7933 => x"00",
          7934 => x"00",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"00",
          7963 => x"00",
          7964 => x"00",
          7965 => x"00",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"01",
          7978 => x"01",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"00",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"dc",
          7992 => x"e4",
          7993 => x"ec",
          7994 => x"80",
          7995 => x"0d",
          7996 => x"f0",
          7997 => x"78",
          7998 => x"70",
          7999 => x"68",
          8000 => x"38",
          8001 => x"2e",
          8002 => x"2f",
          8003 => x"f0",
          8004 => x"f0",
          8005 => x"0d",
          8006 => x"f0",
          8007 => x"58",
          8008 => x"50",
          8009 => x"48",
          8010 => x"38",
          8011 => x"2e",
          8012 => x"2f",
          8013 => x"f0",
          8014 => x"f0",
          8015 => x"0d",
          8016 => x"f0",
          8017 => x"58",
          8018 => x"50",
          8019 => x"48",
          8020 => x"28",
          8021 => x"3e",
          8022 => x"2f",
          8023 => x"f0",
          8024 => x"f0",
          8025 => x"f0",
          8026 => x"f0",
          8027 => x"18",
          8028 => x"10",
          8029 => x"08",
          8030 => x"f0",
          8031 => x"f0",
          8032 => x"1c",
          8033 => x"f0",
          8034 => x"f0",
          8035 => x"cd",
          8036 => x"f0",
          8037 => x"dd",
          8038 => x"b1",
          8039 => x"73",
          8040 => x"a2",
          8041 => x"b9",
          8042 => x"be",
          8043 => x"f0",
          8044 => x"f0",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"f3",
          9081 => x"fb",
          9082 => x"c3",
          9083 => x"e6",
          9084 => x"63",
          9085 => x"6a",
          9086 => x"23",
          9087 => x"2c",
          9088 => x"03",
          9089 => x"0b",
          9090 => x"13",
          9091 => x"52",
          9092 => x"83",
          9093 => x"8b",
          9094 => x"93",
          9095 => x"bc",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"03",
          9112 => x"00",
        others => X"00"
    );

    shared variable RAM5 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"88",
             5 => x"88",
             6 => x"00",
             7 => x"00",
             8 => x"06",
             9 => x"2a",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"05",
            14 => x"ff",
            15 => x"04",
            16 => x"73",
            17 => x"73",
            18 => x"04",
            19 => x"00",
            20 => x"07",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"81",
            25 => x"0a",
            26 => x"81",
            27 => x"00",
            28 => x"07",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"51",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"05",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"06",
            49 => x"ff",
            50 => x"00",
            51 => x"00",
            52 => x"73",
            53 => x"83",
            54 => x"0c",
            55 => x"00",
            56 => x"09",
            57 => x"06",
            58 => x"00",
            59 => x"00",
            60 => x"09",
            61 => x"81",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"53",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"09",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"06",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"83",
            81 => x"05",
            82 => x"04",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"0c",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"0c",
            91 => x"00",
            92 => x"06",
            93 => x"71",
            94 => x"05",
            95 => x"00",
            96 => x"06",
            97 => x"54",
            98 => x"ff",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"05",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"53",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"0b",
           134 => x"a6",
           135 => x"0b",
           136 => x"0b",
           137 => x"e6",
           138 => x"0b",
           139 => x"0b",
           140 => x"a6",
           141 => x"0b",
           142 => x"0b",
           143 => x"e8",
           144 => x"0b",
           145 => x"0b",
           146 => x"ac",
           147 => x"0b",
           148 => x"0b",
           149 => x"f0",
           150 => x"0b",
           151 => x"0b",
           152 => x"b4",
           153 => x"0b",
           154 => x"0b",
           155 => x"f8",
           156 => x"0b",
           157 => x"0b",
           158 => x"bc",
           159 => x"0b",
           160 => x"0b",
           161 => x"80",
           162 => x"0b",
           163 => x"0b",
           164 => x"c4",
           165 => x"0b",
           166 => x"0b",
           167 => x"88",
           168 => x"0b",
           169 => x"0b",
           170 => x"cb",
           171 => x"0b",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"b9",
           193 => x"b9",
           194 => x"84",
           195 => x"b9",
           196 => x"84",
           197 => x"b9",
           198 => x"84",
           199 => x"b9",
           200 => x"84",
           201 => x"b9",
           202 => x"84",
           203 => x"b9",
           204 => x"84",
           205 => x"b9",
           206 => x"84",
           207 => x"b9",
           208 => x"84",
           209 => x"b9",
           210 => x"84",
           211 => x"b9",
           212 => x"84",
           213 => x"b9",
           214 => x"84",
           215 => x"b9",
           216 => x"84",
           217 => x"84",
           218 => x"04",
           219 => x"2d",
           220 => x"90",
           221 => x"a8",
           222 => x"80",
           223 => x"d3",
           224 => x"c0",
           225 => x"82",
           226 => x"80",
           227 => x"0c",
           228 => x"08",
           229 => x"d4",
           230 => x"d4",
           231 => x"b9",
           232 => x"b9",
           233 => x"84",
           234 => x"84",
           235 => x"04",
           236 => x"2d",
           237 => x"90",
           238 => x"87",
           239 => x"80",
           240 => x"f1",
           241 => x"c0",
           242 => x"82",
           243 => x"80",
           244 => x"0c",
           245 => x"08",
           246 => x"d4",
           247 => x"d4",
           248 => x"b9",
           249 => x"b9",
           250 => x"84",
           251 => x"84",
           252 => x"04",
           253 => x"2d",
           254 => x"90",
           255 => x"fd",
           256 => x"80",
           257 => x"95",
           258 => x"c0",
           259 => x"82",
           260 => x"80",
           261 => x"0c",
           262 => x"08",
           263 => x"d4",
           264 => x"d4",
           265 => x"b9",
           266 => x"b9",
           267 => x"84",
           268 => x"84",
           269 => x"04",
           270 => x"2d",
           271 => x"90",
           272 => x"e9",
           273 => x"80",
           274 => x"c6",
           275 => x"c0",
           276 => x"83",
           277 => x"80",
           278 => x"0c",
           279 => x"08",
           280 => x"d4",
           281 => x"d4",
           282 => x"b9",
           283 => x"b9",
           284 => x"84",
           285 => x"84",
           286 => x"04",
           287 => x"2d",
           288 => x"90",
           289 => x"aa",
           290 => x"80",
           291 => x"d1",
           292 => x"c0",
           293 => x"80",
           294 => x"80",
           295 => x"0c",
           296 => x"80",
           297 => x"0c",
           298 => x"08",
           299 => x"d4",
           300 => x"d4",
           301 => x"b9",
           302 => x"b9",
           303 => x"84",
           304 => x"84",
           305 => x"04",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"81",
           311 => x"05",
           312 => x"72",
           313 => x"72",
           314 => x"72",
           315 => x"10",
           316 => x"53",
           317 => x"d5",
           318 => x"84",
           319 => x"ec",
           320 => x"04",
           321 => x"70",
           322 => x"52",
           323 => x"3f",
           324 => x"78",
           325 => x"81",
           326 => x"55",
           327 => x"81",
           328 => x"74",
           329 => x"9f",
           330 => x"74",
           331 => x"38",
           332 => x"c8",
           333 => x"2e",
           334 => x"70",
           335 => x"8a",
           336 => x"2a",
           337 => x"cb",
           338 => x"84",
           339 => x"80",
           340 => x"0d",
           341 => x"02",
           342 => x"fe",
           343 => x"7e",
           344 => x"3f",
           345 => x"3d",
           346 => x"88",
           347 => x"3f",
           348 => x"61",
           349 => x"8c",
           350 => x"2a",
           351 => x"ff",
           352 => x"80",
           353 => x"2e",
           354 => x"06",
           355 => x"38",
           356 => x"a3",
           357 => x"80",
           358 => x"72",
           359 => x"70",
           360 => x"80",
           361 => x"5b",
           362 => x"8c",
           363 => x"0c",
           364 => x"54",
           365 => x"70",
           366 => x"81",
           367 => x"98",
           368 => x"79",
           369 => x"53",
           370 => x"58",
           371 => x"39",
           372 => x"38",
           373 => x"7c",
           374 => x"ff",
           375 => x"af",
           376 => x"38",
           377 => x"81",
           378 => x"70",
           379 => x"e0",
           380 => x"38",
           381 => x"54",
           382 => x"59",
           383 => x"52",
           384 => x"33",
           385 => x"c7",
           386 => x"88",
           387 => x"7d",
           388 => x"54",
           389 => x"51",
           390 => x"81",
           391 => x"df",
           392 => x"38",
           393 => x"74",
           394 => x"52",
           395 => x"c8",
           396 => x"38",
           397 => x"7b",
           398 => x"8f",
           399 => x"80",
           400 => x"7a",
           401 => x"73",
           402 => x"80",
           403 => x"90",
           404 => x"29",
           405 => x"2c",
           406 => x"54",
           407 => x"98",
           408 => x"78",
           409 => x"ff",
           410 => x"2a",
           411 => x"73",
           412 => x"31",
           413 => x"80",
           414 => x"85",
           415 => x"54",
           416 => x"81",
           417 => x"85",
           418 => x"38",
           419 => x"38",
           420 => x"80",
           421 => x"80",
           422 => x"2c",
           423 => x"38",
           424 => x"77",
           425 => x"80",
           426 => x"73",
           427 => x"53",
           428 => x"81",
           429 => x"70",
           430 => x"25",
           431 => x"ef",
           432 => x"81",
           433 => x"55",
           434 => x"87",
           435 => x"80",
           436 => x"2e",
           437 => x"81",
           438 => x"e2",
           439 => x"38",
           440 => x"5e",
           441 => x"2e",
           442 => x"06",
           443 => x"77",
           444 => x"80",
           445 => x"80",
           446 => x"a0",
           447 => x"90",
           448 => x"58",
           449 => x"39",
           450 => x"57",
           451 => x"7e",
           452 => x"55",
           453 => x"05",
           454 => x"33",
           455 => x"80",
           456 => x"90",
           457 => x"5f",
           458 => x"55",
           459 => x"80",
           460 => x"90",
           461 => x"fe",
           462 => x"f7",
           463 => x"ff",
           464 => x"ff",
           465 => x"70",
           466 => x"3f",
           467 => x"ff",
           468 => x"2e",
           469 => x"81",
           470 => x"e2",
           471 => x"0a",
           472 => x"80",
           473 => x"56",
           474 => x"06",
           475 => x"fe",
           476 => x"08",
           477 => x"24",
           478 => x"06",
           479 => x"39",
           480 => x"76",
           481 => x"88",
           482 => x"76",
           483 => x"60",
           484 => x"56",
           485 => x"75",
           486 => x"08",
           487 => x"90",
           488 => x"fe",
           489 => x"33",
           490 => x"ff",
           491 => x"77",
           492 => x"81",
           493 => x"84",
           494 => x"78",
           495 => x"39",
           496 => x"5b",
           497 => x"77",
           498 => x"80",
           499 => x"80",
           500 => x"a0",
           501 => x"52",
           502 => x"2e",
           503 => x"52",
           504 => x"2a",
           505 => x"8c",
           506 => x"78",
           507 => x"7d",
           508 => x"73",
           509 => x"52",
           510 => x"06",
           511 => x"ff",
           512 => x"51",
           513 => x"7a",
           514 => x"39",
           515 => x"2c",
           516 => x"ab",
           517 => x"52",
           518 => x"39",
           519 => x"84",
           520 => x"78",
           521 => x"f3",
           522 => x"83",
           523 => x"99",
           524 => x"08",
           525 => x"3f",
           526 => x"78",
           527 => x"85",
           528 => x"70",
           529 => x"ff",
           530 => x"80",
           531 => x"33",
           532 => x"d5",
           533 => x"08",
           534 => x"80",
           535 => x"81",
           536 => x"88",
           537 => x"39",
           538 => x"ac",
           539 => x"55",
           540 => x"2e",
           541 => x"84",
           542 => x"fa",
           543 => x"0b",
           544 => x"32",
           545 => x"ff",
           546 => x"92",
           547 => x"53",
           548 => x"38",
           549 => x"88",
           550 => x"55",
           551 => x"74",
           552 => x"72",
           553 => x"e3",
           554 => x"33",
           555 => x"ff",
           556 => x"73",
           557 => x"fa",
           558 => x"70",
           559 => x"56",
           560 => x"73",
           561 => x"2e",
           562 => x"88",
           563 => x"56",
           564 => x"75",
           565 => x"8c",
           566 => x"c8",
           567 => x"76",
           568 => x"54",
           569 => x"08",
           570 => x"8c",
           571 => x"3d",
           572 => x"ff",
           573 => x"55",
           574 => x"72",
           575 => x"38",
           576 => x"80",
           577 => x"33",
           578 => x"38",
           579 => x"81",
           580 => x"06",
           581 => x"3d",
           582 => x"72",
           583 => x"05",
           584 => x"b9",
           585 => x"51",
           586 => x"b9",
           587 => x"80",
           588 => x"70",
           589 => x"08",
           590 => x"53",
           591 => x"84",
           592 => x"74",
           593 => x"ff",
           594 => x"77",
           595 => x"05",
           596 => x"12",
           597 => x"51",
           598 => x"70",
           599 => x"85",
           600 => x"79",
           601 => x"80",
           602 => x"38",
           603 => x"81",
           604 => x"55",
           605 => x"73",
           606 => x"04",
           607 => x"38",
           608 => x"ff",
           609 => x"ff",
           610 => x"ff",
           611 => x"73",
           612 => x"c7",
           613 => x"53",
           614 => x"70",
           615 => x"84",
           616 => x"04",
           617 => x"54",
           618 => x"51",
           619 => x"70",
           620 => x"85",
           621 => x"78",
           622 => x"80",
           623 => x"53",
           624 => x"ff",
           625 => x"b9",
           626 => x"3d",
           627 => x"72",
           628 => x"70",
           629 => x"71",
           630 => x"14",
           631 => x"13",
           632 => x"84",
           633 => x"72",
           634 => x"ff",
           635 => x"15",
           636 => x"de",
           637 => x"0c",
           638 => x"c8",
           639 => x"0d",
           640 => x"c1",
           641 => x"c8",
           642 => x"ea",
           643 => x"b9",
           644 => x"b9",
           645 => x"74",
           646 => x"51",
           647 => x"54",
           648 => x"0d",
           649 => x"71",
           650 => x"9f",
           651 => x"51",
           652 => x"52",
           653 => x"38",
           654 => x"70",
           655 => x"04",
           656 => x"55",
           657 => x"38",
           658 => x"ff",
           659 => x"b9",
           660 => x"3d",
           661 => x"76",
           662 => x"f5",
           663 => x"12",
           664 => x"51",
           665 => x"08",
           666 => x"80",
           667 => x"80",
           668 => x"a0",
           669 => x"54",
           670 => x"38",
           671 => x"10",
           672 => x"9f",
           673 => x"75",
           674 => x"52",
           675 => x"73",
           676 => x"c8",
           677 => x"0d",
           678 => x"30",
           679 => x"2b",
           680 => x"83",
           681 => x"25",
           682 => x"2a",
           683 => x"80",
           684 => x"71",
           685 => x"8c",
           686 => x"82",
           687 => x"2a",
           688 => x"82",
           689 => x"b9",
           690 => x"54",
           691 => x"56",
           692 => x"52",
           693 => x"75",
           694 => x"81",
           695 => x"29",
           696 => x"53",
           697 => x"78",
           698 => x"2e",
           699 => x"84",
           700 => x"73",
           701 => x"bd",
           702 => x"52",
           703 => x"38",
           704 => x"81",
           705 => x"76",
           706 => x"56",
           707 => x"74",
           708 => x"78",
           709 => x"81",
           710 => x"ff",
           711 => x"55",
           712 => x"c8",
           713 => x"0d",
           714 => x"9f",
           715 => x"32",
           716 => x"72",
           717 => x"56",
           718 => x"75",
           719 => x"88",
           720 => x"7d",
           721 => x"08",
           722 => x"2e",
           723 => x"70",
           724 => x"a0",
           725 => x"f5",
           726 => x"d0",
           727 => x"80",
           728 => x"74",
           729 => x"27",
           730 => x"06",
           731 => x"06",
           732 => x"f9",
           733 => x"89",
           734 => x"27",
           735 => x"81",
           736 => x"56",
           737 => x"78",
           738 => x"75",
           739 => x"c8",
           740 => x"16",
           741 => x"59",
           742 => x"ff",
           743 => x"33",
           744 => x"38",
           745 => x"38",
           746 => x"d0",
           747 => x"73",
           748 => x"c8",
           749 => x"81",
           750 => x"55",
           751 => x"84",
           752 => x"f7",
           753 => x"70",
           754 => x"56",
           755 => x"8f",
           756 => x"33",
           757 => x"73",
           758 => x"2e",
           759 => x"56",
           760 => x"58",
           761 => x"38",
           762 => x"14",
           763 => x"14",
           764 => x"73",
           765 => x"ff",
           766 => x"89",
           767 => x"77",
           768 => x"0c",
           769 => x"26",
           770 => x"38",
           771 => x"56",
           772 => x"0d",
           773 => x"70",
           774 => x"09",
           775 => x"70",
           776 => x"80",
           777 => x"80",
           778 => x"74",
           779 => x"56",
           780 => x"38",
           781 => x"0d",
           782 => x"0c",
           783 => x"ca",
           784 => x"8b",
           785 => x"84",
           786 => x"b9",
           787 => x"52",
           788 => x"10",
           789 => x"04",
           790 => x"83",
           791 => x"ef",
           792 => x"ce",
           793 => x"0d",
           794 => x"3f",
           795 => x"51",
           796 => x"83",
           797 => x"3d",
           798 => x"fc",
           799 => x"b4",
           800 => x"04",
           801 => x"83",
           802 => x"ee",
           803 => x"d0",
           804 => x"0d",
           805 => x"3f",
           806 => x"51",
           807 => x"83",
           808 => x"3d",
           809 => x"a4",
           810 => x"f8",
           811 => x"04",
           812 => x"83",
           813 => x"ee",
           814 => x"d1",
           815 => x"0d",
           816 => x"3f",
           817 => x"51",
           818 => x"ec",
           819 => x"e3",
           820 => x"30",
           821 => x"57",
           822 => x"83",
           823 => x"81",
           824 => x"80",
           825 => x"3d",
           826 => x"84",
           827 => x"08",
           828 => x"82",
           829 => x"07",
           830 => x"72",
           831 => x"2e",
           832 => x"55",
           833 => x"74",
           834 => x"8e",
           835 => x"d1",
           836 => x"51",
           837 => x"0c",
           838 => x"08",
           839 => x"c8",
           840 => x"84",
           841 => x"9d",
           842 => x"84",
           843 => x"55",
           844 => x"19",
           845 => x"e8",
           846 => x"b9",
           847 => x"3f",
           848 => x"f4",
           849 => x"de",
           850 => x"0d",
           851 => x"58",
           852 => x"7a",
           853 => x"08",
           854 => x"76",
           855 => x"c8",
           856 => x"84",
           857 => x"84",
           858 => x"78",
           859 => x"c8",
           860 => x"0d",
           861 => x"cf",
           862 => x"5f",
           863 => x"2e",
           864 => x"fc",
           865 => x"51",
           866 => x"27",
           867 => x"38",
           868 => x"18",
           869 => x"72",
           870 => x"d1",
           871 => x"53",
           872 => x"74",
           873 => x"dd",
           874 => x"80",
           875 => x"53",
           876 => x"81",
           877 => x"38",
           878 => x"ff",
           879 => x"38",
           880 => x"84",
           881 => x"df",
           882 => x"c2",
           883 => x"3f",
           884 => x"51",
           885 => x"98",
           886 => x"a0",
           887 => x"82",
           888 => x"26",
           889 => x"c8",
           890 => x"98",
           891 => x"d5",
           892 => x"87",
           893 => x"fe",
           894 => x"91",
           895 => x"53",
           896 => x"79",
           897 => x"72",
           898 => x"83",
           899 => x"14",
           900 => x"51",
           901 => x"38",
           902 => x"db",
           903 => x"08",
           904 => x"73",
           905 => x"53",
           906 => x"52",
           907 => x"84",
           908 => x"a0",
           909 => x"dd",
           910 => x"08",
           911 => x"16",
           912 => x"3f",
           913 => x"53",
           914 => x"38",
           915 => x"81",
           916 => x"db",
           917 => x"b9",
           918 => x"70",
           919 => x"70",
           920 => x"06",
           921 => x"72",
           922 => x"9b",
           923 => x"2b",
           924 => x"30",
           925 => x"07",
           926 => x"59",
           927 => x"a9",
           928 => x"b9",
           929 => x"3d",
           930 => x"aa",
           931 => x"83",
           932 => x"51",
           933 => x"81",
           934 => x"72",
           935 => x"71",
           936 => x"81",
           937 => x"72",
           938 => x"71",
           939 => x"81",
           940 => x"72",
           941 => x"71",
           942 => x"81",
           943 => x"88",
           944 => x"a9",
           945 => x"51",
           946 => x"9c",
           947 => x"a9",
           948 => x"51",
           949 => x"9c",
           950 => x"72",
           951 => x"2e",
           952 => x"de",
           953 => x"3f",
           954 => x"2a",
           955 => x"2e",
           956 => x"9b",
           957 => x"ce",
           958 => x"86",
           959 => x"80",
           960 => x"81",
           961 => x"51",
           962 => x"3f",
           963 => x"52",
           964 => x"bd",
           965 => x"d4",
           966 => x"9a",
           967 => x"06",
           968 => x"38",
           969 => x"3f",
           970 => x"80",
           971 => x"70",
           972 => x"fd",
           973 => x"9a",
           974 => x"c6",
           975 => x"82",
           976 => x"80",
           977 => x"ca",
           978 => x"61",
           979 => x"60",
           980 => x"c8",
           981 => x"59",
           982 => x"d5",
           983 => x"43",
           984 => x"7e",
           985 => x"51",
           986 => x"bc",
           987 => x"79",
           988 => x"2e",
           989 => x"5e",
           990 => x"70",
           991 => x"38",
           992 => x"81",
           993 => x"5d",
           994 => x"5c",
           995 => x"29",
           996 => x"5b",
           997 => x"84",
           998 => x"08",
           999 => x"c8",
          1000 => x"7d",
          1001 => x"70",
          1002 => x"27",
          1003 => x"80",
          1004 => x"7e",
          1005 => x"08",
          1006 => x"8d",
          1007 => x"b8",
          1008 => x"3f",
          1009 => x"5c",
          1010 => x"84",
          1011 => x"84",
          1012 => x"38",
          1013 => x"82",
          1014 => x"8c",
          1015 => x"38",
          1016 => x"52",
          1017 => x"84",
          1018 => x"67",
          1019 => x"90",
          1020 => x"3f",
          1021 => x"08",
          1022 => x"25",
          1023 => x"83",
          1024 => x"06",
          1025 => x"1b",
          1026 => x"ff",
          1027 => x"32",
          1028 => x"ff",
          1029 => x"94",
          1030 => x"d1",
          1031 => x"52",
          1032 => x"83",
          1033 => x"5b",
          1034 => x"83",
          1035 => x"82",
          1036 => x"80",
          1037 => x"ee",
          1038 => x"f8",
          1039 => x"84",
          1040 => x"84",
          1041 => x"0b",
          1042 => x"ff",
          1043 => x"81",
          1044 => x"d0",
          1045 => x"0b",
          1046 => x"d5",
          1047 => x"a7",
          1048 => x"fc",
          1049 => x"0c",
          1050 => x"26",
          1051 => x"be",
          1052 => x"53",
          1053 => x"fb",
          1054 => x"f4",
          1055 => x"c8",
          1056 => x"ae",
          1057 => x"41",
          1058 => x"de",
          1059 => x"3f",
          1060 => x"7b",
          1061 => x"83",
          1062 => x"3f",
          1063 => x"fa",
          1064 => x"39",
          1065 => x"fa",
          1066 => x"e8",
          1067 => x"3f",
          1068 => x"51",
          1069 => x"d0",
          1070 => x"ff",
          1071 => x"b9",
          1072 => x"68",
          1073 => x"3f",
          1074 => x"08",
          1075 => x"c8",
          1076 => x"e1",
          1077 => x"84",
          1078 => x"cf",
          1079 => x"f9",
          1080 => x"51",
          1081 => x"b8",
          1082 => x"05",
          1083 => x"08",
          1084 => x"fe",
          1085 => x"e9",
          1086 => x"d0",
          1087 => x"52",
          1088 => x"84",
          1089 => x"7e",
          1090 => x"33",
          1091 => x"78",
          1092 => x"05",
          1093 => x"fe",
          1094 => x"e8",
          1095 => x"2e",
          1096 => x"11",
          1097 => x"3f",
          1098 => x"64",
          1099 => x"d7",
          1100 => x"a8",
          1101 => x"cf",
          1102 => x"78",
          1103 => x"26",
          1104 => x"46",
          1105 => x"11",
          1106 => x"3f",
          1107 => x"a0",
          1108 => x"ff",
          1109 => x"b9",
          1110 => x"b8",
          1111 => x"05",
          1112 => x"08",
          1113 => x"c4",
          1114 => x"59",
          1115 => x"70",
          1116 => x"7d",
          1117 => x"78",
          1118 => x"51",
          1119 => x"81",
          1120 => x"b8",
          1121 => x"05",
          1122 => x"08",
          1123 => x"fe",
          1124 => x"e8",
          1125 => x"2e",
          1126 => x"11",
          1127 => x"3f",
          1128 => x"f8",
          1129 => x"3f",
          1130 => x"38",
          1131 => x"33",
          1132 => x"39",
          1133 => x"80",
          1134 => x"c8",
          1135 => x"3d",
          1136 => x"51",
          1137 => x"b1",
          1138 => x"d7",
          1139 => x"a8",
          1140 => x"cc",
          1141 => x"78",
          1142 => x"26",
          1143 => x"d1",
          1144 => x"33",
          1145 => x"3d",
          1146 => x"51",
          1147 => x"80",
          1148 => x"80",
          1149 => x"05",
          1150 => x"ff",
          1151 => x"b9",
          1152 => x"39",
          1153 => x"80",
          1154 => x"c8",
          1155 => x"3d",
          1156 => x"51",
          1157 => x"80",
          1158 => x"f8",
          1159 => x"c7",
          1160 => x"84",
          1161 => x"51",
          1162 => x"78",
          1163 => x"79",
          1164 => x"26",
          1165 => x"f4",
          1166 => x"51",
          1167 => x"b9",
          1168 => x"f3",
          1169 => x"52",
          1170 => x"c8",
          1171 => x"b9",
          1172 => x"98",
          1173 => x"ff",
          1174 => x"b9",
          1175 => x"33",
          1176 => x"83",
          1177 => x"fc",
          1178 => x"af",
          1179 => x"83",
          1180 => x"83",
          1181 => x"b8",
          1182 => x"05",
          1183 => x"08",
          1184 => x"5c",
          1185 => x"7a",
          1186 => x"9f",
          1187 => x"80",
          1188 => x"38",
          1189 => x"c4",
          1190 => x"66",
          1191 => x"d8",
          1192 => x"39",
          1193 => x"05",
          1194 => x"ff",
          1195 => x"b9",
          1196 => x"64",
          1197 => x"45",
          1198 => x"80",
          1199 => x"c8",
          1200 => x"5e",
          1201 => x"82",
          1202 => x"fe",
          1203 => x"e1",
          1204 => x"2e",
          1205 => x"ce",
          1206 => x"23",
          1207 => x"53",
          1208 => x"84",
          1209 => x"f0",
          1210 => x"ff",
          1211 => x"b9",
          1212 => x"68",
          1213 => x"34",
          1214 => x"b8",
          1215 => x"05",
          1216 => x"08",
          1217 => x"71",
          1218 => x"59",
          1219 => x"81",
          1220 => x"d6",
          1221 => x"52",
          1222 => x"39",
          1223 => x"f3",
          1224 => x"ac",
          1225 => x"f0",
          1226 => x"ab",
          1227 => x"b8",
          1228 => x"22",
          1229 => x"45",
          1230 => x"5c",
          1231 => x"f2",
          1232 => x"f2",
          1233 => x"38",
          1234 => x"39",
          1235 => x"64",
          1236 => x"51",
          1237 => x"39",
          1238 => x"2e",
          1239 => x"fc",
          1240 => x"ac",
          1241 => x"33",
          1242 => x"f2",
          1243 => x"f2",
          1244 => x"38",
          1245 => x"39",
          1246 => x"2e",
          1247 => x"fb",
          1248 => x"7c",
          1249 => x"08",
          1250 => x"33",
          1251 => x"f2",
          1252 => x"f2",
          1253 => x"9c",
          1254 => x"47",
          1255 => x"0b",
          1256 => x"8c",
          1257 => x"52",
          1258 => x"c8",
          1259 => x"87",
          1260 => x"3f",
          1261 => x"0c",
          1262 => x"57",
          1263 => x"a6",
          1264 => x"77",
          1265 => x"75",
          1266 => x"c8",
          1267 => x"0b",
          1268 => x"83",
          1269 => x"bc",
          1270 => x"02",
          1271 => x"84",
          1272 => x"13",
          1273 => x"0c",
          1274 => x"95",
          1275 => x"3f",
          1276 => x"51",
          1277 => x"22",
          1278 => x"bc",
          1279 => x"33",
          1280 => x"3f",
          1281 => x"d0",
          1282 => x"51",
          1283 => x"83",
          1284 => x"e7",
          1285 => x"70",
          1286 => x"74",
          1287 => x"70",
          1288 => x"2e",
          1289 => x"70",
          1290 => x"55",
          1291 => x"ff",
          1292 => x"38",
          1293 => x"38",
          1294 => x"53",
          1295 => x"81",
          1296 => x"80",
          1297 => x"39",
          1298 => x"70",
          1299 => x"81",
          1300 => x"80",
          1301 => x"80",
          1302 => x"05",
          1303 => x"70",
          1304 => x"04",
          1305 => x"2e",
          1306 => x"72",
          1307 => x"54",
          1308 => x"e0",
          1309 => x"53",
          1310 => x"f8",
          1311 => x"53",
          1312 => x"b9",
          1313 => x"3d",
          1314 => x"3f",
          1315 => x"38",
          1316 => x"0d",
          1317 => x"33",
          1318 => x"8b",
          1319 => x"ff",
          1320 => x"81",
          1321 => x"52",
          1322 => x"13",
          1323 => x"80",
          1324 => x"52",
          1325 => x"13",
          1326 => x"26",
          1327 => x"87",
          1328 => x"38",
          1329 => x"72",
          1330 => x"13",
          1331 => x"13",
          1332 => x"13",
          1333 => x"13",
          1334 => x"13",
          1335 => x"87",
          1336 => x"98",
          1337 => x"9c",
          1338 => x"0c",
          1339 => x"7f",
          1340 => x"7d",
          1341 => x"7d",
          1342 => x"5c",
          1343 => x"b4",
          1344 => x"c0",
          1345 => x"34",
          1346 => x"85",
          1347 => x"5c",
          1348 => x"a4",
          1349 => x"c0",
          1350 => x"23",
          1351 => x"06",
          1352 => x"86",
          1353 => x"84",
          1354 => x"82",
          1355 => x"06",
          1356 => x"a1",
          1357 => x"0d",
          1358 => x"2e",
          1359 => x"3f",
          1360 => x"98",
          1361 => x"81",
          1362 => x"38",
          1363 => x"0d",
          1364 => x"84",
          1365 => x"2c",
          1366 => x"06",
          1367 => x"3f",
          1368 => x"98",
          1369 => x"38",
          1370 => x"54",
          1371 => x"80",
          1372 => x"98",
          1373 => x"ff",
          1374 => x"14",
          1375 => x"71",
          1376 => x"04",
          1377 => x"83",
          1378 => x"53",
          1379 => x"38",
          1380 => x"2a",
          1381 => x"80",
          1382 => x"81",
          1383 => x"81",
          1384 => x"8a",
          1385 => x"71",
          1386 => x"87",
          1387 => x"86",
          1388 => x"72",
          1389 => x"3d",
          1390 => x"06",
          1391 => x"32",
          1392 => x"38",
          1393 => x"80",
          1394 => x"08",
          1395 => x"54",
          1396 => x"3d",
          1397 => x"70",
          1398 => x"f2",
          1399 => x"3d",
          1400 => x"56",
          1401 => x"38",
          1402 => x"81",
          1403 => x"2e",
          1404 => x"08",
          1405 => x"54",
          1406 => x"91",
          1407 => x"e3",
          1408 => x"72",
          1409 => x"81",
          1410 => x"ff",
          1411 => x"70",
          1412 => x"90",
          1413 => x"33",
          1414 => x"84",
          1415 => x"71",
          1416 => x"70",
          1417 => x"53",
          1418 => x"2a",
          1419 => x"b5",
          1420 => x"96",
          1421 => x"70",
          1422 => x"87",
          1423 => x"8a",
          1424 => x"ab",
          1425 => x"f2",
          1426 => x"83",
          1427 => x"08",
          1428 => x"98",
          1429 => x"9e",
          1430 => x"c0",
          1431 => x"87",
          1432 => x"0c",
          1433 => x"a0",
          1434 => x"f2",
          1435 => x"83",
          1436 => x"08",
          1437 => x"c0",
          1438 => x"9e",
          1439 => x"c0",
          1440 => x"b8",
          1441 => x"f2",
          1442 => x"83",
          1443 => x"08",
          1444 => x"f2",
          1445 => x"90",
          1446 => x"52",
          1447 => x"f2",
          1448 => x"90",
          1449 => x"52",
          1450 => x"52",
          1451 => x"87",
          1452 => x"0a",
          1453 => x"83",
          1454 => x"34",
          1455 => x"70",
          1456 => x"70",
          1457 => x"83",
          1458 => x"9e",
          1459 => x"51",
          1460 => x"81",
          1461 => x"0b",
          1462 => x"80",
          1463 => x"2e",
          1464 => x"ce",
          1465 => x"08",
          1466 => x"52",
          1467 => x"71",
          1468 => x"c0",
          1469 => x"06",
          1470 => x"38",
          1471 => x"80",
          1472 => x"81",
          1473 => x"80",
          1474 => x"f2",
          1475 => x"90",
          1476 => x"52",
          1477 => x"52",
          1478 => x"87",
          1479 => x"06",
          1480 => x"38",
          1481 => x"87",
          1482 => x"70",
          1483 => x"d4",
          1484 => x"08",
          1485 => x"70",
          1486 => x"83",
          1487 => x"08",
          1488 => x"51",
          1489 => x"87",
          1490 => x"51",
          1491 => x"81",
          1492 => x"c0",
          1493 => x"83",
          1494 => x"81",
          1495 => x"83",
          1496 => x"83",
          1497 => x"38",
          1498 => x"83",
          1499 => x"38",
          1500 => x"c6",
          1501 => x"85",
          1502 => x"74",
          1503 => x"54",
          1504 => x"33",
          1505 => x"d7",
          1506 => x"f2",
          1507 => x"83",
          1508 => x"38",
          1509 => x"a6",
          1510 => x"83",
          1511 => x"75",
          1512 => x"54",
          1513 => x"51",
          1514 => x"52",
          1515 => x"3f",
          1516 => x"e4",
          1517 => x"b4",
          1518 => x"b5",
          1519 => x"f4",
          1520 => x"da",
          1521 => x"f2",
          1522 => x"75",
          1523 => x"08",
          1524 => x"54",
          1525 => x"da",
          1526 => x"f2",
          1527 => x"f2",
          1528 => x"3d",
          1529 => x"bd",
          1530 => x"3f",
          1531 => x"29",
          1532 => x"c8",
          1533 => x"b4",
          1534 => x"f2",
          1535 => x"75",
          1536 => x"08",
          1537 => x"54",
          1538 => x"db",
          1539 => x"f2",
          1540 => x"9e",
          1541 => x"51",
          1542 => x"c0",
          1543 => x"83",
          1544 => x"83",
          1545 => x"51",
          1546 => x"08",
          1547 => x"a9",
          1548 => x"3f",
          1549 => x"bc",
          1550 => x"bc",
          1551 => x"51",
          1552 => x"bd",
          1553 => x"54",
          1554 => x"e4",
          1555 => x"cf",
          1556 => x"38",
          1557 => x"ff",
          1558 => x"54",
          1559 => x"ec",
          1560 => x"ac",
          1561 => x"80",
          1562 => x"dc",
          1563 => x"f2",
          1564 => x"d2",
          1565 => x"ff",
          1566 => x"54",
          1567 => x"39",
          1568 => x"a4",
          1569 => x"c9",
          1570 => x"38",
          1571 => x"83",
          1572 => x"83",
          1573 => x"fb",
          1574 => x"33",
          1575 => x"c9",
          1576 => x"80",
          1577 => x"f2",
          1578 => x"54",
          1579 => x"a9",
          1580 => x"80",
          1581 => x"f2",
          1582 => x"54",
          1583 => x"89",
          1584 => x"80",
          1585 => x"f2",
          1586 => x"54",
          1587 => x"e9",
          1588 => x"80",
          1589 => x"f2",
          1590 => x"54",
          1591 => x"c9",
          1592 => x"80",
          1593 => x"f2",
          1594 => x"54",
          1595 => x"a9",
          1596 => x"80",
          1597 => x"de",
          1598 => x"d9",
          1599 => x"f2",
          1600 => x"d8",
          1601 => x"8e",
          1602 => x"38",
          1603 => x"52",
          1604 => x"ff",
          1605 => x"83",
          1606 => x"83",
          1607 => x"ff",
          1608 => x"83",
          1609 => x"83",
          1610 => x"ff",
          1611 => x"83",
          1612 => x"83",
          1613 => x"04",
          1614 => x"04",
          1615 => x"84",
          1616 => x"08",
          1617 => x"57",
          1618 => x"51",
          1619 => x"08",
          1620 => x"0b",
          1621 => x"f8",
          1622 => x"84",
          1623 => x"76",
          1624 => x"08",
          1625 => x"b9",
          1626 => x"c8",
          1627 => x"80",
          1628 => x"72",
          1629 => x"76",
          1630 => x"83",
          1631 => x"51",
          1632 => x"08",
          1633 => x"77",
          1634 => x"04",
          1635 => x"3f",
          1636 => x"38",
          1637 => x"79",
          1638 => x"08",
          1639 => x"76",
          1640 => x"c1",
          1641 => x"a9",
          1642 => x"3d",
          1643 => x"72",
          1644 => x"2e",
          1645 => x"59",
          1646 => x"bc",
          1647 => x"a9",
          1648 => x"52",
          1649 => x"b9",
          1650 => x"54",
          1651 => x"82",
          1652 => x"ff",
          1653 => x"38",
          1654 => x"aa",
          1655 => x"3d",
          1656 => x"51",
          1657 => x"80",
          1658 => x"52",
          1659 => x"c8",
          1660 => x"2e",
          1661 => x"06",
          1662 => x"38",
          1663 => x"56",
          1664 => x"15",
          1665 => x"a0",
          1666 => x"75",
          1667 => x"3d",
          1668 => x"b9",
          1669 => x"52",
          1670 => x"c8",
          1671 => x"08",
          1672 => x"ce",
          1673 => x"2e",
          1674 => x"3f",
          1675 => x"84",
          1676 => x"b9",
          1677 => x"55",
          1678 => x"81",
          1679 => x"ab",
          1680 => x"06",
          1681 => x"c8",
          1682 => x"0d",
          1683 => x"3d",
          1684 => x"3d",
          1685 => x"b4",
          1686 => x"83",
          1687 => x"2e",
          1688 => x"8d",
          1689 => x"78",
          1690 => x"fd",
          1691 => x"80",
          1692 => x"08",
          1693 => x"79",
          1694 => x"06",
          1695 => x"70",
          1696 => x"98",
          1697 => x"05",
          1698 => x"70",
          1699 => x"5d",
          1700 => x"57",
          1701 => x"75",
          1702 => x"0a",
          1703 => x"2c",
          1704 => x"38",
          1705 => x"57",
          1706 => x"42",
          1707 => x"de",
          1708 => x"41",
          1709 => x"80",
          1710 => x"34",
          1711 => x"38",
          1712 => x"2c",
          1713 => x"70",
          1714 => x"82",
          1715 => x"53",
          1716 => x"78",
          1717 => x"84",
          1718 => x"ff",
          1719 => x"81",
          1720 => x"81",
          1721 => x"26",
          1722 => x"82",
          1723 => x"d4",
          1724 => x"ce",
          1725 => x"70",
          1726 => x"bc",
          1727 => x"fe",
          1728 => x"fe",
          1729 => x"fd",
          1730 => x"38",
          1731 => x"d1",
          1732 => x"0c",
          1733 => x"38",
          1734 => x"57",
          1735 => x"08",
          1736 => x"34",
          1737 => x"39",
          1738 => x"2e",
          1739 => x"52",
          1740 => x"d1",
          1741 => x"d1",
          1742 => x"8c",
          1743 => x"88",
          1744 => x"fc",
          1745 => x"81",
          1746 => x"7b",
          1747 => x"cf",
          1748 => x"8b",
          1749 => x"e4",
          1750 => x"83",
          1751 => x"7c",
          1752 => x"8c",
          1753 => x"38",
          1754 => x"ff",
          1755 => x"52",
          1756 => x"d5",
          1757 => x"ff",
          1758 => x"5b",
          1759 => x"ff",
          1760 => x"ff",
          1761 => x"34",
          1762 => x"f3",
          1763 => x"7c",
          1764 => x"11",
          1765 => x"74",
          1766 => x"38",
          1767 => x"b9",
          1768 => x"b9",
          1769 => x"53",
          1770 => x"3f",
          1771 => x"33",
          1772 => x"38",
          1773 => x"ff",
          1774 => x"52",
          1775 => x"d5",
          1776 => x"e7",
          1777 => x"55",
          1778 => x"ff",
          1779 => x"33",
          1780 => x"33",
          1781 => x"af",
          1782 => x"15",
          1783 => x"16",
          1784 => x"3f",
          1785 => x"06",
          1786 => x"75",
          1787 => x"ac",
          1788 => x"d1",
          1789 => x"55",
          1790 => x"33",
          1791 => x"33",
          1792 => x"a9",
          1793 => x"33",
          1794 => x"76",
          1795 => x"7a",
          1796 => x"70",
          1797 => x"57",
          1798 => x"84",
          1799 => x"b2",
          1800 => x"98",
          1801 => x"33",
          1802 => x"f9",
          1803 => x"88",
          1804 => x"80",
          1805 => x"98",
          1806 => x"5a",
          1807 => x"d5",
          1808 => x"e7",
          1809 => x"80",
          1810 => x"88",
          1811 => x"ff",
          1812 => x"58",
          1813 => x"ac",
          1814 => x"b7",
          1815 => x"80",
          1816 => x"88",
          1817 => x"fe",
          1818 => x"33",
          1819 => x"77",
          1820 => x"81",
          1821 => x"70",
          1822 => x"57",
          1823 => x"fe",
          1824 => x"74",
          1825 => x"ac",
          1826 => x"3f",
          1827 => x"76",
          1828 => x"06",
          1829 => x"7c",
          1830 => x"ac",
          1831 => x"3f",
          1832 => x"8b",
          1833 => x"06",
          1834 => x"88",
          1835 => x"38",
          1836 => x"83",
          1837 => x"56",
          1838 => x"87",
          1839 => x"18",
          1840 => x"3f",
          1841 => x"f3",
          1842 => x"e0",
          1843 => x"8b",
          1844 => x"75",
          1845 => x"33",
          1846 => x"80",
          1847 => x"84",
          1848 => x"0c",
          1849 => x"33",
          1850 => x"d5",
          1851 => x"8f",
          1852 => x"51",
          1853 => x"08",
          1854 => x"84",
          1855 => x"84",
          1856 => x"55",
          1857 => x"ff",
          1858 => x"8c",
          1859 => x"f5",
          1860 => x"81",
          1861 => x"74",
          1862 => x"08",
          1863 => x"84",
          1864 => x"ae",
          1865 => x"88",
          1866 => x"8c",
          1867 => x"8c",
          1868 => x"cc",
          1869 => x"99",
          1870 => x"80",
          1871 => x"b9",
          1872 => x"d1",
          1873 => x"56",
          1874 => x"d1",
          1875 => x"d1",
          1876 => x"d1",
          1877 => x"88",
          1878 => x"8c",
          1879 => x"84",
          1880 => x"76",
          1881 => x"ac",
          1882 => x"3f",
          1883 => x"70",
          1884 => x"57",
          1885 => x"38",
          1886 => x"ff",
          1887 => x"29",
          1888 => x"84",
          1889 => x"79",
          1890 => x"08",
          1891 => x"74",
          1892 => x"05",
          1893 => x"5b",
          1894 => x"38",
          1895 => x"17",
          1896 => x"52",
          1897 => x"75",
          1898 => x"05",
          1899 => x"43",
          1900 => x"38",
          1901 => x"34",
          1902 => x"51",
          1903 => x"0a",
          1904 => x"2c",
          1905 => x"60",
          1906 => x"39",
          1907 => x"06",
          1908 => x"38",
          1909 => x"27",
          1910 => x"2c",
          1911 => x"7b",
          1912 => x"75",
          1913 => x"05",
          1914 => x"52",
          1915 => x"81",
          1916 => x"77",
          1917 => x"3d",
          1918 => x"57",
          1919 => x"56",
          1920 => x"84",
          1921 => x"29",
          1922 => x"79",
          1923 => x"60",
          1924 => x"2b",
          1925 => x"5c",
          1926 => x"38",
          1927 => x"ff",
          1928 => x"29",
          1929 => x"84",
          1930 => x"75",
          1931 => x"08",
          1932 => x"75",
          1933 => x"05",
          1934 => x"57",
          1935 => x"38",
          1936 => x"56",
          1937 => x"51",
          1938 => x"08",
          1939 => x"08",
          1940 => x"52",
          1941 => x"d1",
          1942 => x"56",
          1943 => x"d5",
          1944 => x"a7",
          1945 => x"51",
          1946 => x"08",
          1947 => x"84",
          1948 => x"84",
          1949 => x"55",
          1950 => x"3f",
          1951 => x"0c",
          1952 => x"76",
          1953 => x"38",
          1954 => x"52",
          1955 => x"a8",
          1956 => x"81",
          1957 => x"d1",
          1958 => x"24",
          1959 => x"98",
          1960 => x"06",
          1961 => x"ef",
          1962 => x"b4",
          1963 => x"f2",
          1964 => x"74",
          1965 => x"56",
          1966 => x"83",
          1967 => x"55",
          1968 => x"51",
          1969 => x"08",
          1970 => x"83",
          1971 => x"5f",
          1972 => x"d9",
          1973 => x"84",
          1974 => x"ac",
          1975 => x"aa",
          1976 => x"d1",
          1977 => x"ff",
          1978 => x"51",
          1979 => x"d1",
          1980 => x"57",
          1981 => x"84",
          1982 => x"a6",
          1983 => x"a0",
          1984 => x"ac",
          1985 => x"3f",
          1986 => x"79",
          1987 => x"06",
          1988 => x"0b",
          1989 => x"d1",
          1990 => x"b4",
          1991 => x"e9",
          1992 => x"88",
          1993 => x"06",
          1994 => x"ff",
          1995 => x"ff",
          1996 => x"8c",
          1997 => x"2e",
          1998 => x"52",
          1999 => x"d5",
          2000 => x"e7",
          2001 => x"51",
          2002 => x"33",
          2003 => x"34",
          2004 => x"75",
          2005 => x"c8",
          2006 => x"c8",
          2007 => x"75",
          2008 => x"ff",
          2009 => x"88",
          2010 => x"5e",
          2011 => x"84",
          2012 => x"a5",
          2013 => x"a0",
          2014 => x"ac",
          2015 => x"3f",
          2016 => x"60",
          2017 => x"06",
          2018 => x"fa",
          2019 => x"2b",
          2020 => x"81",
          2021 => x"dc",
          2022 => x"0c",
          2023 => x"83",
          2024 => x"41",
          2025 => x"53",
          2026 => x"3f",
          2027 => x"81",
          2028 => x"82",
          2029 => x"f4",
          2030 => x"54",
          2031 => x"d8",
          2032 => x"8a",
          2033 => x"b4",
          2034 => x"0b",
          2035 => x"d1",
          2036 => x"b4",
          2037 => x"84",
          2038 => x"3f",
          2039 => x"84",
          2040 => x"83",
          2041 => x"7a",
          2042 => x"c8",
          2043 => x"2e",
          2044 => x"b9",
          2045 => x"84",
          2046 => x"b9",
          2047 => x"b9",
          2048 => x"56",
          2049 => x"83",
          2050 => x"f2",
          2051 => x"59",
          2052 => x"87",
          2053 => x"1a",
          2054 => x"3f",
          2055 => x"f3",
          2056 => x"e0",
          2057 => x"a0",
          2058 => x"5e",
          2059 => x"5d",
          2060 => x"df",
          2061 => x"39",
          2062 => x"a5",
          2063 => x"05",
          2064 => x"7a",
          2065 => x"f3",
          2066 => x"80",
          2067 => x"70",
          2068 => x"e0",
          2069 => x"57",
          2070 => x"08",
          2071 => x"10",
          2072 => x"57",
          2073 => x"38",
          2074 => x"34",
          2075 => x"34",
          2076 => x"ff",
          2077 => x"f8",
          2078 => x"c3",
          2079 => x"05",
          2080 => x"8d",
          2081 => x"81",
          2082 => x"2e",
          2083 => x"59",
          2084 => x"80",
          2085 => x"90",
          2086 => x"83",
          2087 => x"23",
          2088 => x"71",
          2089 => x"71",
          2090 => x"78",
          2091 => x"84",
          2092 => x"05",
          2093 => x"75",
          2094 => x"33",
          2095 => x"55",
          2096 => x"34",
          2097 => x"ff",
          2098 => x"0d",
          2099 => x"f8",
          2100 => x"f8",
          2101 => x"05",
          2102 => x"b0",
          2103 => x"81",
          2104 => x"81",
          2105 => x"83",
          2106 => x"59",
          2107 => x"73",
          2108 => x"29",
          2109 => x"ff",
          2110 => x"ff",
          2111 => x"75",
          2112 => x"5c",
          2113 => x"f8",
          2114 => x"29",
          2115 => x"7b",
          2116 => x"55",
          2117 => x"80",
          2118 => x"f8",
          2119 => x"34",
          2120 => x"86",
          2121 => x"33",
          2122 => x"33",
          2123 => x"22",
          2124 => x"5e",
          2125 => x"df",
          2126 => x"ff",
          2127 => x"54",
          2128 => x"0b",
          2129 => x"f8",
          2130 => x"98",
          2131 => x"2b",
          2132 => x"56",
          2133 => x"fd",
          2134 => x"f8",
          2135 => x"10",
          2136 => x"90",
          2137 => x"5e",
          2138 => x"b0",
          2139 => x"70",
          2140 => x"70",
          2141 => x"70",
          2142 => x"60",
          2143 => x"40",
          2144 => x"72",
          2145 => x"57",
          2146 => x"ff",
          2147 => x"ff",
          2148 => x"29",
          2149 => x"78",
          2150 => x"79",
          2151 => x"58",
          2152 => x"5c",
          2153 => x"74",
          2154 => x"39",
          2155 => x"53",
          2156 => x"85",
          2157 => x"80",
          2158 => x"b0",
          2159 => x"80",
          2160 => x"80",
          2161 => x"34",
          2162 => x"51",
          2163 => x"70",
          2164 => x"a0",
          2165 => x"54",
          2166 => x"80",
          2167 => x"72",
          2168 => x"70",
          2169 => x"86",
          2170 => x"f7",
          2171 => x"80",
          2172 => x"0b",
          2173 => x"04",
          2174 => x"0c",
          2175 => x"33",
          2176 => x"b7",
          2177 => x"75",
          2178 => x"bc",
          2179 => x"f8",
          2180 => x"a0",
          2181 => x"51",
          2182 => x"83",
          2183 => x"53",
          2184 => x"c4",
          2185 => x"55",
          2186 => x"f8",
          2187 => x"7a",
          2188 => x"7a",
          2189 => x"72",
          2190 => x"22",
          2191 => x"ba",
          2192 => x"82",
          2193 => x"71",
          2194 => x"9f",
          2195 => x"14",
          2196 => x"e0",
          2197 => x"33",
          2198 => x"14",
          2199 => x"38",
          2200 => x"f8",
          2201 => x"55",
          2202 => x"73",
          2203 => x"54",
          2204 => x"b7",
          2205 => x"f8",
          2206 => x"06",
          2207 => x"73",
          2208 => x"31",
          2209 => x"71",
          2210 => x"a7",
          2211 => x"79",
          2212 => x"71",
          2213 => x"75",
          2214 => x"16",
          2215 => x"b7",
          2216 => x"5a",
          2217 => x"77",
          2218 => x"84",
          2219 => x"71",
          2220 => x"72",
          2221 => x"84",
          2222 => x"74",
          2223 => x"22",
          2224 => x"ba",
          2225 => x"fd",
          2226 => x"38",
          2227 => x"f8",
          2228 => x"09",
          2229 => x"31",
          2230 => x"71",
          2231 => x"59",
          2232 => x"83",
          2233 => x"74",
          2234 => x"e0",
          2235 => x"05",
          2236 => x"2e",
          2237 => x"16",
          2238 => x"34",
          2239 => x"f4",
          2240 => x"55",
          2241 => x"15",
          2242 => x"74",
          2243 => x"a9",
          2244 => x"05",
          2245 => x"26",
          2246 => x"ec",
          2247 => x"bc",
          2248 => x"71",
          2249 => x"b9",
          2250 => x"0b",
          2251 => x"33",
          2252 => x"80",
          2253 => x"83",
          2254 => x"c8",
          2255 => x"f8",
          2256 => x"9f",
          2257 => x"70",
          2258 => x"f8",
          2259 => x"33",
          2260 => x"25",
          2261 => x"f8",
          2262 => x"86",
          2263 => x"70",
          2264 => x"72",
          2265 => x"f8",
          2266 => x"0c",
          2267 => x"33",
          2268 => x"11",
          2269 => x"38",
          2270 => x"80",
          2271 => x"0d",
          2272 => x"83",
          2273 => x"ff",
          2274 => x"b4",
          2275 => x"f8",
          2276 => x"02",
          2277 => x"b3",
          2278 => x"05",
          2279 => x"33",
          2280 => x"80",
          2281 => x"51",
          2282 => x"09",
          2283 => x"83",
          2284 => x"c8",
          2285 => x"f4",
          2286 => x"70",
          2287 => x"b9",
          2288 => x"f8",
          2289 => x"83",
          2290 => x"f4",
          2291 => x"70",
          2292 => x"f1",
          2293 => x"84",
          2294 => x"83",
          2295 => x"07",
          2296 => x"b4",
          2297 => x"51",
          2298 => x"39",
          2299 => x"85",
          2300 => x"ff",
          2301 => x"fb",
          2302 => x"f4",
          2303 => x"33",
          2304 => x"83",
          2305 => x"f8",
          2306 => x"83",
          2307 => x"f8",
          2308 => x"07",
          2309 => x"cc",
          2310 => x"06",
          2311 => x"34",
          2312 => x"81",
          2313 => x"83",
          2314 => x"f8",
          2315 => x"07",
          2316 => x"94",
          2317 => x"06",
          2318 => x"34",
          2319 => x"81",
          2320 => x"34",
          2321 => x"81",
          2322 => x"f8",
          2323 => x"0d",
          2324 => x"80",
          2325 => x"83",
          2326 => x"84",
          2327 => x"5b",
          2328 => x"78",
          2329 => x"81",
          2330 => x"80",
          2331 => x"f8",
          2332 => x"7c",
          2333 => x"04",
          2334 => x"38",
          2335 => x"0b",
          2336 => x"f8",
          2337 => x"34",
          2338 => x"58",
          2339 => x"bb",
          2340 => x"7b",
          2341 => x"bc",
          2342 => x"b7",
          2343 => x"34",
          2344 => x"f8",
          2345 => x"8f",
          2346 => x"be",
          2347 => x"80",
          2348 => x"83",
          2349 => x"f6",
          2350 => x"b8",
          2351 => x"56",
          2352 => x"52",
          2353 => x"3f",
          2354 => x"5a",
          2355 => x"84",
          2356 => x"83",
          2357 => x"81",
          2358 => x"c9",
          2359 => x"dd",
          2360 => x"c1",
          2361 => x"0b",
          2362 => x"f8",
          2363 => x"83",
          2364 => x"80",
          2365 => x"84",
          2366 => x"f8",
          2367 => x"81",
          2368 => x"ac",
          2369 => x"c8",
          2370 => x"ff",
          2371 => x"51",
          2372 => x"c8",
          2373 => x"ac",
          2374 => x"fe",
          2375 => x"ff",
          2376 => x"0d",
          2377 => x"84",
          2378 => x"83",
          2379 => x"86",
          2380 => x"22",
          2381 => x"05",
          2382 => x"ce",
          2383 => x"72",
          2384 => x"2e",
          2385 => x"b9",
          2386 => x"75",
          2387 => x"bc",
          2388 => x"f9",
          2389 => x"54",
          2390 => x"a0",
          2391 => x"83",
          2392 => x"72",
          2393 => x"75",
          2394 => x"f8",
          2395 => x"83",
          2396 => x"18",
          2397 => x"ff",
          2398 => x"f9",
          2399 => x"57",
          2400 => x"98",
          2401 => x"ff",
          2402 => x"99",
          2403 => x"81",
          2404 => x"f8",
          2405 => x"72",
          2406 => x"33",
          2407 => x"80",
          2408 => x"0d",
          2409 => x"8d",
          2410 => x"09",
          2411 => x"81",
          2412 => x"f8",
          2413 => x"fa",
          2414 => x"33",
          2415 => x"06",
          2416 => x"a0",
          2417 => x"81",
          2418 => x"ff",
          2419 => x"a5",
          2420 => x"54",
          2421 => x"fa",
          2422 => x"f2",
          2423 => x"3f",
          2424 => x"3d",
          2425 => x"81",
          2426 => x"33",
          2427 => x"53",
          2428 => x"f8",
          2429 => x"d5",
          2430 => x"ff",
          2431 => x"a5",
          2432 => x"34",
          2433 => x"f9",
          2434 => x"3f",
          2435 => x"ef",
          2436 => x"0d",
          2437 => x"c4",
          2438 => x"b8",
          2439 => x"78",
          2440 => x"24",
          2441 => x"b9",
          2442 => x"84",
          2443 => x"83",
          2444 => x"58",
          2445 => x"86",
          2446 => x"bc",
          2447 => x"f6",
          2448 => x"42",
          2449 => x"83",
          2450 => x"05",
          2451 => x"86",
          2452 => x"bc",
          2453 => x"f6",
          2454 => x"29",
          2455 => x"f8",
          2456 => x"81",
          2457 => x"76",
          2458 => x"bd",
          2459 => x"19",
          2460 => x"0b",
          2461 => x"04",
          2462 => x"79",
          2463 => x"9b",
          2464 => x"cc",
          2465 => x"84",
          2466 => x"83",
          2467 => x"5e",
          2468 => x"86",
          2469 => x"bc",
          2470 => x"f6",
          2471 => x"59",
          2472 => x"83",
          2473 => x"5b",
          2474 => x"b0",
          2475 => x"70",
          2476 => x"83",
          2477 => x"44",
          2478 => x"33",
          2479 => x"1f",
          2480 => x"77",
          2481 => x"f9",
          2482 => x"9c",
          2483 => x"b7",
          2484 => x"78",
          2485 => x"38",
          2486 => x"0b",
          2487 => x"04",
          2488 => x"19",
          2489 => x"84",
          2490 => x"77",
          2491 => x"cc",
          2492 => x"80",
          2493 => x"0b",
          2494 => x"04",
          2495 => x"0b",
          2496 => x"33",
          2497 => x"33",
          2498 => x"84",
          2499 => x"80",
          2500 => x"f8",
          2501 => x"71",
          2502 => x"83",
          2503 => x"33",
          2504 => x"f8",
          2505 => x"34",
          2506 => x"06",
          2507 => x"33",
          2508 => x"58",
          2509 => x"98",
          2510 => x"89",
          2511 => x"3f",
          2512 => x"ae",
          2513 => x"f9",
          2514 => x"f8",
          2515 => x"a0",
          2516 => x"51",
          2517 => x"ff",
          2518 => x"51",
          2519 => x"a4",
          2520 => x"57",
          2521 => x"75",
          2522 => x"80",
          2523 => x"84",
          2524 => x"ca",
          2525 => x"81",
          2526 => x"84",
          2527 => x"83",
          2528 => x"83",
          2529 => x"83",
          2530 => x"80",
          2531 => x"84",
          2532 => x"78",
          2533 => x"a7",
          2534 => x"bc",
          2535 => x"f9",
          2536 => x"29",
          2537 => x"f8",
          2538 => x"05",
          2539 => x"ce",
          2540 => x"5c",
          2541 => x"81",
          2542 => x"83",
          2543 => x"34",
          2544 => x"06",
          2545 => x"05",
          2546 => x"86",
          2547 => x"bc",
          2548 => x"f6",
          2549 => x"42",
          2550 => x"34",
          2551 => x"62",
          2552 => x"86",
          2553 => x"bc",
          2554 => x"f6",
          2555 => x"29",
          2556 => x"f8",
          2557 => x"34",
          2558 => x"58",
          2559 => x"b7",
          2560 => x"ff",
          2561 => x"83",
          2562 => x"58",
          2563 => x"bb",
          2564 => x"83",
          2565 => x"38",
          2566 => x"f9",
          2567 => x"26",
          2568 => x"c5",
          2569 => x"0b",
          2570 => x"51",
          2571 => x"c8",
          2572 => x"f8",
          2573 => x"ff",
          2574 => x"ff",
          2575 => x"a0",
          2576 => x"41",
          2577 => x"ff",
          2578 => x"45",
          2579 => x"82",
          2580 => x"06",
          2581 => x"06",
          2582 => x"84",
          2583 => x"1b",
          2584 => x"f9",
          2585 => x"29",
          2586 => x"83",
          2587 => x"33",
          2588 => x"f8",
          2589 => x"34",
          2590 => x"06",
          2591 => x"33",
          2592 => x"40",
          2593 => x"9a",
          2594 => x"ff",
          2595 => x"ac",
          2596 => x"92",
          2597 => x"f8",
          2598 => x"06",
          2599 => x"38",
          2600 => x"33",
          2601 => x"06",
          2602 => x"06",
          2603 => x"5b",
          2604 => x"a7",
          2605 => x"33",
          2606 => x"22",
          2607 => x"56",
          2608 => x"83",
          2609 => x"5a",
          2610 => x"b0",
          2611 => x"70",
          2612 => x"83",
          2613 => x"5b",
          2614 => x"33",
          2615 => x"05",
          2616 => x"7f",
          2617 => x"f9",
          2618 => x"b8",
          2619 => x"0c",
          2620 => x"17",
          2621 => x"7a",
          2622 => x"ff",
          2623 => x"39",
          2624 => x"0b",
          2625 => x"04",
          2626 => x"b7",
          2627 => x"f8",
          2628 => x"f9",
          2629 => x"f4",
          2630 => x"dc",
          2631 => x"c7",
          2632 => x"fb",
          2633 => x"11",
          2634 => x"79",
          2635 => x"ca",
          2636 => x"23",
          2637 => x"33",
          2638 => x"34",
          2639 => x"33",
          2640 => x"f9",
          2641 => x"f8",
          2642 => x"72",
          2643 => x"c4",
          2644 => x"05",
          2645 => x"f9",
          2646 => x"29",
          2647 => x"f8",
          2648 => x"76",
          2649 => x"f4",
          2650 => x"34",
          2651 => x"06",
          2652 => x"33",
          2653 => x"42",
          2654 => x"9a",
          2655 => x"06",
          2656 => x"38",
          2657 => x"e2",
          2658 => x"f9",
          2659 => x"84",
          2660 => x"f3",
          2661 => x"75",
          2662 => x"ea",
          2663 => x"0c",
          2664 => x"33",
          2665 => x"33",
          2666 => x"33",
          2667 => x"b9",
          2668 => x"b0",
          2669 => x"b1",
          2670 => x"b2",
          2671 => x"33",
          2672 => x"84",
          2673 => x"09",
          2674 => x"f9",
          2675 => x"33",
          2676 => x"84",
          2677 => x"ed",
          2678 => x"3f",
          2679 => x"83",
          2680 => x"60",
          2681 => x"83",
          2682 => x"fe",
          2683 => x"33",
          2684 => x"77",
          2685 => x"84",
          2686 => x"41",
          2687 => x"10",
          2688 => x"08",
          2689 => x"80",
          2690 => x"33",
          2691 => x"70",
          2692 => x"42",
          2693 => x"34",
          2694 => x"56",
          2695 => x"b9",
          2696 => x"06",
          2697 => x"75",
          2698 => x"f8",
          2699 => x"83",
          2700 => x"70",
          2701 => x"2e",
          2702 => x"83",
          2703 => x"0b",
          2704 => x"33",
          2705 => x"57",
          2706 => x"17",
          2707 => x"f9",
          2708 => x"80",
          2709 => x"33",
          2710 => x"70",
          2711 => x"41",
          2712 => x"34",
          2713 => x"5b",
          2714 => x"b9",
          2715 => x"81",
          2716 => x"33",
          2717 => x"33",
          2718 => x"80",
          2719 => x"5a",
          2720 => x"ff",
          2721 => x"ff",
          2722 => x"7e",
          2723 => x"80",
          2724 => x"39",
          2725 => x"2e",
          2726 => x"58",
          2727 => x"d9",
          2728 => x"fb",
          2729 => x"75",
          2730 => x"9d",
          2731 => x"05",
          2732 => x"5e",
          2733 => x"57",
          2734 => x"39",
          2735 => x"2e",
          2736 => x"83",
          2737 => x"b7",
          2738 => x"75",
          2739 => x"83",
          2740 => x"e4",
          2741 => x"0b",
          2742 => x"76",
          2743 => x"b9",
          2744 => x"e3",
          2745 => x"17",
          2746 => x"33",
          2747 => x"84",
          2748 => x"2e",
          2749 => x"75",
          2750 => x"52",
          2751 => x"3f",
          2752 => x"57",
          2753 => x"b9",
          2754 => x"06",
          2755 => x"81",
          2756 => x"81",
          2757 => x"5b",
          2758 => x"38",
          2759 => x"76",
          2760 => x"77",
          2761 => x"83",
          2762 => x"ff",
          2763 => x"b4",
          2764 => x"34",
          2765 => x"5f",
          2766 => x"b9",
          2767 => x"5b",
          2768 => x"f8",
          2769 => x"81",
          2770 => x"74",
          2771 => x"83",
          2772 => x"29",
          2773 => x"f7",
          2774 => x"5d",
          2775 => x"83",
          2776 => x"57",
          2777 => x"b7",
          2778 => x"d6",
          2779 => x"f6",
          2780 => x"31",
          2781 => x"38",
          2782 => x"27",
          2783 => x"83",
          2784 => x"83",
          2785 => x"76",
          2786 => x"81",
          2787 => x"29",
          2788 => x"a0",
          2789 => x"81",
          2790 => x"71",
          2791 => x"7f",
          2792 => x"1a",
          2793 => x"b7",
          2794 => x"5d",
          2795 => x"7c",
          2796 => x"84",
          2797 => x"71",
          2798 => x"77",
          2799 => x"17",
          2800 => x"7b",
          2801 => x"81",
          2802 => x"5e",
          2803 => x"84",
          2804 => x"43",
          2805 => x"99",
          2806 => x"33",
          2807 => x"80",
          2808 => x"b1",
          2809 => x"b7",
          2810 => x"33",
          2811 => x"94",
          2812 => x"78",
          2813 => x"83",
          2814 => x"06",
          2815 => x"5c",
          2816 => x"b7",
          2817 => x"89",
          2818 => x"76",
          2819 => x"61",
          2820 => x"38",
          2821 => x"62",
          2822 => x"1f",
          2823 => x"79",
          2824 => x"ac",
          2825 => x"a4",
          2826 => x"2b",
          2827 => x"07",
          2828 => x"57",
          2829 => x"70",
          2830 => x"84",
          2831 => x"38",
          2832 => x"33",
          2833 => x"81",
          2834 => x"73",
          2835 => x"77",
          2836 => x"1b",
          2837 => x"75",
          2838 => x"f4",
          2839 => x"98",
          2840 => x"e0",
          2841 => x"5a",
          2842 => x"f4",
          2843 => x"34",
          2844 => x"81",
          2845 => x"f4",
          2846 => x"06",
          2847 => x"f4",
          2848 => x"2b",
          2849 => x"58",
          2850 => x"81",
          2851 => x"f8",
          2852 => x"06",
          2853 => x"fa",
          2854 => x"33",
          2855 => x"b7",
          2856 => x"b7",
          2857 => x"ee",
          2858 => x"56",
          2859 => x"70",
          2860 => x"39",
          2861 => x"85",
          2862 => x"e5",
          2863 => x"06",
          2864 => x"34",
          2865 => x"f9",
          2866 => x"f4",
          2867 => x"81",
          2868 => x"f8",
          2869 => x"0b",
          2870 => x"81",
          2871 => x"83",
          2872 => x"75",
          2873 => x"83",
          2874 => x"07",
          2875 => x"fd",
          2876 => x"06",
          2877 => x"f4",
          2878 => x"33",
          2879 => x"75",
          2880 => x"83",
          2881 => x"07",
          2882 => x"c5",
          2883 => x"06",
          2884 => x"34",
          2885 => x"81",
          2886 => x"f8",
          2887 => x"f4",
          2888 => x"75",
          2889 => x"83",
          2890 => x"75",
          2891 => x"83",
          2892 => x"75",
          2893 => x"83",
          2894 => x"75",
          2895 => x"83",
          2896 => x"d0",
          2897 => x"fd",
          2898 => x"bf",
          2899 => x"f4",
          2900 => x"f8",
          2901 => x"c9",
          2902 => x"33",
          2903 => x"33",
          2904 => x"33",
          2905 => x"0b",
          2906 => x"81",
          2907 => x"84",
          2908 => x"77",
          2909 => x"33",
          2910 => x"56",
          2911 => x"9c",
          2912 => x"fe",
          2913 => x"a1",
          2914 => x"c4",
          2915 => x"80",
          2916 => x"0d",
          2917 => x"e9",
          2918 => x"5c",
          2919 => x"10",
          2920 => x"05",
          2921 => x"0b",
          2922 => x"0b",
          2923 => x"51",
          2924 => x"70",
          2925 => x"e6",
          2926 => x"34",
          2927 => x"ef",
          2928 => x"3f",
          2929 => x"ff",
          2930 => x"06",
          2931 => x"52",
          2932 => x"33",
          2933 => x"75",
          2934 => x"83",
          2935 => x"70",
          2936 => x"f0",
          2937 => x"05",
          2938 => x"59",
          2939 => x"75",
          2940 => x"33",
          2941 => x"77",
          2942 => x"33",
          2943 => x"06",
          2944 => x"11",
          2945 => x"f6",
          2946 => x"70",
          2947 => x"33",
          2948 => x"81",
          2949 => x"ff",
          2950 => x"24",
          2951 => x"56",
          2952 => x"16",
          2953 => x"81",
          2954 => x"76",
          2955 => x"33",
          2956 => x"ff",
          2957 => x"7b",
          2958 => x"57",
          2959 => x"38",
          2960 => x"ff",
          2961 => x"79",
          2962 => x"a7",
          2963 => x"81",
          2964 => x"42",
          2965 => x"38",
          2966 => x"17",
          2967 => x"7b",
          2968 => x"81",
          2969 => x"5f",
          2970 => x"84",
          2971 => x"59",
          2972 => x"b1",
          2973 => x"b7",
          2974 => x"5d",
          2975 => x"7d",
          2976 => x"84",
          2977 => x"71",
          2978 => x"75",
          2979 => x"39",
          2980 => x"b7",
          2981 => x"f8",
          2982 => x"f6",
          2983 => x"5f",
          2984 => x"38",
          2985 => x"06",
          2986 => x"27",
          2987 => x"f6",
          2988 => x"58",
          2989 => x"57",
          2990 => x"bc",
          2991 => x"52",
          2992 => x"38",
          2993 => x"eb",
          2994 => x"05",
          2995 => x"40",
          2996 => x"75",
          2997 => x"09",
          2998 => x"f9",
          2999 => x"f8",
          3000 => x"ff",
          3001 => x"f6",
          3002 => x"f8",
          3003 => x"56",
          3004 => x"39",
          3005 => x"f8",
          3006 => x"56",
          3007 => x"76",
          3008 => x"f4",
          3009 => x"75",
          3010 => x"70",
          3011 => x"33",
          3012 => x"76",
          3013 => x"7b",
          3014 => x"f1",
          3015 => x"34",
          3016 => x"23",
          3017 => x"f6",
          3018 => x"f8",
          3019 => x"fa",
          3020 => x"33",
          3021 => x"34",
          3022 => x"97",
          3023 => x"54",
          3024 => x"db",
          3025 => x"0c",
          3026 => x"51",
          3027 => x"c8",
          3028 => x"0d",
          3029 => x"83",
          3030 => x"83",
          3031 => x"59",
          3032 => x"14",
          3033 => x"59",
          3034 => x"0d",
          3035 => x"53",
          3036 => x"32",
          3037 => x"9f",
          3038 => x"f7",
          3039 => x"81",
          3040 => x"54",
          3041 => x"25",
          3042 => x"2e",
          3043 => x"83",
          3044 => x"72",
          3045 => x"05",
          3046 => x"71",
          3047 => x"06",
          3048 => x"58",
          3049 => x"f0",
          3050 => x"80",
          3051 => x"c0",
          3052 => x"f6",
          3053 => x"76",
          3054 => x"70",
          3055 => x"74",
          3056 => x"e8",
          3057 => x"f6",
          3058 => x"76",
          3059 => x"2e",
          3060 => x"15",
          3061 => x"81",
          3062 => x"f7",
          3063 => x"33",
          3064 => x"70",
          3065 => x"27",
          3066 => x"70",
          3067 => x"54",
          3068 => x"ff",
          3069 => x"81",
          3070 => x"85",
          3071 => x"34",
          3072 => x"2e",
          3073 => x"a2",
          3074 => x"83",
          3075 => x"70",
          3076 => x"33",
          3077 => x"83",
          3078 => x"ff",
          3079 => x"33",
          3080 => x"83",
          3081 => x"ff",
          3082 => x"33",
          3083 => x"ff",
          3084 => x"38",
          3085 => x"81",
          3086 => x"06",
          3087 => x"38",
          3088 => x"74",
          3089 => x"08",
          3090 => x"08",
          3091 => x"38",
          3092 => x"83",
          3093 => x"81",
          3094 => x"fe",
          3095 => x"77",
          3096 => x"53",
          3097 => x"10",
          3098 => x"08",
          3099 => x"80",
          3100 => x"c0",
          3101 => x"27",
          3102 => x"ce",
          3103 => x"38",
          3104 => x"87",
          3105 => x"0c",
          3106 => x"2e",
          3107 => x"54",
          3108 => x"81",
          3109 => x"a8",
          3110 => x"38",
          3111 => x"c3",
          3112 => x"39",
          3113 => x"56",
          3114 => x"38",
          3115 => x"b4",
          3116 => x"79",
          3117 => x"ff",
          3118 => x"2b",
          3119 => x"73",
          3120 => x"81",
          3121 => x"87",
          3122 => x"57",
          3123 => x"78",
          3124 => x"11",
          3125 => x"05",
          3126 => x"c0",
          3127 => x"57",
          3128 => x"2e",
          3129 => x"59",
          3130 => x"39",
          3131 => x"0b",
          3132 => x"81",
          3133 => x"70",
          3134 => x"59",
          3135 => x"09",
          3136 => x"2e",
          3137 => x"10",
          3138 => x"5d",
          3139 => x"81",
          3140 => x"93",
          3141 => x"33",
          3142 => x"84",
          3143 => x"38",
          3144 => x"cc",
          3145 => x"8f",
          3146 => x"f0",
          3147 => x"2e",
          3148 => x"81",
          3149 => x"34",
          3150 => x"90",
          3151 => x"15",
          3152 => x"34",
          3153 => x"53",
          3154 => x"83",
          3155 => x"27",
          3156 => x"54",
          3157 => x"fc",
          3158 => x"05",
          3159 => x"74",
          3160 => x"98",
          3161 => x"81",
          3162 => x"0b",
          3163 => x"39",
          3164 => x"81",
          3165 => x"83",
          3166 => x"a1",
          3167 => x"a2",
          3168 => x"f7",
          3169 => x"5e",
          3170 => x"09",
          3171 => x"7a",
          3172 => x"2e",
          3173 => x"93",
          3174 => x"f8",
          3175 => x"33",
          3176 => x"73",
          3177 => x"ac",
          3178 => x"58",
          3179 => x"84",
          3180 => x"39",
          3181 => x"2e",
          3182 => x"a8",
          3183 => x"33",
          3184 => x"5a",
          3185 => x"55",
          3186 => x"ff",
          3187 => x"27",
          3188 => x"f8",
          3189 => x"ff",
          3190 => x"27",
          3191 => x"f9",
          3192 => x"52",
          3193 => x"59",
          3194 => x"39",
          3195 => x"51",
          3196 => x"f7",
          3197 => x"fc",
          3198 => x"f5",
          3199 => x"3d",
          3200 => x"53",
          3201 => x"34",
          3202 => x"71",
          3203 => x"55",
          3204 => x"0b",
          3205 => x"98",
          3206 => x"80",
          3207 => x"9c",
          3208 => x"51",
          3209 => x"33",
          3210 => x"74",
          3211 => x"2e",
          3212 => x"51",
          3213 => x"38",
          3214 => x"38",
          3215 => x"90",
          3216 => x"52",
          3217 => x"72",
          3218 => x"c0",
          3219 => x"27",
          3220 => x"38",
          3221 => x"75",
          3222 => x"ff",
          3223 => x"75",
          3224 => x"06",
          3225 => x"2e",
          3226 => x"88",
          3227 => x"c8",
          3228 => x"0d",
          3229 => x"56",
          3230 => x"73",
          3231 => x"70",
          3232 => x"57",
          3233 => x"51",
          3234 => x"56",
          3235 => x"34",
          3236 => x"13",
          3237 => x"e1",
          3238 => x"08",
          3239 => x"80",
          3240 => x"c0",
          3241 => x"55",
          3242 => x"98",
          3243 => x"08",
          3244 => x"14",
          3245 => x"52",
          3246 => x"fe",
          3247 => x"08",
          3248 => x"c8",
          3249 => x"c0",
          3250 => x"ce",
          3251 => x"08",
          3252 => x"74",
          3253 => x"87",
          3254 => x"73",
          3255 => x"db",
          3256 => x"72",
          3257 => x"55",
          3258 => x"53",
          3259 => x"81",
          3260 => x"74",
          3261 => x"aa",
          3262 => x"11",
          3263 => x"38",
          3264 => x"70",
          3265 => x"f0",
          3266 => x"3d",
          3267 => x"0c",
          3268 => x"39",
          3269 => x"a3",
          3270 => x"f3",
          3271 => x"80",
          3272 => x"51",
          3273 => x"72",
          3274 => x"75",
          3275 => x"72",
          3276 => x"08",
          3277 => x"54",
          3278 => x"70",
          3279 => x"81",
          3280 => x"38",
          3281 => x"15",
          3282 => x"e2",
          3283 => x"08",
          3284 => x"80",
          3285 => x"c0",
          3286 => x"55",
          3287 => x"98",
          3288 => x"08",
          3289 => x"14",
          3290 => x"52",
          3291 => x"fe",
          3292 => x"08",
          3293 => x"c8",
          3294 => x"c0",
          3295 => x"ce",
          3296 => x"08",
          3297 => x"74",
          3298 => x"87",
          3299 => x"73",
          3300 => x"db",
          3301 => x"72",
          3302 => x"55",
          3303 => x"53",
          3304 => x"ff",
          3305 => x"51",
          3306 => x"2e",
          3307 => x"c8",
          3308 => x"e8",
          3309 => x"08",
          3310 => x"83",
          3311 => x"81",
          3312 => x"e8",
          3313 => x"f3",
          3314 => x"54",
          3315 => x"c0",
          3316 => x"f6",
          3317 => x"9c",
          3318 => x"38",
          3319 => x"c0",
          3320 => x"74",
          3321 => x"ff",
          3322 => x"9c",
          3323 => x"c0",
          3324 => x"9c",
          3325 => x"81",
          3326 => x"55",
          3327 => x"81",
          3328 => x"a4",
          3329 => x"ff",
          3330 => x"ff",
          3331 => x"38",
          3332 => x"d5",
          3333 => x"e4",
          3334 => x"3d",
          3335 => x"b8",
          3336 => x"83",
          3337 => x"11",
          3338 => x"2b",
          3339 => x"33",
          3340 => x"90",
          3341 => x"5d",
          3342 => x"71",
          3343 => x"11",
          3344 => x"71",
          3345 => x"81",
          3346 => x"2b",
          3347 => x"52",
          3348 => x"13",
          3349 => x"71",
          3350 => x"2a",
          3351 => x"34",
          3352 => x"13",
          3353 => x"84",
          3354 => x"2b",
          3355 => x"54",
          3356 => x"14",
          3357 => x"80",
          3358 => x"13",
          3359 => x"84",
          3360 => x"b9",
          3361 => x"33",
          3362 => x"07",
          3363 => x"74",
          3364 => x"3d",
          3365 => x"33",
          3366 => x"75",
          3367 => x"71",
          3368 => x"58",
          3369 => x"12",
          3370 => x"b8",
          3371 => x"12",
          3372 => x"07",
          3373 => x"12",
          3374 => x"07",
          3375 => x"77",
          3376 => x"84",
          3377 => x"12",
          3378 => x"ff",
          3379 => x"52",
          3380 => x"84",
          3381 => x"81",
          3382 => x"2b",
          3383 => x"33",
          3384 => x"8f",
          3385 => x"2a",
          3386 => x"54",
          3387 => x"14",
          3388 => x"70",
          3389 => x"71",
          3390 => x"81",
          3391 => x"ff",
          3392 => x"53",
          3393 => x"34",
          3394 => x"08",
          3395 => x"33",
          3396 => x"74",
          3397 => x"98",
          3398 => x"5d",
          3399 => x"25",
          3400 => x"33",
          3401 => x"07",
          3402 => x"75",
          3403 => x"b8",
          3404 => x"33",
          3405 => x"74",
          3406 => x"71",
          3407 => x"5c",
          3408 => x"82",
          3409 => x"3d",
          3410 => x"b9",
          3411 => x"8f",
          3412 => x"51",
          3413 => x"84",
          3414 => x"a0",
          3415 => x"80",
          3416 => x"51",
          3417 => x"08",
          3418 => x"16",
          3419 => x"84",
          3420 => x"84",
          3421 => x"34",
          3422 => x"b8",
          3423 => x"fe",
          3424 => x"06",
          3425 => x"74",
          3426 => x"84",
          3427 => x"84",
          3428 => x"55",
          3429 => x"15",
          3430 => x"7b",
          3431 => x"27",
          3432 => x"05",
          3433 => x"70",
          3434 => x"08",
          3435 => x"88",
          3436 => x"55",
          3437 => x"80",
          3438 => x"70",
          3439 => x"07",
          3440 => x"70",
          3441 => x"56",
          3442 => x"27",
          3443 => x"75",
          3444 => x"13",
          3445 => x"75",
          3446 => x"85",
          3447 => x"83",
          3448 => x"33",
          3449 => x"ff",
          3450 => x"70",
          3451 => x"51",
          3452 => x"51",
          3453 => x"75",
          3454 => x"83",
          3455 => x"07",
          3456 => x"5a",
          3457 => x"84",
          3458 => x"53",
          3459 => x"14",
          3460 => x"70",
          3461 => x"07",
          3462 => x"74",
          3463 => x"88",
          3464 => x"52",
          3465 => x"06",
          3466 => x"b8",
          3467 => x"81",
          3468 => x"19",
          3469 => x"8b",
          3470 => x"58",
          3471 => x"34",
          3472 => x"08",
          3473 => x"33",
          3474 => x"70",
          3475 => x"86",
          3476 => x"b9",
          3477 => x"85",
          3478 => x"2b",
          3479 => x"52",
          3480 => x"34",
          3481 => x"78",
          3482 => x"71",
          3483 => x"5c",
          3484 => x"85",
          3485 => x"84",
          3486 => x"8b",
          3487 => x"15",
          3488 => x"07",
          3489 => x"33",
          3490 => x"5a",
          3491 => x"12",
          3492 => x"b8",
          3493 => x"12",
          3494 => x"07",
          3495 => x"33",
          3496 => x"58",
          3497 => x"70",
          3498 => x"84",
          3499 => x"12",
          3500 => x"ff",
          3501 => x"57",
          3502 => x"84",
          3503 => x"fe",
          3504 => x"b9",
          3505 => x"a0",
          3506 => x"84",
          3507 => x"77",
          3508 => x"08",
          3509 => x"04",
          3510 => x"0c",
          3511 => x"82",
          3512 => x"f4",
          3513 => x"b8",
          3514 => x"81",
          3515 => x"76",
          3516 => x"34",
          3517 => x"17",
          3518 => x"b9",
          3519 => x"05",
          3520 => x"ff",
          3521 => x"56",
          3522 => x"34",
          3523 => x"10",
          3524 => x"55",
          3525 => x"83",
          3526 => x"fe",
          3527 => x"0d",
          3528 => x"b9",
          3529 => x"2e",
          3530 => x"af",
          3531 => x"81",
          3532 => x"fb",
          3533 => x"ff",
          3534 => x"ff",
          3535 => x"83",
          3536 => x"11",
          3537 => x"2b",
          3538 => x"ff",
          3539 => x"73",
          3540 => x"12",
          3541 => x"2b",
          3542 => x"44",
          3543 => x"52",
          3544 => x"fd",
          3545 => x"71",
          3546 => x"19",
          3547 => x"2b",
          3548 => x"56",
          3549 => x"38",
          3550 => x"1b",
          3551 => x"60",
          3552 => x"58",
          3553 => x"18",
          3554 => x"76",
          3555 => x"8b",
          3556 => x"70",
          3557 => x"71",
          3558 => x"53",
          3559 => x"ba",
          3560 => x"12",
          3561 => x"07",
          3562 => x"33",
          3563 => x"7e",
          3564 => x"71",
          3565 => x"57",
          3566 => x"59",
          3567 => x"1d",
          3568 => x"84",
          3569 => x"2b",
          3570 => x"14",
          3571 => x"07",
          3572 => x"40",
          3573 => x"7b",
          3574 => x"16",
          3575 => x"2b",
          3576 => x"2a",
          3577 => x"79",
          3578 => x"70",
          3579 => x"71",
          3580 => x"05",
          3581 => x"2b",
          3582 => x"5d",
          3583 => x"75",
          3584 => x"70",
          3585 => x"8b",
          3586 => x"82",
          3587 => x"2b",
          3588 => x"5d",
          3589 => x"34",
          3590 => x"08",
          3591 => x"33",
          3592 => x"56",
          3593 => x"7e",
          3594 => x"3f",
          3595 => x"61",
          3596 => x"06",
          3597 => x"b6",
          3598 => x"0c",
          3599 => x"0b",
          3600 => x"84",
          3601 => x"60",
          3602 => x"e8",
          3603 => x"7e",
          3604 => x"b9",
          3605 => x"81",
          3606 => x"08",
          3607 => x"87",
          3608 => x"b9",
          3609 => x"07",
          3610 => x"2a",
          3611 => x"34",
          3612 => x"22",
          3613 => x"08",
          3614 => x"15",
          3615 => x"b9",
          3616 => x"76",
          3617 => x"7f",
          3618 => x"f4",
          3619 => x"b9",
          3620 => x"1c",
          3621 => x"71",
          3622 => x"81",
          3623 => x"ff",
          3624 => x"5b",
          3625 => x"1c",
          3626 => x"7c",
          3627 => x"34",
          3628 => x"08",
          3629 => x"71",
          3630 => x"ff",
          3631 => x"ff",
          3632 => x"57",
          3633 => x"34",
          3634 => x"83",
          3635 => x"5b",
          3636 => x"61",
          3637 => x"51",
          3638 => x"39",
          3639 => x"06",
          3640 => x"ff",
          3641 => x"ff",
          3642 => x"71",
          3643 => x"1b",
          3644 => x"2b",
          3645 => x"54",
          3646 => x"f9",
          3647 => x"24",
          3648 => x"8f",
          3649 => x"61",
          3650 => x"39",
          3651 => x"0c",
          3652 => x"82",
          3653 => x"f4",
          3654 => x"b8",
          3655 => x"81",
          3656 => x"7e",
          3657 => x"34",
          3658 => x"19",
          3659 => x"b9",
          3660 => x"05",
          3661 => x"ff",
          3662 => x"44",
          3663 => x"89",
          3664 => x"10",
          3665 => x"f8",
          3666 => x"34",
          3667 => x"39",
          3668 => x"83",
          3669 => x"fb",
          3670 => x"2e",
          3671 => x"3f",
          3672 => x"95",
          3673 => x"33",
          3674 => x"83",
          3675 => x"87",
          3676 => x"2b",
          3677 => x"15",
          3678 => x"2a",
          3679 => x"53",
          3680 => x"34",
          3681 => x"b8",
          3682 => x"12",
          3683 => x"07",
          3684 => x"33",
          3685 => x"5b",
          3686 => x"73",
          3687 => x"05",
          3688 => x"33",
          3689 => x"81",
          3690 => x"5c",
          3691 => x"1e",
          3692 => x"82",
          3693 => x"2b",
          3694 => x"33",
          3695 => x"70",
          3696 => x"57",
          3697 => x"1d",
          3698 => x"70",
          3699 => x"71",
          3700 => x"33",
          3701 => x"70",
          3702 => x"5c",
          3703 => x"83",
          3704 => x"1f",
          3705 => x"88",
          3706 => x"83",
          3707 => x"84",
          3708 => x"b9",
          3709 => x"ff",
          3710 => x"84",
          3711 => x"a0",
          3712 => x"80",
          3713 => x"51",
          3714 => x"08",
          3715 => x"17",
          3716 => x"84",
          3717 => x"84",
          3718 => x"34",
          3719 => x"b8",
          3720 => x"fe",
          3721 => x"06",
          3722 => x"61",
          3723 => x"84",
          3724 => x"84",
          3725 => x"5d",
          3726 => x"1c",
          3727 => x"54",
          3728 => x"1a",
          3729 => x"07",
          3730 => x"33",
          3731 => x"5c",
          3732 => x"84",
          3733 => x"84",
          3734 => x"33",
          3735 => x"83",
          3736 => x"87",
          3737 => x"88",
          3738 => x"59",
          3739 => x"64",
          3740 => x"1d",
          3741 => x"2b",
          3742 => x"2a",
          3743 => x"7f",
          3744 => x"70",
          3745 => x"8b",
          3746 => x"70",
          3747 => x"07",
          3748 => x"77",
          3749 => x"5a",
          3750 => x"17",
          3751 => x"b8",
          3752 => x"33",
          3753 => x"74",
          3754 => x"88",
          3755 => x"88",
          3756 => x"41",
          3757 => x"05",
          3758 => x"fa",
          3759 => x"33",
          3760 => x"79",
          3761 => x"71",
          3762 => x"5e",
          3763 => x"34",
          3764 => x"08",
          3765 => x"33",
          3766 => x"74",
          3767 => x"71",
          3768 => x"56",
          3769 => x"60",
          3770 => x"34",
          3771 => x"81",
          3772 => x"ff",
          3773 => x"58",
          3774 => x"34",
          3775 => x"33",
          3776 => x"83",
          3777 => x"12",
          3778 => x"2b",
          3779 => x"88",
          3780 => x"42",
          3781 => x"83",
          3782 => x"1f",
          3783 => x"2b",
          3784 => x"33",
          3785 => x"81",
          3786 => x"54",
          3787 => x"7c",
          3788 => x"b8",
          3789 => x"12",
          3790 => x"07",
          3791 => x"33",
          3792 => x"78",
          3793 => x"71",
          3794 => x"57",
          3795 => x"5a",
          3796 => x"85",
          3797 => x"17",
          3798 => x"8b",
          3799 => x"86",
          3800 => x"2b",
          3801 => x"52",
          3802 => x"34",
          3803 => x"08",
          3804 => x"88",
          3805 => x"88",
          3806 => x"34",
          3807 => x"08",
          3808 => x"33",
          3809 => x"74",
          3810 => x"88",
          3811 => x"45",
          3812 => x"34",
          3813 => x"08",
          3814 => x"71",
          3815 => x"05",
          3816 => x"88",
          3817 => x"45",
          3818 => x"1a",
          3819 => x"b8",
          3820 => x"12",
          3821 => x"62",
          3822 => x"5d",
          3823 => x"c3",
          3824 => x"05",
          3825 => x"ff",
          3826 => x"86",
          3827 => x"2b",
          3828 => x"1c",
          3829 => x"07",
          3830 => x"41",
          3831 => x"61",
          3832 => x"70",
          3833 => x"71",
          3834 => x"05",
          3835 => x"88",
          3836 => x"5f",
          3837 => x"86",
          3838 => x"84",
          3839 => x"12",
          3840 => x"ff",
          3841 => x"55",
          3842 => x"84",
          3843 => x"81",
          3844 => x"2b",
          3845 => x"33",
          3846 => x"8f",
          3847 => x"2a",
          3848 => x"58",
          3849 => x"1e",
          3850 => x"70",
          3851 => x"71",
          3852 => x"81",
          3853 => x"ff",
          3854 => x"49",
          3855 => x"34",
          3856 => x"ff",
          3857 => x"52",
          3858 => x"08",
          3859 => x"93",
          3860 => x"c8",
          3861 => x"51",
          3862 => x"27",
          3863 => x"3d",
          3864 => x"08",
          3865 => x"77",
          3866 => x"c8",
          3867 => x"e4",
          3868 => x"84",
          3869 => x"77",
          3870 => x"51",
          3871 => x"c8",
          3872 => x"f4",
          3873 => x"0b",
          3874 => x"53",
          3875 => x"b6",
          3876 => x"76",
          3877 => x"84",
          3878 => x"34",
          3879 => x"b8",
          3880 => x"0b",
          3881 => x"84",
          3882 => x"80",
          3883 => x"88",
          3884 => x"17",
          3885 => x"b4",
          3886 => x"b8",
          3887 => x"82",
          3888 => x"77",
          3889 => x"fe",
          3890 => x"05",
          3891 => x"87",
          3892 => x"71",
          3893 => x"04",
          3894 => x"52",
          3895 => x"71",
          3896 => x"08",
          3897 => x"72",
          3898 => x"c4",
          3899 => x"0c",
          3900 => x"7c",
          3901 => x"33",
          3902 => x"74",
          3903 => x"33",
          3904 => x"73",
          3905 => x"c0",
          3906 => x"76",
          3907 => x"08",
          3908 => x"a7",
          3909 => x"73",
          3910 => x"74",
          3911 => x"2e",
          3912 => x"84",
          3913 => x"84",
          3914 => x"06",
          3915 => x"ac",
          3916 => x"7e",
          3917 => x"5a",
          3918 => x"26",
          3919 => x"54",
          3920 => x"bd",
          3921 => x"98",
          3922 => x"51",
          3923 => x"81",
          3924 => x"38",
          3925 => x"e2",
          3926 => x"fc",
          3927 => x"83",
          3928 => x"b9",
          3929 => x"80",
          3930 => x"5a",
          3931 => x"38",
          3932 => x"84",
          3933 => x"9f",
          3934 => x"71",
          3935 => x"12",
          3936 => x"53",
          3937 => x"98",
          3938 => x"96",
          3939 => x"83",
          3940 => x"b9",
          3941 => x"80",
          3942 => x"0c",
          3943 => x"0c",
          3944 => x"3d",
          3945 => x"92",
          3946 => x"71",
          3947 => x"51",
          3948 => x"98",
          3949 => x"c0",
          3950 => x"81",
          3951 => x"52",
          3952 => x"2e",
          3953 => x"54",
          3954 => x"3d",
          3955 => x"33",
          3956 => x"09",
          3957 => x"75",
          3958 => x"80",
          3959 => x"3f",
          3960 => x"38",
          3961 => x"8c",
          3962 => x"08",
          3963 => x"33",
          3964 => x"84",
          3965 => x"06",
          3966 => x"19",
          3967 => x"08",
          3968 => x"08",
          3969 => x"ff",
          3970 => x"82",
          3971 => x"81",
          3972 => x"18",
          3973 => x"33",
          3974 => x"06",
          3975 => x"76",
          3976 => x"38",
          3977 => x"57",
          3978 => x"ff",
          3979 => x"0b",
          3980 => x"84",
          3981 => x"80",
          3982 => x"0b",
          3983 => x"19",
          3984 => x"34",
          3985 => x"80",
          3986 => x"e1",
          3987 => x"08",
          3988 => x"88",
          3989 => x"74",
          3990 => x"34",
          3991 => x"19",
          3992 => x"a4",
          3993 => x"84",
          3994 => x"75",
          3995 => x"55",
          3996 => x"08",
          3997 => x"81",
          3998 => x"33",
          3999 => x"34",
          4000 => x"51",
          4001 => x"80",
          4002 => x"f3",
          4003 => x"56",
          4004 => x"17",
          4005 => x"77",
          4006 => x"04",
          4007 => x"2e",
          4008 => x"a5",
          4009 => x"dd",
          4010 => x"2a",
          4011 => x"5b",
          4012 => x"83",
          4013 => x"81",
          4014 => x"53",
          4015 => x"f8",
          4016 => x"2e",
          4017 => x"b4",
          4018 => x"83",
          4019 => x"1c",
          4020 => x"53",
          4021 => x"2e",
          4022 => x"71",
          4023 => x"81",
          4024 => x"53",
          4025 => x"f8",
          4026 => x"2e",
          4027 => x"b4",
          4028 => x"83",
          4029 => x"88",
          4030 => x"84",
          4031 => x"fe",
          4032 => x"b9",
          4033 => x"88",
          4034 => x"17",
          4035 => x"83",
          4036 => x"7b",
          4037 => x"81",
          4038 => x"17",
          4039 => x"c8",
          4040 => x"81",
          4041 => x"df",
          4042 => x"05",
          4043 => x"71",
          4044 => x"57",
          4045 => x"2e",
          4046 => x"87",
          4047 => x"17",
          4048 => x"83",
          4049 => x"7b",
          4050 => x"81",
          4051 => x"17",
          4052 => x"c8",
          4053 => x"81",
          4054 => x"f7",
          4055 => x"77",
          4056 => x"12",
          4057 => x"07",
          4058 => x"2b",
          4059 => x"80",
          4060 => x"5c",
          4061 => x"04",
          4062 => x"17",
          4063 => x"f6",
          4064 => x"08",
          4065 => x"38",
          4066 => x"b4",
          4067 => x"b9",
          4068 => x"08",
          4069 => x"55",
          4070 => x"f7",
          4071 => x"18",
          4072 => x"33",
          4073 => x"df",
          4074 => x"b8",
          4075 => x"5c",
          4076 => x"7b",
          4077 => x"84",
          4078 => x"17",
          4079 => x"a0",
          4080 => x"33",
          4081 => x"84",
          4082 => x"81",
          4083 => x"70",
          4084 => x"bb",
          4085 => x"7b",
          4086 => x"84",
          4087 => x"17",
          4088 => x"c8",
          4089 => x"27",
          4090 => x"74",
          4091 => x"38",
          4092 => x"08",
          4093 => x"51",
          4094 => x"39",
          4095 => x"17",
          4096 => x"f4",
          4097 => x"08",
          4098 => x"38",
          4099 => x"b4",
          4100 => x"b9",
          4101 => x"08",
          4102 => x"55",
          4103 => x"84",
          4104 => x"18",
          4105 => x"33",
          4106 => x"ec",
          4107 => x"18",
          4108 => x"33",
          4109 => x"81",
          4110 => x"39",
          4111 => x"57",
          4112 => x"38",
          4113 => x"78",
          4114 => x"74",
          4115 => x"2e",
          4116 => x"0c",
          4117 => x"a8",
          4118 => x"1a",
          4119 => x"b6",
          4120 => x"7c",
          4121 => x"38",
          4122 => x"81",
          4123 => x"b9",
          4124 => x"58",
          4125 => x"58",
          4126 => x"fe",
          4127 => x"06",
          4128 => x"88",
          4129 => x"0b",
          4130 => x"0c",
          4131 => x"09",
          4132 => x"2a",
          4133 => x"b4",
          4134 => x"85",
          4135 => x"5d",
          4136 => x"bd",
          4137 => x"52",
          4138 => x"84",
          4139 => x"ff",
          4140 => x"79",
          4141 => x"2b",
          4142 => x"83",
          4143 => x"06",
          4144 => x"5e",
          4145 => x"56",
          4146 => x"5a",
          4147 => x"5b",
          4148 => x"1a",
          4149 => x"16",
          4150 => x"b4",
          4151 => x"2e",
          4152 => x"71",
          4153 => x"81",
          4154 => x"53",
          4155 => x"f0",
          4156 => x"2e",
          4157 => x"b4",
          4158 => x"38",
          4159 => x"81",
          4160 => x"7a",
          4161 => x"84",
          4162 => x"06",
          4163 => x"81",
          4164 => x"a8",
          4165 => x"1a",
          4166 => x"dd",
          4167 => x"70",
          4168 => x"9b",
          4169 => x"7f",
          4170 => x"84",
          4171 => x"19",
          4172 => x"1b",
          4173 => x"56",
          4174 => x"19",
          4175 => x"38",
          4176 => x"19",
          4177 => x"c8",
          4178 => x"81",
          4179 => x"83",
          4180 => x"05",
          4181 => x"38",
          4182 => x"06",
          4183 => x"76",
          4184 => x"cb",
          4185 => x"70",
          4186 => x"8b",
          4187 => x"7c",
          4188 => x"84",
          4189 => x"19",
          4190 => x"1b",
          4191 => x"40",
          4192 => x"82",
          4193 => x"81",
          4194 => x"1e",
          4195 => x"ee",
          4196 => x"81",
          4197 => x"81",
          4198 => x"81",
          4199 => x"09",
          4200 => x"c8",
          4201 => x"70",
          4202 => x"84",
          4203 => x"74",
          4204 => x"33",
          4205 => x"fc",
          4206 => x"76",
          4207 => x"3f",
          4208 => x"76",
          4209 => x"33",
          4210 => x"84",
          4211 => x"06",
          4212 => x"83",
          4213 => x"1b",
          4214 => x"c8",
          4215 => x"27",
          4216 => x"74",
          4217 => x"38",
          4218 => x"81",
          4219 => x"5a",
          4220 => x"53",
          4221 => x"f3",
          4222 => x"76",
          4223 => x"83",
          4224 => x"b8",
          4225 => x"b9",
          4226 => x"fd",
          4227 => x"fc",
          4228 => x"33",
          4229 => x"f0",
          4230 => x"58",
          4231 => x"75",
          4232 => x"79",
          4233 => x"7a",
          4234 => x"3d",
          4235 => x"5a",
          4236 => x"57",
          4237 => x"9c",
          4238 => x"19",
          4239 => x"80",
          4240 => x"38",
          4241 => x"08",
          4242 => x"77",
          4243 => x"51",
          4244 => x"80",
          4245 => x"b9",
          4246 => x"b9",
          4247 => x"07",
          4248 => x"55",
          4249 => x"2e",
          4250 => x"55",
          4251 => x"0d",
          4252 => x"b9",
          4253 => x"79",
          4254 => x"84",
          4255 => x"b9",
          4256 => x"ff",
          4257 => x"b9",
          4258 => x"fe",
          4259 => x"08",
          4260 => x"52",
          4261 => x"84",
          4262 => x"38",
          4263 => x"70",
          4264 => x"84",
          4265 => x"55",
          4266 => x"08",
          4267 => x"54",
          4268 => x"9c",
          4269 => x"70",
          4270 => x"2e",
          4271 => x"78",
          4272 => x"08",
          4273 => x"b9",
          4274 => x"55",
          4275 => x"38",
          4276 => x"fe",
          4277 => x"78",
          4278 => x"0c",
          4279 => x"84",
          4280 => x"c8",
          4281 => x"84",
          4282 => x"84",
          4283 => x"73",
          4284 => x"7a",
          4285 => x"b9",
          4286 => x"b9",
          4287 => x"3d",
          4288 => x"ff",
          4289 => x"f8",
          4290 => x"55",
          4291 => x"df",
          4292 => x"d7",
          4293 => x"08",
          4294 => x"56",
          4295 => x"85",
          4296 => x"5a",
          4297 => x"17",
          4298 => x"0c",
          4299 => x"80",
          4300 => x"98",
          4301 => x"b8",
          4302 => x"84",
          4303 => x"82",
          4304 => x"0d",
          4305 => x"2e",
          4306 => x"89",
          4307 => x"38",
          4308 => x"14",
          4309 => x"8d",
          4310 => x"b0",
          4311 => x"19",
          4312 => x"51",
          4313 => x"55",
          4314 => x"38",
          4315 => x"ff",
          4316 => x"b9",
          4317 => x"73",
          4318 => x"38",
          4319 => x"c8",
          4320 => x"0d",
          4321 => x"05",
          4322 => x"27",
          4323 => x"98",
          4324 => x"2e",
          4325 => x"7a",
          4326 => x"57",
          4327 => x"88",
          4328 => x"81",
          4329 => x"90",
          4330 => x"18",
          4331 => x"0c",
          4332 => x"0c",
          4333 => x"2a",
          4334 => x"76",
          4335 => x"08",
          4336 => x"c8",
          4337 => x"b9",
          4338 => x"19",
          4339 => x"91",
          4340 => x"94",
          4341 => x"3f",
          4342 => x"84",
          4343 => x"38",
          4344 => x"2e",
          4345 => x"c8",
          4346 => x"b9",
          4347 => x"7d",
          4348 => x"08",
          4349 => x"78",
          4350 => x"71",
          4351 => x"7b",
          4352 => x"80",
          4353 => x"05",
          4354 => x"38",
          4355 => x"75",
          4356 => x"1c",
          4357 => x"e4",
          4358 => x"e7",
          4359 => x"98",
          4360 => x"0c",
          4361 => x"19",
          4362 => x"1a",
          4363 => x"b9",
          4364 => x"c8",
          4365 => x"a8",
          4366 => x"08",
          4367 => x"5c",
          4368 => x"db",
          4369 => x"1a",
          4370 => x"33",
          4371 => x"8a",
          4372 => x"06",
          4373 => x"a7",
          4374 => x"9c",
          4375 => x"58",
          4376 => x"19",
          4377 => x"05",
          4378 => x"81",
          4379 => x"0d",
          4380 => x"5c",
          4381 => x"70",
          4382 => x"80",
          4383 => x"75",
          4384 => x"2e",
          4385 => x"58",
          4386 => x"81",
          4387 => x"19",
          4388 => x"3f",
          4389 => x"38",
          4390 => x"0c",
          4391 => x"1c",
          4392 => x"2e",
          4393 => x"06",
          4394 => x"86",
          4395 => x"30",
          4396 => x"25",
          4397 => x"57",
          4398 => x"06",
          4399 => x"38",
          4400 => x"ff",
          4401 => x"3f",
          4402 => x"c8",
          4403 => x"56",
          4404 => x"c8",
          4405 => x"b4",
          4406 => x"33",
          4407 => x"b9",
          4408 => x"fe",
          4409 => x"1a",
          4410 => x"31",
          4411 => x"a0",
          4412 => x"19",
          4413 => x"06",
          4414 => x"08",
          4415 => x"81",
          4416 => x"57",
          4417 => x"81",
          4418 => x"81",
          4419 => x"8d",
          4420 => x"90",
          4421 => x"5e",
          4422 => x"ff",
          4423 => x"56",
          4424 => x"be",
          4425 => x"98",
          4426 => x"94",
          4427 => x"39",
          4428 => x"09",
          4429 => x"9b",
          4430 => x"2b",
          4431 => x"38",
          4432 => x"29",
          4433 => x"5b",
          4434 => x"81",
          4435 => x"07",
          4436 => x"c5",
          4437 => x"38",
          4438 => x"75",
          4439 => x"57",
          4440 => x"70",
          4441 => x"80",
          4442 => x"fe",
          4443 => x"80",
          4444 => x"06",
          4445 => x"ff",
          4446 => x"fe",
          4447 => x"8b",
          4448 => x"29",
          4449 => x"40",
          4450 => x"19",
          4451 => x"7e",
          4452 => x"1d",
          4453 => x"3d",
          4454 => x"08",
          4455 => x"cf",
          4456 => x"b9",
          4457 => x"70",
          4458 => x"b8",
          4459 => x"58",
          4460 => x"38",
          4461 => x"78",
          4462 => x"81",
          4463 => x"1b",
          4464 => x"c8",
          4465 => x"81",
          4466 => x"76",
          4467 => x"33",
          4468 => x"38",
          4469 => x"ff",
          4470 => x"76",
          4471 => x"83",
          4472 => x"81",
          4473 => x"8f",
          4474 => x"78",
          4475 => x"2a",
          4476 => x"81",
          4477 => x"81",
          4478 => x"76",
          4479 => x"38",
          4480 => x"a7",
          4481 => x"78",
          4482 => x"81",
          4483 => x"1a",
          4484 => x"81",
          4485 => x"81",
          4486 => x"80",
          4487 => x"b9",
          4488 => x"80",
          4489 => x"c8",
          4490 => x"b4",
          4491 => x"33",
          4492 => x"b9",
          4493 => x"fe",
          4494 => x"1c",
          4495 => x"31",
          4496 => x"a0",
          4497 => x"1b",
          4498 => x"06",
          4499 => x"08",
          4500 => x"81",
          4501 => x"57",
          4502 => x"39",
          4503 => x"06",
          4504 => x"86",
          4505 => x"93",
          4506 => x"06",
          4507 => x"0c",
          4508 => x"38",
          4509 => x"7b",
          4510 => x"08",
          4511 => x"fc",
          4512 => x"2e",
          4513 => x"0b",
          4514 => x"19",
          4515 => x"06",
          4516 => x"33",
          4517 => x"59",
          4518 => x"33",
          4519 => x"5b",
          4520 => x"c8",
          4521 => x"71",
          4522 => x"57",
          4523 => x"81",
          4524 => x"81",
          4525 => x"7a",
          4526 => x"81",
          4527 => x"75",
          4528 => x"06",
          4529 => x"58",
          4530 => x"33",
          4531 => x"75",
          4532 => x"8d",
          4533 => x"41",
          4534 => x"70",
          4535 => x"39",
          4536 => x"3d",
          4537 => x"ff",
          4538 => x"39",
          4539 => x"ab",
          4540 => x"5d",
          4541 => x"74",
          4542 => x"5d",
          4543 => x"70",
          4544 => x"74",
          4545 => x"40",
          4546 => x"70",
          4547 => x"05",
          4548 => x"38",
          4549 => x"06",
          4550 => x"38",
          4551 => x"0b",
          4552 => x"7b",
          4553 => x"55",
          4554 => x"70",
          4555 => x"74",
          4556 => x"38",
          4557 => x"2e",
          4558 => x"8f",
          4559 => x"76",
          4560 => x"72",
          4561 => x"57",
          4562 => x"a0",
          4563 => x"80",
          4564 => x"ca",
          4565 => x"05",
          4566 => x"55",
          4567 => x"55",
          4568 => x"78",
          4569 => x"38",
          4570 => x"76",
          4571 => x"38",
          4572 => x"38",
          4573 => x"a2",
          4574 => x"74",
          4575 => x"81",
          4576 => x"8e",
          4577 => x"81",
          4578 => x"77",
          4579 => x"7d",
          4580 => x"08",
          4581 => x"7b",
          4582 => x"80",
          4583 => x"c8",
          4584 => x"2e",
          4585 => x"80",
          4586 => x"08",
          4587 => x"57",
          4588 => x"81",
          4589 => x"52",
          4590 => x"84",
          4591 => x"7d",
          4592 => x"08",
          4593 => x"38",
          4594 => x"59",
          4595 => x"18",
          4596 => x"18",
          4597 => x"06",
          4598 => x"b8",
          4599 => x"a4",
          4600 => x"85",
          4601 => x"19",
          4602 => x"1e",
          4603 => x"e5",
          4604 => x"80",
          4605 => x"2e",
          4606 => x"7b",
          4607 => x"51",
          4608 => x"56",
          4609 => x"88",
          4610 => x"89",
          4611 => x"ff",
          4612 => x"1e",
          4613 => x"af",
          4614 => x"7f",
          4615 => x"b8",
          4616 => x"9c",
          4617 => x"85",
          4618 => x"1d",
          4619 => x"a0",
          4620 => x"76",
          4621 => x"55",
          4622 => x"08",
          4623 => x"05",
          4624 => x"34",
          4625 => x"1e",
          4626 => x"5a",
          4627 => x"1d",
          4628 => x"0c",
          4629 => x"70",
          4630 => x"74",
          4631 => x"7d",
          4632 => x"08",
          4633 => x"fd",
          4634 => x"b4",
          4635 => x"33",
          4636 => x"08",
          4637 => x"38",
          4638 => x"b4",
          4639 => x"74",
          4640 => x"18",
          4641 => x"38",
          4642 => x"39",
          4643 => x"31",
          4644 => x"84",
          4645 => x"08",
          4646 => x"08",
          4647 => x"75",
          4648 => x"05",
          4649 => x"ff",
          4650 => x"e4",
          4651 => x"43",
          4652 => x"b4",
          4653 => x"1c",
          4654 => x"06",
          4655 => x"b8",
          4656 => x"dc",
          4657 => x"85",
          4658 => x"1d",
          4659 => x"8c",
          4660 => x"ff",
          4661 => x"34",
          4662 => x"1c",
          4663 => x"1c",
          4664 => x"77",
          4665 => x"2e",
          4666 => x"81",
          4667 => x"18",
          4668 => x"81",
          4669 => x"75",
          4670 => x"ff",
          4671 => x"cb",
          4672 => x"b3",
          4673 => x"58",
          4674 => x"7b",
          4675 => x"52",
          4676 => x"c8",
          4677 => x"f1",
          4678 => x"a9",
          4679 => x"1c",
          4680 => x"1d",
          4681 => x"56",
          4682 => x"84",
          4683 => x"1c",
          4684 => x"c8",
          4685 => x"27",
          4686 => x"61",
          4687 => x"38",
          4688 => x"08",
          4689 => x"51",
          4690 => x"39",
          4691 => x"43",
          4692 => x"06",
          4693 => x"70",
          4694 => x"38",
          4695 => x"5d",
          4696 => x"08",
          4697 => x"cf",
          4698 => x"2e",
          4699 => x"c8",
          4700 => x"a8",
          4701 => x"08",
          4702 => x"7e",
          4703 => x"08",
          4704 => x"41",
          4705 => x"fc",
          4706 => x"39",
          4707 => x"fc",
          4708 => x"b4",
          4709 => x"61",
          4710 => x"3f",
          4711 => x"08",
          4712 => x"81",
          4713 => x"e3",
          4714 => x"08",
          4715 => x"34",
          4716 => x"38",
          4717 => x"38",
          4718 => x"70",
          4719 => x"78",
          4720 => x"70",
          4721 => x"82",
          4722 => x"83",
          4723 => x"ff",
          4724 => x"76",
          4725 => x"79",
          4726 => x"70",
          4727 => x"18",
          4728 => x"34",
          4729 => x"9c",
          4730 => x"58",
          4731 => x"74",
          4732 => x"32",
          4733 => x"55",
          4734 => x"72",
          4735 => x"81",
          4736 => x"77",
          4737 => x"58",
          4738 => x"18",
          4739 => x"34",
          4740 => x"77",
          4741 => x"34",
          4742 => x"80",
          4743 => x"8c",
          4744 => x"73",
          4745 => x"8b",
          4746 => x"08",
          4747 => x"33",
          4748 => x"81",
          4749 => x"75",
          4750 => x"16",
          4751 => x"07",
          4752 => x"55",
          4753 => x"98",
          4754 => x"54",
          4755 => x"04",
          4756 => x"1d",
          4757 => x"5b",
          4758 => x"74",
          4759 => x"b9",
          4760 => x"81",
          4761 => x"27",
          4762 => x"73",
          4763 => x"78",
          4764 => x"56",
          4765 => x"5c",
          4766 => x"ba",
          4767 => x"07",
          4768 => x"55",
          4769 => x"34",
          4770 => x"1f",
          4771 => x"89",
          4772 => x"2e",
          4773 => x"57",
          4774 => x"11",
          4775 => x"9c",
          4776 => x"88",
          4777 => x"53",
          4778 => x"8a",
          4779 => x"06",
          4780 => x"5a",
          4781 => x"71",
          4782 => x"56",
          4783 => x"72",
          4784 => x"30",
          4785 => x"53",
          4786 => x"3d",
          4787 => x"5c",
          4788 => x"74",
          4789 => x"80",
          4790 => x"2e",
          4791 => x"1d",
          4792 => x"41",
          4793 => x"38",
          4794 => x"57",
          4795 => x"55",
          4796 => x"0c",
          4797 => x"ff",
          4798 => x"18",
          4799 => x"73",
          4800 => x"70",
          4801 => x"07",
          4802 => x"38",
          4803 => x"74",
          4804 => x"e4",
          4805 => x"ff",
          4806 => x"81",
          4807 => x"81",
          4808 => x"56",
          4809 => x"ff",
          4810 => x"81",
          4811 => x"18",
          4812 => x"70",
          4813 => x"57",
          4814 => x"cb",
          4815 => x"30",
          4816 => x"58",
          4817 => x"14",
          4818 => x"55",
          4819 => x"dc",
          4820 => x"07",
          4821 => x"88",
          4822 => x"3d",
          4823 => x"90",
          4824 => x"51",
          4825 => x"08",
          4826 => x"8d",
          4827 => x"0c",
          4828 => x"33",
          4829 => x"80",
          4830 => x"80",
          4831 => x"51",
          4832 => x"84",
          4833 => x"81",
          4834 => x"80",
          4835 => x"7d",
          4836 => x"80",
          4837 => x"af",
          4838 => x"70",
          4839 => x"54",
          4840 => x"9f",
          4841 => x"2e",
          4842 => x"d1",
          4843 => x"a7",
          4844 => x"70",
          4845 => x"9f",
          4846 => x"7c",
          4847 => x"ff",
          4848 => x"77",
          4849 => x"2e",
          4850 => x"83",
          4851 => x"56",
          4852 => x"83",
          4853 => x"82",
          4854 => x"77",
          4855 => x"78",
          4856 => x"fe",
          4857 => x"2e",
          4858 => x"54",
          4859 => x"38",
          4860 => x"74",
          4861 => x"53",
          4862 => x"88",
          4863 => x"57",
          4864 => x"38",
          4865 => x"ae",
          4866 => x"5a",
          4867 => x"72",
          4868 => x"26",
          4869 => x"70",
          4870 => x"7c",
          4871 => x"2e",
          4872 => x"83",
          4873 => x"83",
          4874 => x"76",
          4875 => x"81",
          4876 => x"77",
          4877 => x"53",
          4878 => x"57",
          4879 => x"7c",
          4880 => x"06",
          4881 => x"7d",
          4882 => x"e3",
          4883 => x"75",
          4884 => x"80",
          4885 => x"7d",
          4886 => x"2e",
          4887 => x"ab",
          4888 => x"84",
          4889 => x"54",
          4890 => x"ac",
          4891 => x"09",
          4892 => x"2a",
          4893 => x"f0",
          4894 => x"78",
          4895 => x"56",
          4896 => x"57",
          4897 => x"79",
          4898 => x"7c",
          4899 => x"fd",
          4900 => x"8a",
          4901 => x"2e",
          4902 => x"22",
          4903 => x"fc",
          4904 => x"7b",
          4905 => x"ae",
          4906 => x"54",
          4907 => x"81",
          4908 => x"79",
          4909 => x"7b",
          4910 => x"08",
          4911 => x"c8",
          4912 => x"81",
          4913 => x"1c",
          4914 => x"5d",
          4915 => x"1c",
          4916 => x"d3",
          4917 => x"88",
          4918 => x"54",
          4919 => x"88",
          4920 => x"fe",
          4921 => x"2e",
          4922 => x"fb",
          4923 => x"07",
          4924 => x"7d",
          4925 => x"06",
          4926 => x"06",
          4927 => x"fd",
          4928 => x"7c",
          4929 => x"38",
          4930 => x"34",
          4931 => x"3d",
          4932 => x"38",
          4933 => x"ff",
          4934 => x"38",
          4935 => x"5c",
          4936 => x"5a",
          4937 => x"f6",
          4938 => x"ff",
          4939 => x"55",
          4940 => x"ff",
          4941 => x"54",
          4942 => x"74",
          4943 => x"f0",
          4944 => x"ff",
          4945 => x"80",
          4946 => x"81",
          4947 => x"56",
          4948 => x"ff",
          4949 => x"bf",
          4950 => x"7d",
          4951 => x"53",
          4952 => x"93",
          4953 => x"06",
          4954 => x"58",
          4955 => x"59",
          4956 => x"16",
          4957 => x"b3",
          4958 => x"ff",
          4959 => x"ae",
          4960 => x"1d",
          4961 => x"34",
          4962 => x"14",
          4963 => x"2b",
          4964 => x"1f",
          4965 => x"1b",
          4966 => x"72",
          4967 => x"05",
          4968 => x"5b",
          4969 => x"1d",
          4970 => x"09",
          4971 => x"39",
          4972 => x"f6",
          4973 => x"0c",
          4974 => x"67",
          4975 => x"33",
          4976 => x"7e",
          4977 => x"2e",
          4978 => x"5b",
          4979 => x"ba",
          4980 => x"75",
          4981 => x"a4",
          4982 => x"38",
          4983 => x"70",
          4984 => x"2e",
          4985 => x"81",
          4986 => x"80",
          4987 => x"ff",
          4988 => x"81",
          4989 => x"7c",
          4990 => x"34",
          4991 => x"33",
          4992 => x"33",
          4993 => x"c8",
          4994 => x"41",
          4995 => x"78",
          4996 => x"81",
          4997 => x"38",
          4998 => x"0b",
          4999 => x"81",
          5000 => x"81",
          5001 => x"3f",
          5002 => x"38",
          5003 => x"0c",
          5004 => x"17",
          5005 => x"2b",
          5006 => x"d4",
          5007 => x"26",
          5008 => x"42",
          5009 => x"84",
          5010 => x"81",
          5011 => x"33",
          5012 => x"07",
          5013 => x"81",
          5014 => x"33",
          5015 => x"07",
          5016 => x"17",
          5017 => x"90",
          5018 => x"33",
          5019 => x"71",
          5020 => x"56",
          5021 => x"33",
          5022 => x"ff",
          5023 => x"59",
          5024 => x"38",
          5025 => x"80",
          5026 => x"8a",
          5027 => x"87",
          5028 => x"61",
          5029 => x"80",
          5030 => x"56",
          5031 => x"8f",
          5032 => x"98",
          5033 => x"18",
          5034 => x"74",
          5035 => x"33",
          5036 => x"88",
          5037 => x"07",
          5038 => x"44",
          5039 => x"17",
          5040 => x"2b",
          5041 => x"2e",
          5042 => x"2a",
          5043 => x"38",
          5044 => x"ed",
          5045 => x"84",
          5046 => x"38",
          5047 => x"ff",
          5048 => x"83",
          5049 => x"75",
          5050 => x"5d",
          5051 => x"a4",
          5052 => x"0c",
          5053 => x"7c",
          5054 => x"22",
          5055 => x"e0",
          5056 => x"19",
          5057 => x"10",
          5058 => x"05",
          5059 => x"59",
          5060 => x"b8",
          5061 => x"0b",
          5062 => x"18",
          5063 => x"7c",
          5064 => x"05",
          5065 => x"86",
          5066 => x"18",
          5067 => x"58",
          5068 => x"0d",
          5069 => x"97",
          5070 => x"70",
          5071 => x"89",
          5072 => x"ff",
          5073 => x"2e",
          5074 => x"e5",
          5075 => x"5a",
          5076 => x"79",
          5077 => x"12",
          5078 => x"38",
          5079 => x"55",
          5080 => x"89",
          5081 => x"58",
          5082 => x"55",
          5083 => x"38",
          5084 => x"70",
          5085 => x"07",
          5086 => x"98",
          5087 => x"83",
          5088 => x"f9",
          5089 => x"38",
          5090 => x"58",
          5091 => x"c0",
          5092 => x"81",
          5093 => x"81",
          5094 => x"70",
          5095 => x"77",
          5096 => x"83",
          5097 => x"83",
          5098 => x"5b",
          5099 => x"16",
          5100 => x"2b",
          5101 => x"33",
          5102 => x"1b",
          5103 => x"40",
          5104 => x"0c",
          5105 => x"80",
          5106 => x"1d",
          5107 => x"71",
          5108 => x"f0",
          5109 => x"43",
          5110 => x"7a",
          5111 => x"83",
          5112 => x"7a",
          5113 => x"38",
          5114 => x"81",
          5115 => x"84",
          5116 => x"ff",
          5117 => x"84",
          5118 => x"7f",
          5119 => x"83",
          5120 => x"81",
          5121 => x"33",
          5122 => x"b7",
          5123 => x"70",
          5124 => x"7f",
          5125 => x"38",
          5126 => x"80",
          5127 => x"58",
          5128 => x"38",
          5129 => x"38",
          5130 => x"1a",
          5131 => x"fe",
          5132 => x"80",
          5133 => x"58",
          5134 => x"70",
          5135 => x"ff",
          5136 => x"2e",
          5137 => x"38",
          5138 => x"fc",
          5139 => x"5d",
          5140 => x"71",
          5141 => x"40",
          5142 => x"80",
          5143 => x"39",
          5144 => x"84",
          5145 => x"75",
          5146 => x"85",
          5147 => x"40",
          5148 => x"84",
          5149 => x"83",
          5150 => x"5c",
          5151 => x"33",
          5152 => x"71",
          5153 => x"77",
          5154 => x"2e",
          5155 => x"83",
          5156 => x"81",
          5157 => x"5c",
          5158 => x"58",
          5159 => x"38",
          5160 => x"77",
          5161 => x"81",
          5162 => x"33",
          5163 => x"07",
          5164 => x"06",
          5165 => x"5a",
          5166 => x"83",
          5167 => x"81",
          5168 => x"53",
          5169 => x"ff",
          5170 => x"80",
          5171 => x"77",
          5172 => x"79",
          5173 => x"84",
          5174 => x"57",
          5175 => x"81",
          5176 => x"11",
          5177 => x"71",
          5178 => x"72",
          5179 => x"5e",
          5180 => x"84",
          5181 => x"06",
          5182 => x"11",
          5183 => x"71",
          5184 => x"72",
          5185 => x"47",
          5186 => x"86",
          5187 => x"06",
          5188 => x"11",
          5189 => x"71",
          5190 => x"72",
          5191 => x"94",
          5192 => x"11",
          5193 => x"71",
          5194 => x"72",
          5195 => x"62",
          5196 => x"5c",
          5197 => x"77",
          5198 => x"5d",
          5199 => x"18",
          5200 => x"0c",
          5201 => x"39",
          5202 => x"7a",
          5203 => x"54",
          5204 => x"53",
          5205 => x"b3",
          5206 => x"09",
          5207 => x"c8",
          5208 => x"a8",
          5209 => x"08",
          5210 => x"60",
          5211 => x"c8",
          5212 => x"74",
          5213 => x"81",
          5214 => x"58",
          5215 => x"80",
          5216 => x"5f",
          5217 => x"88",
          5218 => x"80",
          5219 => x"33",
          5220 => x"81",
          5221 => x"75",
          5222 => x"7d",
          5223 => x"40",
          5224 => x"2e",
          5225 => x"39",
          5226 => x"3d",
          5227 => x"39",
          5228 => x"bf",
          5229 => x"18",
          5230 => x"33",
          5231 => x"39",
          5232 => x"33",
          5233 => x"5d",
          5234 => x"80",
          5235 => x"33",
          5236 => x"2e",
          5237 => x"ba",
          5238 => x"33",
          5239 => x"73",
          5240 => x"08",
          5241 => x"80",
          5242 => x"86",
          5243 => x"75",
          5244 => x"38",
          5245 => x"05",
          5246 => x"08",
          5247 => x"3d",
          5248 => x"0c",
          5249 => x"11",
          5250 => x"73",
          5251 => x"81",
          5252 => x"79",
          5253 => x"83",
          5254 => x"7e",
          5255 => x"33",
          5256 => x"9f",
          5257 => x"89",
          5258 => x"56",
          5259 => x"26",
          5260 => x"06",
          5261 => x"58",
          5262 => x"85",
          5263 => x"32",
          5264 => x"79",
          5265 => x"92",
          5266 => x"83",
          5267 => x"fe",
          5268 => x"7a",
          5269 => x"e6",
          5270 => x"fb",
          5271 => x"80",
          5272 => x"54",
          5273 => x"84",
          5274 => x"b9",
          5275 => x"80",
          5276 => x"56",
          5277 => x"0d",
          5278 => x"70",
          5279 => x"c8",
          5280 => x"2e",
          5281 => x"7c",
          5282 => x"2e",
          5283 => x"ea",
          5284 => x"bb",
          5285 => x"7a",
          5286 => x"11",
          5287 => x"07",
          5288 => x"56",
          5289 => x"0b",
          5290 => x"34",
          5291 => x"0b",
          5292 => x"8b",
          5293 => x"0b",
          5294 => x"34",
          5295 => x"a9",
          5296 => x"34",
          5297 => x"9e",
          5298 => x"7e",
          5299 => x"80",
          5300 => x"08",
          5301 => x"81",
          5302 => x"7c",
          5303 => x"79",
          5304 => x"05",
          5305 => x"80",
          5306 => x"06",
          5307 => x"fe",
          5308 => x"70",
          5309 => x"82",
          5310 => x"5e",
          5311 => x"06",
          5312 => x"2a",
          5313 => x"38",
          5314 => x"11",
          5315 => x"0c",
          5316 => x"71",
          5317 => x"40",
          5318 => x"38",
          5319 => x"11",
          5320 => x"71",
          5321 => x"72",
          5322 => x"70",
          5323 => x"51",
          5324 => x"1a",
          5325 => x"34",
          5326 => x"9c",
          5327 => x"55",
          5328 => x"80",
          5329 => x"0c",
          5330 => x"52",
          5331 => x"80",
          5332 => x"92",
          5333 => x"7d",
          5334 => x"78",
          5335 => x"c8",
          5336 => x"26",
          5337 => x"08",
          5338 => x"31",
          5339 => x"33",
          5340 => x"82",
          5341 => x"fc",
          5342 => x"fb",
          5343 => x"fb",
          5344 => x"fb",
          5345 => x"84",
          5346 => x"57",
          5347 => x"7a",
          5348 => x"39",
          5349 => x"98",
          5350 => x"5d",
          5351 => x"7c",
          5352 => x"79",
          5353 => x"c8",
          5354 => x"2e",
          5355 => x"81",
          5356 => x"08",
          5357 => x"74",
          5358 => x"84",
          5359 => x"17",
          5360 => x"56",
          5361 => x"81",
          5362 => x"81",
          5363 => x"55",
          5364 => x"d9",
          5365 => x"0b",
          5366 => x"16",
          5367 => x"71",
          5368 => x"5b",
          5369 => x"8f",
          5370 => x"80",
          5371 => x"a0",
          5372 => x"5e",
          5373 => x"9b",
          5374 => x"2e",
          5375 => x"a9",
          5376 => x"57",
          5377 => x"38",
          5378 => x"09",
          5379 => x"53",
          5380 => x"ff",
          5381 => x"80",
          5382 => x"76",
          5383 => x"1d",
          5384 => x"fb",
          5385 => x"39",
          5386 => x"16",
          5387 => x"ff",
          5388 => x"7d",
          5389 => x"84",
          5390 => x"16",
          5391 => x"c8",
          5392 => x"27",
          5393 => x"74",
          5394 => x"38",
          5395 => x"08",
          5396 => x"51",
          5397 => x"ec",
          5398 => x"f8",
          5399 => x"f8",
          5400 => x"79",
          5401 => x"19",
          5402 => x"5a",
          5403 => x"1a",
          5404 => x"05",
          5405 => x"38",
          5406 => x"76",
          5407 => x"0c",
          5408 => x"80",
          5409 => x"c8",
          5410 => x"39",
          5411 => x"f0",
          5412 => x"40",
          5413 => x"79",
          5414 => x"75",
          5415 => x"74",
          5416 => x"84",
          5417 => x"84",
          5418 => x"55",
          5419 => x"55",
          5420 => x"81",
          5421 => x"81",
          5422 => x"08",
          5423 => x"81",
          5424 => x"38",
          5425 => x"7a",
          5426 => x"05",
          5427 => x"38",
          5428 => x"55",
          5429 => x"ff",
          5430 => x"0c",
          5431 => x"9c",
          5432 => x"60",
          5433 => x"70",
          5434 => x"56",
          5435 => x"15",
          5436 => x"2e",
          5437 => x"75",
          5438 => x"77",
          5439 => x"33",
          5440 => x"c8",
          5441 => x"33",
          5442 => x"b4",
          5443 => x"27",
          5444 => x"1e",
          5445 => x"81",
          5446 => x"59",
          5447 => x"77",
          5448 => x"08",
          5449 => x"08",
          5450 => x"5c",
          5451 => x"84",
          5452 => x"74",
          5453 => x"04",
          5454 => x"08",
          5455 => x"71",
          5456 => x"38",
          5457 => x"77",
          5458 => x"33",
          5459 => x"09",
          5460 => x"76",
          5461 => x"51",
          5462 => x"08",
          5463 => x"5b",
          5464 => x"38",
          5465 => x"11",
          5466 => x"59",
          5467 => x"70",
          5468 => x"05",
          5469 => x"2e",
          5470 => x"56",
          5471 => x"ff",
          5472 => x"39",
          5473 => x"19",
          5474 => x"ff",
          5475 => x"c8",
          5476 => x"9c",
          5477 => x"34",
          5478 => x"84",
          5479 => x"1a",
          5480 => x"33",
          5481 => x"fe",
          5482 => x"a0",
          5483 => x"19",
          5484 => x"5b",
          5485 => x"94",
          5486 => x"1a",
          5487 => x"3f",
          5488 => x"39",
          5489 => x"3f",
          5490 => x"74",
          5491 => x"57",
          5492 => x"34",
          5493 => x"3d",
          5494 => x"82",
          5495 => x"0d",
          5496 => x"66",
          5497 => x"89",
          5498 => x"08",
          5499 => x"33",
          5500 => x"16",
          5501 => x"78",
          5502 => x"41",
          5503 => x"1a",
          5504 => x"1a",
          5505 => x"58",
          5506 => x"38",
          5507 => x"7b",
          5508 => x"7a",
          5509 => x"ff",
          5510 => x"8a",
          5511 => x"06",
          5512 => x"9e",
          5513 => x"2e",
          5514 => x"a1",
          5515 => x"74",
          5516 => x"38",
          5517 => x"16",
          5518 => x"38",
          5519 => x"08",
          5520 => x"85",
          5521 => x"29",
          5522 => x"80",
          5523 => x"89",
          5524 => x"98",
          5525 => x"85",
          5526 => x"7b",
          5527 => x"ff",
          5528 => x"85",
          5529 => x"31",
          5530 => x"84",
          5531 => x"1f",
          5532 => x"56",
          5533 => x"ff",
          5534 => x"75",
          5535 => x"7a",
          5536 => x"79",
          5537 => x"94",
          5538 => x"57",
          5539 => x"74",
          5540 => x"85",
          5541 => x"c0",
          5542 => x"56",
          5543 => x"0d",
          5544 => x"3d",
          5545 => x"82",
          5546 => x"60",
          5547 => x"ff",
          5548 => x"7a",
          5549 => x"57",
          5550 => x"80",
          5551 => x"5f",
          5552 => x"d5",
          5553 => x"52",
          5554 => x"3f",
          5555 => x"38",
          5556 => x"0c",
          5557 => x"08",
          5558 => x"05",
          5559 => x"95",
          5560 => x"75",
          5561 => x"56",
          5562 => x"83",
          5563 => x"b4",
          5564 => x"81",
          5565 => x"3f",
          5566 => x"2e",
          5567 => x"b9",
          5568 => x"08",
          5569 => x"08",
          5570 => x"fe",
          5571 => x"82",
          5572 => x"81",
          5573 => x"05",
          5574 => x"ff",
          5575 => x"39",
          5576 => x"77",
          5577 => x"7f",
          5578 => x"0c",
          5579 => x"9c",
          5580 => x"1a",
          5581 => x"3f",
          5582 => x"c8",
          5583 => x"58",
          5584 => x"ff",
          5585 => x"55",
          5586 => x"e4",
          5587 => x"b8",
          5588 => x"57",
          5589 => x"08",
          5590 => x"83",
          5591 => x"08",
          5592 => x"fd",
          5593 => x"82",
          5594 => x"81",
          5595 => x"05",
          5596 => x"ff",
          5597 => x"39",
          5598 => x"3f",
          5599 => x"74",
          5600 => x"57",
          5601 => x"08",
          5602 => x"33",
          5603 => x"b9",
          5604 => x"c8",
          5605 => x"a8",
          5606 => x"08",
          5607 => x"58",
          5608 => x"8b",
          5609 => x"17",
          5610 => x"33",
          5611 => x"b4",
          5612 => x"fd",
          5613 => x"81",
          5614 => x"0d",
          5615 => x"0b",
          5616 => x"04",
          5617 => x"77",
          5618 => x"75",
          5619 => x"74",
          5620 => x"84",
          5621 => x"83",
          5622 => x"56",
          5623 => x"70",
          5624 => x"80",
          5625 => x"08",
          5626 => x"ac",
          5627 => x"bc",
          5628 => x"52",
          5629 => x"3f",
          5630 => x"38",
          5631 => x"0c",
          5632 => x"8b",
          5633 => x"8b",
          5634 => x"70",
          5635 => x"7a",
          5636 => x"79",
          5637 => x"96",
          5638 => x"81",
          5639 => x"7b",
          5640 => x"18",
          5641 => x"18",
          5642 => x"18",
          5643 => x"18",
          5644 => x"cc",
          5645 => x"18",
          5646 => x"5b",
          5647 => x"ff",
          5648 => x"90",
          5649 => x"79",
          5650 => x"0c",
          5651 => x"17",
          5652 => x"18",
          5653 => x"81",
          5654 => x"38",
          5655 => x"b4",
          5656 => x"b9",
          5657 => x"08",
          5658 => x"55",
          5659 => x"81",
          5660 => x"18",
          5661 => x"33",
          5662 => x"fd",
          5663 => x"94",
          5664 => x"95",
          5665 => x"7b",
          5666 => x"18",
          5667 => x"18",
          5668 => x"18",
          5669 => x"18",
          5670 => x"cc",
          5671 => x"18",
          5672 => x"5b",
          5673 => x"ff",
          5674 => x"90",
          5675 => x"79",
          5676 => x"16",
          5677 => x"b9",
          5678 => x"ba",
          5679 => x"b4",
          5680 => x"55",
          5681 => x"54",
          5682 => x"56",
          5683 => x"53",
          5684 => x"52",
          5685 => x"22",
          5686 => x"2e",
          5687 => x"54",
          5688 => x"84",
          5689 => x"81",
          5690 => x"84",
          5691 => x"da",
          5692 => x"39",
          5693 => x"57",
          5694 => x"70",
          5695 => x"52",
          5696 => x"ee",
          5697 => x"d1",
          5698 => x"38",
          5699 => x"84",
          5700 => x"8b",
          5701 => x"0d",
          5702 => x"ff",
          5703 => x"91",
          5704 => x"d0",
          5705 => x"f5",
          5706 => x"58",
          5707 => x"81",
          5708 => x"57",
          5709 => x"70",
          5710 => x"81",
          5711 => x"51",
          5712 => x"70",
          5713 => x"70",
          5714 => x"09",
          5715 => x"38",
          5716 => x"07",
          5717 => x"76",
          5718 => x"1b",
          5719 => x"38",
          5720 => x"24",
          5721 => x"c3",
          5722 => x"3d",
          5723 => x"94",
          5724 => x"b9",
          5725 => x"84",
          5726 => x"7a",
          5727 => x"51",
          5728 => x"55",
          5729 => x"02",
          5730 => x"58",
          5731 => x"02",
          5732 => x"06",
          5733 => x"7a",
          5734 => x"71",
          5735 => x"5b",
          5736 => x"76",
          5737 => x"0c",
          5738 => x"08",
          5739 => x"38",
          5740 => x"3d",
          5741 => x"33",
          5742 => x"79",
          5743 => x"39",
          5744 => x"84",
          5745 => x"ff",
          5746 => x"80",
          5747 => x"34",
          5748 => x"05",
          5749 => x"3f",
          5750 => x"c8",
          5751 => x"3d",
          5752 => x"dd",
          5753 => x"5b",
          5754 => x"80",
          5755 => x"52",
          5756 => x"b9",
          5757 => x"83",
          5758 => x"58",
          5759 => x"38",
          5760 => x"5f",
          5761 => x"76",
          5762 => x"51",
          5763 => x"08",
          5764 => x"59",
          5765 => x"38",
          5766 => x"9a",
          5767 => x"70",
          5768 => x"83",
          5769 => x"3d",
          5770 => x"b7",
          5771 => x"b9",
          5772 => x"7a",
          5773 => x"c8",
          5774 => x"38",
          5775 => x"9a",
          5776 => x"70",
          5777 => x"83",
          5778 => x"a4",
          5779 => x"51",
          5780 => x"08",
          5781 => x"ff",
          5782 => x"38",
          5783 => x"fd",
          5784 => x"89",
          5785 => x"57",
          5786 => x"56",
          5787 => x"57",
          5788 => x"75",
          5789 => x"2e",
          5790 => x"ff",
          5791 => x"19",
          5792 => x"33",
          5793 => x"80",
          5794 => x"7e",
          5795 => x"fd",
          5796 => x"38",
          5797 => x"10",
          5798 => x"70",
          5799 => x"7a",
          5800 => x"70",
          5801 => x"82",
          5802 => x"80",
          5803 => x"16",
          5804 => x"5e",
          5805 => x"ee",
          5806 => x"34",
          5807 => x"df",
          5808 => x"84",
          5809 => x"04",
          5810 => x"98",
          5811 => x"59",
          5812 => x"33",
          5813 => x"90",
          5814 => x"0c",
          5815 => x"a0",
          5816 => x"84",
          5817 => x"38",
          5818 => x"08",
          5819 => x"33",
          5820 => x"59",
          5821 => x"84",
          5822 => x"16",
          5823 => x"c8",
          5824 => x"27",
          5825 => x"74",
          5826 => x"38",
          5827 => x"08",
          5828 => x"51",
          5829 => x"dd",
          5830 => x"11",
          5831 => x"84",
          5832 => x"e5",
          5833 => x"59",
          5834 => x"81",
          5835 => x"80",
          5836 => x"5a",
          5837 => x"34",
          5838 => x"e5",
          5839 => x"79",
          5840 => x"7f",
          5841 => x"82",
          5842 => x"c8",
          5843 => x"3d",
          5844 => x"74",
          5845 => x"73",
          5846 => x"72",
          5847 => x"84",
          5848 => x"83",
          5849 => x"53",
          5850 => x"53",
          5851 => x"56",
          5852 => x"15",
          5853 => x"81",
          5854 => x"89",
          5855 => x"81",
          5856 => x"fd",
          5857 => x"ff",
          5858 => x"fd",
          5859 => x"73",
          5860 => x"06",
          5861 => x"98",
          5862 => x"2e",
          5863 => x"d9",
          5864 => x"17",
          5865 => x"81",
          5866 => x"80",
          5867 => x"51",
          5868 => x"08",
          5869 => x"81",
          5870 => x"81",
          5871 => x"73",
          5872 => x"73",
          5873 => x"0b",
          5874 => x"b9",
          5875 => x"15",
          5876 => x"58",
          5877 => x"08",
          5878 => x"09",
          5879 => x"16",
          5880 => x"27",
          5881 => x"15",
          5882 => x"16",
          5883 => x"80",
          5884 => x"2e",
          5885 => x"0b",
          5886 => x"04",
          5887 => x"08",
          5888 => x"73",
          5889 => x"c2",
          5890 => x"08",
          5891 => x"0c",
          5892 => x"2e",
          5893 => x"08",
          5894 => x"27",
          5895 => x"71",
          5896 => x"2a",
          5897 => x"80",
          5898 => x"e9",
          5899 => x"b7",
          5900 => x"8a",
          5901 => x"a2",
          5902 => x"53",
          5903 => x"54",
          5904 => x"51",
          5905 => x"08",
          5906 => x"98",
          5907 => x"fd",
          5908 => x"16",
          5909 => x"39",
          5910 => x"84",
          5911 => x"f6",
          5912 => x"80",
          5913 => x"fc",
          5914 => x"c5",
          5915 => x"84",
          5916 => x"80",
          5917 => x"c8",
          5918 => x"0c",
          5919 => x"3f",
          5920 => x"c8",
          5921 => x"70",
          5922 => x"af",
          5923 => x"81",
          5924 => x"c5",
          5925 => x"9a",
          5926 => x"70",
          5927 => x"83",
          5928 => x"7a",
          5929 => x"74",
          5930 => x"84",
          5931 => x"8d",
          5932 => x"80",
          5933 => x"80",
          5934 => x"33",
          5935 => x"90",
          5936 => x"5a",
          5937 => x"78",
          5938 => x"38",
          5939 => x"38",
          5940 => x"38",
          5941 => x"52",
          5942 => x"71",
          5943 => x"73",
          5944 => x"04",
          5945 => x"3f",
          5946 => x"71",
          5947 => x"d7",
          5948 => x"55",
          5949 => x"74",
          5950 => x"73",
          5951 => x"86",
          5952 => x"72",
          5953 => x"72",
          5954 => x"76",
          5955 => x"74",
          5956 => x"c8",
          5957 => x"2e",
          5958 => x"38",
          5959 => x"3f",
          5960 => x"3f",
          5961 => x"30",
          5962 => x"c8",
          5963 => x"b9",
          5964 => x"77",
          5965 => x"3f",
          5966 => x"3f",
          5967 => x"30",
          5968 => x"c8",
          5969 => x"75",
          5970 => x"84",
          5971 => x"8a",
          5972 => x"fe",
          5973 => x"81",
          5974 => x"75",
          5975 => x"3d",
          5976 => x"70",
          5977 => x"3f",
          5978 => x"c8",
          5979 => x"b9",
          5980 => x"52",
          5981 => x"b9",
          5982 => x"e5",
          5983 => x"98",
          5984 => x"38",
          5985 => x"75",
          5986 => x"b9",
          5987 => x"0b",
          5988 => x"04",
          5989 => x"80",
          5990 => x"3d",
          5991 => x"08",
          5992 => x"7f",
          5993 => x"fe",
          5994 => x"57",
          5995 => x"0c",
          5996 => x"0d",
          5997 => x"5a",
          5998 => x"77",
          5999 => x"5a",
          6000 => x"81",
          6001 => x"08",
          6002 => x"33",
          6003 => x"81",
          6004 => x"17",
          6005 => x"b9",
          6006 => x"5a",
          6007 => x"7e",
          6008 => x"33",
          6009 => x"77",
          6010 => x"12",
          6011 => x"07",
          6012 => x"2b",
          6013 => x"80",
          6014 => x"63",
          6015 => x"62",
          6016 => x"52",
          6017 => x"f2",
          6018 => x"0c",
          6019 => x"84",
          6020 => x"95",
          6021 => x"08",
          6022 => x"33",
          6023 => x"5e",
          6024 => x"84",
          6025 => x"17",
          6026 => x"c8",
          6027 => x"27",
          6028 => x"74",
          6029 => x"38",
          6030 => x"08",
          6031 => x"51",
          6032 => x"97",
          6033 => x"56",
          6034 => x"3f",
          6035 => x"e8",
          6036 => x"80",
          6037 => x"70",
          6038 => x"7c",
          6039 => x"5c",
          6040 => x"7a",
          6041 => x"17",
          6042 => x"34",
          6043 => x"81",
          6044 => x"07",
          6045 => x"1d",
          6046 => x"5f",
          6047 => x"38",
          6048 => x"39",
          6049 => x"7a",
          6050 => x"07",
          6051 => x"39",
          6052 => x"3d",
          6053 => x"2e",
          6054 => x"2e",
          6055 => x"2e",
          6056 => x"22",
          6057 => x"38",
          6058 => x"38",
          6059 => x"38",
          6060 => x"06",
          6061 => x"80",
          6062 => x"8c",
          6063 => x"d5",
          6064 => x"54",
          6065 => x"08",
          6066 => x"0b",
          6067 => x"18",
          6068 => x"90",
          6069 => x"75",
          6070 => x"b9",
          6071 => x"54",
          6072 => x"52",
          6073 => x"b9",
          6074 => x"80",
          6075 => x"08",
          6076 => x"c8",
          6077 => x"53",
          6078 => x"3f",
          6079 => x"9c",
          6080 => x"57",
          6081 => x"38",
          6082 => x"33",
          6083 => x"78",
          6084 => x"9c",
          6085 => x"e2",
          6086 => x"54",
          6087 => x"55",
          6088 => x"18",
          6089 => x"88",
          6090 => x"08",
          6091 => x"84",
          6092 => x"38",
          6093 => x"be",
          6094 => x"84",
          6095 => x"81",
          6096 => x"18",
          6097 => x"0b",
          6098 => x"38",
          6099 => x"27",
          6100 => x"38",
          6101 => x"83",
          6102 => x"84",
          6103 => x"52",
          6104 => x"b9",
          6105 => x"80",
          6106 => x"08",
          6107 => x"c8",
          6108 => x"53",
          6109 => x"3f",
          6110 => x"9c",
          6111 => x"57",
          6112 => x"81",
          6113 => x"81",
          6114 => x"54",
          6115 => x"55",
          6116 => x"f3",
          6117 => x"0b",
          6118 => x"39",
          6119 => x"18",
          6120 => x"b9",
          6121 => x"fd",
          6122 => x"59",
          6123 => x"08",
          6124 => x"39",
          6125 => x"ff",
          6126 => x"b7",
          6127 => x"84",
          6128 => x"75",
          6129 => x"04",
          6130 => x"3d",
          6131 => x"84",
          6132 => x"08",
          6133 => x"70",
          6134 => x"56",
          6135 => x"80",
          6136 => x"05",
          6137 => x"56",
          6138 => x"08",
          6139 => x"88",
          6140 => x"57",
          6141 => x"76",
          6142 => x"2e",
          6143 => x"08",
          6144 => x"7a",
          6145 => x"3d",
          6146 => x"84",
          6147 => x"08",
          6148 => x"52",
          6149 => x"b9",
          6150 => x"a0",
          6151 => x"a7",
          6152 => x"17",
          6153 => x"07",
          6154 => x"39",
          6155 => x"38",
          6156 => x"78",
          6157 => x"57",
          6158 => x"52",
          6159 => x"b9",
          6160 => x"80",
          6161 => x"07",
          6162 => x"9a",
          6163 => x"79",
          6164 => x"38",
          6165 => x"38",
          6166 => x"51",
          6167 => x"08",
          6168 => x"04",
          6169 => x"80",
          6170 => x"b9",
          6171 => x"74",
          6172 => x"38",
          6173 => x"81",
          6174 => x"84",
          6175 => x"ff",
          6176 => x"77",
          6177 => x"58",
          6178 => x"34",
          6179 => x"38",
          6180 => x"3f",
          6181 => x"c8",
          6182 => x"84",
          6183 => x"82",
          6184 => x"17",
          6185 => x"51",
          6186 => x"b9",
          6187 => x"ff",
          6188 => x"18",
          6189 => x"31",
          6190 => x"a0",
          6191 => x"17",
          6192 => x"06",
          6193 => x"08",
          6194 => x"81",
          6195 => x"79",
          6196 => x"78",
          6197 => x"51",
          6198 => x"08",
          6199 => x"80",
          6200 => x"2e",
          6201 => x"ff",
          6202 => x"52",
          6203 => x"b9",
          6204 => x"fe",
          6205 => x"75",
          6206 => x"94",
          6207 => x"5c",
          6208 => x"7a",
          6209 => x"a2",
          6210 => x"b9",
          6211 => x"56",
          6212 => x"53",
          6213 => x"3d",
          6214 => x"c8",
          6215 => x"2e",
          6216 => x"9f",
          6217 => x"93",
          6218 => x"3f",
          6219 => x"c8",
          6220 => x"c8",
          6221 => x"c8",
          6222 => x"38",
          6223 => x"2a",
          6224 => x"ff",
          6225 => x"3d",
          6226 => x"84",
          6227 => x"b9",
          6228 => x"b9",
          6229 => x"84",
          6230 => x"38",
          6231 => x"c8",
          6232 => x"7a",
          6233 => x"08",
          6234 => x"79",
          6235 => x"71",
          6236 => x"7a",
          6237 => x"80",
          6238 => x"05",
          6239 => x"38",
          6240 => x"75",
          6241 => x"1b",
          6242 => x"fe",
          6243 => x"81",
          6244 => x"82",
          6245 => x"17",
          6246 => x"18",
          6247 => x"81",
          6248 => x"84",
          6249 => x"17",
          6250 => x"a0",
          6251 => x"17",
          6252 => x"06",
          6253 => x"08",
          6254 => x"81",
          6255 => x"fe",
          6256 => x"58",
          6257 => x"7b",
          6258 => x"74",
          6259 => x"84",
          6260 => x"08",
          6261 => x"c8",
          6262 => x"b9",
          6263 => x"80",
          6264 => x"b0",
          6265 => x"38",
          6266 => x"08",
          6267 => x"38",
          6268 => x"33",
          6269 => x"79",
          6270 => x"75",
          6271 => x"04",
          6272 => x"ff",
          6273 => x"09",
          6274 => x"b8",
          6275 => x"05",
          6276 => x"38",
          6277 => x"7d",
          6278 => x"7d",
          6279 => x"80",
          6280 => x"1a",
          6281 => x"34",
          6282 => x"56",
          6283 => x"2a",
          6284 => x"33",
          6285 => x"7d",
          6286 => x"1b",
          6287 => x"56",
          6288 => x"ff",
          6289 => x"ae",
          6290 => x"71",
          6291 => x"78",
          6292 => x"5b",
          6293 => x"55",
          6294 => x"5b",
          6295 => x"ff",
          6296 => x"56",
          6297 => x"69",
          6298 => x"34",
          6299 => x"a1",
          6300 => x"99",
          6301 => x"9a",
          6302 => x"9b",
          6303 => x"2e",
          6304 => x"8b",
          6305 => x"18",
          6306 => x"84",
          6307 => x"c8",
          6308 => x"2a",
          6309 => x"88",
          6310 => x"fe",
          6311 => x"80",
          6312 => x"74",
          6313 => x"0b",
          6314 => x"56",
          6315 => x"77",
          6316 => x"7b",
          6317 => x"8b",
          6318 => x"18",
          6319 => x"84",
          6320 => x"d1",
          6321 => x"70",
          6322 => x"38",
          6323 => x"9f",
          6324 => x"b8",
          6325 => x"81",
          6326 => x"fc",
          6327 => x"b4",
          6328 => x"b9",
          6329 => x"84",
          6330 => x"7f",
          6331 => x"a5",
          6332 => x"3f",
          6333 => x"c8",
          6334 => x"33",
          6335 => x"ce",
          6336 => x"08",
          6337 => x"57",
          6338 => x"ff",
          6339 => x"58",
          6340 => x"70",
          6341 => x"05",
          6342 => x"38",
          6343 => x"9e",
          6344 => x"84",
          6345 => x"a8",
          6346 => x"0b",
          6347 => x"04",
          6348 => x"06",
          6349 => x"38",
          6350 => x"05",
          6351 => x"38",
          6352 => x"08",
          6353 => x"70",
          6354 => x"05",
          6355 => x"56",
          6356 => x"70",
          6357 => x"17",
          6358 => x"17",
          6359 => x"30",
          6360 => x"2e",
          6361 => x"be",
          6362 => x"72",
          6363 => x"55",
          6364 => x"84",
          6365 => x"c2",
          6366 => x"96",
          6367 => x"79",
          6368 => x"fc",
          6369 => x"e4",
          6370 => x"b9",
          6371 => x"39",
          6372 => x"06",
          6373 => x"a8",
          6374 => x"b9",
          6375 => x"93",
          6376 => x"cd",
          6377 => x"05",
          6378 => x"34",
          6379 => x"80",
          6380 => x"18",
          6381 => x"56",
          6382 => x"76",
          6383 => x"83",
          6384 => x"2a",
          6385 => x"81",
          6386 => x"81",
          6387 => x"1a",
          6388 => x"41",
          6389 => x"e0",
          6390 => x"05",
          6391 => x"38",
          6392 => x"19",
          6393 => x"82",
          6394 => x"17",
          6395 => x"33",
          6396 => x"75",
          6397 => x"51",
          6398 => x"08",
          6399 => x"5c",
          6400 => x"80",
          6401 => x"38",
          6402 => x"09",
          6403 => x"ff",
          6404 => x"18",
          6405 => x"f3",
          6406 => x"2e",
          6407 => x"2a",
          6408 => x"88",
          6409 => x"7f",
          6410 => x"08",
          6411 => x"5c",
          6412 => x"52",
          6413 => x"b9",
          6414 => x"80",
          6415 => x"08",
          6416 => x"2e",
          6417 => x"5f",
          6418 => x"a8",
          6419 => x"52",
          6420 => x"3f",
          6421 => x"38",
          6422 => x"0c",
          6423 => x"08",
          6424 => x"17",
          6425 => x"38",
          6426 => x"3f",
          6427 => x"c8",
          6428 => x"56",
          6429 => x"56",
          6430 => x"e5",
          6431 => x"b9",
          6432 => x"0b",
          6433 => x"04",
          6434 => x"98",
          6435 => x"58",
          6436 => x"c8",
          6437 => x"b9",
          6438 => x"75",
          6439 => x"04",
          6440 => x"52",
          6441 => x"3f",
          6442 => x"2e",
          6443 => x"b9",
          6444 => x"08",
          6445 => x"08",
          6446 => x"fe",
          6447 => x"82",
          6448 => x"81",
          6449 => x"05",
          6450 => x"fe",
          6451 => x"39",
          6452 => x"17",
          6453 => x"fe",
          6454 => x"c8",
          6455 => x"08",
          6456 => x"18",
          6457 => x"55",
          6458 => x"38",
          6459 => x"09",
          6460 => x"b4",
          6461 => x"7a",
          6462 => x"eb",
          6463 => x"3d",
          6464 => x"84",
          6465 => x"82",
          6466 => x"3d",
          6467 => x"c8",
          6468 => x"2e",
          6469 => x"96",
          6470 => x"96",
          6471 => x"3f",
          6472 => x"c8",
          6473 => x"33",
          6474 => x"d2",
          6475 => x"8b",
          6476 => x"07",
          6477 => x"34",
          6478 => x"78",
          6479 => x"c8",
          6480 => x"0d",
          6481 => x"53",
          6482 => x"51",
          6483 => x"08",
          6484 => x"8a",
          6485 => x"3d",
          6486 => x"3d",
          6487 => x"84",
          6488 => x"08",
          6489 => x"81",
          6490 => x"38",
          6491 => x"71",
          6492 => x"96",
          6493 => x"97",
          6494 => x"98",
          6495 => x"99",
          6496 => x"18",
          6497 => x"84",
          6498 => x"96",
          6499 => x"6d",
          6500 => x"05",
          6501 => x"3f",
          6502 => x"08",
          6503 => x"80",
          6504 => x"8b",
          6505 => x"78",
          6506 => x"07",
          6507 => x"81",
          6508 => x"58",
          6509 => x"a4",
          6510 => x"16",
          6511 => x"16",
          6512 => x"09",
          6513 => x"76",
          6514 => x"51",
          6515 => x"08",
          6516 => x"59",
          6517 => x"bd",
          6518 => x"c3",
          6519 => x"e4",
          6520 => x"56",
          6521 => x"82",
          6522 => x"2b",
          6523 => x"88",
          6524 => x"5f",
          6525 => x"b9",
          6526 => x"5e",
          6527 => x"52",
          6528 => x"c8",
          6529 => x"2e",
          6530 => x"81",
          6531 => x"80",
          6532 => x"16",
          6533 => x"17",
          6534 => x"77",
          6535 => x"09",
          6536 => x"c8",
          6537 => x"a8",
          6538 => x"5a",
          6539 => x"ad",
          6540 => x"2e",
          6541 => x"54",
          6542 => x"53",
          6543 => x"db",
          6544 => x"53",
          6545 => x"fe",
          6546 => x"80",
          6547 => x"75",
          6548 => x"84",
          6549 => x"08",
          6550 => x"84",
          6551 => x"79",
          6552 => x"56",
          6553 => x"8a",
          6554 => x"57",
          6555 => x"fc",
          6556 => x"33",
          6557 => x"38",
          6558 => x"39",
          6559 => x"ff",
          6560 => x"9c",
          6561 => x"84",
          6562 => x"3d",
          6563 => x"70",
          6564 => x"74",
          6565 => x"33",
          6566 => x"5a",
          6567 => x"3d",
          6568 => x"06",
          6569 => x"38",
          6570 => x"26",
          6571 => x"3f",
          6572 => x"51",
          6573 => x"83",
          6574 => x"81",
          6575 => x"e6",
          6576 => x"56",
          6577 => x"74",
          6578 => x"18",
          6579 => x"57",
          6580 => x"77",
          6581 => x"81",
          6582 => x"81",
          6583 => x"89",
          6584 => x"27",
          6585 => x"7b",
          6586 => x"5a",
          6587 => x"81",
          6588 => x"81",
          6589 => x"9f",
          6590 => x"57",
          6591 => x"38",
          6592 => x"05",
          6593 => x"7a",
          6594 => x"ff",
          6595 => x"80",
          6596 => x"56",
          6597 => x"08",
          6598 => x"b4",
          6599 => x"0c",
          6600 => x"74",
          6601 => x"08",
          6602 => x"f8",
          6603 => x"0c",
          6604 => x"33",
          6605 => x"51",
          6606 => x"08",
          6607 => x"38",
          6608 => x"6c",
          6609 => x"05",
          6610 => x"34",
          6611 => x"5d",
          6612 => x"fe",
          6613 => x"55",
          6614 => x"27",
          6615 => x"39",
          6616 => x"81",
          6617 => x"75",
          6618 => x"53",
          6619 => x"84",
          6620 => x"08",
          6621 => x"38",
          6622 => x"5a",
          6623 => x"18",
          6624 => x"33",
          6625 => x"81",
          6626 => x"18",
          6627 => x"c4",
          6628 => x"85",
          6629 => x"19",
          6630 => x"9c",
          6631 => x"74",
          6632 => x"30",
          6633 => x"74",
          6634 => x"5a",
          6635 => x"75",
          6636 => x"c8",
          6637 => x"2e",
          6638 => x"2e",
          6639 => x"b9",
          6640 => x"70",
          6641 => x"74",
          6642 => x"17",
          6643 => x"76",
          6644 => x"81",
          6645 => x"80",
          6646 => x"05",
          6647 => x"34",
          6648 => x"d6",
          6649 => x"5d",
          6650 => x"fe",
          6651 => x"55",
          6652 => x"39",
          6653 => x"52",
          6654 => x"3f",
          6655 => x"81",
          6656 => x"08",
          6657 => x"19",
          6658 => x"27",
          6659 => x"82",
          6660 => x"59",
          6661 => x"75",
          6662 => x"c8",
          6663 => x"2e",
          6664 => x"70",
          6665 => x"38",
          6666 => x"08",
          6667 => x"81",
          6668 => x"fd",
          6669 => x"02",
          6670 => x"5b",
          6671 => x"38",
          6672 => x"38",
          6673 => x"38",
          6674 => x"59",
          6675 => x"54",
          6676 => x"17",
          6677 => x"80",
          6678 => x"81",
          6679 => x"2a",
          6680 => x"81",
          6681 => x"89",
          6682 => x"59",
          6683 => x"06",
          6684 => x"84",
          6685 => x"79",
          6686 => x"27",
          6687 => x"83",
          6688 => x"80",
          6689 => x"87",
          6690 => x"14",
          6691 => x"84",
          6692 => x"38",
          6693 => x"d8",
          6694 => x"38",
          6695 => x"38",
          6696 => x"38",
          6697 => x"c8",
          6698 => x"84",
          6699 => x"81",
          6700 => x"84",
          6701 => x"fe",
          6702 => x"fe",
          6703 => x"38",
          6704 => x"ab",
          6705 => x"80",
          6706 => x"51",
          6707 => x"08",
          6708 => x"38",
          6709 => x"5e",
          6710 => x"0c",
          6711 => x"7a",
          6712 => x"90",
          6713 => x"90",
          6714 => x"94",
          6715 => x"fe",
          6716 => x"0c",
          6717 => x"84",
          6718 => x"ff",
          6719 => x"59",
          6720 => x"39",
          6721 => x"5e",
          6722 => x"e3",
          6723 => x"08",
          6724 => x"44",
          6725 => x"70",
          6726 => x"8a",
          6727 => x"70",
          6728 => x"85",
          6729 => x"2e",
          6730 => x"56",
          6731 => x"10",
          6732 => x"56",
          6733 => x"75",
          6734 => x"33",
          6735 => x"5d",
          6736 => x"3f",
          6737 => x"70",
          6738 => x"84",
          6739 => x"40",
          6740 => x"3d",
          6741 => x"fe",
          6742 => x"84",
          6743 => x"84",
          6744 => x"84",
          6745 => x"74",
          6746 => x"38",
          6747 => x"7e",
          6748 => x"ff",
          6749 => x"38",
          6750 => x"2a",
          6751 => x"5b",
          6752 => x"30",
          6753 => x"91",
          6754 => x"2e",
          6755 => x"60",
          6756 => x"81",
          6757 => x"38",
          6758 => x"fe",
          6759 => x"56",
          6760 => x"09",
          6761 => x"29",
          6762 => x"58",
          6763 => x"b6",
          6764 => x"71",
          6765 => x"14",
          6766 => x"33",
          6767 => x"33",
          6768 => x"88",
          6769 => x"07",
          6770 => x"a2",
          6771 => x"3d",
          6772 => x"41",
          6773 => x"ff",
          6774 => x"7a",
          6775 => x"81",
          6776 => x"80",
          6777 => x"45",
          6778 => x"06",
          6779 => x"70",
          6780 => x"83",
          6781 => x"78",
          6782 => x"ec",
          6783 => x"38",
          6784 => x"ec",
          6785 => x"57",
          6786 => x"76",
          6787 => x"51",
          6788 => x"08",
          6789 => x"08",
          6790 => x"84",
          6791 => x"08",
          6792 => x"57",
          6793 => x"5d",
          6794 => x"11",
          6795 => x"6b",
          6796 => x"62",
          6797 => x"5d",
          6798 => x"56",
          6799 => x"78",
          6800 => x"68",
          6801 => x"84",
          6802 => x"89",
          6803 => x"06",
          6804 => x"84",
          6805 => x"7a",
          6806 => x"80",
          6807 => x"fe",
          6808 => x"c8",
          6809 => x"0c",
          6810 => x"0b",
          6811 => x"84",
          6812 => x"11",
          6813 => x"74",
          6814 => x"81",
          6815 => x"7a",
          6816 => x"e5",
          6817 => x"5b",
          6818 => x"70",
          6819 => x"45",
          6820 => x"e0",
          6821 => x"ff",
          6822 => x"38",
          6823 => x"46",
          6824 => x"76",
          6825 => x"78",
          6826 => x"30",
          6827 => x"5d",
          6828 => x"38",
          6829 => x"7c",
          6830 => x"e0",
          6831 => x"52",
          6832 => x"57",
          6833 => x"61",
          6834 => x"08",
          6835 => x"6c",
          6836 => x"9c",
          6837 => x"39",
          6838 => x"24",
          6839 => x"0c",
          6840 => x"48",
          6841 => x"38",
          6842 => x"fc",
          6843 => x"f5",
          6844 => x"18",
          6845 => x"38",
          6846 => x"9f",
          6847 => x"80",
          6848 => x"9f",
          6849 => x"06",
          6850 => x"84",
          6851 => x"81",
          6852 => x"f4",
          6853 => x"57",
          6854 => x"76",
          6855 => x"55",
          6856 => x"74",
          6857 => x"77",
          6858 => x"ff",
          6859 => x"6a",
          6860 => x"34",
          6861 => x"32",
          6862 => x"05",
          6863 => x"68",
          6864 => x"83",
          6865 => x"83",
          6866 => x"05",
          6867 => x"94",
          6868 => x"bf",
          6869 => x"05",
          6870 => x"61",
          6871 => x"34",
          6872 => x"05",
          6873 => x"9e",
          6874 => x"d4",
          6875 => x"05",
          6876 => x"80",
          6877 => x"05",
          6878 => x"cc",
          6879 => x"ff",
          6880 => x"74",
          6881 => x"34",
          6882 => x"61",
          6883 => x"83",
          6884 => x"81",
          6885 => x"58",
          6886 => x"60",
          6887 => x"34",
          6888 => x"6b",
          6889 => x"79",
          6890 => x"84",
          6891 => x"17",
          6892 => x"69",
          6893 => x"05",
          6894 => x"38",
          6895 => x"86",
          6896 => x"62",
          6897 => x"61",
          6898 => x"74",
          6899 => x"90",
          6900 => x"46",
          6901 => x"34",
          6902 => x"83",
          6903 => x"60",
          6904 => x"84",
          6905 => x"80",
          6906 => x"05",
          6907 => x"38",
          6908 => x"76",
          6909 => x"80",
          6910 => x"83",
          6911 => x"75",
          6912 => x"54",
          6913 => x"c4",
          6914 => x"9b",
          6915 => x"5b",
          6916 => x"2e",
          6917 => x"ff",
          6918 => x"2e",
          6919 => x"38",
          6920 => x"81",
          6921 => x"80",
          6922 => x"19",
          6923 => x"34",
          6924 => x"05",
          6925 => x"05",
          6926 => x"67",
          6927 => x"34",
          6928 => x"1f",
          6929 => x"85",
          6930 => x"2a",
          6931 => x"34",
          6932 => x"34",
          6933 => x"61",
          6934 => x"c8",
          6935 => x"83",
          6936 => x"05",
          6937 => x"83",
          6938 => x"77",
          6939 => x"2a",
          6940 => x"81",
          6941 => x"fe",
          6942 => x"c8",
          6943 => x"52",
          6944 => x"57",
          6945 => x"84",
          6946 => x"9f",
          6947 => x"62",
          6948 => x"16",
          6949 => x"38",
          6950 => x"e6",
          6951 => x"9d",
          6952 => x"e6",
          6953 => x"22",
          6954 => x"38",
          6955 => x"78",
          6956 => x"c8",
          6957 => x"89",
          6958 => x"84",
          6959 => x"58",
          6960 => x"f5",
          6961 => x"84",
          6962 => x"f8",
          6963 => x"81",
          6964 => x"57",
          6965 => x"63",
          6966 => x"f4",
          6967 => x"75",
          6968 => x"34",
          6969 => x"05",
          6970 => x"a3",
          6971 => x"80",
          6972 => x"05",
          6973 => x"80",
          6974 => x"61",
          6975 => x"7b",
          6976 => x"59",
          6977 => x"2a",
          6978 => x"61",
          6979 => x"34",
          6980 => x"af",
          6981 => x"80",
          6982 => x"05",
          6983 => x"80",
          6984 => x"80",
          6985 => x"05",
          6986 => x"70",
          6987 => x"05",
          6988 => x"2e",
          6989 => x"58",
          6990 => x"ff",
          6991 => x"39",
          6992 => x"51",
          6993 => x"b9",
          6994 => x"29",
          6995 => x"05",
          6996 => x"53",
          6997 => x"3f",
          6998 => x"c8",
          6999 => x"0c",
          7000 => x"6a",
          7001 => x"70",
          7002 => x"ff",
          7003 => x"05",
          7004 => x"61",
          7005 => x"34",
          7006 => x"8a",
          7007 => x"f9",
          7008 => x"60",
          7009 => x"84",
          7010 => x"81",
          7011 => x"f4",
          7012 => x"81",
          7013 => x"75",
          7014 => x"75",
          7015 => x"75",
          7016 => x"34",
          7017 => x"80",
          7018 => x"e1",
          7019 => x"05",
          7020 => x"7a",
          7021 => x"05",
          7022 => x"83",
          7023 => x"7f",
          7024 => x"83",
          7025 => x"05",
          7026 => x"76",
          7027 => x"69",
          7028 => x"87",
          7029 => x"bd",
          7030 => x"60",
          7031 => x"69",
          7032 => x"3d",
          7033 => x"61",
          7034 => x"25",
          7035 => x"f8",
          7036 => x"51",
          7037 => x"09",
          7038 => x"55",
          7039 => x"70",
          7040 => x"74",
          7041 => x"cd",
          7042 => x"83",
          7043 => x"0c",
          7044 => x"7b",
          7045 => x"57",
          7046 => x"17",
          7047 => x"88",
          7048 => x"59",
          7049 => x"bb",
          7050 => x"81",
          7051 => x"04",
          7052 => x"8c",
          7053 => x"d1",
          7054 => x"72",
          7055 => x"0c",
          7056 => x"56",
          7057 => x"94",
          7058 => x"02",
          7059 => x"58",
          7060 => x"70",
          7061 => x"74",
          7062 => x"77",
          7063 => x"80",
          7064 => x"17",
          7065 => x"81",
          7066 => x"74",
          7067 => x"0c",
          7068 => x"9f",
          7069 => x"c0",
          7070 => x"c9",
          7071 => x"7c",
          7072 => x"b9",
          7073 => x"3d",
          7074 => x"05",
          7075 => x"3f",
          7076 => x"07",
          7077 => x"56",
          7078 => x"fd",
          7079 => x"b9",
          7080 => x"3d",
          7081 => x"22",
          7082 => x"26",
          7083 => x"52",
          7084 => x"0d",
          7085 => x"70",
          7086 => x"38",
          7087 => x"8c",
          7088 => x"81",
          7089 => x"54",
          7090 => x"10",
          7091 => x"51",
          7092 => x"ff",
          7093 => x"3d",
          7094 => x"05",
          7095 => x"53",
          7096 => x"8c",
          7097 => x"0c",
          7098 => x"2e",
          7099 => x"ff",
          7100 => x"8c",
          7101 => x"51",
          7102 => x"77",
          7103 => x"e1",
          7104 => x"e9",
          7105 => x"80",
          7106 => x"22",
          7107 => x"7a",
          7108 => x"b7",
          7109 => x"72",
          7110 => x"06",
          7111 => x"b1",
          7112 => x"70",
          7113 => x"30",
          7114 => x"53",
          7115 => x"75",
          7116 => x"3d",
          7117 => x"a2",
          7118 => x"10",
          7119 => x"08",
          7120 => x"ff",
          7121 => x"ff",
          7122 => x"57",
          7123 => x"ff",
          7124 => x"16",
          7125 => x"db",
          7126 => x"06",
          7127 => x"83",
          7128 => x"f0",
          7129 => x"51",
          7130 => x"06",
          7131 => x"06",
          7132 => x"73",
          7133 => x"52",
          7134 => x"ff",
          7135 => x"00",
          7136 => x"19",
          7137 => x"19",
          7138 => x"19",
          7139 => x"19",
          7140 => x"19",
          7141 => x"19",
          7142 => x"19",
          7143 => x"18",
          7144 => x"18",
          7145 => x"18",
          7146 => x"1e",
          7147 => x"1f",
          7148 => x"1f",
          7149 => x"1f",
          7150 => x"1f",
          7151 => x"1f",
          7152 => x"1f",
          7153 => x"1f",
          7154 => x"1f",
          7155 => x"1f",
          7156 => x"1f",
          7157 => x"1f",
          7158 => x"1f",
          7159 => x"1f",
          7160 => x"1f",
          7161 => x"1f",
          7162 => x"1f",
          7163 => x"1f",
          7164 => x"1f",
          7165 => x"1f",
          7166 => x"1f",
          7167 => x"1f",
          7168 => x"1f",
          7169 => x"1f",
          7170 => x"1f",
          7171 => x"1f",
          7172 => x"1f",
          7173 => x"1f",
          7174 => x"1f",
          7175 => x"1f",
          7176 => x"24",
          7177 => x"1f",
          7178 => x"24",
          7179 => x"22",
          7180 => x"1f",
          7181 => x"1f",
          7182 => x"1f",
          7183 => x"1f",
          7184 => x"1f",
          7185 => x"1f",
          7186 => x"1f",
          7187 => x"1f",
          7188 => x"1f",
          7189 => x"1f",
          7190 => x"1f",
          7191 => x"1f",
          7192 => x"1f",
          7193 => x"1f",
          7194 => x"1f",
          7195 => x"1f",
          7196 => x"1f",
          7197 => x"1f",
          7198 => x"1f",
          7199 => x"1f",
          7200 => x"1f",
          7201 => x"1f",
          7202 => x"1f",
          7203 => x"1f",
          7204 => x"1f",
          7205 => x"1f",
          7206 => x"21",
          7207 => x"1f",
          7208 => x"1f",
          7209 => x"1f",
          7210 => x"1f",
          7211 => x"21",
          7212 => x"1f",
          7213 => x"1f",
          7214 => x"21",
          7215 => x"32",
          7216 => x"32",
          7217 => x"32",
          7218 => x"3b",
          7219 => x"39",
          7220 => x"3a",
          7221 => x"37",
          7222 => x"39",
          7223 => x"37",
          7224 => x"34",
          7225 => x"38",
          7226 => x"34",
          7227 => x"37",
          7228 => x"36",
          7229 => x"46",
          7230 => x"46",
          7231 => x"46",
          7232 => x"46",
          7233 => x"47",
          7234 => x"47",
          7235 => x"47",
          7236 => x"47",
          7237 => x"47",
          7238 => x"47",
          7239 => x"47",
          7240 => x"47",
          7241 => x"47",
          7242 => x"47",
          7243 => x"47",
          7244 => x"47",
          7245 => x"47",
          7246 => x"47",
          7247 => x"47",
          7248 => x"48",
          7249 => x"48",
          7250 => x"48",
          7251 => x"47",
          7252 => x"47",
          7253 => x"48",
          7254 => x"47",
          7255 => x"47",
          7256 => x"47",
          7257 => x"47",
          7258 => x"55",
          7259 => x"54",
          7260 => x"54",
          7261 => x"56",
          7262 => x"55",
          7263 => x"52",
          7264 => x"52",
          7265 => x"52",
          7266 => x"55",
          7267 => x"56",
          7268 => x"52",
          7269 => x"52",
          7270 => x"52",
          7271 => x"52",
          7272 => x"52",
          7273 => x"52",
          7274 => x"52",
          7275 => x"52",
          7276 => x"52",
          7277 => x"55",
          7278 => x"52",
          7279 => x"54",
          7280 => x"53",
          7281 => x"52",
          7282 => x"52",
          7283 => x"52",
          7284 => x"59",
          7285 => x"59",
          7286 => x"59",
          7287 => x"59",
          7288 => x"59",
          7289 => x"59",
          7290 => x"59",
          7291 => x"59",
          7292 => x"59",
          7293 => x"59",
          7294 => x"59",
          7295 => x"59",
          7296 => x"59",
          7297 => x"59",
          7298 => x"59",
          7299 => x"59",
          7300 => x"59",
          7301 => x"59",
          7302 => x"5a",
          7303 => x"59",
          7304 => x"5a",
          7305 => x"5a",
          7306 => x"59",
          7307 => x"59",
          7308 => x"59",
          7309 => x"63",
          7310 => x"61",
          7311 => x"61",
          7312 => x"61",
          7313 => x"61",
          7314 => x"61",
          7315 => x"61",
          7316 => x"5e",
          7317 => x"61",
          7318 => x"61",
          7319 => x"61",
          7320 => x"61",
          7321 => x"63",
          7322 => x"63",
          7323 => x"63",
          7324 => x"de",
          7325 => x"de",
          7326 => x"de",
          7327 => x"de",
          7328 => x"0e",
          7329 => x"0b",
          7330 => x"0b",
          7331 => x"0b",
          7332 => x"0b",
          7333 => x"0b",
          7334 => x"0b",
          7335 => x"0f",
          7336 => x"0b",
          7337 => x"0b",
          7338 => x"0b",
          7339 => x"0b",
          7340 => x"0b",
          7341 => x"0b",
          7342 => x"0b",
          7343 => x"0b",
          7344 => x"0b",
          7345 => x"0b",
          7346 => x"0b",
          7347 => x"0b",
          7348 => x"0b",
          7349 => x"0b",
          7350 => x"0b",
          7351 => x"0b",
          7352 => x"0b",
          7353 => x"0b",
          7354 => x"0b",
          7355 => x"0b",
          7356 => x"0e",
          7357 => x"0b",
          7358 => x"0b",
          7359 => x"0b",
          7360 => x"0b",
          7361 => x"0b",
          7362 => x"0e",
          7363 => x"0e",
          7364 => x"0b",
          7365 => x"0b",
          7366 => x"0e",
          7367 => x"0b",
          7368 => x"0e",
          7369 => x"0b",
          7370 => x"0b",
          7371 => x"0b",
          7372 => x"0e",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"68",
          7383 => x"64",
          7384 => x"64",
          7385 => x"6c",
          7386 => x"70",
          7387 => x"74",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"30",
          7392 => x"00",
          7393 => x"00",
          7394 => x"00",
          7395 => x"6b",
          7396 => x"72",
          7397 => x"72",
          7398 => x"20",
          7399 => x"63",
          7400 => x"6f",
          7401 => x"70",
          7402 => x"73",
          7403 => x"73",
          7404 => x"6e",
          7405 => x"79",
          7406 => x"6c",
          7407 => x"63",
          7408 => x"6d",
          7409 => x"70",
          7410 => x"20",
          7411 => x"65",
          7412 => x"72",
          7413 => x"72",
          7414 => x"20",
          7415 => x"62",
          7416 => x"73",
          7417 => x"6f",
          7418 => x"64",
          7419 => x"73",
          7420 => x"6e",
          7421 => x"00",
          7422 => x"6e",
          7423 => x"73",
          7424 => x"64",
          7425 => x"20",
          7426 => x"65",
          7427 => x"74",
          7428 => x"6c",
          7429 => x"65",
          7430 => x"64",
          7431 => x"6c",
          7432 => x"64",
          7433 => x"73",
          7434 => x"63",
          7435 => x"69",
          7436 => x"76",
          7437 => x"6c",
          7438 => x"00",
          7439 => x"68",
          7440 => x"00",
          7441 => x"65",
          7442 => x"00",
          7443 => x"6f",
          7444 => x"2e",
          7445 => x"61",
          7446 => x"2e",
          7447 => x"72",
          7448 => x"63",
          7449 => x"00",
          7450 => x"79",
          7451 => x"61",
          7452 => x"79",
          7453 => x"2e",
          7454 => x"61",
          7455 => x"38",
          7456 => x"20",
          7457 => x"00",
          7458 => x"00",
          7459 => x"34",
          7460 => x"20",
          7461 => x"00",
          7462 => x"20",
          7463 => x"2f",
          7464 => x"00",
          7465 => x"00",
          7466 => x"72",
          7467 => x"29",
          7468 => x"2a",
          7469 => x"3a",
          7470 => x"73",
          7471 => x"73",
          7472 => x"20",
          7473 => x"20",
          7474 => x"00",
          7475 => x"70",
          7476 => x"73",
          7477 => x"20",
          7478 => x"20",
          7479 => x"00",
          7480 => x"74",
          7481 => x"48",
          7482 => x"00",
          7483 => x"54",
          7484 => x"72",
          7485 => x"52",
          7486 => x"6e",
          7487 => x"00",
          7488 => x"54",
          7489 => x"72",
          7490 => x"52",
          7491 => x"6e",
          7492 => x"00",
          7493 => x"57",
          7494 => x"72",
          7495 => x"43",
          7496 => x"6e",
          7497 => x"00",
          7498 => x"74",
          7499 => x"00",
          7500 => x"69",
          7501 => x"74",
          7502 => x"67",
          7503 => x"65",
          7504 => x"61",
          7505 => x"69",
          7506 => x"00",
          7507 => x"65",
          7508 => x"00",
          7509 => x"75",
          7510 => x"69",
          7511 => x"69",
          7512 => x"73",
          7513 => x"72",
          7514 => x"65",
          7515 => x"74",
          7516 => x"6c",
          7517 => x"00",
          7518 => x"00",
          7519 => x"64",
          7520 => x"64",
          7521 => x"55",
          7522 => x"3a",
          7523 => x"25",
          7524 => x"6c",
          7525 => x"74",
          7526 => x"00",
          7527 => x"74",
          7528 => x"6c",
          7529 => x"2e",
          7530 => x"6c",
          7531 => x"64",
          7532 => x"6c",
          7533 => x"00",
          7534 => x"65",
          7535 => x"63",
          7536 => x"29",
          7537 => x"65",
          7538 => x"63",
          7539 => x"30",
          7540 => x"0a",
          7541 => x"25",
          7542 => x"00",
          7543 => x"25",
          7544 => x"6d",
          7545 => x"2e",
          7546 => x"38",
          7547 => x"29",
          7548 => x"28",
          7549 => x"00",
          7550 => x"67",
          7551 => x"38",
          7552 => x"2d",
          7553 => x"6e",
          7554 => x"00",
          7555 => x"65",
          7556 => x"6f",
          7557 => x"00",
          7558 => x"5c",
          7559 => x"6d",
          7560 => x"61",
          7561 => x"63",
          7562 => x"72",
          7563 => x"6f",
          7564 => x"00",
          7565 => x"2f",
          7566 => x"64",
          7567 => x"25",
          7568 => x"43",
          7569 => x"75",
          7570 => x"00",
          7571 => x"63",
          7572 => x"65",
          7573 => x"00",
          7574 => x"73",
          7575 => x"20",
          7576 => x"73",
          7577 => x"6f",
          7578 => x"73",
          7579 => x"58",
          7580 => x"20",
          7581 => x"6d",
          7582 => x"72",
          7583 => x"73",
          7584 => x"58",
          7585 => x"20",
          7586 => x"53",
          7587 => x"64",
          7588 => x"20",
          7589 => x"58",
          7590 => x"73",
          7591 => x"20",
          7592 => x"20",
          7593 => x"20",
          7594 => x"20",
          7595 => x"58",
          7596 => x"20",
          7597 => x"20",
          7598 => x"72",
          7599 => x"20",
          7600 => x"25",
          7601 => x"00",
          7602 => x"73",
          7603 => x"44",
          7604 => x"63",
          7605 => x"20",
          7606 => x"4d",
          7607 => x"20",
          7608 => x"43",
          7609 => x"65",
          7610 => x"20",
          7611 => x"25",
          7612 => x"00",
          7613 => x"49",
          7614 => x"32",
          7615 => x"43",
          7616 => x"20",
          7617 => x"00",
          7618 => x"53",
          7619 => x"55",
          7620 => x"20",
          7621 => x"54",
          7622 => x"6e",
          7623 => x"32",
          7624 => x"20",
          7625 => x"20",
          7626 => x"65",
          7627 => x"32",
          7628 => x"20",
          7629 => x"44",
          7630 => x"69",
          7631 => x"32",
          7632 => x"20",
          7633 => x"20",
          7634 => x"58",
          7635 => x"0a",
          7636 => x"41",
          7637 => x"28",
          7638 => x"38",
          7639 => x"20",
          7640 => x"52",
          7641 => x"58",
          7642 => x"0a",
          7643 => x"52",
          7644 => x"28",
          7645 => x"38",
          7646 => x"20",
          7647 => x"41",
          7648 => x"58",
          7649 => x"0a",
          7650 => x"20",
          7651 => x"66",
          7652 => x"6b",
          7653 => x"4f",
          7654 => x"61",
          7655 => x"64",
          7656 => x"65",
          7657 => x"4f",
          7658 => x"00",
          7659 => x"f0",
          7660 => x"00",
          7661 => x"00",
          7662 => x"f0",
          7663 => x"00",
          7664 => x"00",
          7665 => x"f0",
          7666 => x"00",
          7667 => x"00",
          7668 => x"f0",
          7669 => x"00",
          7670 => x"00",
          7671 => x"f0",
          7672 => x"00",
          7673 => x"00",
          7674 => x"f0",
          7675 => x"00",
          7676 => x"00",
          7677 => x"f0",
          7678 => x"00",
          7679 => x"00",
          7680 => x"f0",
          7681 => x"00",
          7682 => x"00",
          7683 => x"f0",
          7684 => x"00",
          7685 => x"00",
          7686 => x"f0",
          7687 => x"00",
          7688 => x"00",
          7689 => x"f0",
          7690 => x"00",
          7691 => x"43",
          7692 => x"41",
          7693 => x"35",
          7694 => x"46",
          7695 => x"32",
          7696 => x"00",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"20",
          7703 => x"65",
          7704 => x"74",
          7705 => x"65",
          7706 => x"6c",
          7707 => x"73",
          7708 => x"73",
          7709 => x"00",
          7710 => x"20",
          7711 => x"69",
          7712 => x"72",
          7713 => x"65",
          7714 => x"79",
          7715 => x"6f",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"42",
          7720 => x"44",
          7721 => x"00",
          7722 => x"00",
          7723 => x"00",
          7724 => x"00",
          7725 => x"00",
          7726 => x"00",
          7727 => x"00",
          7728 => x"00",
          7729 => x"00",
          7730 => x"00",
          7731 => x"00",
          7732 => x"00",
          7733 => x"35",
          7734 => x"36",
          7735 => x"25",
          7736 => x"2c",
          7737 => x"64",
          7738 => x"00",
          7739 => x"64",
          7740 => x"25",
          7741 => x"3a",
          7742 => x"25",
          7743 => x"32",
          7744 => x"5b",
          7745 => x"00",
          7746 => x"20",
          7747 => x"00",
          7748 => x"78",
          7749 => x"00",
          7750 => x"78",
          7751 => x"00",
          7752 => x"78",
          7753 => x"20",
          7754 => x"66",
          7755 => x"00",
          7756 => x"3a",
          7757 => x"00",
          7758 => x"00",
          7759 => x"54",
          7760 => x"90",
          7761 => x"30",
          7762 => x"45",
          7763 => x"20",
          7764 => x"20",
          7765 => x"20",
          7766 => x"20",
          7767 => x"00",
          7768 => x"00",
          7769 => x"10",
          7770 => x"00",
          7771 => x"8f",
          7772 => x"8e",
          7773 => x"55",
          7774 => x"9e",
          7775 => x"a6",
          7776 => x"ae",
          7777 => x"b6",
          7778 => x"be",
          7779 => x"c6",
          7780 => x"ce",
          7781 => x"d6",
          7782 => x"de",
          7783 => x"e6",
          7784 => x"ee",
          7785 => x"f6",
          7786 => x"fe",
          7787 => x"5d",
          7788 => x"3f",
          7789 => x"00",
          7790 => x"02",
          7791 => x"00",
          7792 => x"00",
          7793 => x"00",
          7794 => x"00",
          7795 => x"00",
          7796 => x"00",
          7797 => x"00",
          7798 => x"00",
          7799 => x"00",
          7800 => x"00",
          7801 => x"00",
          7802 => x"00",
          7803 => x"23",
          7804 => x"00",
          7805 => x"25",
          7806 => x"25",
          7807 => x"25",
          7808 => x"25",
          7809 => x"25",
          7810 => x"25",
          7811 => x"25",
          7812 => x"25",
          7813 => x"25",
          7814 => x"25",
          7815 => x"25",
          7816 => x"25",
          7817 => x"00",
          7818 => x"03",
          7819 => x"03",
          7820 => x"03",
          7821 => x"00",
          7822 => x"23",
          7823 => x"22",
          7824 => x"00",
          7825 => x"03",
          7826 => x"03",
          7827 => x"01",
          7828 => x"01",
          7829 => x"01",
          7830 => x"02",
          7831 => x"01",
          7832 => x"01",
          7833 => x"01",
          7834 => x"01",
          7835 => x"01",
          7836 => x"01",
          7837 => x"01",
          7838 => x"01",
          7839 => x"01",
          7840 => x"01",
          7841 => x"01",
          7842 => x"01",
          7843 => x"01",
          7844 => x"01",
          7845 => x"01",
          7846 => x"01",
          7847 => x"01",
          7848 => x"01",
          7849 => x"01",
          7850 => x"00",
          7851 => x"01",
          7852 => x"01",
          7853 => x"01",
          7854 => x"02",
          7855 => x"02",
          7856 => x"02",
          7857 => x"01",
          7858 => x"01",
          7859 => x"01",
          7860 => x"02",
          7861 => x"01",
          7862 => x"02",
          7863 => x"2c",
          7864 => x"01",
          7865 => x"02",
          7866 => x"02",
          7867 => x"02",
          7868 => x"02",
          7869 => x"01",
          7870 => x"02",
          7871 => x"01",
          7872 => x"02",
          7873 => x"03",
          7874 => x"03",
          7875 => x"03",
          7876 => x"03",
          7877 => x"03",
          7878 => x"00",
          7879 => x"03",
          7880 => x"03",
          7881 => x"03",
          7882 => x"03",
          7883 => x"04",
          7884 => x"04",
          7885 => x"04",
          7886 => x"01",
          7887 => x"00",
          7888 => x"1e",
          7889 => x"1f",
          7890 => x"1f",
          7891 => x"1f",
          7892 => x"1f",
          7893 => x"1f",
          7894 => x"06",
          7895 => x"1f",
          7896 => x"1f",
          7897 => x"1f",
          7898 => x"1f",
          7899 => x"06",
          7900 => x"00",
          7901 => x"1f",
          7902 => x"1f",
          7903 => x"1f",
          7904 => x"00",
          7905 => x"21",
          7906 => x"00",
          7907 => x"2c",
          7908 => x"2c",
          7909 => x"2c",
          7910 => x"ff",
          7911 => x"00",
          7912 => x"01",
          7913 => x"00",
          7914 => x"01",
          7915 => x"00",
          7916 => x"03",
          7917 => x"00",
          7918 => x"03",
          7919 => x"00",
          7920 => x"03",
          7921 => x"00",
          7922 => x"04",
          7923 => x"00",
          7924 => x"04",
          7925 => x"00",
          7926 => x"04",
          7927 => x"00",
          7928 => x"04",
          7929 => x"00",
          7930 => x"04",
          7931 => x"00",
          7932 => x"04",
          7933 => x"00",
          7934 => x"04",
          7935 => x"00",
          7936 => x"05",
          7937 => x"00",
          7938 => x"05",
          7939 => x"00",
          7940 => x"05",
          7941 => x"00",
          7942 => x"05",
          7943 => x"00",
          7944 => x"07",
          7945 => x"00",
          7946 => x"07",
          7947 => x"00",
          7948 => x"08",
          7949 => x"00",
          7950 => x"08",
          7951 => x"00",
          7952 => x"08",
          7953 => x"00",
          7954 => x"08",
          7955 => x"00",
          7956 => x"08",
          7957 => x"00",
          7958 => x"08",
          7959 => x"00",
          7960 => x"09",
          7961 => x"00",
          7962 => x"09",
          7963 => x"00",
          7964 => x"09",
          7965 => x"00",
          7966 => x"09",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"78",
          7975 => x"e1",
          7976 => x"e1",
          7977 => x"01",
          7978 => x"10",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"00",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"f0",
          7992 => x"f0",
          7993 => x"f0",
          7994 => x"fd",
          7995 => x"3a",
          7996 => x"f0",
          7997 => x"77",
          7998 => x"6f",
          7999 => x"67",
          8000 => x"37",
          8001 => x"2c",
          8002 => x"3f",
          8003 => x"f0",
          8004 => x"f0",
          8005 => x"3b",
          8006 => x"f0",
          8007 => x"57",
          8008 => x"4f",
          8009 => x"47",
          8010 => x"37",
          8011 => x"2c",
          8012 => x"3f",
          8013 => x"f0",
          8014 => x"f0",
          8015 => x"2a",
          8016 => x"f0",
          8017 => x"57",
          8018 => x"4f",
          8019 => x"47",
          8020 => x"27",
          8021 => x"3c",
          8022 => x"3f",
          8023 => x"f0",
          8024 => x"f0",
          8025 => x"f0",
          8026 => x"f0",
          8027 => x"17",
          8028 => x"0f",
          8029 => x"07",
          8030 => x"f0",
          8031 => x"f0",
          8032 => x"f0",
          8033 => x"f0",
          8034 => x"f0",
          8035 => x"4d",
          8036 => x"f0",
          8037 => x"78",
          8038 => x"d5",
          8039 => x"4c",
          8040 => x"5f",
          8041 => x"d0",
          8042 => x"bb",
          8043 => x"f0",
          8044 => x"f0",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"01",
          9080 => x"f2",
          9081 => x"fa",
          9082 => x"c2",
          9083 => x"e5",
          9084 => x"62",
          9085 => x"6b",
          9086 => x"22",
          9087 => x"4f",
          9088 => x"02",
          9089 => x"0a",
          9090 => x"12",
          9091 => x"1a",
          9092 => x"82",
          9093 => x"8a",
          9094 => x"92",
          9095 => x"9a",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
        others => X"00"
    );

    shared variable RAM6 : ramArray :=
    (
             0 => x"0d",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"83",
             9 => x"2b",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"82",
            14 => x"83",
            15 => x"a5",
            16 => x"05",
            17 => x"09",
            18 => x"51",
            19 => x"00",
            20 => x"2e",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"10",
            26 => x"0a",
            27 => x"00",
            28 => x"2e",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"04",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"53",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"81",
            45 => x"04",
            46 => x"00",
            47 => x"00",
            48 => x"9f",
            49 => x"06",
            50 => x"00",
            51 => x"00",
            52 => x"06",
            53 => x"05",
            54 => x"06",
            55 => x"00",
            56 => x"05",
            57 => x"81",
            58 => x"00",
            59 => x"00",
            60 => x"05",
            61 => x"09",
            62 => x"00",
            63 => x"00",
            64 => x"04",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"83",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"b5",
            83 => x"00",
            84 => x"08",
            85 => x"2d",
            86 => x"8c",
            87 => x"00",
            88 => x"08",
            89 => x"2d",
            90 => x"8c",
            91 => x"00",
            92 => x"09",
            93 => x"54",
            94 => x"ff",
            95 => x"00",
            96 => x"09",
            97 => x"70",
            98 => x"05",
            99 => x"04",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"04",
           133 => x"0b",
           134 => x"8c",
           135 => x"04",
           136 => x"0b",
           137 => x"8c",
           138 => x"04",
           139 => x"0b",
           140 => x"8d",
           141 => x"04",
           142 => x"0b",
           143 => x"8d",
           144 => x"04",
           145 => x"0b",
           146 => x"8e",
           147 => x"04",
           148 => x"0b",
           149 => x"8e",
           150 => x"04",
           151 => x"0b",
           152 => x"8f",
           153 => x"04",
           154 => x"0b",
           155 => x"8f",
           156 => x"04",
           157 => x"0b",
           158 => x"90",
           159 => x"04",
           160 => x"0b",
           161 => x"91",
           162 => x"04",
           163 => x"0b",
           164 => x"91",
           165 => x"04",
           166 => x"0b",
           167 => x"92",
           168 => x"04",
           169 => x"0b",
           170 => x"92",
           171 => x"04",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"84",
           193 => x"84",
           194 => x"04",
           195 => x"84",
           196 => x"04",
           197 => x"84",
           198 => x"04",
           199 => x"84",
           200 => x"04",
           201 => x"84",
           202 => x"04",
           203 => x"84",
           204 => x"04",
           205 => x"84",
           206 => x"04",
           207 => x"84",
           208 => x"04",
           209 => x"84",
           210 => x"04",
           211 => x"84",
           212 => x"04",
           213 => x"84",
           214 => x"04",
           215 => x"84",
           216 => x"04",
           217 => x"2d",
           218 => x"90",
           219 => x"d1",
           220 => x"80",
           221 => x"d2",
           222 => x"c0",
           223 => x"80",
           224 => x"80",
           225 => x"0c",
           226 => x"08",
           227 => x"d4",
           228 => x"d4",
           229 => x"b9",
           230 => x"b9",
           231 => x"84",
           232 => x"84",
           233 => x"04",
           234 => x"2d",
           235 => x"90",
           236 => x"a5",
           237 => x"80",
           238 => x"df",
           239 => x"c0",
           240 => x"82",
           241 => x"80",
           242 => x"0c",
           243 => x"08",
           244 => x"d4",
           245 => x"d4",
           246 => x"b9",
           247 => x"b9",
           248 => x"84",
           249 => x"84",
           250 => x"04",
           251 => x"2d",
           252 => x"90",
           253 => x"bd",
           254 => x"80",
           255 => x"93",
           256 => x"c0",
           257 => x"83",
           258 => x"80",
           259 => x"0c",
           260 => x"08",
           261 => x"d4",
           262 => x"d4",
           263 => x"b9",
           264 => x"b9",
           265 => x"84",
           266 => x"84",
           267 => x"04",
           268 => x"2d",
           269 => x"90",
           270 => x"f7",
           271 => x"80",
           272 => x"a0",
           273 => x"c0",
           274 => x"82",
           275 => x"80",
           276 => x"0c",
           277 => x"08",
           278 => x"d4",
           279 => x"d4",
           280 => x"b9",
           281 => x"b9",
           282 => x"84",
           283 => x"84",
           284 => x"04",
           285 => x"2d",
           286 => x"90",
           287 => x"e1",
           288 => x"80",
           289 => x"d0",
           290 => x"c0",
           291 => x"80",
           292 => x"80",
           293 => x"0c",
           294 => x"08",
           295 => x"d4",
           296 => x"08",
           297 => x"d4",
           298 => x"d4",
           299 => x"b9",
           300 => x"b9",
           301 => x"84",
           302 => x"84",
           303 => x"04",
           304 => x"2d",
           305 => x"90",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"73",
           311 => x"81",
           312 => x"07",
           313 => x"72",
           314 => x"09",
           315 => x"0a",
           316 => x"51",
           317 => x"84",
           318 => x"70",
           319 => x"93",
           320 => x"ba",
           321 => x"70",
           322 => x"74",
           323 => x"c5",
           324 => x"0d",
           325 => x"32",
           326 => x"58",
           327 => x"09",
           328 => x"77",
           329 => x"07",
           330 => x"80",
           331 => x"b2",
           332 => x"b9",
           333 => x"ff",
           334 => x"75",
           335 => x"73",
           336 => x"9f",
           337 => x"24",
           338 => x"71",
           339 => x"04",
           340 => x"3d",
           341 => x"86",
           342 => x"56",
           343 => x"53",
           344 => x"9d",
           345 => x"8d",
           346 => x"3d",
           347 => x"85",
           348 => x"0d",
           349 => x"70",
           350 => x"81",
           351 => x"5b",
           352 => x"06",
           353 => x"7b",
           354 => x"81",
           355 => x"81",
           356 => x"81",
           357 => x"70",
           358 => x"38",
           359 => x"2a",
           360 => x"7e",
           361 => x"07",
           362 => x"38",
           363 => x"c8",
           364 => x"2a",
           365 => x"05",
           366 => x"70",
           367 => x"70",
           368 => x"80",
           369 => x"06",
           370 => x"33",
           371 => x"b8",
           372 => x"93",
           373 => x"8a",
           374 => x"38",
           375 => x"8b",
           376 => x"cc",
           377 => x"70",
           378 => x"81",
           379 => x"38",
           380 => x"97",
           381 => x"05",
           382 => x"54",
           383 => x"7c",
           384 => x"7c",
           385 => x"fe",
           386 => x"39",
           387 => x"08",
           388 => x"41",
           389 => x"75",
           390 => x"08",
           391 => x"18",
           392 => x"88",
           393 => x"55",
           394 => x"79",
           395 => x"b9",
           396 => x"c5",
           397 => x"2b",
           398 => x"2e",
           399 => x"fc",
           400 => x"55",
           401 => x"5f",
           402 => x"80",
           403 => x"79",
           404 => x"80",
           405 => x"90",
           406 => x"06",
           407 => x"75",
           408 => x"54",
           409 => x"83",
           410 => x"86",
           411 => x"54",
           412 => x"79",
           413 => x"83",
           414 => x"2e",
           415 => x"06",
           416 => x"2a",
           417 => x"7a",
           418 => x"97",
           419 => x"8f",
           420 => x"7e",
           421 => x"80",
           422 => x"90",
           423 => x"9d",
           424 => x"3f",
           425 => x"80",
           426 => x"54",
           427 => x"06",
           428 => x"79",
           429 => x"05",
           430 => x"75",
           431 => x"87",
           432 => x"29",
           433 => x"5b",
           434 => x"7a",
           435 => x"7a",
           436 => x"e3",
           437 => x"2e",
           438 => x"81",
           439 => x"96",
           440 => x"52",
           441 => x"d8",
           442 => x"81",
           443 => x"38",
           444 => x"80",
           445 => x"55",
           446 => x"52",
           447 => x"7a",
           448 => x"33",
           449 => x"c8",
           450 => x"f8",
           451 => x"08",
           452 => x"42",
           453 => x"84",
           454 => x"13",
           455 => x"84",
           456 => x"70",
           457 => x"41",
           458 => x"5c",
           459 => x"84",
           460 => x"70",
           461 => x"25",
           462 => x"85",
           463 => x"83",
           464 => x"ff",
           465 => x"75",
           466 => x"d8",
           467 => x"ff",
           468 => x"ff",
           469 => x"70",
           470 => x"3f",
           471 => x"fc",
           472 => x"fc",
           473 => x"58",
           474 => x"81",
           475 => x"38",
           476 => x"71",
           477 => x"7e",
           478 => x"bf",
           479 => x"ad",
           480 => x"5b",
           481 => x"7a",
           482 => x"59",
           483 => x"7f",
           484 => x"06",
           485 => x"38",
           486 => x"c8",
           487 => x"31",
           488 => x"58",
           489 => x"7c",
           490 => x"f7",
           491 => x"08",
           492 => x"79",
           493 => x"3f",
           494 => x"06",
           495 => x"c4",
           496 => x"58",
           497 => x"39",
           498 => x"80",
           499 => x"54",
           500 => x"52",
           501 => x"7c",
           502 => x"90",
           503 => x"7c",
           504 => x"88",
           505 => x"fb",
           506 => x"2c",
           507 => x"2c",
           508 => x"53",
           509 => x"7c",
           510 => x"81",
           511 => x"38",
           512 => x"2a",
           513 => x"5b",
           514 => x"c8",
           515 => x"98",
           516 => x"52",
           517 => x"7c",
           518 => x"be",
           519 => x"3f",
           520 => x"06",
           521 => x"fd",
           522 => x"71",
           523 => x"fd",
           524 => x"a8",
           525 => x"b5",
           526 => x"0d",
           527 => x"08",
           528 => x"32",
           529 => x"57",
           530 => x"06",
           531 => x"56",
           532 => x"84",
           533 => x"14",
           534 => x"08",
           535 => x"70",
           536 => x"2e",
           537 => x"d7",
           538 => x"d5",
           539 => x"08",
           540 => x"80",
           541 => x"75",
           542 => x"04",
           543 => x"80",
           544 => x"81",
           545 => x"57",
           546 => x"06",
           547 => x"33",
           548 => x"98",
           549 => x"0c",
           550 => x"05",
           551 => x"38",
           552 => x"53",
           553 => x"2e",
           554 => x"56",
           555 => x"39",
           556 => x"52",
           557 => x"04",
           558 => x"33",
           559 => x"56",
           560 => x"38",
           561 => x"80",
           562 => x"72",
           563 => x"08",
           564 => x"05",
           565 => x"13",
           566 => x"b9",
           567 => x"52",
           568 => x"08",
           569 => x"c8",
           570 => x"05",
           571 => x"fb",
           572 => x"81",
           573 => x"55",
           574 => x"38",
           575 => x"b3",
           576 => x"71",
           577 => x"70",
           578 => x"f0",
           579 => x"08",
           580 => x"ff",
           581 => x"87",
           582 => x"53",
           583 => x"81",
           584 => x"84",
           585 => x"75",
           586 => x"84",
           587 => x"08",
           588 => x"33",
           589 => x"c8",
           590 => x"07",
           591 => x"73",
           592 => x"04",
           593 => x"34",
           594 => x"75",
           595 => x"81",
           596 => x"ff",
           597 => x"33",
           598 => x"34",
           599 => x"0c",
           600 => x"76",
           601 => x"70",
           602 => x"a1",
           603 => x"70",
           604 => x"05",
           605 => x"38",
           606 => x"0d",
           607 => x"d9",
           608 => x"13",
           609 => x"34",
           610 => x"38",
           611 => x"33",
           612 => x"38",
           613 => x"53",
           614 => x"51",
           615 => x"31",
           616 => x"0d",
           617 => x"54",
           618 => x"33",
           619 => x"34",
           620 => x"0c",
           621 => x"75",
           622 => x"70",
           623 => x"05",
           624 => x"34",
           625 => x"84",
           626 => x"fc",
           627 => x"54",
           628 => x"75",
           629 => x"71",
           630 => x"81",
           631 => x"ff",
           632 => x"70",
           633 => x"04",
           634 => x"53",
           635 => x"ff",
           636 => x"2e",
           637 => x"c8",
           638 => x"b9",
           639 => x"3d",
           640 => x"80",
           641 => x"b9",
           642 => x"b2",
           643 => x"84",
           644 => x"84",
           645 => x"34",
           646 => x"08",
           647 => x"08",
           648 => x"3d",
           649 => x"71",
           650 => x"2e",
           651 => x"33",
           652 => x"12",
           653 => x"ea",
           654 => x"52",
           655 => x"0d",
           656 => x"72",
           657 => x"8e",
           658 => x"34",
           659 => x"84",
           660 => x"fa",
           661 => x"52",
           662 => x"80",
           663 => x"e0",
           664 => x"73",
           665 => x"c8",
           666 => x"26",
           667 => x"2e",
           668 => x"2a",
           669 => x"54",
           670 => x"a8",
           671 => x"74",
           672 => x"11",
           673 => x"06",
           674 => x"52",
           675 => x"38",
           676 => x"b9",
           677 => x"3d",
           678 => x"70",
           679 => x"84",
           680 => x"70",
           681 => x"80",
           682 => x"71",
           683 => x"70",
           684 => x"74",
           685 => x"73",
           686 => x"10",
           687 => x"81",
           688 => x"30",
           689 => x"84",
           690 => x"51",
           691 => x"51",
           692 => x"54",
           693 => x"0d",
           694 => x"54",
           695 => x"73",
           696 => x"0c",
           697 => x"0d",
           698 => x"80",
           699 => x"3f",
           700 => x"52",
           701 => x"fe",
           702 => x"31",
           703 => x"c5",
           704 => x"38",
           705 => x"31",
           706 => x"80",
           707 => x"10",
           708 => x"07",
           709 => x"70",
           710 => x"31",
           711 => x"58",
           712 => x"b9",
           713 => x"3d",
           714 => x"7a",
           715 => x"7d",
           716 => x"57",
           717 => x"55",
           718 => x"08",
           719 => x"0c",
           720 => x"7b",
           721 => x"77",
           722 => x"a0",
           723 => x"15",
           724 => x"73",
           725 => x"80",
           726 => x"38",
           727 => x"26",
           728 => x"a0",
           729 => x"74",
           730 => x"ff",
           731 => x"ff",
           732 => x"38",
           733 => x"54",
           734 => x"78",
           735 => x"13",
           736 => x"56",
           737 => x"38",
           738 => x"56",
           739 => x"b9",
           740 => x"70",
           741 => x"56",
           742 => x"fe",
           743 => x"70",
           744 => x"a6",
           745 => x"a0",
           746 => x"38",
           747 => x"89",
           748 => x"b9",
           749 => x"58",
           750 => x"55",
           751 => x"0b",
           752 => x"04",
           753 => x"80",
           754 => x"56",
           755 => x"06",
           756 => x"70",
           757 => x"38",
           758 => x"b0",
           759 => x"80",
           760 => x"8a",
           761 => x"c4",
           762 => x"e0",
           763 => x"d0",
           764 => x"90",
           765 => x"81",
           766 => x"81",
           767 => x"38",
           768 => x"79",
           769 => x"a0",
           770 => x"84",
           771 => x"81",
           772 => x"3d",
           773 => x"0c",
           774 => x"2e",
           775 => x"15",
           776 => x"73",
           777 => x"73",
           778 => x"a0",
           779 => x"80",
           780 => x"e1",
           781 => x"3d",
           782 => x"78",
           783 => x"fe",
           784 => x"0c",
           785 => x"3f",
           786 => x"84",
           787 => x"73",
           788 => x"10",
           789 => x"08",
           790 => x"3f",
           791 => x"51",
           792 => x"83",
           793 => x"3d",
           794 => x"9d",
           795 => x"f4",
           796 => x"04",
           797 => x"83",
           798 => x"ee",
           799 => x"cf",
           800 => x"0d",
           801 => x"3f",
           802 => x"51",
           803 => x"83",
           804 => x"3d",
           805 => x"c5",
           806 => x"bc",
           807 => x"04",
           808 => x"83",
           809 => x"ee",
           810 => x"d0",
           811 => x"0d",
           812 => x"3f",
           813 => x"51",
           814 => x"83",
           815 => x"3d",
           816 => x"ed",
           817 => x"c4",
           818 => x"04",
           819 => x"80",
           820 => x"79",
           821 => x"57",
           822 => x"26",
           823 => x"70",
           824 => x"74",
           825 => x"8c",
           826 => x"3f",
           827 => x"c8",
           828 => x"51",
           829 => x"78",
           830 => x"2a",
           831 => x"80",
           832 => x"08",
           833 => x"38",
           834 => x"f5",
           835 => x"83",
           836 => x"d0",
           837 => x"c8",
           838 => x"c8",
           839 => x"b9",
           840 => x"54",
           841 => x"82",
           842 => x"57",
           843 => x"7a",
           844 => x"74",
           845 => x"87",
           846 => x"84",
           847 => x"a7",
           848 => x"d1",
           849 => x"51",
           850 => x"3d",
           851 => x"33",
           852 => x"52",
           853 => x"c8",
           854 => x"38",
           855 => x"b9",
           856 => x"04",
           857 => x"54",
           858 => x"51",
           859 => x"b9",
           860 => x"3d",
           861 => x"80",
           862 => x"41",
           863 => x"80",
           864 => x"d1",
           865 => x"84",
           866 => x"79",
           867 => x"ed",
           868 => x"73",
           869 => x"38",
           870 => x"dd",
           871 => x"08",
           872 => x"78",
           873 => x"51",
           874 => x"27",
           875 => x"55",
           876 => x"38",
           877 => x"83",
           878 => x"81",
           879 => x"88",
           880 => x"38",
           881 => x"eb",
           882 => x"26",
           883 => x"d5",
           884 => x"80",
           885 => x"08",
           886 => x"76",
           887 => x"2e",
           888 => x"78",
           889 => x"b9",
           890 => x"d2",
           891 => x"84",
           892 => x"eb",
           893 => x"38",
           894 => x"dc",
           895 => x"08",
           896 => x"73",
           897 => x"53",
           898 => x"52",
           899 => x"82",
           900 => x"a0",
           901 => x"dd",
           902 => x"51",
           903 => x"ac",
           904 => x"3f",
           905 => x"18",
           906 => x"08",
           907 => x"3f",
           908 => x"54",
           909 => x"26",
           910 => x"ac",
           911 => x"81",
           912 => x"e9",
           913 => x"06",
           914 => x"ec",
           915 => x"09",
           916 => x"fc",
           917 => x"84",
           918 => x"2c",
           919 => x"32",
           920 => x"07",
           921 => x"53",
           922 => x"51",
           923 => x"98",
           924 => x"70",
           925 => x"72",
           926 => x"58",
           927 => x"ff",
           928 => x"84",
           929 => x"fe",
           930 => x"53",
           931 => x"3f",
           932 => x"80",
           933 => x"70",
           934 => x"38",
           935 => x"52",
           936 => x"70",
           937 => x"38",
           938 => x"52",
           939 => x"70",
           940 => x"38",
           941 => x"52",
           942 => x"70",
           943 => x"72",
           944 => x"38",
           945 => x"81",
           946 => x"51",
           947 => x"3f",
           948 => x"81",
           949 => x"51",
           950 => x"3f",
           951 => x"80",
           952 => x"9b",
           953 => x"ef",
           954 => x"87",
           955 => x"80",
           956 => x"51",
           957 => x"9b",
           958 => x"72",
           959 => x"71",
           960 => x"39",
           961 => x"a8",
           962 => x"8f",
           963 => x"51",
           964 => x"ff",
           965 => x"83",
           966 => x"51",
           967 => x"81",
           968 => x"94",
           969 => x"d7",
           970 => x"3f",
           971 => x"2a",
           972 => x"2e",
           973 => x"51",
           974 => x"9a",
           975 => x"72",
           976 => x"71",
           977 => x"39",
           978 => x"ff",
           979 => x"52",
           980 => x"b9",
           981 => x"40",
           982 => x"83",
           983 => x"3d",
           984 => x"3f",
           985 => x"7e",
           986 => x"ee",
           987 => x"59",
           988 => x"81",
           989 => x"06",
           990 => x"67",
           991 => x"dc",
           992 => x"09",
           993 => x"33",
           994 => x"80",
           995 => x"90",
           996 => x"52",
           997 => x"08",
           998 => x"7b",
           999 => x"b9",
          1000 => x"5e",
          1001 => x"1c",
          1002 => x"7c",
          1003 => x"7b",
          1004 => x"52",
          1005 => x"c8",
          1006 => x"2e",
          1007 => x"48",
          1008 => x"a4",
          1009 => x"06",
          1010 => x"38",
          1011 => x"3f",
          1012 => x"f3",
          1013 => x"7a",
          1014 => x"24",
          1015 => x"e4",
          1016 => x"f0",
          1017 => x"f2",
          1018 => x"56",
          1019 => x"53",
          1020 => x"ae",
          1021 => x"c8",
          1022 => x"80",
          1023 => x"7a",
          1024 => x"7a",
          1025 => x"81",
          1026 => x"7a",
          1027 => x"81",
          1028 => x"61",
          1029 => x"81",
          1030 => x"d3",
          1031 => x"80",
          1032 => x"0b",
          1033 => x"06",
          1034 => x"53",
          1035 => x"51",
          1036 => x"08",
          1037 => x"83",
          1038 => x"80",
          1039 => x"3f",
          1040 => x"38",
          1041 => x"3f",
          1042 => x"81",
          1043 => x"09",
          1044 => x"84",
          1045 => x"82",
          1046 => x"83",
          1047 => x"51",
          1048 => x"79",
          1049 => x"63",
          1050 => x"89",
          1051 => x"83",
          1052 => x"83",
          1053 => x"e4",
          1054 => x"ba",
          1055 => x"b9",
          1056 => x"fb",
          1057 => x"41",
          1058 => x"51",
          1059 => x"f3",
          1060 => x"56",
          1061 => x"53",
          1062 => x"f2",
          1063 => x"3f",
          1064 => x"f9",
          1065 => x"3f",
          1066 => x"fa",
          1067 => x"95",
          1068 => x"b8",
          1069 => x"fa",
          1070 => x"53",
          1071 => x"84",
          1072 => x"38",
          1073 => x"fa",
          1074 => x"c8",
          1075 => x"b9",
          1076 => x"d0",
          1077 => x"ff",
          1078 => x"eb",
          1079 => x"2e",
          1080 => x"8c",
          1081 => x"04",
          1082 => x"80",
          1083 => x"c8",
          1084 => x"3d",
          1085 => x"51",
          1086 => x"86",
          1087 => x"78",
          1088 => x"3f",
          1089 => x"52",
          1090 => x"7e",
          1091 => x"38",
          1092 => x"84",
          1093 => x"3d",
          1094 => x"51",
          1095 => x"80",
          1096 => x"f0",
          1097 => x"b4",
          1098 => x"38",
          1099 => x"83",
          1100 => x"d5",
          1101 => x"51",
          1102 => x"59",
          1103 => x"9f",
          1104 => x"70",
          1105 => x"84",
          1106 => x"f0",
          1107 => x"f8",
          1108 => x"53",
          1109 => x"84",
          1110 => x"38",
          1111 => x"80",
          1112 => x"c8",
          1113 => x"d7",
          1114 => x"5d",
          1115 => x"65",
          1116 => x"7a",
          1117 => x"54",
          1118 => x"d4",
          1119 => x"5c",
          1120 => x"39",
          1121 => x"80",
          1122 => x"c8",
          1123 => x"3d",
          1124 => x"51",
          1125 => x"80",
          1126 => x"f8",
          1127 => x"c8",
          1128 => x"f6",
          1129 => x"ba",
          1130 => x"93",
          1131 => x"5b",
          1132 => x"eb",
          1133 => x"ff",
          1134 => x"b9",
          1135 => x"b8",
          1136 => x"05",
          1137 => x"08",
          1138 => x"83",
          1139 => x"d5",
          1140 => x"51",
          1141 => x"59",
          1142 => x"9f",
          1143 => x"49",
          1144 => x"05",
          1145 => x"b8",
          1146 => x"05",
          1147 => x"08",
          1148 => x"02",
          1149 => x"81",
          1150 => x"53",
          1151 => x"84",
          1152 => x"b9",
          1153 => x"ff",
          1154 => x"b9",
          1155 => x"b8",
          1156 => x"05",
          1157 => x"08",
          1158 => x"fe",
          1159 => x"e6",
          1160 => x"38",
          1161 => x"88",
          1162 => x"59",
          1163 => x"7a",
          1164 => x"79",
          1165 => x"3f",
          1166 => x"05",
          1167 => x"08",
          1168 => x"88",
          1169 => x"08",
          1170 => x"b9",
          1171 => x"84",
          1172 => x"f4",
          1173 => x"53",
          1174 => x"84",
          1175 => x"cc",
          1176 => x"38",
          1177 => x"fe",
          1178 => x"e5",
          1179 => x"38",
          1180 => x"2e",
          1181 => x"47",
          1182 => x"80",
          1183 => x"c8",
          1184 => x"5c",
          1185 => x"5c",
          1186 => x"07",
          1187 => x"79",
          1188 => x"83",
          1189 => x"d6",
          1190 => x"53",
          1191 => x"83",
          1192 => x"f9",
          1193 => x"84",
          1194 => x"53",
          1195 => x"84",
          1196 => x"38",
          1197 => x"05",
          1198 => x"ff",
          1199 => x"b9",
          1200 => x"64",
          1201 => x"70",
          1202 => x"3d",
          1203 => x"51",
          1204 => x"80",
          1205 => x"80",
          1206 => x"40",
          1207 => x"11",
          1208 => x"3f",
          1209 => x"f1",
          1210 => x"53",
          1211 => x"84",
          1212 => x"38",
          1213 => x"7c",
          1214 => x"39",
          1215 => x"80",
          1216 => x"c8",
          1217 => x"64",
          1218 => x"46",
          1219 => x"09",
          1220 => x"83",
          1221 => x"b0",
          1222 => x"96",
          1223 => x"3f",
          1224 => x"d4",
          1225 => x"fe",
          1226 => x"e0",
          1227 => x"2e",
          1228 => x"05",
          1229 => x"78",
          1230 => x"33",
          1231 => x"83",
          1232 => x"83",
          1233 => x"a1",
          1234 => x"b5",
          1235 => x"3f",
          1236 => x"e8",
          1237 => x"cc",
          1238 => x"80",
          1239 => x"49",
          1240 => x"d3",
          1241 => x"ce",
          1242 => x"83",
          1243 => x"83",
          1244 => x"9b",
          1245 => x"dd",
          1246 => x"80",
          1247 => x"47",
          1248 => x"5d",
          1249 => x"a4",
          1250 => x"ca",
          1251 => x"83",
          1252 => x"83",
          1253 => x"fb",
          1254 => x"05",
          1255 => x"80",
          1256 => x"94",
          1257 => x"80",
          1258 => x"b9",
          1259 => x"55",
          1260 => x"bf",
          1261 => x"77",
          1262 => x"56",
          1263 => x"da",
          1264 => x"2b",
          1265 => x"52",
          1266 => x"b9",
          1267 => x"83",
          1268 => x"80",
          1269 => x"81",
          1270 => x"83",
          1271 => x"5e",
          1272 => x"88",
          1273 => x"ac",
          1274 => x"3f",
          1275 => x"8c",
          1276 => x"b4",
          1277 => x"70",
          1278 => x"d2",
          1279 => x"15",
          1280 => x"82",
          1281 => x"51",
          1282 => x"f0",
          1283 => x"52",
          1284 => x"ec",
          1285 => x"77",
          1286 => x"53",
          1287 => x"33",
          1288 => x"a0",
          1289 => x"15",
          1290 => x"53",
          1291 => x"81",
          1292 => x"82",
          1293 => x"e7",
          1294 => x"06",
          1295 => x"38",
          1296 => x"73",
          1297 => x"e1",
          1298 => x"54",
          1299 => x"38",
          1300 => x"70",
          1301 => x"72",
          1302 => x"81",
          1303 => x"51",
          1304 => x"0d",
          1305 => x"80",
          1306 => x"80",
          1307 => x"54",
          1308 => x"54",
          1309 => x"53",
          1310 => x"fe",
          1311 => x"76",
          1312 => x"84",
          1313 => x"86",
          1314 => x"ec",
          1315 => x"e5",
          1316 => x"3d",
          1317 => x"11",
          1318 => x"70",
          1319 => x"33",
          1320 => x"26",
          1321 => x"83",
          1322 => x"85",
          1323 => x"26",
          1324 => x"85",
          1325 => x"88",
          1326 => x"e7",
          1327 => x"54",
          1328 => x"cc",
          1329 => x"0c",
          1330 => x"82",
          1331 => x"83",
          1332 => x"84",
          1333 => x"85",
          1334 => x"86",
          1335 => x"74",
          1336 => x"c0",
          1337 => x"98",
          1338 => x"c8",
          1339 => x"0d",
          1340 => x"81",
          1341 => x"5e",
          1342 => x"08",
          1343 => x"98",
          1344 => x"87",
          1345 => x"1c",
          1346 => x"79",
          1347 => x"08",
          1348 => x"98",
          1349 => x"87",
          1350 => x"1c",
          1351 => x"ff",
          1352 => x"58",
          1353 => x"56",
          1354 => x"54",
          1355 => x"ff",
          1356 => x"bf",
          1357 => x"3d",
          1358 => x"81",
          1359 => x"a6",
          1360 => x"70",
          1361 => x"09",
          1362 => x"e3",
          1363 => x"3d",
          1364 => x"3f",
          1365 => x"98",
          1366 => x"81",
          1367 => x"e6",
          1368 => x"70",
          1369 => x"d2",
          1370 => x"70",
          1371 => x"51",
          1372 => x"08",
          1373 => x"71",
          1374 => x"81",
          1375 => x"38",
          1376 => x"0d",
          1377 => x"33",
          1378 => x"06",
          1379 => x"f4",
          1380 => x"96",
          1381 => x"70",
          1382 => x"70",
          1383 => x"72",
          1384 => x"2e",
          1385 => x"52",
          1386 => x"51",
          1387 => x"2e",
          1388 => x"74",
          1389 => x"86",
          1390 => x"81",
          1391 => x"81",
          1392 => x"cb",
          1393 => x"71",
          1394 => x"84",
          1395 => x"53",
          1396 => x"ff",
          1397 => x"30",
          1398 => x"83",
          1399 => x"fa",
          1400 => x"70",
          1401 => x"e7",
          1402 => x"70",
          1403 => x"80",
          1404 => x"94",
          1405 => x"53",
          1406 => x"71",
          1407 => x"70",
          1408 => x"53",
          1409 => x"2a",
          1410 => x"81",
          1411 => x"52",
          1412 => x"94",
          1413 => x"75",
          1414 => x"76",
          1415 => x"04",
          1416 => x"51",
          1417 => x"06",
          1418 => x"93",
          1419 => x"ff",
          1420 => x"70",
          1421 => x"52",
          1422 => x"0d",
          1423 => x"2a",
          1424 => x"84",
          1425 => x"83",
          1426 => x"08",
          1427 => x"94",
          1428 => x"9e",
          1429 => x"c0",
          1430 => x"87",
          1431 => x"0c",
          1432 => x"9c",
          1433 => x"f2",
          1434 => x"83",
          1435 => x"08",
          1436 => x"bc",
          1437 => x"9e",
          1438 => x"c0",
          1439 => x"87",
          1440 => x"f2",
          1441 => x"83",
          1442 => x"08",
          1443 => x"8c",
          1444 => x"83",
          1445 => x"9e",
          1446 => x"51",
          1447 => x"83",
          1448 => x"9e",
          1449 => x"51",
          1450 => x"81",
          1451 => x"0b",
          1452 => x"80",
          1453 => x"2e",
          1454 => x"cb",
          1455 => x"08",
          1456 => x"52",
          1457 => x"71",
          1458 => x"c0",
          1459 => x"06",
          1460 => x"38",
          1461 => x"80",
          1462 => x"90",
          1463 => x"80",
          1464 => x"f2",
          1465 => x"90",
          1466 => x"52",
          1467 => x"52",
          1468 => x"87",
          1469 => x"80",
          1470 => x"83",
          1471 => x"34",
          1472 => x"70",
          1473 => x"70",
          1474 => x"83",
          1475 => x"9e",
          1476 => x"51",
          1477 => x"81",
          1478 => x"0b",
          1479 => x"80",
          1480 => x"83",
          1481 => x"34",
          1482 => x"06",
          1483 => x"f2",
          1484 => x"90",
          1485 => x"52",
          1486 => x"71",
          1487 => x"90",
          1488 => x"53",
          1489 => x"0b",
          1490 => x"06",
          1491 => x"38",
          1492 => x"87",
          1493 => x"70",
          1494 => x"04",
          1495 => x"0d",
          1496 => x"3f",
          1497 => x"9f",
          1498 => x"3f",
          1499 => x"ef",
          1500 => x"85",
          1501 => x"75",
          1502 => x"55",
          1503 => x"33",
          1504 => x"d3",
          1505 => x"f2",
          1506 => x"83",
          1507 => x"38",
          1508 => x"c4",
          1509 => x"83",
          1510 => x"74",
          1511 => x"56",
          1512 => x"33",
          1513 => x"b0",
          1514 => x"08",
          1515 => x"aa",
          1516 => x"d9",
          1517 => x"f2",
          1518 => x"ff",
          1519 => x"c1",
          1520 => x"83",
          1521 => x"83",
          1522 => x"52",
          1523 => x"c8",
          1524 => x"31",
          1525 => x"83",
          1526 => x"83",
          1527 => x"83",
          1528 => x"87",
          1529 => x"56",
          1530 => x"cf",
          1531 => x"c0",
          1532 => x"b9",
          1533 => x"ff",
          1534 => x"83",
          1535 => x"52",
          1536 => x"c8",
          1537 => x"31",
          1538 => x"83",
          1539 => x"83",
          1540 => x"ff",
          1541 => x"e8",
          1542 => x"51",
          1543 => x"52",
          1544 => x"3f",
          1545 => x"e4",
          1546 => x"b4",
          1547 => x"b3",
          1548 => x"8d",
          1549 => x"da",
          1550 => x"f2",
          1551 => x"75",
          1552 => x"08",
          1553 => x"54",
          1554 => x"da",
          1555 => x"f2",
          1556 => x"97",
          1557 => x"51",
          1558 => x"33",
          1559 => x"fe",
          1560 => x"bf",
          1561 => x"75",
          1562 => x"83",
          1563 => x"83",
          1564 => x"fc",
          1565 => x"51",
          1566 => x"33",
          1567 => x"d7",
          1568 => x"dc",
          1569 => x"f2",
          1570 => x"91",
          1571 => x"52",
          1572 => x"3f",
          1573 => x"2e",
          1574 => x"d4",
          1575 => x"b1",
          1576 => x"73",
          1577 => x"83",
          1578 => x"11",
          1579 => x"b1",
          1580 => x"75",
          1581 => x"83",
          1582 => x"11",
          1583 => x"b1",
          1584 => x"73",
          1585 => x"83",
          1586 => x"11",
          1587 => x"b0",
          1588 => x"74",
          1589 => x"83",
          1590 => x"11",
          1591 => x"b0",
          1592 => x"75",
          1593 => x"83",
          1594 => x"11",
          1595 => x"b0",
          1596 => x"73",
          1597 => x"83",
          1598 => x"83",
          1599 => x"83",
          1600 => x"f9",
          1601 => x"02",
          1602 => x"8c",
          1603 => x"05",
          1604 => x"51",
          1605 => x"04",
          1606 => x"3f",
          1607 => x"51",
          1608 => x"04",
          1609 => x"3f",
          1610 => x"51",
          1611 => x"04",
          1612 => x"3f",
          1613 => x"0c",
          1614 => x"0c",
          1615 => x"96",
          1616 => x"3d",
          1617 => x"70",
          1618 => x"08",
          1619 => x"c8",
          1620 => x"ff",
          1621 => x"80",
          1622 => x"3f",
          1623 => x"38",
          1624 => x"c8",
          1625 => x"84",
          1626 => x"b9",
          1627 => x"55",
          1628 => x"70",
          1629 => x"78",
          1630 => x"38",
          1631 => x"53",
          1632 => x"c8",
          1633 => x"38",
          1634 => x"0d",
          1635 => x"ea",
          1636 => x"e8",
          1637 => x"3f",
          1638 => x"3d",
          1639 => x"34",
          1640 => x"ad",
          1641 => x"0c",
          1642 => x"ab",
          1643 => x"5d",
          1644 => x"a0",
          1645 => x"3d",
          1646 => x"f3",
          1647 => x"bf",
          1648 => x"79",
          1649 => x"84",
          1650 => x"33",
          1651 => x"73",
          1652 => x"81",
          1653 => x"c2",
          1654 => x"0c",
          1655 => x"aa",
          1656 => x"05",
          1657 => x"08",
          1658 => x"78",
          1659 => x"b9",
          1660 => x"80",
          1661 => x"ff",
          1662 => x"fa",
          1663 => x"05",
          1664 => x"81",
          1665 => x"73",
          1666 => x"38",
          1667 => x"8d",
          1668 => x"84",
          1669 => x"08",
          1670 => x"b9",
          1671 => x"b4",
          1672 => x"82",
          1673 => x"80",
          1674 => x"d2",
          1675 => x"0b",
          1676 => x"84",
          1677 => x"58",
          1678 => x"52",
          1679 => x"ff",
          1680 => x"81",
          1681 => x"b9",
          1682 => x"3d",
          1683 => x"b9",
          1684 => x"b4",
          1685 => x"f3",
          1686 => x"74",
          1687 => x"80",
          1688 => x"91",
          1689 => x"57",
          1690 => x"90",
          1691 => x"5f",
          1692 => x"c8",
          1693 => x"56",
          1694 => x"ff",
          1695 => x"2b",
          1696 => x"70",
          1697 => x"2c",
          1698 => x"05",
          1699 => x"5c",
          1700 => x"81",
          1701 => x"78",
          1702 => x"80",
          1703 => x"98",
          1704 => x"cb",
          1705 => x"56",
          1706 => x"33",
          1707 => x"83",
          1708 => x"56",
          1709 => x"76",
          1710 => x"80",
          1711 => x"99",
          1712 => x"98",
          1713 => x"2b",
          1714 => x"70",
          1715 => x"5f",
          1716 => x"7a",
          1717 => x"d1",
          1718 => x"76",
          1719 => x"29",
          1720 => x"70",
          1721 => x"95",
          1722 => x"70",
          1723 => x"de",
          1724 => x"25",
          1725 => x"18",
          1726 => x"ff",
          1727 => x"38",
          1728 => x"2e",
          1729 => x"56",
          1730 => x"e9",
          1731 => x"84",
          1732 => x"7f",
          1733 => x"b0",
          1734 => x"05",
          1735 => x"15",
          1736 => x"84",
          1737 => x"d9",
          1738 => x"80",
          1739 => x"08",
          1740 => x"84",
          1741 => x"84",
          1742 => x"d1",
          1743 => x"d1",
          1744 => x"27",
          1745 => x"52",
          1746 => x"34",
          1747 => x"b5",
          1748 => x"2e",
          1749 => x"f2",
          1750 => x"8f",
          1751 => x"75",
          1752 => x"d1",
          1753 => x"b6",
          1754 => x"51",
          1755 => x"08",
          1756 => x"84",
          1757 => x"b4",
          1758 => x"05",
          1759 => x"81",
          1760 => x"51",
          1761 => x"8c",
          1762 => x"83",
          1763 => x"38",
          1764 => x"fc",
          1765 => x"38",
          1766 => x"a8",
          1767 => x"84",
          1768 => x"84",
          1769 => x"05",
          1770 => x"94",
          1771 => x"8c",
          1772 => x"9e",
          1773 => x"51",
          1774 => x"08",
          1775 => x"84",
          1776 => x"b3",
          1777 => x"05",
          1778 => x"81",
          1779 => x"8c",
          1780 => x"88",
          1781 => x"fa",
          1782 => x"81",
          1783 => x"7b",
          1784 => x"a8",
          1785 => x"ff",
          1786 => x"55",
          1787 => x"d5",
          1788 => x"84",
          1789 => x"52",
          1790 => x"8c",
          1791 => x"88",
          1792 => x"ff",
          1793 => x"8c",
          1794 => x"74",
          1795 => x"5b",
          1796 => x"2b",
          1797 => x"43",
          1798 => x"38",
          1799 => x"ff",
          1800 => x"70",
          1801 => x"88",
          1802 => x"24",
          1803 => x"52",
          1804 => x"81",
          1805 => x"70",
          1806 => x"56",
          1807 => x"84",
          1808 => x"b1",
          1809 => x"81",
          1810 => x"d1",
          1811 => x"25",
          1812 => x"16",
          1813 => x"d5",
          1814 => x"b1",
          1815 => x"81",
          1816 => x"d1",
          1817 => x"25",
          1818 => x"18",
          1819 => x"52",
          1820 => x"75",
          1821 => x"05",
          1822 => x"5b",
          1823 => x"38",
          1824 => x"55",
          1825 => x"d5",
          1826 => x"d8",
          1827 => x"57",
          1828 => x"ff",
          1829 => x"33",
          1830 => x"d5",
          1831 => x"b0",
          1832 => x"f4",
          1833 => x"ff",
          1834 => x"d1",
          1835 => x"d8",
          1836 => x"10",
          1837 => x"5e",
          1838 => x"2b",
          1839 => x"81",
          1840 => x"fb",
          1841 => x"83",
          1842 => x"f2",
          1843 => x"74",
          1844 => x"56",
          1845 => x"b0",
          1846 => x"38",
          1847 => x"0b",
          1848 => x"c8",
          1849 => x"8c",
          1850 => x"84",
          1851 => x"af",
          1852 => x"a0",
          1853 => x"ac",
          1854 => x"3f",
          1855 => x"75",
          1856 => x"06",
          1857 => x"51",
          1858 => x"d1",
          1859 => x"34",
          1860 => x"0b",
          1861 => x"55",
          1862 => x"ac",
          1863 => x"3f",
          1864 => x"ff",
          1865 => x"52",
          1866 => x"d1",
          1867 => x"d1",
          1868 => x"74",
          1869 => x"9f",
          1870 => x"34",
          1871 => x"84",
          1872 => x"84",
          1873 => x"5c",
          1874 => x"84",
          1875 => x"84",
          1876 => x"84",
          1877 => x"52",
          1878 => x"d1",
          1879 => x"2c",
          1880 => x"56",
          1881 => x"d5",
          1882 => x"98",
          1883 => x"2b",
          1884 => x"5d",
          1885 => x"f0",
          1886 => x"51",
          1887 => x"0a",
          1888 => x"2c",
          1889 => x"74",
          1890 => x"ac",
          1891 => x"3f",
          1892 => x"0a",
          1893 => x"33",
          1894 => x"b9",
          1895 => x"81",
          1896 => x"08",
          1897 => x"3f",
          1898 => x"0a",
          1899 => x"33",
          1900 => x"e6",
          1901 => x"77",
          1902 => x"33",
          1903 => x"80",
          1904 => x"98",
          1905 => x"5b",
          1906 => x"b6",
          1907 => x"ff",
          1908 => x"b8",
          1909 => x"75",
          1910 => x"98",
          1911 => x"38",
          1912 => x"34",
          1913 => x"0a",
          1914 => x"33",
          1915 => x"38",
          1916 => x"34",
          1917 => x"b3",
          1918 => x"33",
          1919 => x"17",
          1920 => x"57",
          1921 => x"0a",
          1922 => x"2c",
          1923 => x"58",
          1924 => x"98",
          1925 => x"06",
          1926 => x"a8",
          1927 => x"51",
          1928 => x"0a",
          1929 => x"2c",
          1930 => x"75",
          1931 => x"ac",
          1932 => x"3f",
          1933 => x"0a",
          1934 => x"33",
          1935 => x"b9",
          1936 => x"08",
          1937 => x"75",
          1938 => x"c8",
          1939 => x"c8",
          1940 => x"75",
          1941 => x"84",
          1942 => x"56",
          1943 => x"84",
          1944 => x"a9",
          1945 => x"a0",
          1946 => x"ac",
          1947 => x"3f",
          1948 => x"7a",
          1949 => x"06",
          1950 => x"8b",
          1951 => x"b4",
          1952 => x"38",
          1953 => x"ca",
          1954 => x"08",
          1955 => x"ff",
          1956 => x"29",
          1957 => x"84",
          1958 => x"76",
          1959 => x"70",
          1960 => x"ff",
          1961 => x"25",
          1962 => x"f3",
          1963 => x"83",
          1964 => x"55",
          1965 => x"58",
          1966 => x"0b",
          1967 => x"08",
          1968 => x"74",
          1969 => x"b4",
          1970 => x"0b",
          1971 => x"3d",
          1972 => x"80",
          1973 => x"16",
          1974 => x"ff",
          1975 => x"ff",
          1976 => x"84",
          1977 => x"81",
          1978 => x"7b",
          1979 => x"84",
          1980 => x"57",
          1981 => x"38",
          1982 => x"ff",
          1983 => x"52",
          1984 => x"d5",
          1985 => x"e0",
          1986 => x"5a",
          1987 => x"ff",
          1988 => x"80",
          1989 => x"84",
          1990 => x"0c",
          1991 => x"a9",
          1992 => x"d1",
          1993 => x"ff",
          1994 => x"51",
          1995 => x"81",
          1996 => x"d1",
          1997 => x"80",
          1998 => x"08",
          1999 => x"84",
          2000 => x"a5",
          2001 => x"88",
          2002 => x"8c",
          2003 => x"8c",
          2004 => x"39",
          2005 => x"b9",
          2006 => x"b9",
          2007 => x"53",
          2008 => x"3f",
          2009 => x"d1",
          2010 => x"58",
          2011 => x"38",
          2012 => x"ff",
          2013 => x"52",
          2014 => x"d5",
          2015 => x"f0",
          2016 => x"41",
          2017 => x"ff",
          2018 => x"d6",
          2019 => x"82",
          2020 => x"05",
          2021 => x"80",
          2022 => x"7b",
          2023 => x"10",
          2024 => x"41",
          2025 => x"75",
          2026 => x"94",
          2027 => x"70",
          2028 => x"27",
          2029 => x"34",
          2030 => x"05",
          2031 => x"81",
          2032 => x"52",
          2033 => x"f3",
          2034 => x"80",
          2035 => x"84",
          2036 => x"0c",
          2037 => x"52",
          2038 => x"f8",
          2039 => x"38",
          2040 => x"5d",
          2041 => x"52",
          2042 => x"b9",
          2043 => x"7b",
          2044 => x"84",
          2045 => x"3f",
          2046 => x"84",
          2047 => x"84",
          2048 => x"58",
          2049 => x"06",
          2050 => x"83",
          2051 => x"58",
          2052 => x"2b",
          2053 => x"81",
          2054 => x"cb",
          2055 => x"83",
          2056 => x"f2",
          2057 => x"74",
          2058 => x"06",
          2059 => x"80",
          2060 => x"fe",
          2061 => x"e6",
          2062 => x"ff",
          2063 => x"81",
          2064 => x"93",
          2065 => x"83",
          2066 => x"51",
          2067 => x"33",
          2068 => x"f2",
          2069 => x"56",
          2070 => x"c8",
          2071 => x"70",
          2072 => x"08",
          2073 => x"82",
          2074 => x"b8",
          2075 => x"b8",
          2076 => x"51",
          2077 => x"38",
          2078 => x"80",
          2079 => x"c7",
          2080 => x"81",
          2081 => x"38",
          2082 => x"82",
          2083 => x"80",
          2084 => x"57",
          2085 => x"2e",
          2086 => x"75",
          2087 => x"f6",
          2088 => x"2b",
          2089 => x"07",
          2090 => x"5b",
          2091 => x"70",
          2092 => x"84",
          2093 => x"38",
          2094 => x"f4",
          2095 => x"31",
          2096 => x"15",
          2097 => x"34",
          2098 => x"3d",
          2099 => x"83",
          2100 => x"83",
          2101 => x"74",
          2102 => x"a7",
          2103 => x"70",
          2104 => x"70",
          2105 => x"70",
          2106 => x"5d",
          2107 => x"73",
          2108 => x"75",
          2109 => x"81",
          2110 => x"83",
          2111 => x"70",
          2112 => x"5b",
          2113 => x"f8",
          2114 => x"7d",
          2115 => x"5c",
          2116 => x"7d",
          2117 => x"38",
          2118 => x"83",
          2119 => x"56",
          2120 => x"59",
          2121 => x"bc",
          2122 => x"bb",
          2123 => x"f6",
          2124 => x"57",
          2125 => x"81",
          2126 => x"81",
          2127 => x"54",
          2128 => x"80",
          2129 => x"83",
          2130 => x"70",
          2131 => x"88",
          2132 => x"56",
          2133 => x"38",
          2134 => x"83",
          2135 => x"70",
          2136 => x"71",
          2137 => x"11",
          2138 => x"a7",
          2139 => x"33",
          2140 => x"33",
          2141 => x"22",
          2142 => x"29",
          2143 => x"5f",
          2144 => x"38",
          2145 => x"19",
          2146 => x"81",
          2147 => x"ff",
          2148 => x"75",
          2149 => x"7b",
          2150 => x"53",
          2151 => x"5b",
          2152 => x"06",
          2153 => x"39",
          2154 => x"9a",
          2155 => x"8c",
          2156 => x"34",
          2157 => x"ee",
          2158 => x"ff",
          2159 => x"56",
          2160 => x"ee",
          2161 => x"74",
          2162 => x"83",
          2163 => x"e0",
          2164 => x"86",
          2165 => x"07",
          2166 => x"70",
          2167 => x"53",
          2168 => x"08",
          2169 => x"72",
          2170 => x"81",
          2171 => x"34",
          2172 => x"80",
          2173 => x"0d",
          2174 => x"c8",
          2175 => x"05",
          2176 => x"84",
          2177 => x"53",
          2178 => x"b7",
          2179 => x"f8",
          2180 => x"a7",
          2181 => x"5f",
          2182 => x"70",
          2183 => x"33",
          2184 => x"83",
          2185 => x"05",
          2186 => x"f8",
          2187 => x"06",
          2188 => x"72",
          2189 => x"53",
          2190 => x"f6",
          2191 => x"b7",
          2192 => x"26",
          2193 => x"76",
          2194 => x"9f",
          2195 => x"70",
          2196 => x"e0",
          2197 => x"54",
          2198 => x"81",
          2199 => x"e3",
          2200 => x"83",
          2201 => x"54",
          2202 => x"74",
          2203 => x"14",
          2204 => x"84",
          2205 => x"83",
          2206 => x"ff",
          2207 => x"54",
          2208 => x"74",
          2209 => x"71",
          2210 => x"86",
          2211 => x"80",
          2212 => x"06",
          2213 => x"57",
          2214 => x"9a",
          2215 => x"84",
          2216 => x"05",
          2217 => x"33",
          2218 => x"15",
          2219 => x"33",
          2220 => x"55",
          2221 => x"72",
          2222 => x"04",
          2223 => x"f6",
          2224 => x"b7",
          2225 => x"27",
          2226 => x"dd",
          2227 => x"83",
          2228 => x"2e",
          2229 => x"76",
          2230 => x"71",
          2231 => x"52",
          2232 => x"38",
          2233 => x"15",
          2234 => x"0b",
          2235 => x"81",
          2236 => x"80",
          2237 => x"e0",
          2238 => x"57",
          2239 => x"fd",
          2240 => x"33",
          2241 => x"fa",
          2242 => x"33",
          2243 => x"fc",
          2244 => x"84",
          2245 => x"86",
          2246 => x"c3",
          2247 => x"b7",
          2248 => x"38",
          2249 => x"84",
          2250 => x"80",
          2251 => x"f8",
          2252 => x"72",
          2253 => x"70",
          2254 => x"b9",
          2255 => x"f8",
          2256 => x"70",
          2257 => x"54",
          2258 => x"83",
          2259 => x"bb",
          2260 => x"75",
          2261 => x"f8",
          2262 => x"0c",
          2263 => x"33",
          2264 => x"2c",
          2265 => x"83",
          2266 => x"c8",
          2267 => x"f9",
          2268 => x"ff",
          2269 => x"83",
          2270 => x"34",
          2271 => x"3d",
          2272 => x"34",
          2273 => x"33",
          2274 => x"fe",
          2275 => x"f8",
          2276 => x"0d",
          2277 => x"26",
          2278 => x"88",
          2279 => x"f4",
          2280 => x"2b",
          2281 => x"07",
          2282 => x"2e",
          2283 => x"0b",
          2284 => x"b9",
          2285 => x"f8",
          2286 => x"51",
          2287 => x"84",
          2288 => x"83",
          2289 => x"70",
          2290 => x"f8",
          2291 => x"51",
          2292 => x"80",
          2293 => x"0b",
          2294 => x"04",
          2295 => x"84",
          2296 => x"ff",
          2297 => x"07",
          2298 => x"a5",
          2299 => x"06",
          2300 => x"34",
          2301 => x"81",
          2302 => x"f8",
          2303 => x"f4",
          2304 => x"70",
          2305 => x"83",
          2306 => x"70",
          2307 => x"83",
          2308 => x"d0",
          2309 => x"fe",
          2310 => x"bf",
          2311 => x"f4",
          2312 => x"33",
          2313 => x"70",
          2314 => x"83",
          2315 => x"c0",
          2316 => x"fe",
          2317 => x"af",
          2318 => x"f4",
          2319 => x"33",
          2320 => x"f4",
          2321 => x"33",
          2322 => x"83",
          2323 => x"3d",
          2324 => x"05",
          2325 => x"33",
          2326 => x"33",
          2327 => x"5d",
          2328 => x"38",
          2329 => x"2e",
          2330 => x"34",
          2331 => x"83",
          2332 => x"23",
          2333 => x"0d",
          2334 => x"db",
          2335 => x"81",
          2336 => x"83",
          2337 => x"f9",
          2338 => x"79",
          2339 => x"b7",
          2340 => x"55",
          2341 => x"e3",
          2342 => x"84",
          2343 => x"c0",
          2344 => x"83",
          2345 => x"34",
          2346 => x"b7",
          2347 => x"34",
          2348 => x"0b",
          2349 => x"f8",
          2350 => x"84",
          2351 => x"33",
          2352 => x"7a",
          2353 => x"fa",
          2354 => x"5a",
          2355 => x"10",
          2356 => x"59",
          2357 => x"3f",
          2358 => x"b8",
          2359 => x"26",
          2360 => x"80",
          2361 => x"80",
          2362 => x"f8",
          2363 => x"7c",
          2364 => x"04",
          2365 => x"0b",
          2366 => x"f8",
          2367 => x"34",
          2368 => x"f7",
          2369 => x"b9",
          2370 => x"fe",
          2371 => x"ac",
          2372 => x"b9",
          2373 => x"f7",
          2374 => x"51",
          2375 => x"81",
          2376 => x"3d",
          2377 => x"33",
          2378 => x"33",
          2379 => x"12",
          2380 => x"f6",
          2381 => x"29",
          2382 => x"f7",
          2383 => x"57",
          2384 => x"89",
          2385 => x"81",
          2386 => x"38",
          2387 => x"b7",
          2388 => x"f8",
          2389 => x"56",
          2390 => x"a7",
          2391 => x"33",
          2392 => x"22",
          2393 => x"53",
          2394 => x"f8",
          2395 => x"54",
          2396 => x"80",
          2397 => x"81",
          2398 => x"f8",
          2399 => x"5b",
          2400 => x"84",
          2401 => x"81",
          2402 => x"81",
          2403 => x"77",
          2404 => x"83",
          2405 => x"53",
          2406 => x"c0",
          2407 => x"38",
          2408 => x"3d",
          2409 => x"75",
          2410 => x"2e",
          2411 => x"52",
          2412 => x"83",
          2413 => x"f8",
          2414 => x"13",
          2415 => x"81",
          2416 => x"52",
          2417 => x"70",
          2418 => x"26",
          2419 => x"fd",
          2420 => x"06",
          2421 => x"fe",
          2422 => x"fe",
          2423 => x"de",
          2424 => x"89",
          2425 => x"09",
          2426 => x"f9",
          2427 => x"05",
          2428 => x"83",
          2429 => x"fc",
          2430 => x"81",
          2431 => x"fe",
          2432 => x"f9",
          2433 => x"f8",
          2434 => x"e2",
          2435 => x"51",
          2436 => x"3d",
          2437 => x"b8",
          2438 => x"81",
          2439 => x"38",
          2440 => x"8a",
          2441 => x"84",
          2442 => x"38",
          2443 => x"33",
          2444 => x"05",
          2445 => x"33",
          2446 => x"b7",
          2447 => x"f8",
          2448 => x"5a",
          2449 => x"34",
          2450 => x"62",
          2451 => x"7f",
          2452 => x"b7",
          2453 => x"f8",
          2454 => x"72",
          2455 => x"83",
          2456 => x"34",
          2457 => x"58",
          2458 => x"b7",
          2459 => x"ff",
          2460 => x"80",
          2461 => x"0d",
          2462 => x"b7",
          2463 => x"2e",
          2464 => x"89",
          2465 => x"0c",
          2466 => x"33",
          2467 => x"05",
          2468 => x"33",
          2469 => x"b7",
          2470 => x"f8",
          2471 => x"5f",
          2472 => x"34",
          2473 => x"19",
          2474 => x"a7",
          2475 => x"33",
          2476 => x"22",
          2477 => x"11",
          2478 => x"f4",
          2479 => x"81",
          2480 => x"60",
          2481 => x"f8",
          2482 => x"0c",
          2483 => x"82",
          2484 => x"38",
          2485 => x"a8",
          2486 => x"80",
          2487 => x"0d",
          2488 => x"d0",
          2489 => x"38",
          2490 => x"57",
          2491 => x"b8",
          2492 => x"59",
          2493 => x"80",
          2494 => x"0d",
          2495 => x"80",
          2496 => x"bc",
          2497 => x"f9",
          2498 => x"40",
          2499 => x"a0",
          2500 => x"83",
          2501 => x"72",
          2502 => x"78",
          2503 => x"f8",
          2504 => x"83",
          2505 => x"1b",
          2506 => x"ff",
          2507 => x"f9",
          2508 => x"43",
          2509 => x"84",
          2510 => x"fe",
          2511 => x"fa",
          2512 => x"fe",
          2513 => x"f8",
          2514 => x"f8",
          2515 => x"a7",
          2516 => x"40",
          2517 => x"83",
          2518 => x"5a",
          2519 => x"86",
          2520 => x"1a",
          2521 => x"56",
          2522 => x"39",
          2523 => x"0b",
          2524 => x"b8",
          2525 => x"34",
          2526 => x"0b",
          2527 => x"04",
          2528 => x"34",
          2529 => x"34",
          2530 => x"34",
          2531 => x"0b",
          2532 => x"04",
          2533 => x"fa",
          2534 => x"b7",
          2535 => x"f8",
          2536 => x"75",
          2537 => x"83",
          2538 => x"29",
          2539 => x"f7",
          2540 => x"5b",
          2541 => x"78",
          2542 => x"75",
          2543 => x"f9",
          2544 => x"ff",
          2545 => x"29",
          2546 => x"33",
          2547 => x"b7",
          2548 => x"f8",
          2549 => x"5e",
          2550 => x"18",
          2551 => x"29",
          2552 => x"33",
          2553 => x"b7",
          2554 => x"f8",
          2555 => x"72",
          2556 => x"83",
          2557 => x"05",
          2558 => x"5c",
          2559 => x"84",
          2560 => x"38",
          2561 => x"34",
          2562 => x"06",
          2563 => x"78",
          2564 => x"2e",
          2565 => x"a8",
          2566 => x"83",
          2567 => x"b4",
          2568 => x"83",
          2569 => x"80",
          2570 => x"81",
          2571 => x"b9",
          2572 => x"f8",
          2573 => x"81",
          2574 => x"81",
          2575 => x"a7",
          2576 => x"5c",
          2577 => x"ff",
          2578 => x"53",
          2579 => x"2e",
          2580 => x"ff",
          2581 => x"ff",
          2582 => x"40",
          2583 => x"80",
          2584 => x"f8",
          2585 => x"71",
          2586 => x"0b",
          2587 => x"f8",
          2588 => x"83",
          2589 => x"1a",
          2590 => x"ff",
          2591 => x"f9",
          2592 => x"5a",
          2593 => x"98",
          2594 => x"81",
          2595 => x"81",
          2596 => x"77",
          2597 => x"83",
          2598 => x"ff",
          2599 => x"a7",
          2600 => x"bc",
          2601 => x"ff",
          2602 => x"ff",
          2603 => x"43",
          2604 => x"86",
          2605 => x"bc",
          2606 => x"f6",
          2607 => x"5e",
          2608 => x"34",
          2609 => x"1e",
          2610 => x"a7",
          2611 => x"33",
          2612 => x"22",
          2613 => x"11",
          2614 => x"f4",
          2615 => x"81",
          2616 => x"79",
          2617 => x"f8",
          2618 => x"84",
          2619 => x"c8",
          2620 => x"fa",
          2621 => x"33",
          2622 => x"81",
          2623 => x"ca",
          2624 => x"80",
          2625 => x"0d",
          2626 => x"84",
          2627 => x"f8",
          2628 => x"f8",
          2629 => x"fc",
          2630 => x"3d",
          2631 => x"8a",
          2632 => x"2e",
          2633 => x"81",
          2634 => x"34",
          2635 => x"80",
          2636 => x"05",
          2637 => x"17",
          2638 => x"7b",
          2639 => x"bc",
          2640 => x"5c",
          2641 => x"83",
          2642 => x"72",
          2643 => x"b7",
          2644 => x"80",
          2645 => x"f8",
          2646 => x"71",
          2647 => x"83",
          2648 => x"33",
          2649 => x"f8",
          2650 => x"05",
          2651 => x"ff",
          2652 => x"f9",
          2653 => x"5a",
          2654 => x"98",
          2655 => x"ff",
          2656 => x"a2",
          2657 => x"90",
          2658 => x"f8",
          2659 => x"0c",
          2660 => x"2e",
          2661 => x"56",
          2662 => x"51",
          2663 => x"c8",
          2664 => x"b0",
          2665 => x"b1",
          2666 => x"b2",
          2667 => x"ff",
          2668 => x"b9",
          2669 => x"b9",
          2670 => x"b9",
          2671 => x"c9",
          2672 => x"38",
          2673 => x"2e",
          2674 => x"f8",
          2675 => x"f8",
          2676 => x"e4",
          2677 => x"fe",
          2678 => x"f2",
          2679 => x"06",
          2680 => x"41",
          2681 => x"52",
          2682 => x"3f",
          2683 => x"c9",
          2684 => x"5b",
          2685 => x"10",
          2686 => x"57",
          2687 => x"75",
          2688 => x"7e",
          2689 => x"7d",
          2690 => x"f8",
          2691 => x"31",
          2692 => x"5a",
          2693 => x"f8",
          2694 => x"33",
          2695 => x"84",
          2696 => x"ff",
          2697 => x"5f",
          2698 => x"83",
          2699 => x"0b",
          2700 => x"33",
          2701 => x"80",
          2702 => x"75",
          2703 => x"80",
          2704 => x"f8",
          2705 => x"57",
          2706 => x"81",
          2707 => x"fc",
          2708 => x"7f",
          2709 => x"f9",
          2710 => x"31",
          2711 => x"5a",
          2712 => x"f9",
          2713 => x"33",
          2714 => x"84",
          2715 => x"09",
          2716 => x"bc",
          2717 => x"f8",
          2718 => x"a0",
          2719 => x"51",
          2720 => x"83",
          2721 => x"87",
          2722 => x"5d",
          2723 => x"38",
          2724 => x"f2",
          2725 => x"80",
          2726 => x"22",
          2727 => x"fb",
          2728 => x"34",
          2729 => x"56",
          2730 => x"b9",
          2731 => x"7c",
          2732 => x"59",
          2733 => x"75",
          2734 => x"a2",
          2735 => x"80",
          2736 => x"33",
          2737 => x"84",
          2738 => x"56",
          2739 => x"76",
          2740 => x"83",
          2741 => x"80",
          2742 => x"76",
          2743 => x"84",
          2744 => x"83",
          2745 => x"81",
          2746 => x"c9",
          2747 => x"0b",
          2748 => x"80",
          2749 => x"56",
          2750 => x"81",
          2751 => x"f3",
          2752 => x"33",
          2753 => x"84",
          2754 => x"ff",
          2755 => x"70",
          2756 => x"70",
          2757 => x"52",
          2758 => x"83",
          2759 => x"23",
          2760 => x"5f",
          2761 => x"76",
          2762 => x"33",
          2763 => x"f9",
          2764 => x"f9",
          2765 => x"33",
          2766 => x"84",
          2767 => x"40",
          2768 => x"83",
          2769 => x"70",
          2770 => x"71",
          2771 => x"05",
          2772 => x"7e",
          2773 => x"83",
          2774 => x"5f",
          2775 => x"79",
          2776 => x"5d",
          2777 => x"84",
          2778 => x"8e",
          2779 => x"f8",
          2780 => x"7c",
          2781 => x"e5",
          2782 => x"76",
          2783 => x"75",
          2784 => x"06",
          2785 => x"5a",
          2786 => x"31",
          2787 => x"71",
          2788 => x"a7",
          2789 => x"7f",
          2790 => x"71",
          2791 => x"79",
          2792 => x"9a",
          2793 => x"84",
          2794 => x"05",
          2795 => x"33",
          2796 => x"18",
          2797 => x"33",
          2798 => x"58",
          2799 => x"e0",
          2800 => x"33",
          2801 => x"70",
          2802 => x"05",
          2803 => x"33",
          2804 => x"1d",
          2805 => x"ff",
          2806 => x"c9",
          2807 => x"38",
          2808 => x"d8",
          2809 => x"84",
          2810 => x"c9",
          2811 => x"2e",
          2812 => x"75",
          2813 => x"38",
          2814 => x"ff",
          2815 => x"5c",
          2816 => x"84",
          2817 => x"f6",
          2818 => x"60",
          2819 => x"26",
          2820 => x"f2",
          2821 => x"29",
          2822 => x"70",
          2823 => x"05",
          2824 => x"8b",
          2825 => x"8b",
          2826 => x"98",
          2827 => x"2b",
          2828 => x"5f",
          2829 => x"77",
          2830 => x"70",
          2831 => x"ee",
          2832 => x"bb",
          2833 => x"60",
          2834 => x"7d",
          2835 => x"5a",
          2836 => x"31",
          2837 => x"40",
          2838 => x"26",
          2839 => x"84",
          2840 => x"e0",
          2841 => x"05",
          2842 => x"26",
          2843 => x"19",
          2844 => x"34",
          2845 => x"38",
          2846 => x"ff",
          2847 => x"f8",
          2848 => x"84",
          2849 => x"07",
          2850 => x"09",
          2851 => x"83",
          2852 => x"ff",
          2853 => x"f8",
          2854 => x"1e",
          2855 => x"84",
          2856 => x"84",
          2857 => x"fa",
          2858 => x"07",
          2859 => x"18",
          2860 => x"fb",
          2861 => x"06",
          2862 => x"34",
          2863 => x"fb",
          2864 => x"f4",
          2865 => x"81",
          2866 => x"f8",
          2867 => x"33",
          2868 => x"83",
          2869 => x"f1",
          2870 => x"70",
          2871 => x"39",
          2872 => x"56",
          2873 => x"39",
          2874 => x"90",
          2875 => x"fe",
          2876 => x"ef",
          2877 => x"f8",
          2878 => x"f4",
          2879 => x"56",
          2880 => x"39",
          2881 => x"a0",
          2882 => x"fe",
          2883 => x"fe",
          2884 => x"f4",
          2885 => x"33",
          2886 => x"83",
          2887 => x"f8",
          2888 => x"56",
          2889 => x"39",
          2890 => x"56",
          2891 => x"39",
          2892 => x"56",
          2893 => x"39",
          2894 => x"56",
          2895 => x"39",
          2896 => x"80",
          2897 => x"34",
          2898 => x"81",
          2899 => x"f8",
          2900 => x"83",
          2901 => x"d2",
          2902 => x"b0",
          2903 => x"b1",
          2904 => x"b2",
          2905 => x"80",
          2906 => x"39",
          2907 => x"0b",
          2908 => x"04",
          2909 => x"f9",
          2910 => x"05",
          2911 => x"42",
          2912 => x"51",
          2913 => x"08",
          2914 => x"b8",
          2915 => x"34",
          2916 => x"3d",
          2917 => x"ef",
          2918 => x"11",
          2919 => x"7b",
          2920 => x"ca",
          2921 => x"80",
          2922 => x"80",
          2923 => x"81",
          2924 => x"33",
          2925 => x"56",
          2926 => x"f9",
          2927 => x"3f",
          2928 => x"d8",
          2929 => x"33",
          2930 => x"72",
          2931 => x"75",
          2932 => x"bc",
          2933 => x"38",
          2934 => x"39",
          2935 => x"09",
          2936 => x"57",
          2937 => x"81",
          2938 => x"59",
          2939 => x"38",
          2940 => x"bb",
          2941 => x"81",
          2942 => x"f8",
          2943 => x"ff",
          2944 => x"29",
          2945 => x"f8",
          2946 => x"05",
          2947 => x"ce",
          2948 => x"77",
          2949 => x"ff",
          2950 => x"7b",
          2951 => x"33",
          2952 => x"ff",
          2953 => x"7c",
          2954 => x"80",
          2955 => x"bb",
          2956 => x"38",
          2957 => x"34",
          2958 => x"22",
          2959 => x"90",
          2960 => x"81",
          2961 => x"5f",
          2962 => x"86",
          2963 => x"7f",
          2964 => x"41",
          2965 => x"ea",
          2966 => x"e0",
          2967 => x"33",
          2968 => x"70",
          2969 => x"05",
          2970 => x"33",
          2971 => x"1d",
          2972 => x"ec",
          2973 => x"84",
          2974 => x"05",
          2975 => x"33",
          2976 => x"18",
          2977 => x"33",
          2978 => x"58",
          2979 => x"fa",
          2980 => x"84",
          2981 => x"f8",
          2982 => x"f8",
          2983 => x"5c",
          2984 => x"d2",
          2985 => x"ff",
          2986 => x"61",
          2987 => x"f8",
          2988 => x"19",
          2989 => x"80",
          2990 => x"b7",
          2991 => x"12",
          2992 => x"8d",
          2993 => x"34",
          2994 => x"81",
          2995 => x"59",
          2996 => x"38",
          2997 => x"2e",
          2998 => x"f8",
          2999 => x"f8",
          3000 => x"76",
          3001 => x"38",
          3002 => x"83",
          3003 => x"1a",
          3004 => x"e7",
          3005 => x"f8",
          3006 => x"58",
          3007 => x"80",
          3008 => x"f8",
          3009 => x"34",
          3010 => x"76",
          3011 => x"f4",
          3012 => x"79",
          3013 => x"79",
          3014 => x"23",
          3015 => x"f8",
          3016 => x"f6",
          3017 => x"f8",
          3018 => x"83",
          3019 => x"f8",
          3020 => x"1a",
          3021 => x"cd",
          3022 => x"02",
          3023 => x"54",
          3024 => x"51",
          3025 => x"c8",
          3026 => x"73",
          3027 => x"b9",
          3028 => x"3d",
          3029 => x"0b",
          3030 => x"06",
          3031 => x"55",
          3032 => x"81",
          3033 => x"74",
          3034 => x"3d",
          3035 => x"82",
          3036 => x"73",
          3037 => x"70",
          3038 => x"83",
          3039 => x"7b",
          3040 => x"7b",
          3041 => x"80",
          3042 => x"80",
          3043 => x"33",
          3044 => x"33",
          3045 => x"80",
          3046 => x"5d",
          3047 => x"ff",
          3048 => x"55",
          3049 => x"81",
          3050 => x"34",
          3051 => x"87",
          3052 => x"2e",
          3053 => x"57",
          3054 => x"14",
          3055 => x"f9",
          3056 => x"f6",
          3057 => x"83",
          3058 => x"72",
          3059 => x"ff",
          3060 => x"fc",
          3061 => x"79",
          3062 => x"83",
          3063 => x"14",
          3064 => x"14",
          3065 => x"74",
          3066 => x"33",
          3067 => x"56",
          3068 => x"81",
          3069 => x"70",
          3070 => x"2e",
          3071 => x"a1",
          3072 => x"80",
          3073 => x"f7",
          3074 => x"33",
          3075 => x"33",
          3076 => x"a3",
          3077 => x"56",
          3078 => x"81",
          3079 => x"16",
          3080 => x"38",
          3081 => x"81",
          3082 => x"16",
          3083 => x"81",
          3084 => x"8d",
          3085 => x"72",
          3086 => x"ff",
          3087 => x"8c",
          3088 => x"81",
          3089 => x"9c",
          3090 => x"9c",
          3091 => x"ec",
          3092 => x"08",
          3093 => x"70",
          3094 => x"27",
          3095 => x"34",
          3096 => x"19",
          3097 => x"72",
          3098 => x"79",
          3099 => x"73",
          3100 => x"87",
          3101 => x"7d",
          3102 => x"f7",
          3103 => x"83",
          3104 => x"34",
          3105 => x"d0",
          3106 => x"81",
          3107 => x"33",
          3108 => x"34",
          3109 => x"f7",
          3110 => x"9c",
          3111 => x"80",
          3112 => x"8a",
          3113 => x"74",
          3114 => x"9b",
          3115 => x"83",
          3116 => x"38",
          3117 => x"81",
          3118 => x"98",
          3119 => x"38",
          3120 => x"70",
          3121 => x"06",
          3122 => x"53",
          3123 => x"38",
          3124 => x"76",
          3125 => x"d8",
          3126 => x"87",
          3127 => x"0c",
          3128 => x"81",
          3129 => x"06",
          3130 => x"9b",
          3131 => x"80",
          3132 => x"72",
          3133 => x"32",
          3134 => x"40",
          3135 => x"2e",
          3136 => x"ff",
          3137 => x"10",
          3138 => x"33",
          3139 => x"38",
          3140 => x"57",
          3141 => x"bf",
          3142 => x"38",
          3143 => x"91",
          3144 => x"51",
          3145 => x"0c",
          3146 => x"81",
          3147 => x"ff",
          3148 => x"33",
          3149 => x"15",
          3150 => x"f7",
          3151 => x"fc",
          3152 => x"15",
          3153 => x"06",
          3154 => x"38",
          3155 => x"75",
          3156 => x"06",
          3157 => x"fb",
          3158 => x"fa",
          3159 => x"55",
          3160 => x"c0",
          3161 => x"76",
          3162 => x"ff",
          3163 => x"ca",
          3164 => x"09",
          3165 => x"72",
          3166 => x"f7",
          3167 => x"f7",
          3168 => x"83",
          3169 => x"5c",
          3170 => x"2e",
          3171 => x"59",
          3172 => x"81",
          3173 => x"fd",
          3174 => x"54",
          3175 => x"bf",
          3176 => x"54",
          3177 => x"f7",
          3178 => x"33",
          3179 => x"73",
          3180 => x"95",
          3181 => x"84",
          3182 => x"f7",
          3183 => x"bb",
          3184 => x"57",
          3185 => x"80",
          3186 => x"81",
          3187 => x"73",
          3188 => x"f8",
          3189 => x"81",
          3190 => x"75",
          3191 => x"f8",
          3192 => x"81",
          3193 => x"ff",
          3194 => x"95",
          3195 => x"ac",
          3196 => x"83",
          3197 => x"59",
          3198 => x"51",
          3199 => x"fa",
          3200 => x"08",
          3201 => x"13",
          3202 => x"e0",
          3203 => x"08",
          3204 => x"80",
          3205 => x"c0",
          3206 => x"55",
          3207 => x"98",
          3208 => x"08",
          3209 => x"14",
          3210 => x"52",
          3211 => x"fe",
          3212 => x"08",
          3213 => x"c8",
          3214 => x"c0",
          3215 => x"ce",
          3216 => x"08",
          3217 => x"74",
          3218 => x"87",
          3219 => x"73",
          3220 => x"db",
          3221 => x"72",
          3222 => x"55",
          3223 => x"53",
          3224 => x"ff",
          3225 => x"ff",
          3226 => x"0c",
          3227 => x"b9",
          3228 => x"3d",
          3229 => x"33",
          3230 => x"08",
          3231 => x"06",
          3232 => x"55",
          3233 => x"2a",
          3234 => x"2a",
          3235 => x"15",
          3236 => x"82",
          3237 => x"80",
          3238 => x"d4",
          3239 => x"34",
          3240 => x"87",
          3241 => x"08",
          3242 => x"c0",
          3243 => x"9c",
          3244 => x"81",
          3245 => x"56",
          3246 => x"81",
          3247 => x"a4",
          3248 => x"80",
          3249 => x"80",
          3250 => x"80",
          3251 => x"9c",
          3252 => x"55",
          3253 => x"33",
          3254 => x"70",
          3255 => x"2e",
          3256 => x"55",
          3257 => x"71",
          3258 => x"57",
          3259 => x"74",
          3260 => x"38",
          3261 => x"75",
          3262 => x"80",
          3263 => x"92",
          3264 => x"71",
          3265 => x"26",
          3266 => x"88",
          3267 => x"c8",
          3268 => x"c2",
          3269 => x"05",
          3270 => x"83",
          3271 => x"fc",
          3272 => x"07",
          3273 => x"34",
          3274 => x"34",
          3275 => x"34",
          3276 => x"d4",
          3277 => x"56",
          3278 => x"38",
          3279 => x"70",
          3280 => x"f0",
          3281 => x"82",
          3282 => x"80",
          3283 => x"d4",
          3284 => x"34",
          3285 => x"87",
          3286 => x"08",
          3287 => x"c0",
          3288 => x"9c",
          3289 => x"81",
          3290 => x"56",
          3291 => x"81",
          3292 => x"a4",
          3293 => x"80",
          3294 => x"80",
          3295 => x"80",
          3296 => x"9c",
          3297 => x"55",
          3298 => x"33",
          3299 => x"70",
          3300 => x"2e",
          3301 => x"55",
          3302 => x"71",
          3303 => x"57",
          3304 => x"81",
          3305 => x"74",
          3306 => x"80",
          3307 => x"b9",
          3308 => x"51",
          3309 => x"d4",
          3310 => x"0b",
          3311 => x"0b",
          3312 => x"80",
          3313 => x"83",
          3314 => x"05",
          3315 => x"87",
          3316 => x"2e",
          3317 => x"98",
          3318 => x"87",
          3319 => x"87",
          3320 => x"70",
          3321 => x"71",
          3322 => x"98",
          3323 => x"87",
          3324 => x"98",
          3325 => x"38",
          3326 => x"08",
          3327 => x"71",
          3328 => x"98",
          3329 => x"38",
          3330 => x"81",
          3331 => x"8a",
          3332 => x"fe",
          3333 => x"83",
          3334 => x"82",
          3335 => x"b9",
          3336 => x"70",
          3337 => x"73",
          3338 => x"8b",
          3339 => x"70",
          3340 => x"71",
          3341 => x"53",
          3342 => x"80",
          3343 => x"82",
          3344 => x"2b",
          3345 => x"33",
          3346 => x"90",
          3347 => x"56",
          3348 => x"84",
          3349 => x"2b",
          3350 => x"88",
          3351 => x"13",
          3352 => x"87",
          3353 => x"17",
          3354 => x"88",
          3355 => x"59",
          3356 => x"85",
          3357 => x"52",
          3358 => x"87",
          3359 => x"74",
          3360 => x"84",
          3361 => x"12",
          3362 => x"80",
          3363 => x"52",
          3364 => x"89",
          3365 => x"13",
          3366 => x"07",
          3367 => x"33",
          3368 => x"58",
          3369 => x"84",
          3370 => x"b9",
          3371 => x"85",
          3372 => x"2b",
          3373 => x"86",
          3374 => x"2b",
          3375 => x"52",
          3376 => x"34",
          3377 => x"81",
          3378 => x"ff",
          3379 => x"54",
          3380 => x"34",
          3381 => x"33",
          3382 => x"83",
          3383 => x"12",
          3384 => x"2b",
          3385 => x"88",
          3386 => x"57",
          3387 => x"83",
          3388 => x"17",
          3389 => x"2b",
          3390 => x"33",
          3391 => x"81",
          3392 => x"52",
          3393 => x"73",
          3394 => x"b8",
          3395 => x"12",
          3396 => x"07",
          3397 => x"71",
          3398 => x"53",
          3399 => x"80",
          3400 => x"13",
          3401 => x"80",
          3402 => x"76",
          3403 => x"b9",
          3404 => x"12",
          3405 => x"07",
          3406 => x"33",
          3407 => x"57",
          3408 => x"72",
          3409 => x"89",
          3410 => x"84",
          3411 => x"2e",
          3412 => x"77",
          3413 => x"04",
          3414 => x"0c",
          3415 => x"82",
          3416 => x"f4",
          3417 => x"b8",
          3418 => x"81",
          3419 => x"76",
          3420 => x"34",
          3421 => x"17",
          3422 => x"b9",
          3423 => x"05",
          3424 => x"ff",
          3425 => x"56",
          3426 => x"34",
          3427 => x"10",
          3428 => x"55",
          3429 => x"83",
          3430 => x"0d",
          3431 => x"72",
          3432 => x"82",
          3433 => x"51",
          3434 => x"b8",
          3435 => x"71",
          3436 => x"58",
          3437 => x"2e",
          3438 => x"17",
          3439 => x"2b",
          3440 => x"31",
          3441 => x"27",
          3442 => x"74",
          3443 => x"38",
          3444 => x"85",
          3445 => x"5a",
          3446 => x"2e",
          3447 => x"76",
          3448 => x"12",
          3449 => x"ff",
          3450 => x"59",
          3451 => x"80",
          3452 => x"78",
          3453 => x"72",
          3454 => x"70",
          3455 => x"80",
          3456 => x"56",
          3457 => x"34",
          3458 => x"2a",
          3459 => x"83",
          3460 => x"19",
          3461 => x"2b",
          3462 => x"06",
          3463 => x"70",
          3464 => x"52",
          3465 => x"ff",
          3466 => x"b9",
          3467 => x"72",
          3468 => x"70",
          3469 => x"71",
          3470 => x"05",
          3471 => x"15",
          3472 => x"b8",
          3473 => x"11",
          3474 => x"07",
          3475 => x"70",
          3476 => x"84",
          3477 => x"33",
          3478 => x"83",
          3479 => x"5a",
          3480 => x"15",
          3481 => x"55",
          3482 => x"33",
          3483 => x"54",
          3484 => x"79",
          3485 => x"18",
          3486 => x"0c",
          3487 => x"87",
          3488 => x"2b",
          3489 => x"18",
          3490 => x"2a",
          3491 => x"84",
          3492 => x"b9",
          3493 => x"85",
          3494 => x"2b",
          3495 => x"15",
          3496 => x"2a",
          3497 => x"52",
          3498 => x"34",
          3499 => x"81",
          3500 => x"ff",
          3501 => x"54",
          3502 => x"34",
          3503 => x"51",
          3504 => x"84",
          3505 => x"2e",
          3506 => x"73",
          3507 => x"04",
          3508 => x"c8",
          3509 => x"0d",
          3510 => x"b8",
          3511 => x"23",
          3512 => x"ff",
          3513 => x"b9",
          3514 => x"0b",
          3515 => x"54",
          3516 => x"15",
          3517 => x"86",
          3518 => x"84",
          3519 => x"ff",
          3520 => x"ff",
          3521 => x"55",
          3522 => x"17",
          3523 => x"10",
          3524 => x"05",
          3525 => x"0b",
          3526 => x"2e",
          3527 => x"3d",
          3528 => x"84",
          3529 => x"61",
          3530 => x"85",
          3531 => x"38",
          3532 => x"7f",
          3533 => x"83",
          3534 => x"ff",
          3535 => x"70",
          3536 => x"7a",
          3537 => x"88",
          3538 => x"ff",
          3539 => x"05",
          3540 => x"81",
          3541 => x"90",
          3542 => x"46",
          3543 => x"59",
          3544 => x"85",
          3545 => x"33",
          3546 => x"10",
          3547 => x"98",
          3548 => x"53",
          3549 => x"c9",
          3550 => x"63",
          3551 => x"38",
          3552 => x"1b",
          3553 => x"63",
          3554 => x"38",
          3555 => x"71",
          3556 => x"11",
          3557 => x"2b",
          3558 => x"52",
          3559 => x"8c",
          3560 => x"83",
          3561 => x"2b",
          3562 => x"12",
          3563 => x"07",
          3564 => x"33",
          3565 => x"59",
          3566 => x"5c",
          3567 => x"85",
          3568 => x"17",
          3569 => x"8b",
          3570 => x"86",
          3571 => x"2b",
          3572 => x"52",
          3573 => x"34",
          3574 => x"08",
          3575 => x"88",
          3576 => x"88",
          3577 => x"34",
          3578 => x"08",
          3579 => x"33",
          3580 => x"74",
          3581 => x"88",
          3582 => x"45",
          3583 => x"34",
          3584 => x"08",
          3585 => x"71",
          3586 => x"05",
          3587 => x"88",
          3588 => x"45",
          3589 => x"1a",
          3590 => x"b8",
          3591 => x"12",
          3592 => x"62",
          3593 => x"5d",
          3594 => x"ec",
          3595 => x"05",
          3596 => x"ff",
          3597 => x"81",
          3598 => x"c8",
          3599 => x"f4",
          3600 => x"0b",
          3601 => x"53",
          3602 => x"c7",
          3603 => x"60",
          3604 => x"84",
          3605 => x"34",
          3606 => x"b8",
          3607 => x"0b",
          3608 => x"84",
          3609 => x"80",
          3610 => x"88",
          3611 => x"18",
          3612 => x"b4",
          3613 => x"b8",
          3614 => x"82",
          3615 => x"84",
          3616 => x"38",
          3617 => x"54",
          3618 => x"51",
          3619 => x"84",
          3620 => x"61",
          3621 => x"2b",
          3622 => x"33",
          3623 => x"81",
          3624 => x"44",
          3625 => x"81",
          3626 => x"05",
          3627 => x"19",
          3628 => x"b8",
          3629 => x"33",
          3630 => x"8f",
          3631 => x"ff",
          3632 => x"47",
          3633 => x"05",
          3634 => x"63",
          3635 => x"1e",
          3636 => x"34",
          3637 => x"05",
          3638 => x"bc",
          3639 => x"ff",
          3640 => x"81",
          3641 => x"ff",
          3642 => x"33",
          3643 => x"10",
          3644 => x"98",
          3645 => x"53",
          3646 => x"25",
          3647 => x"78",
          3648 => x"8b",
          3649 => x"5b",
          3650 => x"8f",
          3651 => x"b8",
          3652 => x"23",
          3653 => x"ff",
          3654 => x"b9",
          3655 => x"0b",
          3656 => x"59",
          3657 => x"1a",
          3658 => x"86",
          3659 => x"84",
          3660 => x"ff",
          3661 => x"ff",
          3662 => x"57",
          3663 => x"64",
          3664 => x"70",
          3665 => x"05",
          3666 => x"05",
          3667 => x"ee",
          3668 => x"61",
          3669 => x"27",
          3670 => x"80",
          3671 => x"fb",
          3672 => x"0c",
          3673 => x"11",
          3674 => x"71",
          3675 => x"33",
          3676 => x"83",
          3677 => x"85",
          3678 => x"88",
          3679 => x"58",
          3680 => x"05",
          3681 => x"b9",
          3682 => x"85",
          3683 => x"2b",
          3684 => x"15",
          3685 => x"2a",
          3686 => x"41",
          3687 => x"87",
          3688 => x"70",
          3689 => x"07",
          3690 => x"5f",
          3691 => x"81",
          3692 => x"1f",
          3693 => x"8b",
          3694 => x"73",
          3695 => x"07",
          3696 => x"43",
          3697 => x"81",
          3698 => x"1f",
          3699 => x"2b",
          3700 => x"14",
          3701 => x"07",
          3702 => x"40",
          3703 => x"60",
          3704 => x"70",
          3705 => x"71",
          3706 => x"70",
          3707 => x"05",
          3708 => x"84",
          3709 => x"83",
          3710 => x"39",
          3711 => x"0c",
          3712 => x"82",
          3713 => x"f4",
          3714 => x"b8",
          3715 => x"81",
          3716 => x"7f",
          3717 => x"34",
          3718 => x"15",
          3719 => x"b9",
          3720 => x"05",
          3721 => x"ff",
          3722 => x"5e",
          3723 => x"34",
          3724 => x"10",
          3725 => x"5c",
          3726 => x"83",
          3727 => x"7f",
          3728 => x"87",
          3729 => x"2b",
          3730 => x"1d",
          3731 => x"2a",
          3732 => x"61",
          3733 => x"34",
          3734 => x"11",
          3735 => x"71",
          3736 => x"33",
          3737 => x"70",
          3738 => x"56",
          3739 => x"78",
          3740 => x"08",
          3741 => x"88",
          3742 => x"88",
          3743 => x"34",
          3744 => x"08",
          3745 => x"71",
          3746 => x"05",
          3747 => x"2b",
          3748 => x"06",
          3749 => x"5d",
          3750 => x"82",
          3751 => x"b9",
          3752 => x"12",
          3753 => x"07",
          3754 => x"71",
          3755 => x"70",
          3756 => x"5a",
          3757 => x"81",
          3758 => x"5b",
          3759 => x"16",
          3760 => x"07",
          3761 => x"33",
          3762 => x"5e",
          3763 => x"1e",
          3764 => x"b8",
          3765 => x"12",
          3766 => x"07",
          3767 => x"33",
          3768 => x"44",
          3769 => x"7c",
          3770 => x"05",
          3771 => x"33",
          3772 => x"81",
          3773 => x"5b",
          3774 => x"16",
          3775 => x"70",
          3776 => x"71",
          3777 => x"81",
          3778 => x"83",
          3779 => x"63",
          3780 => x"59",
          3781 => x"7b",
          3782 => x"70",
          3783 => x"8b",
          3784 => x"70",
          3785 => x"07",
          3786 => x"5d",
          3787 => x"75",
          3788 => x"b9",
          3789 => x"83",
          3790 => x"2b",
          3791 => x"12",
          3792 => x"07",
          3793 => x"33",
          3794 => x"59",
          3795 => x"5d",
          3796 => x"79",
          3797 => x"70",
          3798 => x"71",
          3799 => x"05",
          3800 => x"88",
          3801 => x"5e",
          3802 => x"16",
          3803 => x"b8",
          3804 => x"71",
          3805 => x"70",
          3806 => x"79",
          3807 => x"b8",
          3808 => x"12",
          3809 => x"07",
          3810 => x"71",
          3811 => x"5c",
          3812 => x"79",
          3813 => x"b8",
          3814 => x"33",
          3815 => x"74",
          3816 => x"71",
          3817 => x"5c",
          3818 => x"82",
          3819 => x"b9",
          3820 => x"83",
          3821 => x"57",
          3822 => x"5a",
          3823 => x"b6",
          3824 => x"84",
          3825 => x"ff",
          3826 => x"39",
          3827 => x"8b",
          3828 => x"84",
          3829 => x"2b",
          3830 => x"43",
          3831 => x"63",
          3832 => x"08",
          3833 => x"33",
          3834 => x"74",
          3835 => x"71",
          3836 => x"41",
          3837 => x"64",
          3838 => x"34",
          3839 => x"81",
          3840 => x"ff",
          3841 => x"42",
          3842 => x"34",
          3843 => x"33",
          3844 => x"83",
          3845 => x"12",
          3846 => x"2b",
          3847 => x"88",
          3848 => x"45",
          3849 => x"83",
          3850 => x"1f",
          3851 => x"2b",
          3852 => x"33",
          3853 => x"81",
          3854 => x"5f",
          3855 => x"7d",
          3856 => x"ff",
          3857 => x"60",
          3858 => x"c8",
          3859 => x"2e",
          3860 => x"b9",
          3861 => x"73",
          3862 => x"7b",
          3863 => x"f9",
          3864 => x"b8",
          3865 => x"38",
          3866 => x"b9",
          3867 => x"51",
          3868 => x"54",
          3869 => x"38",
          3870 => x"08",
          3871 => x"b9",
          3872 => x"ff",
          3873 => x"80",
          3874 => x"80",
          3875 => x"fe",
          3876 => x"55",
          3877 => x"34",
          3878 => x"15",
          3879 => x"b9",
          3880 => x"81",
          3881 => x"08",
          3882 => x"80",
          3883 => x"70",
          3884 => x"88",
          3885 => x"b9",
          3886 => x"b9",
          3887 => x"76",
          3888 => x"34",
          3889 => x"38",
          3890 => x"8f",
          3891 => x"26",
          3892 => x"52",
          3893 => x"0d",
          3894 => x"33",
          3895 => x"38",
          3896 => x"c8",
          3897 => x"38",
          3898 => x"b9",
          3899 => x"c8",
          3900 => x"0d",
          3901 => x"05",
          3902 => x"76",
          3903 => x"17",
          3904 => x"55",
          3905 => x"87",
          3906 => x"52",
          3907 => x"c8",
          3908 => x"2e",
          3909 => x"54",
          3910 => x"38",
          3911 => x"80",
          3912 => x"74",
          3913 => x"04",
          3914 => x"ff",
          3915 => x"ff",
          3916 => x"7c",
          3917 => x"33",
          3918 => x"74",
          3919 => x"33",
          3920 => x"73",
          3921 => x"c0",
          3922 => x"76",
          3923 => x"08",
          3924 => x"a7",
          3925 => x"73",
          3926 => x"74",
          3927 => x"2e",
          3928 => x"84",
          3929 => x"84",
          3930 => x"06",
          3931 => x"ac",
          3932 => x"02",
          3933 => x"05",
          3934 => x"53",
          3935 => x"c4",
          3936 => x"83",
          3937 => x"c0",
          3938 => x"2e",
          3939 => x"70",
          3940 => x"84",
          3941 => x"88",
          3942 => x"c8",
          3943 => x"75",
          3944 => x"86",
          3945 => x"c0",
          3946 => x"38",
          3947 => x"51",
          3948 => x"c0",
          3949 => x"87",
          3950 => x"38",
          3951 => x"14",
          3952 => x"80",
          3953 => x"06",
          3954 => x"f6",
          3955 => x"19",
          3956 => x"2e",
          3957 => x"56",
          3958 => x"53",
          3959 => x"a3",
          3960 => x"83",
          3961 => x"0c",
          3962 => x"18",
          3963 => x"19",
          3964 => x"59",
          3965 => x"81",
          3966 => x"83",
          3967 => x"1a",
          3968 => x"c8",
          3969 => x"27",
          3970 => x"74",
          3971 => x"38",
          3972 => x"81",
          3973 => x"78",
          3974 => x"81",
          3975 => x"57",
          3976 => x"ee",
          3977 => x"56",
          3978 => x"34",
          3979 => x"d5",
          3980 => x"0b",
          3981 => x"34",
          3982 => x"e1",
          3983 => x"bb",
          3984 => x"19",
          3985 => x"34",
          3986 => x"80",
          3987 => x"18",
          3988 => x"74",
          3989 => x"34",
          3990 => x"19",
          3991 => x"a3",
          3992 => x"84",
          3993 => x"74",
          3994 => x"56",
          3995 => x"2a",
          3996 => x"18",
          3997 => x"5b",
          3998 => x"18",
          3999 => x"19",
          4000 => x"33",
          4001 => x"08",
          4002 => x"39",
          4003 => x"59",
          4004 => x"9c",
          4005 => x"58",
          4006 => x"0d",
          4007 => x"82",
          4008 => x"82",
          4009 => x"06",
          4010 => x"89",
          4011 => x"80",
          4012 => x"38",
          4013 => x"09",
          4014 => x"78",
          4015 => x"51",
          4016 => x"80",
          4017 => x"78",
          4018 => x"79",
          4019 => x"81",
          4020 => x"05",
          4021 => x"79",
          4022 => x"33",
          4023 => x"09",
          4024 => x"78",
          4025 => x"51",
          4026 => x"80",
          4027 => x"78",
          4028 => x"7a",
          4029 => x"70",
          4030 => x"71",
          4031 => x"79",
          4032 => x"84",
          4033 => x"75",
          4034 => x"b4",
          4035 => x"0b",
          4036 => x"7b",
          4037 => x"38",
          4038 => x"81",
          4039 => x"b9",
          4040 => x"59",
          4041 => x"fd",
          4042 => x"77",
          4043 => x"33",
          4044 => x"0c",
          4045 => x"83",
          4046 => x"75",
          4047 => x"b4",
          4048 => x"0b",
          4049 => x"7c",
          4050 => x"38",
          4051 => x"81",
          4052 => x"b9",
          4053 => x"59",
          4054 => x"fc",
          4055 => x"06",
          4056 => x"82",
          4057 => x"2b",
          4058 => x"88",
          4059 => x"fe",
          4060 => x"41",
          4061 => x"0d",
          4062 => x"b8",
          4063 => x"5c",
          4064 => x"c8",
          4065 => x"be",
          4066 => x"34",
          4067 => x"84",
          4068 => x"18",
          4069 => x"33",
          4070 => x"fd",
          4071 => x"a0",
          4072 => x"17",
          4073 => x"fd",
          4074 => x"53",
          4075 => x"52",
          4076 => x"08",
          4077 => x"38",
          4078 => x"b4",
          4079 => x"7c",
          4080 => x"17",
          4081 => x"38",
          4082 => x"39",
          4083 => x"17",
          4084 => x"f5",
          4085 => x"08",
          4086 => x"38",
          4087 => x"b4",
          4088 => x"b9",
          4089 => x"08",
          4090 => x"55",
          4091 => x"b8",
          4092 => x"18",
          4093 => x"33",
          4094 => x"a0",
          4095 => x"b8",
          4096 => x"5e",
          4097 => x"c8",
          4098 => x"cb",
          4099 => x"34",
          4100 => x"84",
          4101 => x"18",
          4102 => x"33",
          4103 => x"fb",
          4104 => x"a0",
          4105 => x"17",
          4106 => x"fa",
          4107 => x"a0",
          4108 => x"17",
          4109 => x"39",
          4110 => x"9f",
          4111 => x"5d",
          4112 => x"9c",
          4113 => x"38",
          4114 => x"38",
          4115 => x"81",
          4116 => x"c8",
          4117 => x"2a",
          4118 => x"b4",
          4119 => x"86",
          4120 => x"5d",
          4121 => x"fa",
          4122 => x"52",
          4123 => x"84",
          4124 => x"ff",
          4125 => x"79",
          4126 => x"83",
          4127 => x"ff",
          4128 => x"76",
          4129 => x"81",
          4130 => x"c8",
          4131 => x"2e",
          4132 => x"87",
          4133 => x"0b",
          4134 => x"2e",
          4135 => x"5b",
          4136 => x"84",
          4137 => x"19",
          4138 => x"3f",
          4139 => x"38",
          4140 => x"0c",
          4141 => x"82",
          4142 => x"11",
          4143 => x"0a",
          4144 => x"57",
          4145 => x"2a",
          4146 => x"2a",
          4147 => x"2a",
          4148 => x"83",
          4149 => x"2a",
          4150 => x"05",
          4151 => x"78",
          4152 => x"33",
          4153 => x"09",
          4154 => x"77",
          4155 => x"51",
          4156 => x"80",
          4157 => x"77",
          4158 => x"ac",
          4159 => x"05",
          4160 => x"57",
          4161 => x"7a",
          4162 => x"8f",
          4163 => x"34",
          4164 => x"2a",
          4165 => x"b4",
          4166 => x"83",
          4167 => x"19",
          4168 => x"f0",
          4169 => x"08",
          4170 => x"38",
          4171 => x"b4",
          4172 => x"a0",
          4173 => x"5c",
          4174 => x"82",
          4175 => x"e4",
          4176 => x"81",
          4177 => x"b9",
          4178 => x"56",
          4179 => x"fc",
          4180 => x"b8",
          4181 => x"8f",
          4182 => x"f0",
          4183 => x"74",
          4184 => x"fc",
          4185 => x"19",
          4186 => x"ef",
          4187 => x"08",
          4188 => x"38",
          4189 => x"b4",
          4190 => x"a0",
          4191 => x"59",
          4192 => x"38",
          4193 => x"09",
          4194 => x"76",
          4195 => x"51",
          4196 => x"39",
          4197 => x"53",
          4198 => x"3f",
          4199 => x"2e",
          4200 => x"b9",
          4201 => x"08",
          4202 => x"08",
          4203 => x"5f",
          4204 => x"19",
          4205 => x"06",
          4206 => x"53",
          4207 => x"e4",
          4208 => x"54",
          4209 => x"1a",
          4210 => x"5a",
          4211 => x"81",
          4212 => x"08",
          4213 => x"a8",
          4214 => x"b9",
          4215 => x"7d",
          4216 => x"55",
          4217 => x"fa",
          4218 => x"52",
          4219 => x"7b",
          4220 => x"1c",
          4221 => x"ec",
          4222 => x"7b",
          4223 => x"7c",
          4224 => x"76",
          4225 => x"79",
          4226 => x"58",
          4227 => x"83",
          4228 => x"11",
          4229 => x"7f",
          4230 => x"5d",
          4231 => x"56",
          4232 => x"5a",
          4233 => x"5b",
          4234 => x"f6",
          4235 => x"5c",
          4236 => x"08",
          4237 => x"76",
          4238 => x"94",
          4239 => x"2e",
          4240 => x"93",
          4241 => x"19",
          4242 => x"75",
          4243 => x"79",
          4244 => x"08",
          4245 => x"84",
          4246 => x"84",
          4247 => x"72",
          4248 => x"51",
          4249 => x"77",
          4250 => x"73",
          4251 => x"3d",
          4252 => x"84",
          4253 => x"52",
          4254 => x"74",
          4255 => x"84",
          4256 => x"08",
          4257 => x"84",
          4258 => x"57",
          4259 => x"19",
          4260 => x"75",
          4261 => x"58",
          4262 => x"a0",
          4263 => x"30",
          4264 => x"07",
          4265 => x"55",
          4266 => x"c8",
          4267 => x"08",
          4268 => x"73",
          4269 => x"73",
          4270 => x"80",
          4271 => x"52",
          4272 => x"c8",
          4273 => x"84",
          4274 => x"58",
          4275 => x"e3",
          4276 => x"08",
          4277 => x"74",
          4278 => x"1a",
          4279 => x"79",
          4280 => x"b9",
          4281 => x"0b",
          4282 => x"04",
          4283 => x"39",
          4284 => x"53",
          4285 => x"84",
          4286 => x"84",
          4287 => x"8c",
          4288 => x"2e",
          4289 => x"39",
          4290 => x"59",
          4291 => x"80",
          4292 => x"80",
          4293 => x"18",
          4294 => x"33",
          4295 => x"73",
          4296 => x"22",
          4297 => x"ac",
          4298 => x"19",
          4299 => x"72",
          4300 => x"13",
          4301 => x"17",
          4302 => x"75",
          4303 => x"04",
          4304 => x"3d",
          4305 => x"80",
          4306 => x"70",
          4307 => x"a5",
          4308 => x"fe",
          4309 => x"27",
          4310 => x"29",
          4311 => x"98",
          4312 => x"77",
          4313 => x"08",
          4314 => x"a4",
          4315 => x"27",
          4316 => x"84",
          4317 => x"38",
          4318 => x"cd",
          4319 => x"b9",
          4320 => x"3d",
          4321 => x"a0",
          4322 => x"7a",
          4323 => x"0c",
          4324 => x"80",
          4325 => x"5b",
          4326 => x"08",
          4327 => x"2a",
          4328 => x"27",
          4329 => x"79",
          4330 => x"9c",
          4331 => x"c8",
          4332 => x"18",
          4333 => x"89",
          4334 => x"52",
          4335 => x"c8",
          4336 => x"b9",
          4337 => x"84",
          4338 => x"9c",
          4339 => x"82",
          4340 => x"38",
          4341 => x"a7",
          4342 => x"56",
          4343 => x"9c",
          4344 => x"81",
          4345 => x"b9",
          4346 => x"84",
          4347 => x"58",
          4348 => x"1a",
          4349 => x"75",
          4350 => x"76",
          4351 => x"5e",
          4352 => x"84",
          4353 => x"81",
          4354 => x"f4",
          4355 => x"75",
          4356 => x"75",
          4357 => x"51",
          4358 => x"80",
          4359 => x"7a",
          4360 => x"c8",
          4361 => x"b4",
          4362 => x"81",
          4363 => x"84",
          4364 => x"b9",
          4365 => x"08",
          4366 => x"1a",
          4367 => x"33",
          4368 => x"fe",
          4369 => x"a0",
          4370 => x"19",
          4371 => x"39",
          4372 => x"ff",
          4373 => x"06",
          4374 => x"1d",
          4375 => x"80",
          4376 => x"8a",
          4377 => x"08",
          4378 => x"39",
          4379 => x"3d",
          4380 => x"41",
          4381 => x"ff",
          4382 => x"75",
          4383 => x"5f",
          4384 => x"76",
          4385 => x"78",
          4386 => x"06",
          4387 => x"b8",
          4388 => x"bd",
          4389 => x"85",
          4390 => x"1a",
          4391 => x"9c",
          4392 => x"80",
          4393 => x"bf",
          4394 => x"60",
          4395 => x"70",
          4396 => x"80",
          4397 => x"45",
          4398 => x"df",
          4399 => x"bf",
          4400 => x"81",
          4401 => x"f6",
          4402 => x"b9",
          4403 => x"08",
          4404 => x"b9",
          4405 => x"54",
          4406 => x"19",
          4407 => x"84",
          4408 => x"06",
          4409 => x"83",
          4410 => x"08",
          4411 => x"7a",
          4412 => x"82",
          4413 => x"81",
          4414 => x"19",
          4415 => x"52",
          4416 => x"77",
          4417 => x"09",
          4418 => x"2a",
          4419 => x"38",
          4420 => x"70",
          4421 => x"59",
          4422 => x"81",
          4423 => x"81",
          4424 => x"fe",
          4425 => x"0b",
          4426 => x"0c",
          4427 => x"df",
          4428 => x"2e",
          4429 => x"08",
          4430 => x"88",
          4431 => x"b7",
          4432 => x"8d",
          4433 => x"58",
          4434 => x"05",
          4435 => x"2b",
          4436 => x"80",
          4437 => x"87",
          4438 => x"42",
          4439 => x"17",
          4440 => x"33",
          4441 => x"77",
          4442 => x"26",
          4443 => x"43",
          4444 => x"ff",
          4445 => x"83",
          4446 => x"55",
          4447 => x"55",
          4448 => x"80",
          4449 => x"33",
          4450 => x"ff",
          4451 => x"74",
          4452 => x"ac",
          4453 => x"94",
          4454 => x"70",
          4455 => x"f5",
          4456 => x"84",
          4457 => x"ff",
          4458 => x"0c",
          4459 => x"80",
          4460 => x"cc",
          4461 => x"74",
          4462 => x"38",
          4463 => x"81",
          4464 => x"b9",
          4465 => x"56",
          4466 => x"5a",
          4467 => x"70",
          4468 => x"99",
          4469 => x"81",
          4470 => x"34",
          4471 => x"75",
          4472 => x"2e",
          4473 => x"75",
          4474 => x"38",
          4475 => x"81",
          4476 => x"70",
          4477 => x"70",
          4478 => x"5d",
          4479 => x"cd",
          4480 => x"76",
          4481 => x"57",
          4482 => x"70",
          4483 => x"ff",
          4484 => x"2e",
          4485 => x"38",
          4486 => x"0c",
          4487 => x"84",
          4488 => x"08",
          4489 => x"b9",
          4490 => x"54",
          4491 => x"1b",
          4492 => x"84",
          4493 => x"06",
          4494 => x"83",
          4495 => x"08",
          4496 => x"78",
          4497 => x"82",
          4498 => x"81",
          4499 => x"1b",
          4500 => x"52",
          4501 => x"77",
          4502 => x"e4",
          4503 => x"81",
          4504 => x"76",
          4505 => x"2e",
          4506 => x"bf",
          4507 => x"05",
          4508 => x"af",
          4509 => x"52",
          4510 => x"c8",
          4511 => x"2e",
          4512 => x"80",
          4513 => x"ff",
          4514 => x"8d",
          4515 => x"81",
          4516 => x"1a",
          4517 => x"07",
          4518 => x"78",
          4519 => x"05",
          4520 => x"e5",
          4521 => x"33",
          4522 => x"42",
          4523 => x"79",
          4524 => x"51",
          4525 => x"08",
          4526 => x"43",
          4527 => x"3f",
          4528 => x"81",
          4529 => x"18",
          4530 => x"78",
          4531 => x"59",
          4532 => x"2e",
          4533 => x"22",
          4534 => x"1d",
          4535 => x"ae",
          4536 => x"93",
          4537 => x"2e",
          4538 => x"94",
          4539 => x"70",
          4540 => x"5a",
          4541 => x"38",
          4542 => x"57",
          4543 => x"1d",
          4544 => x"5d",
          4545 => x"5b",
          4546 => x"75",
          4547 => x"81",
          4548 => x"ef",
          4549 => x"81",
          4550 => x"aa",
          4551 => x"81",
          4552 => x"08",
          4553 => x"57",
          4554 => x"76",
          4555 => x"55",
          4556 => x"c2",
          4557 => x"80",
          4558 => x"56",
          4559 => x"07",
          4560 => x"06",
          4561 => x"56",
          4562 => x"84",
          4563 => x"77",
          4564 => x"74",
          4565 => x"cf",
          4566 => x"06",
          4567 => x"15",
          4568 => x"19",
          4569 => x"e3",
          4570 => x"34",
          4571 => x"a0",
          4572 => x"98",
          4573 => x"88",
          4574 => x"57",
          4575 => x"38",
          4576 => x"26",
          4577 => x"05",
          4578 => x"74",
          4579 => x"38",
          4580 => x"c8",
          4581 => x"e3",
          4582 => x"7a",
          4583 => x"b9",
          4584 => x"84",
          4585 => x"02",
          4586 => x"7d",
          4587 => x"33",
          4588 => x"5f",
          4589 => x"8d",
          4590 => x"3f",
          4591 => x"52",
          4592 => x"c8",
          4593 => x"82",
          4594 => x"5e",
          4595 => x"b4",
          4596 => x"83",
          4597 => x"81",
          4598 => x"53",
          4599 => x"d4",
          4600 => x"2e",
          4601 => x"b4",
          4602 => x"9c",
          4603 => x"81",
          4604 => x"70",
          4605 => x"80",
          4606 => x"78",
          4607 => x"7d",
          4608 => x"08",
          4609 => x"ff",
          4610 => x"81",
          4611 => x"38",
          4612 => x"98",
          4613 => x"2e",
          4614 => x"40",
          4615 => x"53",
          4616 => x"d3",
          4617 => x"2e",
          4618 => x"b4",
          4619 => x"38",
          4620 => x"80",
          4621 => x"15",
          4622 => x"1f",
          4623 => x"81",
          4624 => x"59",
          4625 => x"9c",
          4626 => x"5e",
          4627 => x"83",
          4628 => x"c8",
          4629 => x"30",
          4630 => x"57",
          4631 => x"52",
          4632 => x"c8",
          4633 => x"2e",
          4634 => x"54",
          4635 => x"18",
          4636 => x"c8",
          4637 => x"bf",
          4638 => x"34",
          4639 => x"55",
          4640 => x"82",
          4641 => x"ac",
          4642 => x"9c",
          4643 => x"71",
          4644 => x"3f",
          4645 => x"c8",
          4646 => x"c8",
          4647 => x"2a",
          4648 => x"81",
          4649 => x"81",
          4650 => x"76",
          4651 => x"1d",
          4652 => x"56",
          4653 => x"83",
          4654 => x"81",
          4655 => x"53",
          4656 => x"d0",
          4657 => x"2e",
          4658 => x"b4",
          4659 => x"38",
          4660 => x"81",
          4661 => x"1c",
          4662 => x"8c",
          4663 => x"9b",
          4664 => x"76",
          4665 => x"ff",
          4666 => x"22",
          4667 => x"c8",
          4668 => x"70",
          4669 => x"56",
          4670 => x"ff",
          4671 => x"27",
          4672 => x"81",
          4673 => x"58",
          4674 => x"7c",
          4675 => x"80",
          4676 => x"b9",
          4677 => x"fc",
          4678 => x"fe",
          4679 => x"b4",
          4680 => x"81",
          4681 => x"81",
          4682 => x"38",
          4683 => x"b4",
          4684 => x"b9",
          4685 => x"08",
          4686 => x"42",
          4687 => x"bc",
          4688 => x"1d",
          4689 => x"33",
          4690 => x"a4",
          4691 => x"57",
          4692 => x"81",
          4693 => x"81",
          4694 => x"9f",
          4695 => x"07",
          4696 => x"1c",
          4697 => x"51",
          4698 => x"76",
          4699 => x"b9",
          4700 => x"08",
          4701 => x"1d",
          4702 => x"5f",
          4703 => x"c8",
          4704 => x"1c",
          4705 => x"38",
          4706 => x"e8",
          4707 => x"2e",
          4708 => x"54",
          4709 => x"53",
          4710 => x"ac",
          4711 => x"18",
          4712 => x"52",
          4713 => x"f8",
          4714 => x"71",
          4715 => x"1e",
          4716 => x"b5",
          4717 => x"d9",
          4718 => x"08",
          4719 => x"72",
          4720 => x"14",
          4721 => x"7a",
          4722 => x"70",
          4723 => x"8f",
          4724 => x"1a",
          4725 => x"5b",
          4726 => x"25",
          4727 => x"7c",
          4728 => x"18",
          4729 => x"58",
          4730 => x"18",
          4731 => x"38",
          4732 => x"89",
          4733 => x"25",
          4734 => x"38",
          4735 => x"70",
          4736 => x"74",
          4737 => x"18",
          4738 => x"7c",
          4739 => x"16",
          4740 => x"38",
          4741 => x"1e",
          4742 => x"56",
          4743 => x"08",
          4744 => x"38",
          4745 => x"53",
          4746 => x"1c",
          4747 => x"12",
          4748 => x"07",
          4749 => x"2b",
          4750 => x"97",
          4751 => x"2b",
          4752 => x"5b",
          4753 => x"33",
          4754 => x"5d",
          4755 => x"0d",
          4756 => x"77",
          4757 => x"58",
          4758 => x"2b",
          4759 => x"84",
          4760 => x"55",
          4761 => x"76",
          4762 => x"54",
          4763 => x"82",
          4764 => x"08",
          4765 => x"22",
          4766 => x"fd",
          4767 => x"78",
          4768 => x"58",
          4769 => x"7a",
          4770 => x"8c",
          4771 => x"73",
          4772 => x"80",
          4773 => x"7e",
          4774 => x"bf",
          4775 => x"38",
          4776 => x"5b",
          4777 => x"2a",
          4778 => x"2e",
          4779 => x"ff",
          4780 => x"05",
          4781 => x"19",
          4782 => x"56",
          4783 => x"39",
          4784 => x"7b",
          4785 => x"06",
          4786 => x"ef",
          4787 => x"57",
          4788 => x"53",
          4789 => x"74",
          4790 => x"80",
          4791 => x"88",
          4792 => x"3d",
          4793 => x"a7",
          4794 => x"80",
          4795 => x"33",
          4796 => x"7f",
          4797 => x"83",
          4798 => x"10",
          4799 => x"57",
          4800 => x"32",
          4801 => x"25",
          4802 => x"90",
          4803 => x"38",
          4804 => x"e4",
          4805 => x"81",
          4806 => x"2e",
          4807 => x"38",
          4808 => x"06",
          4809 => x"81",
          4810 => x"76",
          4811 => x"10",
          4812 => x"62",
          4813 => x"54",
          4814 => x"80",
          4815 => x"70",
          4816 => x"55",
          4817 => x"81",
          4818 => x"54",
          4819 => x"80",
          4820 => x"77",
          4821 => x"72",
          4822 => x"94",
          4823 => x"fe",
          4824 => x"73",
          4825 => x"c8",
          4826 => x"fe",
          4827 => x"c8",
          4828 => x"e4",
          4829 => x"7a",
          4830 => x"ff",
          4831 => x"7b",
          4832 => x"08",
          4833 => x"04",
          4834 => x"70",
          4835 => x"56",
          4836 => x"42",
          4837 => x"72",
          4838 => x"32",
          4839 => x"40",
          4840 => x"0c",
          4841 => x"81",
          4842 => x"83",
          4843 => x"2e",
          4844 => x"05",
          4845 => x"70",
          4846 => x"59",
          4847 => x"38",
          4848 => x"59",
          4849 => x"80",
          4850 => x"70",
          4851 => x"55",
          4852 => x"73",
          4853 => x"2e",
          4854 => x"38",
          4855 => x"54",
          4856 => x"18",
          4857 => x"80",
          4858 => x"5e",
          4859 => x"eb",
          4860 => x"a0",
          4861 => x"13",
          4862 => x"5e",
          4863 => x"59",
          4864 => x"ed",
          4865 => x"74",
          4866 => x"55",
          4867 => x"38",
          4868 => x"7b",
          4869 => x"32",
          4870 => x"70",
          4871 => x"80",
          4872 => x"86",
          4873 => x"79",
          4874 => x"38",
          4875 => x"2b",
          4876 => x"5d",
          4877 => x"56",
          4878 => x"33",
          4879 => x"38",
          4880 => x"8c",
          4881 => x"38",
          4882 => x"82",
          4883 => x"56",
          4884 => x"7c",
          4885 => x"5a",
          4886 => x"80",
          4887 => x"79",
          4888 => x"3f",
          4889 => x"56",
          4890 => x"81",
          4891 => x"2e",
          4892 => x"85",
          4893 => x"84",
          4894 => x"59",
          4895 => x"55",
          4896 => x"80",
          4897 => x"11",
          4898 => x"56",
          4899 => x"2e",
          4900 => x"fd",
          4901 => x"ae",
          4902 => x"77",
          4903 => x"06",
          4904 => x"80",
          4905 => x"53",
          4906 => x"a0",
          4907 => x"34",
          4908 => x"38",
          4909 => x"34",
          4910 => x"c8",
          4911 => x"b9",
          4912 => x"2a",
          4913 => x"86",
          4914 => x"56",
          4915 => x"90",
          4916 => x"80",
          4917 => x"71",
          4918 => x"54",
          4919 => x"74",
          4920 => x"56",
          4921 => x"ae",
          4922 => x"76",
          4923 => x"83",
          4924 => x"39",
          4925 => x"8c",
          4926 => x"81",
          4927 => x"5a",
          4928 => x"34",
          4929 => x"f6",
          4930 => x"1d",
          4931 => x"93",
          4932 => x"9d",
          4933 => x"38",
          4934 => x"f7",
          4935 => x"57",
          4936 => x"07",
          4937 => x"85",
          4938 => x"ff",
          4939 => x"5a",
          4940 => x"80",
          4941 => x"56",
          4942 => x"38",
          4943 => x"e4",
          4944 => x"81",
          4945 => x"2e",
          4946 => x"38",
          4947 => x"06",
          4948 => x"81",
          4949 => x"ff",
          4950 => x"38",
          4951 => x"5f",
          4952 => x"26",
          4953 => x"ff",
          4954 => x"06",
          4955 => x"05",
          4956 => x"75",
          4957 => x"fa",
          4958 => x"81",
          4959 => x"ff",
          4960 => x"7d",
          4961 => x"79",
          4962 => x"cd",
          4963 => x"98",
          4964 => x"88",
          4965 => x"7b",
          4966 => x"54",
          4967 => x"a0",
          4968 => x"1b",
          4969 => x"a0",
          4970 => x"2e",
          4971 => x"a3",
          4972 => x"7b",
          4973 => x"c8",
          4974 => x"0d",
          4975 => x"05",
          4976 => x"ff",
          4977 => x"80",
          4978 => x"05",
          4979 => x"75",
          4980 => x"38",
          4981 => x"d1",
          4982 => x"b2",
          4983 => x"05",
          4984 => x"80",
          4985 => x"7f",
          4986 => x"7b",
          4987 => x"51",
          4988 => x"08",
          4989 => x"58",
          4990 => x"77",
          4991 => x"1d",
          4992 => x"17",
          4993 => x"b9",
          4994 => x"06",
          4995 => x"38",
          4996 => x"2a",
          4997 => x"b1",
          4998 => x"ff",
          4999 => x"55",
          5000 => x"53",
          5001 => x"95",
          5002 => x"85",
          5003 => x"18",
          5004 => x"b7",
          5005 => x"88",
          5006 => x"82",
          5007 => x"81",
          5008 => x"33",
          5009 => x"75",
          5010 => x"75",
          5011 => x"17",
          5012 => x"2b",
          5013 => x"09",
          5014 => x"17",
          5015 => x"2b",
          5016 => x"dc",
          5017 => x"71",
          5018 => x"14",
          5019 => x"33",
          5020 => x"5f",
          5021 => x"17",
          5022 => x"33",
          5023 => x"40",
          5024 => x"d9",
          5025 => x"29",
          5026 => x"77",
          5027 => x"2e",
          5028 => x"42",
          5029 => x"33",
          5030 => x"07",
          5031 => x"75",
          5032 => x"82",
          5033 => x"cb",
          5034 => x"5c",
          5035 => x"11",
          5036 => x"71",
          5037 => x"72",
          5038 => x"53",
          5039 => x"c7",
          5040 => x"88",
          5041 => x"80",
          5042 => x"84",
          5043 => x"c1",
          5044 => x"fd",
          5045 => x"56",
          5046 => x"a9",
          5047 => x"ff",
          5048 => x"75",
          5049 => x"5d",
          5050 => x"81",
          5051 => x"7b",
          5052 => x"1a",
          5053 => x"59",
          5054 => x"17",
          5055 => x"80",
          5056 => x"78",
          5057 => x"78",
          5058 => x"06",
          5059 => x"2a",
          5060 => x"26",
          5061 => x"ff",
          5062 => x"84",
          5063 => x"38",
          5064 => x"81",
          5065 => x"7c",
          5066 => x"8c",
          5067 => x"80",
          5068 => x"3d",
          5069 => x"0c",
          5070 => x"11",
          5071 => x"74",
          5072 => x"81",
          5073 => x"7a",
          5074 => x"83",
          5075 => x"7f",
          5076 => x"33",
          5077 => x"9f",
          5078 => x"89",
          5079 => x"57",
          5080 => x"26",
          5081 => x"06",
          5082 => x"59",
          5083 => x"85",
          5084 => x"32",
          5085 => x"7a",
          5086 => x"87",
          5087 => x"5c",
          5088 => x"56",
          5089 => x"cf",
          5090 => x"8a",
          5091 => x"fe",
          5092 => x"75",
          5093 => x"38",
          5094 => x"30",
          5095 => x"5c",
          5096 => x"2e",
          5097 => x"5a",
          5098 => x"59",
          5099 => x"81",
          5100 => x"90",
          5101 => x"19",
          5102 => x"fe",
          5103 => x"40",
          5104 => x"5c",
          5105 => x"78",
          5106 => x"bd",
          5107 => x"72",
          5108 => x"05",
          5109 => x"52",
          5110 => x"56",
          5111 => x"0b",
          5112 => x"0c",
          5113 => x"a5",
          5114 => x"52",
          5115 => x"3f",
          5116 => x"38",
          5117 => x"0c",
          5118 => x"33",
          5119 => x"5e",
          5120 => x"09",
          5121 => x"18",
          5122 => x"82",
          5123 => x"30",
          5124 => x"42",
          5125 => x"b6",
          5126 => x"56",
          5127 => x"5d",
          5128 => x"83",
          5129 => x"bd",
          5130 => x"81",
          5131 => x"27",
          5132 => x"0b",
          5133 => x"5d",
          5134 => x"7e",
          5135 => x"31",
          5136 => x"80",
          5137 => x"e1",
          5138 => x"e4",
          5139 => x"05",
          5140 => x"33",
          5141 => x"42",
          5142 => x"75",
          5143 => x"f3",
          5144 => x"77",
          5145 => x"04",
          5146 => x"38",
          5147 => x"fc",
          5148 => x"0b",
          5149 => x"04",
          5150 => x"f8",
          5151 => x"5a",
          5152 => x"71",
          5153 => x"5f",
          5154 => x"80",
          5155 => x"18",
          5156 => x"70",
          5157 => x"05",
          5158 => x"5b",
          5159 => x"91",
          5160 => x"3d",
          5161 => x"39",
          5162 => x"17",
          5163 => x"2b",
          5164 => x"81",
          5165 => x"80",
          5166 => x"38",
          5167 => x"09",
          5168 => x"77",
          5169 => x"51",
          5170 => x"08",
          5171 => x"5a",
          5172 => x"38",
          5173 => x"33",
          5174 => x"07",
          5175 => x"09",
          5176 => x"83",
          5177 => x"2b",
          5178 => x"70",
          5179 => x"07",
          5180 => x"77",
          5181 => x"81",
          5182 => x"83",
          5183 => x"2b",
          5184 => x"70",
          5185 => x"07",
          5186 => x"60",
          5187 => x"81",
          5188 => x"83",
          5189 => x"2b",
          5190 => x"70",
          5191 => x"07",
          5192 => x"83",
          5193 => x"2b",
          5194 => x"70",
          5195 => x"07",
          5196 => x"46",
          5197 => x"7c",
          5198 => x"05",
          5199 => x"86",
          5200 => x"18",
          5201 => x"cf",
          5202 => x"7b",
          5203 => x"75",
          5204 => x"70",
          5205 => x"af",
          5206 => x"2e",
          5207 => x"b9",
          5208 => x"08",
          5209 => x"18",
          5210 => x"41",
          5211 => x"b9",
          5212 => x"56",
          5213 => x"0b",
          5214 => x"5a",
          5215 => x"33",
          5216 => x"07",
          5217 => x"38",
          5218 => x"38",
          5219 => x"12",
          5220 => x"07",
          5221 => x"2b",
          5222 => x"5a",
          5223 => x"59",
          5224 => x"80",
          5225 => x"e3",
          5226 => x"93",
          5227 => x"f2",
          5228 => x"fc",
          5229 => x"a0",
          5230 => x"17",
          5231 => x"85",
          5232 => x"05",
          5233 => x"57",
          5234 => x"2e",
          5235 => x"5a",
          5236 => x"ba",
          5237 => x"74",
          5238 => x"a4",
          5239 => x"38",
          5240 => x"70",
          5241 => x"38",
          5242 => x"2e",
          5243 => x"73",
          5244 => x"92",
          5245 => x"84",
          5246 => x"c8",
          5247 => x"92",
          5248 => x"c8",
          5249 => x"d0",
          5250 => x"57",
          5251 => x"77",
          5252 => x"77",
          5253 => x"08",
          5254 => x"08",
          5255 => x"5b",
          5256 => x"ff",
          5257 => x"26",
          5258 => x"06",
          5259 => x"99",
          5260 => x"ff",
          5261 => x"2a",
          5262 => x"06",
          5263 => x"79",
          5264 => x"2a",
          5265 => x"2e",
          5266 => x"5b",
          5267 => x"54",
          5268 => x"38",
          5269 => x"39",
          5270 => x"80",
          5271 => x"78",
          5272 => x"70",
          5273 => x"3d",
          5274 => x"84",
          5275 => x"08",
          5276 => x"76",
          5277 => x"3d",
          5278 => x"3d",
          5279 => x"b9",
          5280 => x"80",
          5281 => x"5d",
          5282 => x"80",
          5283 => x"83",
          5284 => x"ff",
          5285 => x"5b",
          5286 => x"9b",
          5287 => x"2b",
          5288 => x"5e",
          5289 => x"80",
          5290 => x"17",
          5291 => x"cc",
          5292 => x"0b",
          5293 => x"80",
          5294 => x"17",
          5295 => x"84",
          5296 => x"1c",
          5297 => x"0b",
          5298 => x"34",
          5299 => x"7b",
          5300 => x"11",
          5301 => x"57",
          5302 => x"08",
          5303 => x"80",
          5304 => x"e7",
          5305 => x"7b",
          5306 => x"9c",
          5307 => x"76",
          5308 => x"33",
          5309 => x"7b",
          5310 => x"06",
          5311 => x"81",
          5312 => x"83",
          5313 => x"86",
          5314 => x"b4",
          5315 => x"1b",
          5316 => x"33",
          5317 => x"5e",
          5318 => x"f1",
          5319 => x"83",
          5320 => x"2b",
          5321 => x"70",
          5322 => x"07",
          5323 => x"0c",
          5324 => x"86",
          5325 => x"1a",
          5326 => x"0b",
          5327 => x"06",
          5328 => x"75",
          5329 => x"1a",
          5330 => x"7c",
          5331 => x"07",
          5332 => x"84",
          5333 => x"5b",
          5334 => x"52",
          5335 => x"b9",
          5336 => x"81",
          5337 => x"c8",
          5338 => x"7a",
          5339 => x"05",
          5340 => x"77",
          5341 => x"2e",
          5342 => x"0c",
          5343 => x"0c",
          5344 => x"0c",
          5345 => x"3f",
          5346 => x"59",
          5347 => x"39",
          5348 => x"f3",
          5349 => x"71",
          5350 => x"07",
          5351 => x"55",
          5352 => x"52",
          5353 => x"b9",
          5354 => x"80",
          5355 => x"08",
          5356 => x"c8",
          5357 => x"53",
          5358 => x"3f",
          5359 => x"9c",
          5360 => x"58",
          5361 => x"38",
          5362 => x"33",
          5363 => x"7c",
          5364 => x"80",
          5365 => x"80",
          5366 => x"95",
          5367 => x"2b",
          5368 => x"56",
          5369 => x"0b",
          5370 => x"34",
          5371 => x"56",
          5372 => x"57",
          5373 => x"0b",
          5374 => x"83",
          5375 => x"ff",
          5376 => x"59",
          5377 => x"ae",
          5378 => x"2e",
          5379 => x"7d",
          5380 => x"51",
          5381 => x"08",
          5382 => x"5b",
          5383 => x"ff",
          5384 => x"2e",
          5385 => x"97",
          5386 => x"b8",
          5387 => x"5a",
          5388 => x"08",
          5389 => x"38",
          5390 => x"b4",
          5391 => x"b9",
          5392 => x"08",
          5393 => x"55",
          5394 => x"85",
          5395 => x"17",
          5396 => x"33",
          5397 => x"fe",
          5398 => x"56",
          5399 => x"76",
          5400 => x"5a",
          5401 => x"fe",
          5402 => x"59",
          5403 => x"8a",
          5404 => x"08",
          5405 => x"cd",
          5406 => x"0c",
          5407 => x"1a",
          5408 => x"57",
          5409 => x"b9",
          5410 => x"cf",
          5411 => x"39",
          5412 => x"40",
          5413 => x"57",
          5414 => x"56",
          5415 => x"55",
          5416 => x"22",
          5417 => x"2e",
          5418 => x"76",
          5419 => x"33",
          5420 => x"33",
          5421 => x"2e",
          5422 => x"1b",
          5423 => x"26",
          5424 => x"d5",
          5425 => x"5b",
          5426 => x"ff",
          5427 => x"9b",
          5428 => x"08",
          5429 => x"74",
          5430 => x"1b",
          5431 => x"05",
          5432 => x"76",
          5433 => x"22",
          5434 => x"56",
          5435 => x"7a",
          5436 => x"80",
          5437 => x"75",
          5438 => x"58",
          5439 => x"19",
          5440 => x"b9",
          5441 => x"11",
          5442 => x"38",
          5443 => x"78",
          5444 => x"29",
          5445 => x"70",
          5446 => x"05",
          5447 => x"38",
          5448 => x"7e",
          5449 => x"1c",
          5450 => x"5e",
          5451 => x"75",
          5452 => x"04",
          5453 => x"0d",
          5454 => x"1a",
          5455 => x"80",
          5456 => x"83",
          5457 => x"08",
          5458 => x"1a",
          5459 => x"2e",
          5460 => x"54",
          5461 => x"33",
          5462 => x"c8",
          5463 => x"81",
          5464 => x"dc",
          5465 => x"06",
          5466 => x"56",
          5467 => x"74",
          5468 => x"81",
          5469 => x"80",
          5470 => x"05",
          5471 => x"34",
          5472 => x"bc",
          5473 => x"b8",
          5474 => x"40",
          5475 => x"b9",
          5476 => x"ff",
          5477 => x"1a",
          5478 => x"31",
          5479 => x"a0",
          5480 => x"19",
          5481 => x"06",
          5482 => x"08",
          5483 => x"81",
          5484 => x"7e",
          5485 => x"0c",
          5486 => x"98",
          5487 => x"98",
          5488 => x"a1",
          5489 => x"83",
          5490 => x"55",
          5491 => x"56",
          5492 => x"1b",
          5493 => x"92",
          5494 => x"34",
          5495 => x"3d",
          5496 => x"67",
          5497 => x"0c",
          5498 => x"79",
          5499 => x"75",
          5500 => x"86",
          5501 => x"78",
          5502 => x"74",
          5503 => x"91",
          5504 => x"90",
          5505 => x"58",
          5506 => x"a1",
          5507 => x"57",
          5508 => x"5b",
          5509 => x"83",
          5510 => x"60",
          5511 => x"2a",
          5512 => x"84",
          5513 => x"80",
          5514 => x"86",
          5515 => x"38",
          5516 => x"85",
          5517 => x"b4",
          5518 => x"d3",
          5519 => x"17",
          5520 => x"27",
          5521 => x"79",
          5522 => x"74",
          5523 => x"7b",
          5524 => x"83",
          5525 => x"27",
          5526 => x"54",
          5527 => x"51",
          5528 => x"08",
          5529 => x"7d",
          5530 => x"38",
          5531 => x"29",
          5532 => x"05",
          5533 => x"34",
          5534 => x"59",
          5535 => x"59",
          5536 => x"0c",
          5537 => x"71",
          5538 => x"5a",
          5539 => x"38",
          5540 => x"fe",
          5541 => x"80",
          5542 => x"80",
          5543 => x"3d",
          5544 => x"92",
          5545 => x"74",
          5546 => x"39",
          5547 => x"83",
          5548 => x"5c",
          5549 => x"77",
          5550 => x"38",
          5551 => x"41",
          5552 => x"80",
          5553 => x"16",
          5554 => x"cd",
          5555 => x"85",
          5556 => x"17",
          5557 => x"1b",
          5558 => x"b8",
          5559 => x"2e",
          5560 => x"33",
          5561 => x"16",
          5562 => x"0b",
          5563 => x"54",
          5564 => x"53",
          5565 => x"f4",
          5566 => x"7f",
          5567 => x"84",
          5568 => x"16",
          5569 => x"c8",
          5570 => x"27",
          5571 => x"74",
          5572 => x"38",
          5573 => x"08",
          5574 => x"51",
          5575 => x"ca",
          5576 => x"08",
          5577 => x"40",
          5578 => x"12",
          5579 => x"7c",
          5580 => x"98",
          5581 => x"e7",
          5582 => x"b9",
          5583 => x"33",
          5584 => x"51",
          5585 => x"08",
          5586 => x"38",
          5587 => x"53",
          5588 => x"52",
          5589 => x"c8",
          5590 => x"08",
          5591 => x"17",
          5592 => x"27",
          5593 => x"7b",
          5594 => x"38",
          5595 => x"08",
          5596 => x"51",
          5597 => x"89",
          5598 => x"9b",
          5599 => x"55",
          5600 => x"56",
          5601 => x"16",
          5602 => x"17",
          5603 => x"84",
          5604 => x"b9",
          5605 => x"08",
          5606 => x"17",
          5607 => x"33",
          5608 => x"fe",
          5609 => x"a0",
          5610 => x"16",
          5611 => x"7c",
          5612 => x"56",
          5613 => x"34",
          5614 => x"3d",
          5615 => x"82",
          5616 => x"0d",
          5617 => x"5a",
          5618 => x"56",
          5619 => x"55",
          5620 => x"22",
          5621 => x"2e",
          5622 => x"79",
          5623 => x"33",
          5624 => x"7a",
          5625 => x"19",
          5626 => x"2e",
          5627 => x"81",
          5628 => x"17",
          5629 => x"f5",
          5630 => x"85",
          5631 => x"18",
          5632 => x"08",
          5633 => x"78",
          5634 => x"08",
          5635 => x"56",
          5636 => x"5a",
          5637 => x"33",
          5638 => x"2e",
          5639 => x"74",
          5640 => x"9d",
          5641 => x"9e",
          5642 => x"9f",
          5643 => x"97",
          5644 => x"80",
          5645 => x"92",
          5646 => x"7b",
          5647 => x"51",
          5648 => x"08",
          5649 => x"56",
          5650 => x"c8",
          5651 => x"b4",
          5652 => x"81",
          5653 => x"3f",
          5654 => x"c9",
          5655 => x"34",
          5656 => x"84",
          5657 => x"18",
          5658 => x"33",
          5659 => x"fe",
          5660 => x"a0",
          5661 => x"17",
          5662 => x"56",
          5663 => x"74",
          5664 => x"75",
          5665 => x"74",
          5666 => x"9d",
          5667 => x"9e",
          5668 => x"9f",
          5669 => x"97",
          5670 => x"80",
          5671 => x"92",
          5672 => x"7b",
          5673 => x"51",
          5674 => x"08",
          5675 => x"56",
          5676 => x"81",
          5677 => x"84",
          5678 => x"fc",
          5679 => x"fc",
          5680 => x"52",
          5681 => x"08",
          5682 => x"89",
          5683 => x"08",
          5684 => x"33",
          5685 => x"13",
          5686 => x"77",
          5687 => x"75",
          5688 => x"73",
          5689 => x"04",
          5690 => x"3f",
          5691 => x"72",
          5692 => x"d5",
          5693 => x"5b",
          5694 => x"75",
          5695 => x"26",
          5696 => x"70",
          5697 => x"84",
          5698 => x"90",
          5699 => x"0b",
          5700 => x"04",
          5701 => x"3d",
          5702 => x"81",
          5703 => x"26",
          5704 => x"06",
          5705 => x"80",
          5706 => x"5b",
          5707 => x"70",
          5708 => x"05",
          5709 => x"52",
          5710 => x"70",
          5711 => x"13",
          5712 => x"13",
          5713 => x"30",
          5714 => x"2e",
          5715 => x"be",
          5716 => x"72",
          5717 => x"52",
          5718 => x"84",
          5719 => x"99",
          5720 => x"83",
          5721 => x"fe",
          5722 => x"98",
          5723 => x"d1",
          5724 => x"84",
          5725 => x"74",
          5726 => x"04",
          5727 => x"05",
          5728 => x"08",
          5729 => x"38",
          5730 => x"2b",
          5731 => x"38",
          5732 => x"81",
          5733 => x"38",
          5734 => x"33",
          5735 => x"5a",
          5736 => x"38",
          5737 => x"c8",
          5738 => x"c8",
          5739 => x"8f",
          5740 => x"98",
          5741 => x"17",
          5742 => x"07",
          5743 => x"cc",
          5744 => x"74",
          5745 => x"04",
          5746 => x"08",
          5747 => x"7c",
          5748 => x"b4",
          5749 => x"c5",
          5750 => x"b9",
          5751 => x"d9",
          5752 => x"80",
          5753 => x"08",
          5754 => x"38",
          5755 => x"a0",
          5756 => x"84",
          5757 => x"08",
          5758 => x"08",
          5759 => x"b1",
          5760 => x"33",
          5761 => x"54",
          5762 => x"33",
          5763 => x"c8",
          5764 => x"81",
          5765 => x"d4",
          5766 => x"33",
          5767 => x"63",
          5768 => x"78",
          5769 => x"db",
          5770 => x"a3",
          5771 => x"84",
          5772 => x"52",
          5773 => x"b9",
          5774 => x"bb",
          5775 => x"33",
          5776 => x"63",
          5777 => x"7d",
          5778 => x"2e",
          5779 => x"7a",
          5780 => x"c8",
          5781 => x"2e",
          5782 => x"d8",
          5783 => x"3d",
          5784 => x"bd",
          5785 => x"5b",
          5786 => x"1f",
          5787 => x"5f",
          5788 => x"56",
          5789 => x"80",
          5790 => x"56",
          5791 => x"ff",
          5792 => x"75",
          5793 => x"18",
          5794 => x"af",
          5795 => x"79",
          5796 => x"8a",
          5797 => x"70",
          5798 => x"08",
          5799 => x"7e",
          5800 => x"17",
          5801 => x"38",
          5802 => x"38",
          5803 => x"76",
          5804 => x"05",
          5805 => x"26",
          5806 => x"5e",
          5807 => x"81",
          5808 => x"78",
          5809 => x"0d",
          5810 => x"71",
          5811 => x"07",
          5812 => x"16",
          5813 => x"71",
          5814 => x"3d",
          5815 => x"ff",
          5816 => x"59",
          5817 => x"96",
          5818 => x"16",
          5819 => x"17",
          5820 => x"81",
          5821 => x"38",
          5822 => x"b4",
          5823 => x"b9",
          5824 => x"08",
          5825 => x"55",
          5826 => x"f6",
          5827 => x"17",
          5828 => x"33",
          5829 => x"fb",
          5830 => x"08",
          5831 => x"0b",
          5832 => x"83",
          5833 => x"43",
          5834 => x"09",
          5835 => x"39",
          5836 => x"59",
          5837 => x"5e",
          5838 => x"80",
          5839 => x"5a",
          5840 => x"34",
          5841 => x"39",
          5842 => x"b9",
          5843 => x"f7",
          5844 => x"56",
          5845 => x"54",
          5846 => x"53",
          5847 => x"22",
          5848 => x"2e",
          5849 => x"75",
          5850 => x"33",
          5851 => x"08",
          5852 => x"94",
          5853 => x"2e",
          5854 => x"70",
          5855 => x"2e",
          5856 => x"51",
          5857 => x"08",
          5858 => x"53",
          5859 => x"08",
          5860 => x"74",
          5861 => x"31",
          5862 => x"80",
          5863 => x"81",
          5864 => x"08",
          5865 => x"70",
          5866 => x"78",
          5867 => x"74",
          5868 => x"c8",
          5869 => x"2e",
          5870 => x"38",
          5871 => x"53",
          5872 => x"38",
          5873 => x"81",
          5874 => x"84",
          5875 => x"90",
          5876 => x"55",
          5877 => x"16",
          5878 => x"2e",
          5879 => x"94",
          5880 => x"74",
          5881 => x"90",
          5882 => x"90",
          5883 => x"78",
          5884 => x"78",
          5885 => x"80",
          5886 => x"0d",
          5887 => x"15",
          5888 => x"38",
          5889 => x"80",
          5890 => x"c8",
          5891 => x"16",
          5892 => x"80",
          5893 => x"12",
          5894 => x"78",
          5895 => x"74",
          5896 => x"89",
          5897 => x"2e",
          5898 => x"fe",
          5899 => x"89",
          5900 => x"fe",
          5901 => x"82",
          5902 => x"06",
          5903 => x"08",
          5904 => x"74",
          5905 => x"c8",
          5906 => x"2e",
          5907 => x"2e",
          5908 => x"88",
          5909 => x"dc",
          5910 => x"0b",
          5911 => x"04",
          5912 => x"75",
          5913 => x"3d",
          5914 => x"51",
          5915 => x"55",
          5916 => x"38",
          5917 => x"b9",
          5918 => x"76",
          5919 => x"97",
          5920 => x"b9",
          5921 => x"33",
          5922 => x"24",
          5923 => x"2a",
          5924 => x"80",
          5925 => x"33",
          5926 => x"7d",
          5927 => x"78",
          5928 => x"0c",
          5929 => x"23",
          5930 => x"3f",
          5931 => x"2e",
          5932 => x"38",
          5933 => x"55",
          5934 => x"17",
          5935 => x"71",
          5936 => x"0c",
          5937 => x"0d",
          5938 => x"9e",
          5939 => x"96",
          5940 => x"8e",
          5941 => x"57",
          5942 => x"52",
          5943 => x"0c",
          5944 => x"0d",
          5945 => x"c3",
          5946 => x"52",
          5947 => x"54",
          5948 => x"58",
          5949 => x"38",
          5950 => x"38",
          5951 => x"38",
          5952 => x"53",
          5953 => x"53",
          5954 => x"38",
          5955 => x"52",
          5956 => x"b9",
          5957 => x"84",
          5958 => x"a6",
          5959 => x"92",
          5960 => x"be",
          5961 => x"70",
          5962 => x"b9",
          5963 => x"84",
          5964 => x"75",
          5965 => x"e2",
          5966 => x"8e",
          5967 => x"70",
          5968 => x"b9",
          5969 => x"39",
          5970 => x"3f",
          5971 => x"0c",
          5972 => x"51",
          5973 => x"08",
          5974 => x"72",
          5975 => x"ed",
          5976 => x"3d",
          5977 => x"a5",
          5978 => x"b9",
          5979 => x"84",
          5980 => x"65",
          5981 => x"84",
          5982 => x"08",
          5983 => x"70",
          5984 => x"97",
          5985 => x"52",
          5986 => x"84",
          5987 => x"86",
          5988 => x"0d",
          5989 => x"5f",
          5990 => x"96",
          5991 => x"c8",
          5992 => x"38",
          5993 => x"08",
          5994 => x"59",
          5995 => x"7f",
          5996 => x"3d",
          5997 => x"33",
          5998 => x"38",
          5999 => x"08",
          6000 => x"7b",
          6001 => x"17",
          6002 => x"17",
          6003 => x"38",
          6004 => x"81",
          6005 => x"84",
          6006 => x"ff",
          6007 => x"7f",
          6008 => x"76",
          6009 => x"38",
          6010 => x"82",
          6011 => x"2b",
          6012 => x"88",
          6013 => x"fe",
          6014 => x"25",
          6015 => x"06",
          6016 => x"54",
          6017 => x"fe",
          6018 => x"18",
          6019 => x"77",
          6020 => x"0c",
          6021 => x"17",
          6022 => x"18",
          6023 => x"81",
          6024 => x"38",
          6025 => x"b4",
          6026 => x"b9",
          6027 => x"08",
          6028 => x"55",
          6029 => x"b0",
          6030 => x"18",
          6031 => x"33",
          6032 => x"fe",
          6033 => x"59",
          6034 => x"80",
          6035 => x"80",
          6036 => x"2e",
          6037 => x"30",
          6038 => x"25",
          6039 => x"5c",
          6040 => x"38",
          6041 => x"84",
          6042 => x"18",
          6043 => x"05",
          6044 => x"2b",
          6045 => x"82",
          6046 => x"5d",
          6047 => x"83",
          6048 => x"bf",
          6049 => x"0c",
          6050 => x"81",
          6051 => x"83",
          6052 => x"f7",
          6053 => x"80",
          6054 => x"80",
          6055 => x"80",
          6056 => x"18",
          6057 => x"da",
          6058 => x"dc",
          6059 => x"d4",
          6060 => x"81",
          6061 => x"2e",
          6062 => x"73",
          6063 => x"81",
          6064 => x"57",
          6065 => x"16",
          6066 => x"80",
          6067 => x"8c",
          6068 => x"78",
          6069 => x"38",
          6070 => x"84",
          6071 => x"78",
          6072 => x"73",
          6073 => x"84",
          6074 => x"08",
          6075 => x"c8",
          6076 => x"b9",
          6077 => x"80",
          6078 => x"81",
          6079 => x"38",
          6080 => x"08",
          6081 => x"af",
          6082 => x"16",
          6083 => x"34",
          6084 => x"38",
          6085 => x"f6",
          6086 => x"06",
          6087 => x"08",
          6088 => x"90",
          6089 => x"0b",
          6090 => x"17",
          6091 => x"3f",
          6092 => x"c2",
          6093 => x"81",
          6094 => x"58",
          6095 => x"27",
          6096 => x"98",
          6097 => x"81",
          6098 => x"a1",
          6099 => x"08",
          6100 => x"97",
          6101 => x"ff",
          6102 => x"55",
          6103 => x"73",
          6104 => x"84",
          6105 => x"08",
          6106 => x"c8",
          6107 => x"b9",
          6108 => x"80",
          6109 => x"89",
          6110 => x"38",
          6111 => x"08",
          6112 => x"38",
          6113 => x"33",
          6114 => x"78",
          6115 => x"80",
          6116 => x"fc",
          6117 => x"82",
          6118 => x"e4",
          6119 => x"90",
          6120 => x"84",
          6121 => x"54",
          6122 => x"33",
          6123 => x"c8",
          6124 => x"bb",
          6125 => x"3d",
          6126 => x"ff",
          6127 => x"56",
          6128 => x"38",
          6129 => x"0d",
          6130 => x"9b",
          6131 => x"3f",
          6132 => x"c8",
          6133 => x"33",
          6134 => x"86",
          6135 => x"5b",
          6136 => x"ee",
          6137 => x"87",
          6138 => x"3d",
          6139 => x"71",
          6140 => x"5c",
          6141 => x"38",
          6142 => x"80",
          6143 => x"18",
          6144 => x"5f",
          6145 => x"8f",
          6146 => x"3f",
          6147 => x"c8",
          6148 => x"08",
          6149 => x"84",
          6150 => x"08",
          6151 => x"0c",
          6152 => x"94",
          6153 => x"2b",
          6154 => x"98",
          6155 => x"88",
          6156 => x"38",
          6157 => x"5d",
          6158 => x"74",
          6159 => x"84",
          6160 => x"08",
          6161 => x"77",
          6162 => x"2e",
          6163 => x"7a",
          6164 => x"89",
          6165 => x"fd",
          6166 => x"7d",
          6167 => x"c8",
          6168 => x"0d",
          6169 => x"56",
          6170 => x"82",
          6171 => x"55",
          6172 => x"dd",
          6173 => x"52",
          6174 => x"3f",
          6175 => x"38",
          6176 => x"0c",
          6177 => x"08",
          6178 => x"18",
          6179 => x"ec",
          6180 => x"de",
          6181 => x"b9",
          6182 => x"75",
          6183 => x"38",
          6184 => x"b4",
          6185 => x"33",
          6186 => x"84",
          6187 => x"06",
          6188 => x"83",
          6189 => x"08",
          6190 => x"74",
          6191 => x"82",
          6192 => x"81",
          6193 => x"17",
          6194 => x"52",
          6195 => x"3f",
          6196 => x"79",
          6197 => x"78",
          6198 => x"c8",
          6199 => x"2e",
          6200 => x"81",
          6201 => x"08",
          6202 => x"74",
          6203 => x"84",
          6204 => x"08",
          6205 => x"58",
          6206 => x"16",
          6207 => x"07",
          6208 => x"77",
          6209 => x"fd",
          6210 => x"84",
          6211 => x"81",
          6212 => x"82",
          6213 => x"a0",
          6214 => x"b9",
          6215 => x"80",
          6216 => x"0c",
          6217 => x"52",
          6218 => x"bf",
          6219 => x"b9",
          6220 => x"b9",
          6221 => x"b9",
          6222 => x"cb",
          6223 => x"85",
          6224 => x"74",
          6225 => x"8f",
          6226 => x"3f",
          6227 => x"84",
          6228 => x"84",
          6229 => x"38",
          6230 => x"cb",
          6231 => x"b9",
          6232 => x"57",
          6233 => x"18",
          6234 => x"75",
          6235 => x"76",
          6236 => x"58",
          6237 => x"84",
          6238 => x"81",
          6239 => x"f4",
          6240 => x"77",
          6241 => x"77",
          6242 => x"51",
          6243 => x"08",
          6244 => x"39",
          6245 => x"b4",
          6246 => x"81",
          6247 => x"3f",
          6248 => x"38",
          6249 => x"b4",
          6250 => x"74",
          6251 => x"82",
          6252 => x"81",
          6253 => x"17",
          6254 => x"52",
          6255 => x"3f",
          6256 => x"08",
          6257 => x"38",
          6258 => x"38",
          6259 => x"3f",
          6260 => x"c8",
          6261 => x"b9",
          6262 => x"84",
          6263 => x"38",
          6264 => x"f9",
          6265 => x"f3",
          6266 => x"19",
          6267 => x"90",
          6268 => x"17",
          6269 => x"34",
          6270 => x"38",
          6271 => x"0d",
          6272 => x"ff",
          6273 => x"2e",
          6274 => x"0b",
          6275 => x"81",
          6276 => x"f4",
          6277 => x"34",
          6278 => x"34",
          6279 => x"75",
          6280 => x"d0",
          6281 => x"1a",
          6282 => x"59",
          6283 => x"88",
          6284 => x"75",
          6285 => x"38",
          6286 => x"b8",
          6287 => x"05",
          6288 => x"34",
          6289 => x"56",
          6290 => x"7e",
          6291 => x"57",
          6292 => x"2a",
          6293 => x"33",
          6294 => x"7d",
          6295 => x"51",
          6296 => x"08",
          6297 => x"38",
          6298 => x"17",
          6299 => x"34",
          6300 => x"0b",
          6301 => x"77",
          6302 => x"78",
          6303 => x"83",
          6304 => x"0b",
          6305 => x"83",
          6306 => x"3f",
          6307 => x"b9",
          6308 => x"90",
          6309 => x"74",
          6310 => x"34",
          6311 => x"7a",
          6312 => x"55",
          6313 => x"a0",
          6314 => x"58",
          6315 => x"58",
          6316 => x"5c",
          6317 => x"0b",
          6318 => x"83",
          6319 => x"3f",
          6320 => x"39",
          6321 => x"08",
          6322 => x"9b",
          6323 => x"70",
          6324 => x"81",
          6325 => x"2e",
          6326 => x"fe",
          6327 => x"ab",
          6328 => x"84",
          6329 => x"75",
          6330 => x"04",
          6331 => x"52",
          6332 => x"af",
          6333 => x"b9",
          6334 => x"05",
          6335 => x"7c",
          6336 => x"3d",
          6337 => x"05",
          6338 => x"34",
          6339 => x"3d",
          6340 => x"75",
          6341 => x"81",
          6342 => x"ef",
          6343 => x"ff",
          6344 => x"56",
          6345 => x"6a",
          6346 => x"88",
          6347 => x"0d",
          6348 => x"ff",
          6349 => x"91",
          6350 => x"d0",
          6351 => x"fa",
          6352 => x"70",
          6353 => x"7a",
          6354 => x"81",
          6355 => x"58",
          6356 => x"16",
          6357 => x"9f",
          6358 => x"e0",
          6359 => x"75",
          6360 => x"77",
          6361 => x"ff",
          6362 => x"70",
          6363 => x"58",
          6364 => x"1c",
          6365 => x"fd",
          6366 => x"ff",
          6367 => x"38",
          6368 => x"fe",
          6369 => x"a8",
          6370 => x"84",
          6371 => x"b8",
          6372 => x"81",
          6373 => x"8d",
          6374 => x"84",
          6375 => x"58",
          6376 => x"80",
          6377 => x"81",
          6378 => x"57",
          6379 => x"02",
          6380 => x"8b",
          6381 => x"40",
          6382 => x"57",
          6383 => x"0b",
          6384 => x"84",
          6385 => x"2e",
          6386 => x"2e",
          6387 => x"9a",
          6388 => x"33",
          6389 => x"82",
          6390 => x"fe",
          6391 => x"c7",
          6392 => x"b0",
          6393 => x"2e",
          6394 => x"b4",
          6395 => x"17",
          6396 => x"54",
          6397 => x"33",
          6398 => x"c8",
          6399 => x"81",
          6400 => x"7b",
          6401 => x"bf",
          6402 => x"2e",
          6403 => x"83",
          6404 => x"f2",
          6405 => x"80",
          6406 => x"83",
          6407 => x"90",
          6408 => x"7d",
          6409 => x"34",
          6410 => x"78",
          6411 => x"57",
          6412 => x"74",
          6413 => x"84",
          6414 => x"08",
          6415 => x"19",
          6416 => x"77",
          6417 => x"59",
          6418 => x"81",
          6419 => x"16",
          6420 => x"bd",
          6421 => x"85",
          6422 => x"17",
          6423 => x"19",
          6424 => x"83",
          6425 => x"a5",
          6426 => x"ae",
          6427 => x"b9",
          6428 => x"82",
          6429 => x"74",
          6430 => x"fe",
          6431 => x"84",
          6432 => x"82",
          6433 => x"0d",
          6434 => x"71",
          6435 => x"07",
          6436 => x"b9",
          6437 => x"84",
          6438 => x"38",
          6439 => x"0d",
          6440 => x"7b",
          6441 => x"94",
          6442 => x"7a",
          6443 => x"84",
          6444 => x"16",
          6445 => x"c8",
          6446 => x"27",
          6447 => x"7c",
          6448 => x"38",
          6449 => x"08",
          6450 => x"51",
          6451 => x"fa",
          6452 => x"b8",
          6453 => x"5b",
          6454 => x"b9",
          6455 => x"c8",
          6456 => x"a8",
          6457 => x"5d",
          6458 => x"8e",
          6459 => x"2e",
          6460 => x"54",
          6461 => x"53",
          6462 => x"e0",
          6463 => x"ec",
          6464 => x"02",
          6465 => x"57",
          6466 => x"97",
          6467 => x"b9",
          6468 => x"80",
          6469 => x"0c",
          6470 => x"52",
          6471 => x"d7",
          6472 => x"b9",
          6473 => x"05",
          6474 => x"73",
          6475 => x"09",
          6476 => x"06",
          6477 => x"17",
          6478 => x"34",
          6479 => x"b9",
          6480 => x"3d",
          6481 => x"82",
          6482 => x"3d",
          6483 => x"c8",
          6484 => x"2e",
          6485 => x"96",
          6486 => x"96",
          6487 => x"3f",
          6488 => x"c8",
          6489 => x"33",
          6490 => x"d2",
          6491 => x"22",
          6492 => x"76",
          6493 => x"74",
          6494 => x"77",
          6495 => x"73",
          6496 => x"83",
          6497 => x"3f",
          6498 => x"0c",
          6499 => x"6b",
          6500 => x"cc",
          6501 => x"c5",
          6502 => x"c8",
          6503 => x"07",
          6504 => x"2e",
          6505 => x"56",
          6506 => x"78",
          6507 => x"2e",
          6508 => x"5a",
          6509 => x"7c",
          6510 => x"b4",
          6511 => x"83",
          6512 => x"2e",
          6513 => x"54",
          6514 => x"33",
          6515 => x"c8",
          6516 => x"81",
          6517 => x"78",
          6518 => x"80",
          6519 => x"80",
          6520 => x"a7",
          6521 => x"33",
          6522 => x"88",
          6523 => x"07",
          6524 => x"0c",
          6525 => x"84",
          6526 => x"7c",
          6527 => x"70",
          6528 => x"b9",
          6529 => x"80",
          6530 => x"09",
          6531 => x"34",
          6532 => x"b4",
          6533 => x"81",
          6534 => x"3f",
          6535 => x"2e",
          6536 => x"b9",
          6537 => x"08",
          6538 => x"08",
          6539 => x"fe",
          6540 => x"82",
          6541 => x"77",
          6542 => x"05",
          6543 => x"fe",
          6544 => x"76",
          6545 => x"51",
          6546 => x"08",
          6547 => x"39",
          6548 => x"3f",
          6549 => x"c8",
          6550 => x"08",
          6551 => x"59",
          6552 => x"59",
          6553 => x"59",
          6554 => x"1c",
          6555 => x"2e",
          6556 => x"70",
          6557 => x"ea",
          6558 => x"ba",
          6559 => x"3d",
          6560 => x"ff",
          6561 => x"56",
          6562 => x"8f",
          6563 => x"76",
          6564 => x"55",
          6565 => x"70",
          6566 => x"58",
          6567 => x"a2",
          6568 => x"ff",
          6569 => x"f5",
          6570 => x"ff",
          6571 => x"95",
          6572 => x"08",
          6573 => x"08",
          6574 => x"2e",
          6575 => x"83",
          6576 => x"5b",
          6577 => x"38",
          6578 => x"81",
          6579 => x"57",
          6580 => x"74",
          6581 => x"75",
          6582 => x"38",
          6583 => x"79",
          6584 => x"77",
          6585 => x"74",
          6586 => x"1a",
          6587 => x"34",
          6588 => x"70",
          6589 => x"77",
          6590 => x"33",
          6591 => x"bc",
          6592 => x"b7",
          6593 => x"5c",
          6594 => x"38",
          6595 => x"45",
          6596 => x"52",
          6597 => x"c8",
          6598 => x"2e",
          6599 => x"c8",
          6600 => x"52",
          6601 => x"c8",
          6602 => x"fd",
          6603 => x"c8",
          6604 => x"d8",
          6605 => x"75",
          6606 => x"c8",
          6607 => x"c1",
          6608 => x"8b",
          6609 => x"81",
          6610 => x"58",
          6611 => x"7d",
          6612 => x"51",
          6613 => x"08",
          6614 => x"7a",
          6615 => x"9c",
          6616 => x"09",
          6617 => x"79",
          6618 => x"75",
          6619 => x"3f",
          6620 => x"c8",
          6621 => x"84",
          6622 => x"5c",
          6623 => x"b4",
          6624 => x"18",
          6625 => x"06",
          6626 => x"b8",
          6627 => x"d5",
          6628 => x"2e",
          6629 => x"b4",
          6630 => x"78",
          6631 => x"57",
          6632 => x"74",
          6633 => x"5c",
          6634 => x"1a",
          6635 => x"52",
          6636 => x"b9",
          6637 => x"80",
          6638 => x"84",
          6639 => x"fd",
          6640 => x"76",
          6641 => x"55",
          6642 => x"8b",
          6643 => x"55",
          6644 => x"70",
          6645 => x"74",
          6646 => x"81",
          6647 => x"58",
          6648 => x"fd",
          6649 => x"7d",
          6650 => x"51",
          6651 => x"08",
          6652 => x"df",
          6653 => x"7a",
          6654 => x"ec",
          6655 => x"09",
          6656 => x"c8",
          6657 => x"a8",
          6658 => x"08",
          6659 => x"74",
          6660 => x"08",
          6661 => x"52",
          6662 => x"b9",
          6663 => x"80",
          6664 => x"81",
          6665 => x"e7",
          6666 => x"18",
          6667 => x"52",
          6668 => x"3f",
          6669 => x"62",
          6670 => x"5e",
          6671 => x"9f",
          6672 => x"97",
          6673 => x"8f",
          6674 => x"59",
          6675 => x"80",
          6676 => x"91",
          6677 => x"79",
          6678 => x"08",
          6679 => x"81",
          6680 => x"2e",
          6681 => x"70",
          6682 => x"5c",
          6683 => x"7a",
          6684 => x"2a",
          6685 => x"08",
          6686 => x"78",
          6687 => x"26",
          6688 => x"5b",
          6689 => x"d8",
          6690 => x"9c",
          6691 => x"55",
          6692 => x"dc",
          6693 => x"81",
          6694 => x"c5",
          6695 => x"bb",
          6696 => x"c2",
          6697 => x"b9",
          6698 => x"0b",
          6699 => x"04",
          6700 => x"3f",
          6701 => x"73",
          6702 => x"56",
          6703 => x"8e",
          6704 => x"2e",
          6705 => x"2e",
          6706 => x"7e",
          6707 => x"c8",
          6708 => x"a3",
          6709 => x"59",
          6710 => x"12",
          6711 => x"38",
          6712 => x"0c",
          6713 => x"7b",
          6714 => x"05",
          6715 => x"26",
          6716 => x"16",
          6717 => x"7c",
          6718 => x"39",
          6719 => x"80",
          6720 => x"c5",
          6721 => x"1b",
          6722 => x"08",
          6723 => x"3d",
          6724 => x"33",
          6725 => x"08",
          6726 => x"85",
          6727 => x"33",
          6728 => x"2e",
          6729 => x"ba",
          6730 => x"33",
          6731 => x"75",
          6732 => x"08",
          6733 => x"80",
          6734 => x"11",
          6735 => x"5b",
          6736 => x"a9",
          6737 => x"06",
          6738 => x"7b",
          6739 => x"06",
          6740 => x"9f",
          6741 => x"51",
          6742 => x"08",
          6743 => x"2e",
          6744 => x"26",
          6745 => x"55",
          6746 => x"88",
          6747 => x"38",
          6748 => x"38",
          6749 => x"e7",
          6750 => x"89",
          6751 => x"47",
          6752 => x"65",
          6753 => x"5f",
          6754 => x"80",
          6755 => x"53",
          6756 => x"3f",
          6757 => x"95",
          6758 => x"83",
          6759 => x"59",
          6760 => x"2e",
          6761 => x"90",
          6762 => x"44",
          6763 => x"83",
          6764 => x"33",
          6765 => x"81",
          6766 => x"75",
          6767 => x"11",
          6768 => x"71",
          6769 => x"72",
          6770 => x"5c",
          6771 => x"a3",
          6772 => x"4f",
          6773 => x"80",
          6774 => x"57",
          6775 => x"61",
          6776 => x"63",
          6777 => x"06",
          6778 => x"81",
          6779 => x"6e",
          6780 => x"62",
          6781 => x"38",
          6782 => x"e6",
          6783 => x"9d",
          6784 => x"e6",
          6785 => x"22",
          6786 => x"38",
          6787 => x"78",
          6788 => x"c8",
          6789 => x"c8",
          6790 => x"0b",
          6791 => x"c8",
          6792 => x"05",
          6793 => x"2a",
          6794 => x"7d",
          6795 => x"70",
          6796 => x"44",
          6797 => x"1d",
          6798 => x"31",
          6799 => x"38",
          6800 => x"70",
          6801 => x"3f",
          6802 => x"2e",
          6803 => x"81",
          6804 => x"0b",
          6805 => x"38",
          6806 => x"74",
          6807 => x"5b",
          6808 => x"b9",
          6809 => x"d4",
          6810 => x"93",
          6811 => x"0d",
          6812 => x"d0",
          6813 => x"57",
          6814 => x"77",
          6815 => x"77",
          6816 => x"83",
          6817 => x"57",
          6818 => x"76",
          6819 => x"12",
          6820 => x"38",
          6821 => x"44",
          6822 => x"89",
          6823 => x"59",
          6824 => x"47",
          6825 => x"38",
          6826 => x"70",
          6827 => x"07",
          6828 => x"ce",
          6829 => x"83",
          6830 => x"f9",
          6831 => x"81",
          6832 => x"81",
          6833 => x"38",
          6834 => x"c8",
          6835 => x"5f",
          6836 => x"fe",
          6837 => x"fb",
          6838 => x"83",
          6839 => x"3d",
          6840 => x"06",
          6841 => x"f5",
          6842 => x"43",
          6843 => x"9f",
          6844 => x"77",
          6845 => x"f5",
          6846 => x"0c",
          6847 => x"04",
          6848 => x"38",
          6849 => x"81",
          6850 => x"38",
          6851 => x"70",
          6852 => x"74",
          6853 => x"59",
          6854 => x"33",
          6855 => x"15",
          6856 => x"45",
          6857 => x"34",
          6858 => x"ff",
          6859 => x"34",
          6860 => x"05",
          6861 => x"83",
          6862 => x"91",
          6863 => x"49",
          6864 => x"75",
          6865 => x"75",
          6866 => x"93",
          6867 => x"61",
          6868 => x"34",
          6869 => x"99",
          6870 => x"80",
          6871 => x"05",
          6872 => x"9d",
          6873 => x"61",
          6874 => x"b9",
          6875 => x"9f",
          6876 => x"38",
          6877 => x"a8",
          6878 => x"80",
          6879 => x"ff",
          6880 => x"34",
          6881 => x"05",
          6882 => x"a9",
          6883 => x"05",
          6884 => x"70",
          6885 => x"05",
          6886 => x"38",
          6887 => x"69",
          6888 => x"aa",
          6889 => x"52",
          6890 => x"57",
          6891 => x"60",
          6892 => x"38",
          6893 => x"81",
          6894 => x"f4",
          6895 => x"2e",
          6896 => x"57",
          6897 => x"76",
          6898 => x"55",
          6899 => x"76",
          6900 => x"05",
          6901 => x"64",
          6902 => x"26",
          6903 => x"53",
          6904 => x"3f",
          6905 => x"84",
          6906 => x"81",
          6907 => x"f4",
          6908 => x"5b",
          6909 => x"7f",
          6910 => x"62",
          6911 => x"55",
          6912 => x"74",
          6913 => x"fe",
          6914 => x"85",
          6915 => x"57",
          6916 => x"83",
          6917 => x"ff",
          6918 => x"82",
          6919 => x"c1",
          6920 => x"7d",
          6921 => x"59",
          6922 => x"ff",
          6923 => x"69",
          6924 => x"be",
          6925 => x"81",
          6926 => x"78",
          6927 => x"05",
          6928 => x"62",
          6929 => x"67",
          6930 => x"82",
          6931 => x"05",
          6932 => x"05",
          6933 => x"67",
          6934 => x"83",
          6935 => x"61",
          6936 => x"ca",
          6937 => x"61",
          6938 => x"58",
          6939 => x"98",
          6940 => x"34",
          6941 => x"51",
          6942 => x"b9",
          6943 => x"80",
          6944 => x"81",
          6945 => x"38",
          6946 => x"0c",
          6947 => x"04",
          6948 => x"64",
          6949 => x"ae",
          6950 => x"83",
          6951 => x"2e",
          6952 => x"83",
          6953 => x"70",
          6954 => x"86",
          6955 => x"52",
          6956 => x"b9",
          6957 => x"70",
          6958 => x"0b",
          6959 => x"05",
          6960 => x"27",
          6961 => x"39",
          6962 => x"26",
          6963 => x"77",
          6964 => x"8e",
          6965 => x"44",
          6966 => x"43",
          6967 => x"34",
          6968 => x"05",
          6969 => x"a2",
          6970 => x"61",
          6971 => x"61",
          6972 => x"c4",
          6973 => x"34",
          6974 => x"7c",
          6975 => x"5c",
          6976 => x"2a",
          6977 => x"98",
          6978 => x"82",
          6979 => x"05",
          6980 => x"61",
          6981 => x"34",
          6982 => x"b2",
          6983 => x"ff",
          6984 => x"61",
          6985 => x"c7",
          6986 => x"76",
          6987 => x"81",
          6988 => x"80",
          6989 => x"05",
          6990 => x"34",
          6991 => x"b8",
          6992 => x"79",
          6993 => x"84",
          6994 => x"90",
          6995 => x"b2",
          6996 => x"08",
          6997 => x"b4",
          6998 => x"b9",
          6999 => x"d4",
          7000 => x"ff",
          7001 => x"6a",
          7002 => x"34",
          7003 => x"85",
          7004 => x"ff",
          7005 => x"05",
          7006 => x"61",
          7007 => x"57",
          7008 => x"53",
          7009 => x"3f",
          7010 => x"70",
          7011 => x"76",
          7012 => x"70",
          7013 => x"d2",
          7014 => x"e1",
          7015 => x"c1",
          7016 => x"05",
          7017 => x"34",
          7018 => x"80",
          7019 => x"ff",
          7020 => x"34",
          7021 => x"e9",
          7022 => x"61",
          7023 => x"40",
          7024 => x"61",
          7025 => x"ed",
          7026 => x"34",
          7027 => x"d5",
          7028 => x"54",
          7029 => x"fe",
          7030 => x"53",
          7031 => x"3f",
          7032 => x"f4",
          7033 => x"7b",
          7034 => x"78",
          7035 => x"3d",
          7036 => x"79",
          7037 => x"2e",
          7038 => x"33",
          7039 => x"76",
          7040 => x"57",
          7041 => x"24",
          7042 => x"76",
          7043 => x"c8",
          7044 => x"0d",
          7045 => x"59",
          7046 => x"84",
          7047 => x"38",
          7048 => x"56",
          7049 => x"74",
          7050 => x"0c",
          7051 => x"0d",
          7052 => x"53",
          7053 => x"9e",
          7054 => x"70",
          7055 => x"1b",
          7056 => x"56",
          7057 => x"ff",
          7058 => x"0d",
          7059 => x"58",
          7060 => x"76",
          7061 => x"55",
          7062 => x"0c",
          7063 => x"56",
          7064 => x"77",
          7065 => x"34",
          7066 => x"38",
          7067 => x"18",
          7068 => x"38",
          7069 => x"54",
          7070 => x"9d",
          7071 => x"38",
          7072 => x"84",
          7073 => x"9f",
          7074 => x"c0",
          7075 => x"a2",
          7076 => x"72",
          7077 => x"56",
          7078 => x"51",
          7079 => x"84",
          7080 => x"fd",
          7081 => x"05",
          7082 => x"ff",
          7083 => x"06",
          7084 => x"3d",
          7085 => x"54",
          7086 => x"e9",
          7087 => x"e7",
          7088 => x"38",
          7089 => x"53",
          7090 => x"71",
          7091 => x"51",
          7092 => x"81",
          7093 => x"85",
          7094 => x"92",
          7095 => x"22",
          7096 => x"26",
          7097 => x"c8",
          7098 => x"b5",
          7099 => x"81",
          7100 => x"e5",
          7101 => x"0c",
          7102 => x"0d",
          7103 => x"80",
          7104 => x"83",
          7105 => x"26",
          7106 => x"56",
          7107 => x"73",
          7108 => x"70",
          7109 => x"22",
          7110 => x"ff",
          7111 => x"24",
          7112 => x"15",
          7113 => x"73",
          7114 => x"07",
          7115 => x"38",
          7116 => x"87",
          7117 => x"ff",
          7118 => x"71",
          7119 => x"73",
          7120 => x"ff",
          7121 => x"39",
          7122 => x"06",
          7123 => x"83",
          7124 => x"e6",
          7125 => x"51",
          7126 => x"ff",
          7127 => x"70",
          7128 => x"39",
          7129 => x"57",
          7130 => x"81",
          7131 => x"ff",
          7132 => x"75",
          7133 => x"52",
          7134 => x"ff",
          7135 => x"ff",
          7136 => x"00",
          7137 => x"00",
          7138 => x"00",
          7139 => x"00",
          7140 => x"00",
          7141 => x"00",
          7142 => x"00",
          7143 => x"00",
          7144 => x"00",
          7145 => x"00",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"00",
          7374 => x"6c",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"72",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"65",
          7383 => x"69",
          7384 => x"66",
          7385 => x"61",
          7386 => x"6d",
          7387 => x"72",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"38",
          7392 => x"63",
          7393 => x"63",
          7394 => x"00",
          7395 => x"6e",
          7396 => x"72",
          7397 => x"61",
          7398 => x"73",
          7399 => x"65",
          7400 => x"6f",
          7401 => x"6f",
          7402 => x"65",
          7403 => x"6e",
          7404 => x"65",
          7405 => x"72",
          7406 => x"69",
          7407 => x"6f",
          7408 => x"69",
          7409 => x"6f",
          7410 => x"6e",
          7411 => x"6c",
          7412 => x"6f",
          7413 => x"6f",
          7414 => x"6f",
          7415 => x"69",
          7416 => x"65",
          7417 => x"66",
          7418 => x"20",
          7419 => x"69",
          7420 => x"65",
          7421 => x"00",
          7422 => x"20",
          7423 => x"69",
          7424 => x"69",
          7425 => x"44",
          7426 => x"74",
          7427 => x"63",
          7428 => x"69",
          7429 => x"6c",
          7430 => x"69",
          7431 => x"69",
          7432 => x"61",
          7433 => x"74",
          7434 => x"63",
          7435 => x"6e",
          7436 => x"6e",
          7437 => x"69",
          7438 => x"00",
          7439 => x"74",
          7440 => x"2e",
          7441 => x"6c",
          7442 => x"2e",
          7443 => x"6e",
          7444 => x"79",
          7445 => x"6e",
          7446 => x"72",
          7447 => x"45",
          7448 => x"75",
          7449 => x"00",
          7450 => x"62",
          7451 => x"20",
          7452 => x"62",
          7453 => x"63",
          7454 => x"65",
          7455 => x"30",
          7456 => x"20",
          7457 => x"00",
          7458 => x"00",
          7459 => x"30",
          7460 => x"20",
          7461 => x"00",
          7462 => x"2a",
          7463 => x"37",
          7464 => x"31",
          7465 => x"00",
          7466 => x"20",
          7467 => x"78",
          7468 => x"20",
          7469 => x"53",
          7470 => x"61",
          7471 => x"65",
          7472 => x"20",
          7473 => x"3d",
          7474 => x"00",
          7475 => x"70",
          7476 => x"73",
          7477 => x"20",
          7478 => x"3d",
          7479 => x"00",
          7480 => x"6e",
          7481 => x"20",
          7482 => x"00",
          7483 => x"20",
          7484 => x"72",
          7485 => x"41",
          7486 => x"69",
          7487 => x"74",
          7488 => x"20",
          7489 => x"72",
          7490 => x"41",
          7491 => x"69",
          7492 => x"74",
          7493 => x"20",
          7494 => x"72",
          7495 => x"4f",
          7496 => x"69",
          7497 => x"74",
          7498 => x"6e",
          7499 => x"00",
          7500 => x"20",
          7501 => x"70",
          7502 => x"6e",
          7503 => x"6d",
          7504 => x"6e",
          7505 => x"74",
          7506 => x"00",
          7507 => x"78",
          7508 => x"00",
          7509 => x"70",
          7510 => x"61",
          7511 => x"20",
          7512 => x"69",
          7513 => x"61",
          7514 => x"6c",
          7515 => x"69",
          7516 => x"6c",
          7517 => x"20",
          7518 => x"73",
          7519 => x"61",
          7520 => x"6e",
          7521 => x"50",
          7522 => x"64",
          7523 => x"2e",
          7524 => x"6f",
          7525 => x"6f",
          7526 => x"00",
          7527 => x"72",
          7528 => x"70",
          7529 => x"6e",
          7530 => x"61",
          7531 => x"6f",
          7532 => x"38",
          7533 => x"00",
          7534 => x"72",
          7535 => x"20",
          7536 => x"64",
          7537 => x"78",
          7538 => x"20",
          7539 => x"25",
          7540 => x"2e",
          7541 => x"20",
          7542 => x"00",
          7543 => x"20",
          7544 => x"6f",
          7545 => x"2e",
          7546 => x"30",
          7547 => x"78",
          7548 => x"78",
          7549 => x"00",
          7550 => x"6e",
          7551 => x"30",
          7552 => x"58",
          7553 => x"69",
          7554 => x"00",
          7555 => x"4d",
          7556 => x"43",
          7557 => x"2e",
          7558 => x"73",
          7559 => x"65",
          7560 => x"68",
          7561 => x"20",
          7562 => x"70",
          7563 => x"63",
          7564 => x"00",
          7565 => x"64",
          7566 => x"25",
          7567 => x"2e",
          7568 => x"6f",
          7569 => x"67",
          7570 => x"00",
          7571 => x"69",
          7572 => x"6c",
          7573 => x"3a",
          7574 => x"73",
          7575 => x"20",
          7576 => x"65",
          7577 => x"74",
          7578 => x"65",
          7579 => x"38",
          7580 => x"20",
          7581 => x"65",
          7582 => x"61",
          7583 => x"65",
          7584 => x"38",
          7585 => x"20",
          7586 => x"20",
          7587 => x"64",
          7588 => x"20",
          7589 => x"38",
          7590 => x"69",
          7591 => x"20",
          7592 => x"64",
          7593 => x"20",
          7594 => x"20",
          7595 => x"34",
          7596 => x"20",
          7597 => x"6d",
          7598 => x"46",
          7599 => x"20",
          7600 => x"2e",
          7601 => x"0a",
          7602 => x"69",
          7603 => x"53",
          7604 => x"6f",
          7605 => x"3d",
          7606 => x"64",
          7607 => x"20",
          7608 => x"20",
          7609 => x"72",
          7610 => x"20",
          7611 => x"2e",
          7612 => x"0a",
          7613 => x"50",
          7614 => x"53",
          7615 => x"4f",
          7616 => x"20",
          7617 => x"43",
          7618 => x"49",
          7619 => x"42",
          7620 => x"20",
          7621 => x"43",
          7622 => x"61",
          7623 => x"30",
          7624 => x"20",
          7625 => x"31",
          7626 => x"6d",
          7627 => x"30",
          7628 => x"20",
          7629 => x"52",
          7630 => x"76",
          7631 => x"30",
          7632 => x"20",
          7633 => x"20",
          7634 => x"38",
          7635 => x"2e",
          7636 => x"52",
          7637 => x"20",
          7638 => x"30",
          7639 => x"20",
          7640 => x"42",
          7641 => x"38",
          7642 => x"2e",
          7643 => x"44",
          7644 => x"20",
          7645 => x"30",
          7646 => x"20",
          7647 => x"52",
          7648 => x"38",
          7649 => x"2e",
          7650 => x"6d",
          7651 => x"6e",
          7652 => x"6e",
          7653 => x"56",
          7654 => x"6d",
          7655 => x"65",
          7656 => x"6c",
          7657 => x"56",
          7658 => x"00",
          7659 => x"00",
          7660 => x"00",
          7661 => x"00",
          7662 => x"00",
          7663 => x"00",
          7664 => x"00",
          7665 => x"00",
          7666 => x"00",
          7667 => x"00",
          7668 => x"00",
          7669 => x"00",
          7670 => x"00",
          7671 => x"00",
          7672 => x"00",
          7673 => x"00",
          7674 => x"00",
          7675 => x"00",
          7676 => x"00",
          7677 => x"00",
          7678 => x"00",
          7679 => x"00",
          7680 => x"00",
          7681 => x"00",
          7682 => x"00",
          7683 => x"00",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"00",
          7690 => x"00",
          7691 => x"5b",
          7692 => x"5b",
          7693 => x"5b",
          7694 => x"30",
          7695 => x"5b",
          7696 => x"00",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"74",
          7703 => x"72",
          7704 => x"73",
          7705 => x"6c",
          7706 => x"62",
          7707 => x"69",
          7708 => x"69",
          7709 => x"00",
          7710 => x"20",
          7711 => x"61",
          7712 => x"20",
          7713 => x"68",
          7714 => x"72",
          7715 => x"74",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"5b",
          7720 => x"5b",
          7721 => x"00",
          7722 => x"00",
          7723 => x"00",
          7724 => x"00",
          7725 => x"00",
          7726 => x"00",
          7727 => x"00",
          7728 => x"00",
          7729 => x"00",
          7730 => x"00",
          7731 => x"00",
          7732 => x"00",
          7733 => x"5b",
          7734 => x"5b",
          7735 => x"3a",
          7736 => x"64",
          7737 => x"25",
          7738 => x"00",
          7739 => x"25",
          7740 => x"3a",
          7741 => x"64",
          7742 => x"3a",
          7743 => x"30",
          7744 => x"63",
          7745 => x"00",
          7746 => x"74",
          7747 => x"3a",
          7748 => x"32",
          7749 => x"00",
          7750 => x"32",
          7751 => x"00",
          7752 => x"32",
          7753 => x"6f",
          7754 => x"65",
          7755 => x"00",
          7756 => x"2a",
          7757 => x"00",
          7758 => x"5d",
          7759 => x"41",
          7760 => x"fe",
          7761 => x"2e",
          7762 => x"4d",
          7763 => x"54",
          7764 => x"4f",
          7765 => x"20",
          7766 => x"20",
          7767 => x"00",
          7768 => x"00",
          7769 => x"0e",
          7770 => x"00",
          7771 => x"41",
          7772 => x"49",
          7773 => x"4f",
          7774 => x"9d",
          7775 => x"a5",
          7776 => x"ad",
          7777 => x"b5",
          7778 => x"bd",
          7779 => x"c5",
          7780 => x"cd",
          7781 => x"d5",
          7782 => x"dd",
          7783 => x"e5",
          7784 => x"ed",
          7785 => x"f5",
          7786 => x"fd",
          7787 => x"5b",
          7788 => x"3e",
          7789 => x"01",
          7790 => x"00",
          7791 => x"01",
          7792 => x"10",
          7793 => x"c7",
          7794 => x"e4",
          7795 => x"ea",
          7796 => x"ee",
          7797 => x"c9",
          7798 => x"f6",
          7799 => x"ff",
          7800 => x"a3",
          7801 => x"e1",
          7802 => x"f1",
          7803 => x"bf",
          7804 => x"bc",
          7805 => x"91",
          7806 => x"24",
          7807 => x"55",
          7808 => x"5d",
          7809 => x"14",
          7810 => x"00",
          7811 => x"5a",
          7812 => x"60",
          7813 => x"68",
          7814 => x"58",
          7815 => x"6a",
          7816 => x"84",
          7817 => x"b1",
          7818 => x"a3",
          7819 => x"a6",
          7820 => x"1e",
          7821 => x"61",
          7822 => x"20",
          7823 => x"b0",
          7824 => x"7f",
          7825 => x"61",
          7826 => x"f8",
          7827 => x"78",
          7828 => x"06",
          7829 => x"2e",
          7830 => x"4d",
          7831 => x"82",
          7832 => x"87",
          7833 => x"8b",
          7834 => x"8f",
          7835 => x"93",
          7836 => x"97",
          7837 => x"9b",
          7838 => x"9f",
          7839 => x"a2",
          7840 => x"a7",
          7841 => x"ab",
          7842 => x"af",
          7843 => x"b3",
          7844 => x"b7",
          7845 => x"bb",
          7846 => x"f7",
          7847 => x"c3",
          7848 => x"c7",
          7849 => x"cb",
          7850 => x"dd",
          7851 => x"12",
          7852 => x"f4",
          7853 => x"22",
          7854 => x"65",
          7855 => x"66",
          7856 => x"41",
          7857 => x"40",
          7858 => x"89",
          7859 => x"5a",
          7860 => x"5e",
          7861 => x"62",
          7862 => x"66",
          7863 => x"6a",
          7864 => x"6e",
          7865 => x"9d",
          7866 => x"76",
          7867 => x"7a",
          7868 => x"7e",
          7869 => x"82",
          7870 => x"86",
          7871 => x"b1",
          7872 => x"8e",
          7873 => x"b7",
          7874 => x"fe",
          7875 => x"86",
          7876 => x"b1",
          7877 => x"a3",
          7878 => x"cc",
          7879 => x"8f",
          7880 => x"0a",
          7881 => x"f5",
          7882 => x"f9",
          7883 => x"20",
          7884 => x"22",
          7885 => x"0e",
          7886 => x"d0",
          7887 => x"00",
          7888 => x"63",
          7889 => x"5a",
          7890 => x"06",
          7891 => x"08",
          7892 => x"07",
          7893 => x"54",
          7894 => x"60",
          7895 => x"ba",
          7896 => x"ca",
          7897 => x"f8",
          7898 => x"fa",
          7899 => x"90",
          7900 => x"b0",
          7901 => x"b2",
          7902 => x"c3",
          7903 => x"02",
          7904 => x"f3",
          7905 => x"01",
          7906 => x"84",
          7907 => x"1a",
          7908 => x"02",
          7909 => x"02",
          7910 => x"26",
          7911 => x"00",
          7912 => x"02",
          7913 => x"00",
          7914 => x"04",
          7915 => x"00",
          7916 => x"14",
          7917 => x"00",
          7918 => x"2b",
          7919 => x"00",
          7920 => x"30",
          7921 => x"00",
          7922 => x"3c",
          7923 => x"00",
          7924 => x"3d",
          7925 => x"00",
          7926 => x"3f",
          7927 => x"00",
          7928 => x"40",
          7929 => x"00",
          7930 => x"41",
          7931 => x"00",
          7932 => x"42",
          7933 => x"00",
          7934 => x"43",
          7935 => x"00",
          7936 => x"50",
          7937 => x"00",
          7938 => x"51",
          7939 => x"00",
          7940 => x"54",
          7941 => x"00",
          7942 => x"55",
          7943 => x"00",
          7944 => x"79",
          7945 => x"00",
          7946 => x"78",
          7947 => x"00",
          7948 => x"82",
          7949 => x"00",
          7950 => x"83",
          7951 => x"00",
          7952 => x"85",
          7953 => x"00",
          7954 => x"87",
          7955 => x"00",
          7956 => x"88",
          7957 => x"00",
          7958 => x"89",
          7959 => x"00",
          7960 => x"8c",
          7961 => x"00",
          7962 => x"8d",
          7963 => x"00",
          7964 => x"8e",
          7965 => x"00",
          7966 => x"8f",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"01",
          7971 => x"01",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"f5",
          7976 => x"f5",
          7977 => x"01",
          7978 => x"01",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"00",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"01",
          7995 => x"3b",
          7996 => x"f0",
          7997 => x"76",
          7998 => x"6e",
          7999 => x"66",
          8000 => x"36",
          8001 => x"39",
          8002 => x"f2",
          8003 => x"f0",
          8004 => x"f0",
          8005 => x"3a",
          8006 => x"f0",
          8007 => x"56",
          8008 => x"4e",
          8009 => x"46",
          8010 => x"36",
          8011 => x"39",
          8012 => x"f2",
          8013 => x"f0",
          8014 => x"f0",
          8015 => x"2b",
          8016 => x"f0",
          8017 => x"56",
          8018 => x"4e",
          8019 => x"46",
          8020 => x"26",
          8021 => x"29",
          8022 => x"f8",
          8023 => x"f0",
          8024 => x"f0",
          8025 => x"f0",
          8026 => x"f0",
          8027 => x"16",
          8028 => x"0e",
          8029 => x"06",
          8030 => x"f0",
          8031 => x"1f",
          8032 => x"f0",
          8033 => x"f0",
          8034 => x"f0",
          8035 => x"b5",
          8036 => x"f0",
          8037 => x"a6",
          8038 => x"33",
          8039 => x"43",
          8040 => x"1e",
          8041 => x"a3",
          8042 => x"c4",
          8043 => x"f0",
          8044 => x"f0",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"01",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"e0",
          9081 => x"f9",
          9082 => x"c1",
          9083 => x"e4",
          9084 => x"61",
          9085 => x"69",
          9086 => x"21",
          9087 => x"29",
          9088 => x"01",
          9089 => x"09",
          9090 => x"11",
          9091 => x"19",
          9092 => x"81",
          9093 => x"89",
          9094 => x"91",
          9095 => x"99",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"02",
          9112 => x"00",
        others => X"00"
    );

    shared variable RAM7 : ramArray :=
    (
             0 => x"f8",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"90",
             5 => x"8c",
             6 => x"00",
             7 => x"00",
             8 => x"72",
             9 => x"83",
            10 => x"04",
            11 => x"00",
            12 => x"83",
            13 => x"05",
            14 => x"73",
            15 => x"83",
            16 => x"72",
            17 => x"73",
            18 => x"53",
            19 => x"00",
            20 => x"73",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"0a",
            26 => x"05",
            27 => x"04",
            28 => x"73",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"cd",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"0a",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"09",
            45 => x"05",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"81",
            50 => x"04",
            51 => x"00",
            52 => x"04",
            53 => x"82",
            54 => x"fc",
            55 => x"00",
            56 => x"72",
            57 => x"0a",
            58 => x"00",
            59 => x"00",
            60 => x"72",
            61 => x"0a",
            62 => x"00",
            63 => x"00",
            64 => x"52",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"72",
            77 => x"10",
            78 => x"04",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"93",
            83 => x"00",
            84 => x"90",
            85 => x"cc",
            86 => x"0c",
            87 => x"00",
            88 => x"90",
            89 => x"ab",
            90 => x"0c",
            91 => x"00",
            92 => x"05",
            93 => x"70",
            94 => x"05",
            95 => x"04",
            96 => x"05",
            97 => x"05",
            98 => x"74",
            99 => x"51",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"04",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"05",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"81",
           133 => x"0b",
           134 => x"0b",
           135 => x"b6",
           136 => x"0b",
           137 => x"0b",
           138 => x"f6",
           139 => x"0b",
           140 => x"0b",
           141 => x"b6",
           142 => x"0b",
           143 => x"0b",
           144 => x"f9",
           145 => x"0b",
           146 => x"0b",
           147 => x"bd",
           148 => x"0b",
           149 => x"0b",
           150 => x"81",
           151 => x"0b",
           152 => x"0b",
           153 => x"c5",
           154 => x"0b",
           155 => x"0b",
           156 => x"89",
           157 => x"0b",
           158 => x"0b",
           159 => x"cd",
           160 => x"0b",
           161 => x"0b",
           162 => x"91",
           163 => x"0b",
           164 => x"0b",
           165 => x"d5",
           166 => x"0b",
           167 => x"0b",
           168 => x"99",
           169 => x"0b",
           170 => x"0b",
           171 => x"dc",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"04",
           193 => x"2d",
           194 => x"90",
           195 => x"2d",
           196 => x"90",
           197 => x"2d",
           198 => x"90",
           199 => x"2d",
           200 => x"90",
           201 => x"2d",
           202 => x"90",
           203 => x"2d",
           204 => x"90",
           205 => x"2d",
           206 => x"90",
           207 => x"2d",
           208 => x"90",
           209 => x"2d",
           210 => x"90",
           211 => x"2d",
           212 => x"90",
           213 => x"2d",
           214 => x"90",
           215 => x"2d",
           216 => x"90",
           217 => x"ec",
           218 => x"80",
           219 => x"d5",
           220 => x"c0",
           221 => x"80",
           222 => x"80",
           223 => x"0c",
           224 => x"08",
           225 => x"d4",
           226 => x"d4",
           227 => x"b9",
           228 => x"b9",
           229 => x"84",
           230 => x"84",
           231 => x"04",
           232 => x"2d",
           233 => x"90",
           234 => x"9d",
           235 => x"80",
           236 => x"fa",
           237 => x"c0",
           238 => x"82",
           239 => x"80",
           240 => x"0c",
           241 => x"08",
           242 => x"d4",
           243 => x"d4",
           244 => x"b9",
           245 => x"b9",
           246 => x"84",
           247 => x"84",
           248 => x"04",
           249 => x"2d",
           250 => x"90",
           251 => x"86",
           252 => x"80",
           253 => x"f5",
           254 => x"c0",
           255 => x"83",
           256 => x"80",
           257 => x"0c",
           258 => x"08",
           259 => x"d4",
           260 => x"d4",
           261 => x"b9",
           262 => x"b9",
           263 => x"84",
           264 => x"84",
           265 => x"04",
           266 => x"2d",
           267 => x"90",
           268 => x"9a",
           269 => x"80",
           270 => x"99",
           271 => x"c0",
           272 => x"83",
           273 => x"80",
           274 => x"0c",
           275 => x"08",
           276 => x"d4",
           277 => x"d4",
           278 => x"b9",
           279 => x"b9",
           280 => x"84",
           281 => x"84",
           282 => x"04",
           283 => x"2d",
           284 => x"90",
           285 => x"e2",
           286 => x"80",
           287 => x"f5",
           288 => x"c0",
           289 => x"80",
           290 => x"80",
           291 => x"0c",
           292 => x"08",
           293 => x"d4",
           294 => x"d4",
           295 => x"b9",
           296 => x"d4",
           297 => x"b9",
           298 => x"b9",
           299 => x"84",
           300 => x"84",
           301 => x"04",
           302 => x"2d",
           303 => x"90",
           304 => x"91",
           305 => x"80",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"00",
           311 => x"09",
           312 => x"2b",
           313 => x"04",
           314 => x"05",
           315 => x"72",
           316 => x"51",
           317 => x"70",
           318 => x"71",
           319 => x"0b",
           320 => x"ce",
           321 => x"3d",
           322 => x"53",
           323 => x"81",
           324 => x"3d",
           325 => x"81",
           326 => x"56",
           327 => x"2e",
           328 => x"14",
           329 => x"72",
           330 => x"54",
           331 => x"2e",
           332 => x"84",
           333 => x"08",
           334 => x"08",
           335 => x"14",
           336 => x"07",
           337 => x"80",
           338 => x"52",
           339 => x"0d",
           340 => x"88",
           341 => x"54",
           342 => x"73",
           343 => x"05",
           344 => x"51",
           345 => x"34",
           346 => x"86",
           347 => x"51",
           348 => x"3d",
           349 => x"80",
           350 => x"70",
           351 => x"55",
           352 => x"81",
           353 => x"76",
           354 => x"7b",
           355 => x"81",
           356 => x"26",
           357 => x"30",
           358 => x"ae",
           359 => x"83",
           360 => x"54",
           361 => x"80",
           362 => x"bd",
           363 => x"b9",
           364 => x"83",
           365 => x"10",
           366 => x"19",
           367 => x"05",
           368 => x"5f",
           369 => x"81",
           370 => x"7c",
           371 => x"ff",
           372 => x"06",
           373 => x"5b",
           374 => x"dd",
           375 => x"51",
           376 => x"fe",
           377 => x"2a",
           378 => x"38",
           379 => x"95",
           380 => x"26",
           381 => x"84",
           382 => x"18",
           383 => x"38",
           384 => x"80",
           385 => x"38",
           386 => x"f6",
           387 => x"71",
           388 => x"58",
           389 => x"52",
           390 => x"c8",
           391 => x"08",
           392 => x"26",
           393 => x"05",
           394 => x"34",
           395 => x"84",
           396 => x"08",
           397 => x"98",
           398 => x"80",
           399 => x"29",
           400 => x"59",
           401 => x"55",
           402 => x"84",
           403 => x"53",
           404 => x"80",
           405 => x"72",
           406 => x"81",
           407 => x"38",
           408 => x"54",
           409 => x"7a",
           410 => x"71",
           411 => x"06",
           412 => x"77",
           413 => x"7c",
           414 => x"80",
           415 => x"81",
           416 => x"84",
           417 => x"38",
           418 => x"86",
           419 => x"85",
           420 => x"5f",
           421 => x"84",
           422 => x"70",
           423 => x"25",
           424 => x"a9",
           425 => x"fc",
           426 => x"40",
           427 => x"81",
           428 => x"78",
           429 => x"0a",
           430 => x"80",
           431 => x"51",
           432 => x"0a",
           433 => x"2c",
           434 => x"38",
           435 => x"55",
           436 => x"80",
           437 => x"f3",
           438 => x"2e",
           439 => x"2e",
           440 => x"33",
           441 => x"b9",
           442 => x"74",
           443 => x"a7",
           444 => x"fc",
           445 => x"40",
           446 => x"7c",
           447 => x"39",
           448 => x"7c",
           449 => x"fa",
           450 => x"80",
           451 => x"71",
           452 => x"59",
           453 => x"60",
           454 => x"83",
           455 => x"7c",
           456 => x"05",
           457 => x"57",
           458 => x"06",
           459 => x"78",
           460 => x"05",
           461 => x"7f",
           462 => x"51",
           463 => x"70",
           464 => x"83",
           465 => x"52",
           466 => x"85",
           467 => x"83",
           468 => x"ff",
           469 => x"75",
           470 => x"b9",
           471 => x"81",
           472 => x"29",
           473 => x"5a",
           474 => x"70",
           475 => x"c6",
           476 => x"05",
           477 => x"80",
           478 => x"ff",
           479 => x"fa",
           480 => x"58",
           481 => x"39",
           482 => x"58",
           483 => x"39",
           484 => x"81",
           485 => x"8a",
           486 => x"b9",
           487 => x"71",
           488 => x"2c",
           489 => x"07",
           490 => x"38",
           491 => x"71",
           492 => x"54",
           493 => x"bb",
           494 => x"ff",
           495 => x"5a",
           496 => x"33",
           497 => x"c9",
           498 => x"fc",
           499 => x"54",
           500 => x"7c",
           501 => x"39",
           502 => x"79",
           503 => x"38",
           504 => x"7a",
           505 => x"2e",
           506 => x"98",
           507 => x"90",
           508 => x"51",
           509 => x"39",
           510 => x"7e",
           511 => x"a2",
           512 => x"98",
           513 => x"06",
           514 => x"fb",
           515 => x"70",
           516 => x"7c",
           517 => x"39",
           518 => x"ff",
           519 => x"8b",
           520 => x"ff",
           521 => x"5a",
           522 => x"30",
           523 => x"5b",
           524 => x"d5",
           525 => x"f3",
           526 => x"3d",
           527 => x"ac",
           528 => x"81",
           529 => x"55",
           530 => x"81",
           531 => x"05",
           532 => x"38",
           533 => x"90",
           534 => x"c8",
           535 => x"74",
           536 => x"80",
           537 => x"54",
           538 => x"84",
           539 => x"14",
           540 => x"08",
           541 => x"56",
           542 => x"0d",
           543 => x"54",
           544 => x"2a",
           545 => x"57",
           546 => x"81",
           547 => x"55",
           548 => x"06",
           549 => x"c8",
           550 => x"81",
           551 => x"ea",
           552 => x"08",
           553 => x"80",
           554 => x"05",
           555 => x"ca",
           556 => x"08",
           557 => x"0d",
           558 => x"11",
           559 => x"06",
           560 => x"ae",
           561 => x"73",
           562 => x"53",
           563 => x"74",
           564 => x"81",
           565 => x"81",
           566 => x"84",
           567 => x"74",
           568 => x"15",
           569 => x"b9",
           570 => x"81",
           571 => x"39",
           572 => x"70",
           573 => x"06",
           574 => x"b3",
           575 => x"71",
           576 => x"52",
           577 => x"08",
           578 => x"80",
           579 => x"16",
           580 => x"81",
           581 => x"0c",
           582 => x"06",
           583 => x"08",
           584 => x"33",
           585 => x"04",
           586 => x"2d",
           587 => x"c8",
           588 => x"16",
           589 => x"b9",
           590 => x"a0",
           591 => x"54",
           592 => x"0d",
           593 => x"17",
           594 => x"0d",
           595 => x"70",
           596 => x"38",
           597 => x"54",
           598 => x"54",
           599 => x"c8",
           600 => x"0d",
           601 => x"54",
           602 => x"27",
           603 => x"71",
           604 => x"81",
           605 => x"ef",
           606 => x"3d",
           607 => x"27",
           608 => x"ff",
           609 => x"73",
           610 => x"d9",
           611 => x"71",
           612 => x"df",
           613 => x"70",
           614 => x"33",
           615 => x"74",
           616 => x"3d",
           617 => x"71",
           618 => x"54",
           619 => x"54",
           620 => x"c8",
           621 => x"0d",
           622 => x"54",
           623 => x"81",
           624 => x"55",
           625 => x"73",
           626 => x"04",
           627 => x"56",
           628 => x"33",
           629 => x"52",
           630 => x"38",
           631 => x"38",
           632 => x"51",
           633 => x"0d",
           634 => x"33",
           635 => x"38",
           636 => x"80",
           637 => x"b9",
           638 => x"84",
           639 => x"fb",
           640 => x"56",
           641 => x"84",
           642 => x"81",
           643 => x"54",
           644 => x"38",
           645 => x"74",
           646 => x"c8",
           647 => x"c8",
           648 => x"87",
           649 => x"77",
           650 => x"80",
           651 => x"54",
           652 => x"ff",
           653 => x"06",
           654 => x"52",
           655 => x"3d",
           656 => x"79",
           657 => x"2e",
           658 => x"54",
           659 => x"73",
           660 => x"04",
           661 => x"a0",
           662 => x"51",
           663 => x"52",
           664 => x"38",
           665 => x"b9",
           666 => x"9f",
           667 => x"9f",
           668 => x"71",
           669 => x"57",
           670 => x"2e",
           671 => x"07",
           672 => x"ff",
           673 => x"72",
           674 => x"56",
           675 => x"da",
           676 => x"84",
           677 => x"fc",
           678 => x"06",
           679 => x"70",
           680 => x"2a",
           681 => x"70",
           682 => x"74",
           683 => x"30",
           684 => x"31",
           685 => x"05",
           686 => x"25",
           687 => x"70",
           688 => x"70",
           689 => x"05",
           690 => x"55",
           691 => x"55",
           692 => x"56",
           693 => x"3d",
           694 => x"54",
           695 => x"08",
           696 => x"c8",
           697 => x"3d",
           698 => x"76",
           699 => x"cf",
           700 => x"13",
           701 => x"51",
           702 => x"08",
           703 => x"80",
           704 => x"be",
           705 => x"72",
           706 => x"55",
           707 => x"72",
           708 => x"77",
           709 => x"2c",
           710 => x"71",
           711 => x"55",
           712 => x"84",
           713 => x"fa",
           714 => x"2c",
           715 => x"2c",
           716 => x"31",
           717 => x"59",
           718 => x"c8",
           719 => x"c8",
           720 => x"0d",
           721 => x"0c",
           722 => x"73",
           723 => x"81",
           724 => x"55",
           725 => x"2e",
           726 => x"83",
           727 => x"89",
           728 => x"56",
           729 => x"e0",
           730 => x"81",
           731 => x"81",
           732 => x"8f",
           733 => x"54",
           734 => x"72",
           735 => x"29",
           736 => x"33",
           737 => x"be",
           738 => x"30",
           739 => x"84",
           740 => x"81",
           741 => x"56",
           742 => x"06",
           743 => x"0c",
           744 => x"2e",
           745 => x"2e",
           746 => x"c6",
           747 => x"58",
           748 => x"84",
           749 => x"82",
           750 => x"33",
           751 => x"80",
           752 => x"0d",
           753 => x"57",
           754 => x"33",
           755 => x"81",
           756 => x"0c",
           757 => x"f3",
           758 => x"73",
           759 => x"58",
           760 => x"38",
           761 => x"80",
           762 => x"38",
           763 => x"53",
           764 => x"53",
           765 => x"70",
           766 => x"27",
           767 => x"83",
           768 => x"70",
           769 => x"73",
           770 => x"2e",
           771 => x"0c",
           772 => x"8b",
           773 => x"79",
           774 => x"b0",
           775 => x"81",
           776 => x"55",
           777 => x"58",
           778 => x"56",
           779 => x"53",
           780 => x"fe",
           781 => x"8b",
           782 => x"70",
           783 => x"56",
           784 => x"c8",
           785 => x"e2",
           786 => x"06",
           787 => x"0d",
           788 => x"71",
           789 => x"71",
           790 => x"be",
           791 => x"ac",
           792 => x"04",
           793 => x"83",
           794 => x"ef",
           795 => x"ce",
           796 => x"0d",
           797 => x"3f",
           798 => x"51",
           799 => x"83",
           800 => x"3d",
           801 => x"e6",
           802 => x"f0",
           803 => x"04",
           804 => x"83",
           805 => x"ee",
           806 => x"d0",
           807 => x"0d",
           808 => x"3f",
           809 => x"51",
           810 => x"83",
           811 => x"3d",
           812 => x"8e",
           813 => x"98",
           814 => x"04",
           815 => x"83",
           816 => x"ed",
           817 => x"d1",
           818 => x"0d",
           819 => x"05",
           820 => x"68",
           821 => x"51",
           822 => x"ff",
           823 => x"07",
           824 => x"57",
           825 => x"52",
           826 => x"d9",
           827 => x"b9",
           828 => x"77",
           829 => x"70",
           830 => x"9f",
           831 => x"77",
           832 => x"88",
           833 => x"e0",
           834 => x"51",
           835 => x"54",
           836 => x"d1",
           837 => x"b9",
           838 => x"b9",
           839 => x"84",
           840 => x"05",
           841 => x"51",
           842 => x"08",
           843 => x"38",
           844 => x"38",
           845 => x"39",
           846 => x"3f",
           847 => x"f4",
           848 => x"83",
           849 => x"d0",
           850 => x"f8",
           851 => x"05",
           852 => x"7b",
           853 => x"b9",
           854 => x"91",
           855 => x"84",
           856 => x"78",
           857 => x"60",
           858 => x"7e",
           859 => x"84",
           860 => x"f3",
           861 => x"05",
           862 => x"68",
           863 => x"78",
           864 => x"83",
           865 => x"d2",
           866 => x"73",
           867 => x"81",
           868 => x"38",
           869 => x"a7",
           870 => x"51",
           871 => x"ac",
           872 => x"3f",
           873 => x"90",
           874 => x"79",
           875 => x"33",
           876 => x"83",
           877 => x"27",
           878 => x"70",
           879 => x"2e",
           880 => x"ee",
           881 => x"51",
           882 => x"76",
           883 => x"e9",
           884 => x"58",
           885 => x"c8",
           886 => x"54",
           887 => x"9b",
           888 => x"76",
           889 => x"84",
           890 => x"83",
           891 => x"14",
           892 => x"51",
           893 => x"b8",
           894 => x"51",
           895 => x"ac",
           896 => x"3f",
           897 => x"18",
           898 => x"22",
           899 => x"3f",
           900 => x"54",
           901 => x"26",
           902 => x"a4",
           903 => x"d5",
           904 => x"a9",
           905 => x"73",
           906 => x"72",
           907 => x"ab",
           908 => x"53",
           909 => x"74",
           910 => x"d5",
           911 => x"3f",
           912 => x"ce",
           913 => x"ff",
           914 => x"fc",
           915 => x"2e",
           916 => x"59",
           917 => x"3f",
           918 => x"98",
           919 => x"9b",
           920 => x"75",
           921 => x"58",
           922 => x"80",
           923 => x"08",
           924 => x"32",
           925 => x"70",
           926 => x"55",
           927 => x"24",
           928 => x"0b",
           929 => x"04",
           930 => x"08",
           931 => x"88",
           932 => x"3f",
           933 => x"2a",
           934 => x"b7",
           935 => x"51",
           936 => x"2a",
           937 => x"db",
           938 => x"51",
           939 => x"2a",
           940 => x"ff",
           941 => x"51",
           942 => x"2a",
           943 => x"38",
           944 => x"88",
           945 => x"04",
           946 => x"d8",
           947 => x"88",
           948 => x"04",
           949 => x"ec",
           950 => x"f0",
           951 => x"72",
           952 => x"51",
           953 => x"9b",
           954 => x"72",
           955 => x"71",
           956 => x"81",
           957 => x"51",
           958 => x"3f",
           959 => x"52",
           960 => x"be",
           961 => x"d4",
           962 => x"9b",
           963 => x"06",
           964 => x"38",
           965 => x"3f",
           966 => x"80",
           967 => x"70",
           968 => x"fe",
           969 => x"9a",
           970 => x"e8",
           971 => x"83",
           972 => x"80",
           973 => x"81",
           974 => x"51",
           975 => x"3f",
           976 => x"52",
           977 => x"bd",
           978 => x"41",
           979 => x"81",
           980 => x"84",
           981 => x"3d",
           982 => x"38",
           983 => x"98",
           984 => x"c3",
           985 => x"52",
           986 => x"83",
           987 => x"5b",
           988 => x"79",
           989 => x"ff",
           990 => x"38",
           991 => x"83",
           992 => x"2e",
           993 => x"70",
           994 => x"38",
           995 => x"7b",
           996 => x"08",
           997 => x"c8",
           998 => x"53",
           999 => x"84",
          1000 => x"33",
          1001 => x"81",
          1002 => x"9b",
          1003 => x"5c",
          1004 => x"f8",
          1005 => x"b9",
          1006 => x"80",
          1007 => x"08",
          1008 => x"91",
          1009 => x"62",
          1010 => x"84",
          1011 => x"8b",
          1012 => x"80",
          1013 => x"5b",
          1014 => x"82",
          1015 => x"82",
          1016 => x"d5",
          1017 => x"83",
          1018 => x"7d",
          1019 => x"0a",
          1020 => x"f5",
          1021 => x"b9",
          1022 => x"07",
          1023 => x"5a",
          1024 => x"78",
          1025 => x"38",
          1026 => x"5a",
          1027 => x"61",
          1028 => x"38",
          1029 => x"51",
          1030 => x"51",
          1031 => x"53",
          1032 => x"0b",
          1033 => x"ff",
          1034 => x"81",
          1035 => x"d8",
          1036 => x"c8",
          1037 => x"0b",
          1038 => x"53",
          1039 => x"c8",
          1040 => x"a0",
          1041 => x"e6",
          1042 => x"70",
          1043 => x"2e",
          1044 => x"39",
          1045 => x"3f",
          1046 => x"34",
          1047 => x"7e",
          1048 => x"5a",
          1049 => x"1a",
          1050 => x"81",
          1051 => x"10",
          1052 => x"04",
          1053 => x"51",
          1054 => x"84",
          1055 => x"84",
          1056 => x"06",
          1057 => x"45",
          1058 => x"fc",
          1059 => x"92",
          1060 => x"8c",
          1061 => x"80",
          1062 => x"d2",
          1063 => x"ab",
          1064 => x"fa",
          1065 => x"a4",
          1066 => x"3f",
          1067 => x"de",
          1068 => x"d6",
          1069 => x"3f",
          1070 => x"11",
          1071 => x"3f",
          1072 => x"ba",
          1073 => x"d0",
          1074 => x"b9",
          1075 => x"84",
          1076 => x"51",
          1077 => x"3d",
          1078 => x"51",
          1079 => x"80",
          1080 => x"d7",
          1081 => x"78",
          1082 => x"ff",
          1083 => x"b9",
          1084 => x"b8",
          1085 => x"05",
          1086 => x"08",
          1087 => x"53",
          1088 => x"83",
          1089 => x"f8",
          1090 => x"48",
          1091 => x"a2",
          1092 => x"64",
          1093 => x"b8",
          1094 => x"05",
          1095 => x"08",
          1096 => x"fe",
          1097 => x"e8",
          1098 => x"b0",
          1099 => x"52",
          1100 => x"84",
          1101 => x"7e",
          1102 => x"33",
          1103 => x"78",
          1104 => x"05",
          1105 => x"ff",
          1106 => x"e9",
          1107 => x"2e",
          1108 => x"11",
          1109 => x"3f",
          1110 => x"8a",
          1111 => x"ff",
          1112 => x"b9",
          1113 => x"83",
          1114 => x"67",
          1115 => x"38",
          1116 => x"5a",
          1117 => x"79",
          1118 => x"d7",
          1119 => x"5b",
          1120 => x"d2",
          1121 => x"ff",
          1122 => x"b9",
          1123 => x"b8",
          1124 => x"05",
          1125 => x"08",
          1126 => x"fe",
          1127 => x"e8",
          1128 => x"2e",
          1129 => x"cd",
          1130 => x"82",
          1131 => x"05",
          1132 => x"46",
          1133 => x"53",
          1134 => x"84",
          1135 => x"38",
          1136 => x"80",
          1137 => x"c8",
          1138 => x"52",
          1139 => x"84",
          1140 => x"7e",
          1141 => x"33",
          1142 => x"78",
          1143 => x"05",
          1144 => x"db",
          1145 => x"49",
          1146 => x"80",
          1147 => x"c8",
          1148 => x"59",
          1149 => x"68",
          1150 => x"11",
          1151 => x"3f",
          1152 => x"f5",
          1153 => x"53",
          1154 => x"84",
          1155 => x"38",
          1156 => x"80",
          1157 => x"c8",
          1158 => x"3d",
          1159 => x"51",
          1160 => x"86",
          1161 => x"d8",
          1162 => x"5b",
          1163 => x"5b",
          1164 => x"79",
          1165 => x"f1",
          1166 => x"80",
          1167 => x"c8",
          1168 => x"59",
          1169 => x"c8",
          1170 => x"84",
          1171 => x"38",
          1172 => x"3f",
          1173 => x"11",
          1174 => x"3f",
          1175 => x"f2",
          1176 => x"c0",
          1177 => x"3d",
          1178 => x"51",
          1179 => x"91",
          1180 => x"80",
          1181 => x"08",
          1182 => x"ff",
          1183 => x"b9",
          1184 => x"66",
          1185 => x"81",
          1186 => x"72",
          1187 => x"5d",
          1188 => x"2e",
          1189 => x"51",
          1190 => x"65",
          1191 => x"3f",
          1192 => x"f2",
          1193 => x"64",
          1194 => x"11",
          1195 => x"3f",
          1196 => x"da",
          1197 => x"84",
          1198 => x"53",
          1199 => x"84",
          1200 => x"39",
          1201 => x"7e",
          1202 => x"b8",
          1203 => x"05",
          1204 => x"08",
          1205 => x"02",
          1206 => x"05",
          1207 => x"f0",
          1208 => x"bd",
          1209 => x"38",
          1210 => x"11",
          1211 => x"3f",
          1212 => x"dc",
          1213 => x"33",
          1214 => x"9b",
          1215 => x"ff",
          1216 => x"b9",
          1217 => x"64",
          1218 => x"70",
          1219 => x"2e",
          1220 => x"55",
          1221 => x"d8",
          1222 => x"f3",
          1223 => x"8a",
          1224 => x"51",
          1225 => x"3d",
          1226 => x"51",
          1227 => x"80",
          1228 => x"ce",
          1229 => x"23",
          1230 => x"cd",
          1231 => x"38",
          1232 => x"39",
          1233 => x"2e",
          1234 => x"fc",
          1235 => x"d6",
          1236 => x"d8",
          1237 => x"f6",
          1238 => x"78",
          1239 => x"08",
          1240 => x"51",
          1241 => x"f2",
          1242 => x"38",
          1243 => x"39",
          1244 => x"2e",
          1245 => x"fb",
          1246 => x"7d",
          1247 => x"08",
          1248 => x"33",
          1249 => x"f2",
          1250 => x"f2",
          1251 => x"38",
          1252 => x"39",
          1253 => x"49",
          1254 => x"88",
          1255 => x"0d",
          1256 => x"c0",
          1257 => x"84",
          1258 => x"84",
          1259 => x"57",
          1260 => x"da",
          1261 => x"07",
          1262 => x"08",
          1263 => x"51",
          1264 => x"90",
          1265 => x"80",
          1266 => x"84",
          1267 => x"80",
          1268 => x"8c",
          1269 => x"0c",
          1270 => x"5d",
          1271 => x"80",
          1272 => x"70",
          1273 => x"d5",
          1274 => x"9e",
          1275 => x"95",
          1276 => x"d2",
          1277 => x"b8",
          1278 => x"83",
          1279 => x"81",
          1280 => x"c4",
          1281 => x"ec",
          1282 => x"d2",
          1283 => x"0a",
          1284 => x"3f",
          1285 => x"0d",
          1286 => x"52",
          1287 => x"74",
          1288 => x"70",
          1289 => x"81",
          1290 => x"53",
          1291 => x"71",
          1292 => x"81",
          1293 => x"80",
          1294 => x"ff",
          1295 => x"83",
          1296 => x"38",
          1297 => x"52",
          1298 => x"52",
          1299 => x"83",
          1300 => x"30",
          1301 => x"53",
          1302 => x"70",
          1303 => x"74",
          1304 => x"3d",
          1305 => x"73",
          1306 => x"52",
          1307 => x"53",
          1308 => x"81",
          1309 => x"75",
          1310 => x"06",
          1311 => x"0d",
          1312 => x"0b",
          1313 => x"04",
          1314 => x"da",
          1315 => x"2e",
          1316 => x"86",
          1317 => x"82",
          1318 => x"52",
          1319 => x"13",
          1320 => x"9e",
          1321 => x"51",
          1322 => x"38",
          1323 => x"bb",
          1324 => x"55",
          1325 => x"38",
          1326 => x"87",
          1327 => x"22",
          1328 => x"80",
          1329 => x"9c",
          1330 => x"0c",
          1331 => x"0c",
          1332 => x"0c",
          1333 => x"0c",
          1334 => x"0c",
          1335 => x"0c",
          1336 => x"87",
          1337 => x"c0",
          1338 => x"b9",
          1339 => x"3d",
          1340 => x"5d",
          1341 => x"08",
          1342 => x"b8",
          1343 => x"c0",
          1344 => x"34",
          1345 => x"84",
          1346 => x"5a",
          1347 => x"a8",
          1348 => x"c0",
          1349 => x"23",
          1350 => x"8a",
          1351 => x"ff",
          1352 => x"06",
          1353 => x"33",
          1354 => x"33",
          1355 => x"ff",
          1356 => x"ff",
          1357 => x"fe",
          1358 => x"72",
          1359 => x"e8",
          1360 => x"2b",
          1361 => x"2e",
          1362 => x"2e",
          1363 => x"84",
          1364 => x"ff",
          1365 => x"70",
          1366 => x"09",
          1367 => x"e7",
          1368 => x"2b",
          1369 => x"2e",
          1370 => x"80",
          1371 => x"81",
          1372 => x"c8",
          1373 => x"52",
          1374 => x"07",
          1375 => x"db",
          1376 => x"3d",
          1377 => x"05",
          1378 => x"ff",
          1379 => x"80",
          1380 => x"70",
          1381 => x"52",
          1382 => x"2a",
          1383 => x"38",
          1384 => x"80",
          1385 => x"06",
          1386 => x"06",
          1387 => x"80",
          1388 => x"52",
          1389 => x"0c",
          1390 => x"70",
          1391 => x"72",
          1392 => x"2e",
          1393 => x"52",
          1394 => x"94",
          1395 => x"06",
          1396 => x"39",
          1397 => x"70",
          1398 => x"70",
          1399 => x"04",
          1400 => x"33",
          1401 => x"80",
          1402 => x"33",
          1403 => x"71",
          1404 => x"94",
          1405 => x"06",
          1406 => x"38",
          1407 => x"51",
          1408 => x"06",
          1409 => x"93",
          1410 => x"75",
          1411 => x"80",
          1412 => x"c0",
          1413 => x"17",
          1414 => x"38",
          1415 => x"0d",
          1416 => x"51",
          1417 => x"81",
          1418 => x"71",
          1419 => x"2e",
          1420 => x"08",
          1421 => x"54",
          1422 => x"3d",
          1423 => x"9c",
          1424 => x"2e",
          1425 => x"08",
          1426 => x"a8",
          1427 => x"9e",
          1428 => x"c0",
          1429 => x"87",
          1430 => x"0c",
          1431 => x"98",
          1432 => x"f2",
          1433 => x"83",
          1434 => x"08",
          1435 => x"b8",
          1436 => x"9e",
          1437 => x"c0",
          1438 => x"87",
          1439 => x"0c",
          1440 => x"83",
          1441 => x"08",
          1442 => x"88",
          1443 => x"9e",
          1444 => x"0b",
          1445 => x"c0",
          1446 => x"06",
          1447 => x"71",
          1448 => x"c0",
          1449 => x"06",
          1450 => x"38",
          1451 => x"80",
          1452 => x"90",
          1453 => x"80",
          1454 => x"f2",
          1455 => x"90",
          1456 => x"52",
          1457 => x"52",
          1458 => x"87",
          1459 => x"80",
          1460 => x"83",
          1461 => x"34",
          1462 => x"70",
          1463 => x"70",
          1464 => x"83",
          1465 => x"9e",
          1466 => x"51",
          1467 => x"81",
          1468 => x"0b",
          1469 => x"80",
          1470 => x"2e",
          1471 => x"d0",
          1472 => x"08",
          1473 => x"52",
          1474 => x"71",
          1475 => x"c0",
          1476 => x"06",
          1477 => x"38",
          1478 => x"80",
          1479 => x"a0",
          1480 => x"2e",
          1481 => x"d3",
          1482 => x"80",
          1483 => x"83",
          1484 => x"9e",
          1485 => x"52",
          1486 => x"52",
          1487 => x"9e",
          1488 => x"2a",
          1489 => x"80",
          1490 => x"88",
          1491 => x"83",
          1492 => x"34",
          1493 => x"51",
          1494 => x"0d",
          1495 => x"3d",
          1496 => x"c3",
          1497 => x"86",
          1498 => x"9e",
          1499 => x"85",
          1500 => x"73",
          1501 => x"56",
          1502 => x"33",
          1503 => x"ce",
          1504 => x"f2",
          1505 => x"83",
          1506 => x"38",
          1507 => x"e2",
          1508 => x"83",
          1509 => x"73",
          1510 => x"55",
          1511 => x"33",
          1512 => x"d2",
          1513 => x"d9",
          1514 => x"ac",
          1515 => x"b5",
          1516 => x"83",
          1517 => x"83",
          1518 => x"51",
          1519 => x"51",
          1520 => x"52",
          1521 => x"3f",
          1522 => x"c0",
          1523 => x"b9",
          1524 => x"71",
          1525 => x"52",
          1526 => x"3f",
          1527 => x"38",
          1528 => x"38",
          1529 => x"08",
          1530 => x"c9",
          1531 => x"84",
          1532 => x"84",
          1533 => x"51",
          1534 => x"04",
          1535 => x"c0",
          1536 => x"b9",
          1537 => x"71",
          1538 => x"52",
          1539 => x"3f",
          1540 => x"2e",
          1541 => x"db",
          1542 => x"b0",
          1543 => x"08",
          1544 => x"c3",
          1545 => x"d9",
          1546 => x"f2",
          1547 => x"ff",
          1548 => x"c0",
          1549 => x"83",
          1550 => x"83",
          1551 => x"52",
          1552 => x"c8",
          1553 => x"31",
          1554 => x"83",
          1555 => x"83",
          1556 => x"fe",
          1557 => x"f0",
          1558 => x"d2",
          1559 => x"38",
          1560 => x"ff",
          1561 => x"56",
          1562 => x"39",
          1563 => x"3f",
          1564 => x"2e",
          1565 => x"90",
          1566 => x"cb",
          1567 => x"38",
          1568 => x"83",
          1569 => x"83",
          1570 => x"fc",
          1571 => x"33",
          1572 => x"e3",
          1573 => x"80",
          1574 => x"f2",
          1575 => x"ff",
          1576 => x"54",
          1577 => x"39",
          1578 => x"08",
          1579 => x"ff",
          1580 => x"56",
          1581 => x"39",
          1582 => x"08",
          1583 => x"ff",
          1584 => x"54",
          1585 => x"39",
          1586 => x"08",
          1587 => x"ff",
          1588 => x"55",
          1589 => x"39",
          1590 => x"08",
          1591 => x"ff",
          1592 => x"56",
          1593 => x"39",
          1594 => x"08",
          1595 => x"ff",
          1596 => x"54",
          1597 => x"39",
          1598 => x"3f",
          1599 => x"3f",
          1600 => x"2e",
          1601 => x"0d",
          1602 => x"26",
          1603 => x"fc",
          1604 => x"a4",
          1605 => x"0d",
          1606 => x"d3",
          1607 => x"b4",
          1608 => x"0d",
          1609 => x"bb",
          1610 => x"c4",
          1611 => x"0d",
          1612 => x"a3",
          1613 => x"80",
          1614 => x"84",
          1615 => x"c0",
          1616 => x"aa",
          1617 => x"81",
          1618 => x"b4",
          1619 => x"b9",
          1620 => x"57",
          1621 => x"55",
          1622 => x"90",
          1623 => x"a4",
          1624 => x"b9",
          1625 => x"0b",
          1626 => x"84",
          1627 => x"55",
          1628 => x"30",
          1629 => x"55",
          1630 => x"b0",
          1631 => x"08",
          1632 => x"b9",
          1633 => x"9a",
          1634 => x"3d",
          1635 => x"ad",
          1636 => x"06",
          1637 => x"9a",
          1638 => x"ab",
          1639 => x"76",
          1640 => x"ff",
          1641 => x"c8",
          1642 => x"0d",
          1643 => x"72",
          1644 => x"73",
          1645 => x"8d",
          1646 => x"83",
          1647 => x"ff",
          1648 => x"53",
          1649 => x"3f",
          1650 => x"14",
          1651 => x"38",
          1652 => x"70",
          1653 => x"27",
          1654 => x"c8",
          1655 => x"5a",
          1656 => x"80",
          1657 => x"c8",
          1658 => x"53",
          1659 => x"84",
          1660 => x"73",
          1661 => x"81",
          1662 => x"fe",
          1663 => x"77",
          1664 => x"38",
          1665 => x"55",
          1666 => x"d5",
          1667 => x"0b",
          1668 => x"73",
          1669 => x"b4",
          1670 => x"84",
          1671 => x"f3",
          1672 => x"51",
          1673 => x"08",
          1674 => x"bd",
          1675 => x"80",
          1676 => x"38",
          1677 => x"19",
          1678 => x"75",
          1679 => x"56",
          1680 => x"09",
          1681 => x"84",
          1682 => x"ce",
          1683 => x"08",
          1684 => x"0b",
          1685 => x"83",
          1686 => x"38",
          1687 => x"74",
          1688 => x"2e",
          1689 => x"5a",
          1690 => x"2e",
          1691 => x"5f",
          1692 => x"b9",
          1693 => x"5b",
          1694 => x"81",
          1695 => x"98",
          1696 => x"33",
          1697 => x"98",
          1698 => x"d0",
          1699 => x"53",
          1700 => x"59",
          1701 => x"38",
          1702 => x"81",
          1703 => x"70",
          1704 => x"81",
          1705 => x"2b",
          1706 => x"16",
          1707 => x"38",
          1708 => x"33",
          1709 => x"38",
          1710 => x"d1",
          1711 => x"81",
          1712 => x"70",
          1713 => x"98",
          1714 => x"05",
          1715 => x"33",
          1716 => x"57",
          1717 => x"84",
          1718 => x"57",
          1719 => x"0a",
          1720 => x"2c",
          1721 => x"76",
          1722 => x"16",
          1723 => x"83",
          1724 => x"61",
          1725 => x"08",
          1726 => x"2e",
          1727 => x"bc",
          1728 => x"80",
          1729 => x"81",
          1730 => x"fe",
          1731 => x"76",
          1732 => x"76",
          1733 => x"fd",
          1734 => x"94",
          1735 => x"d8",
          1736 => x"d1",
          1737 => x"34",
          1738 => x"75",
          1739 => x"ac",
          1740 => x"3f",
          1741 => x"76",
          1742 => x"84",
          1743 => x"84",
          1744 => x"79",
          1745 => x"08",
          1746 => x"8c",
          1747 => x"ff",
          1748 => x"93",
          1749 => x"83",
          1750 => x"75",
          1751 => x"34",
          1752 => x"84",
          1753 => x"2e",
          1754 => x"88",
          1755 => x"ac",
          1756 => x"3f",
          1757 => x"ff",
          1758 => x"ff",
          1759 => x"7a",
          1760 => x"7b",
          1761 => x"d1",
          1762 => x"38",
          1763 => x"9e",
          1764 => x"05",
          1765 => x"f9",
          1766 => x"fb",
          1767 => x"3f",
          1768 => x"34",
          1769 => x"81",
          1770 => x"b8",
          1771 => x"d1",
          1772 => x"ff",
          1773 => x"88",
          1774 => x"ac",
          1775 => x"3f",
          1776 => x"ff",
          1777 => x"ff",
          1778 => x"74",
          1779 => x"d1",
          1780 => x"d1",
          1781 => x"27",
          1782 => x"52",
          1783 => x"34",
          1784 => x"b3",
          1785 => x"81",
          1786 => x"57",
          1787 => x"84",
          1788 => x"76",
          1789 => x"33",
          1790 => x"d1",
          1791 => x"d1",
          1792 => x"26",
          1793 => x"d1",
          1794 => x"56",
          1795 => x"15",
          1796 => x"98",
          1797 => x"06",
          1798 => x"ef",
          1799 => x"51",
          1800 => x"33",
          1801 => x"d1",
          1802 => x"77",
          1803 => x"08",
          1804 => x"74",
          1805 => x"05",
          1806 => x"5d",
          1807 => x"38",
          1808 => x"ff",
          1809 => x"29",
          1810 => x"84",
          1811 => x"75",
          1812 => x"7b",
          1813 => x"84",
          1814 => x"ff",
          1815 => x"29",
          1816 => x"84",
          1817 => x"79",
          1818 => x"81",
          1819 => x"08",
          1820 => x"3f",
          1821 => x"0a",
          1822 => x"33",
          1823 => x"a7",
          1824 => x"33",
          1825 => x"84",
          1826 => x"b0",
          1827 => x"05",
          1828 => x"81",
          1829 => x"88",
          1830 => x"84",
          1831 => x"b0",
          1832 => x"51",
          1833 => x"81",
          1834 => x"84",
          1835 => x"80",
          1836 => x"10",
          1837 => x"57",
          1838 => x"82",
          1839 => x"05",
          1840 => x"e7",
          1841 => x"0c",
          1842 => x"83",
          1843 => x"41",
          1844 => x"08",
          1845 => x"f3",
          1846 => x"bc",
          1847 => x"80",
          1848 => x"b9",
          1849 => x"d1",
          1850 => x"38",
          1851 => x"ff",
          1852 => x"52",
          1853 => x"d5",
          1854 => x"f9",
          1855 => x"56",
          1856 => x"ff",
          1857 => x"f0",
          1858 => x"84",
          1859 => x"88",
          1860 => x"80",
          1861 => x"33",
          1862 => x"d5",
          1863 => x"b1",
          1864 => x"51",
          1865 => x"08",
          1866 => x"84",
          1867 => x"84",
          1868 => x"55",
          1869 => x"ff",
          1870 => x"8c",
          1871 => x"7b",
          1872 => x"04",
          1873 => x"06",
          1874 => x"38",
          1875 => x"78",
          1876 => x"77",
          1877 => x"08",
          1878 => x"84",
          1879 => x"98",
          1880 => x"5b",
          1881 => x"84",
          1882 => x"ad",
          1883 => x"98",
          1884 => x"33",
          1885 => x"f3",
          1886 => x"88",
          1887 => x"80",
          1888 => x"98",
          1889 => x"55",
          1890 => x"d5",
          1891 => x"d1",
          1892 => x"80",
          1893 => x"88",
          1894 => x"ff",
          1895 => x"57",
          1896 => x"ac",
          1897 => x"a1",
          1898 => x"80",
          1899 => x"88",
          1900 => x"fe",
          1901 => x"33",
          1902 => x"76",
          1903 => x"81",
          1904 => x"70",
          1905 => x"57",
          1906 => x"fe",
          1907 => x"81",
          1908 => x"f2",
          1909 => x"76",
          1910 => x"70",
          1911 => x"a1",
          1912 => x"1c",
          1913 => x"ff",
          1914 => x"8c",
          1915 => x"e1",
          1916 => x"8c",
          1917 => x"5a",
          1918 => x"88",
          1919 => x"81",
          1920 => x"75",
          1921 => x"80",
          1922 => x"98",
          1923 => x"5c",
          1924 => x"77",
          1925 => x"ff",
          1926 => x"f1",
          1927 => x"88",
          1928 => x"80",
          1929 => x"98",
          1930 => x"41",
          1931 => x"d5",
          1932 => x"89",
          1933 => x"80",
          1934 => x"88",
          1935 => x"ff",
          1936 => x"e0",
          1937 => x"38",
          1938 => x"b9",
          1939 => x"b9",
          1940 => x"53",
          1941 => x"3f",
          1942 => x"33",
          1943 => x"38",
          1944 => x"ff",
          1945 => x"52",
          1946 => x"d5",
          1947 => x"91",
          1948 => x"5b",
          1949 => x"ff",
          1950 => x"e1",
          1951 => x"f3",
          1952 => x"a5",
          1953 => x"ef",
          1954 => x"ac",
          1955 => x"58",
          1956 => x"0a",
          1957 => x"2c",
          1958 => x"76",
          1959 => x"33",
          1960 => x"81",
          1961 => x"7a",
          1962 => x"83",
          1963 => x"38",
          1964 => x"08",
          1965 => x"18",
          1966 => x"80",
          1967 => x"b4",
          1968 => x"38",
          1969 => x"f3",
          1970 => x"80",
          1971 => x"b4",
          1972 => x"51",
          1973 => x"ff",
          1974 => x"25",
          1975 => x"51",
          1976 => x"08",
          1977 => x"08",
          1978 => x"52",
          1979 => x"0b",
          1980 => x"33",
          1981 => x"97",
          1982 => x"51",
          1983 => x"08",
          1984 => x"84",
          1985 => x"a6",
          1986 => x"05",
          1987 => x"81",
          1988 => x"34",
          1989 => x"0b",
          1990 => x"c8",
          1991 => x"ff",
          1992 => x"84",
          1993 => x"81",
          1994 => x"7b",
          1995 => x"70",
          1996 => x"84",
          1997 => x"74",
          1998 => x"ac",
          1999 => x"3f",
          2000 => x"ff",
          2001 => x"52",
          2002 => x"d1",
          2003 => x"d1",
          2004 => x"c7",
          2005 => x"84",
          2006 => x"84",
          2007 => x"05",
          2008 => x"a5",
          2009 => x"84",
          2010 => x"58",
          2011 => x"a7",
          2012 => x"51",
          2013 => x"08",
          2014 => x"84",
          2015 => x"a4",
          2016 => x"05",
          2017 => x"81",
          2018 => x"80",
          2019 => x"70",
          2020 => x"e0",
          2021 => x"56",
          2022 => x"08",
          2023 => x"10",
          2024 => x"57",
          2025 => x"38",
          2026 => x"a8",
          2027 => x"05",
          2028 => x"79",
          2029 => x"b8",
          2030 => x"f8",
          2031 => x"51",
          2032 => x"08",
          2033 => x"83",
          2034 => x"3f",
          2035 => x"0b",
          2036 => x"c8",
          2037 => x"77",
          2038 => x"c9",
          2039 => x"a5",
          2040 => x"5c",
          2041 => x"f8",
          2042 => x"84",
          2043 => x"08",
          2044 => x"38",
          2045 => x"bb",
          2046 => x"0b",
          2047 => x"38",
          2048 => x"1b",
          2049 => x"ff",
          2050 => x"10",
          2051 => x"40",
          2052 => x"82",
          2053 => x"05",
          2054 => x"da",
          2055 => x"0c",
          2056 => x"83",
          2057 => x"41",
          2058 => x"ff",
          2059 => x"38",
          2060 => x"06",
          2061 => x"f9",
          2062 => x"51",
          2063 => x"33",
          2064 => x"57",
          2065 => x"0b",
          2066 => x"74",
          2067 => x"b8",
          2068 => x"83",
          2069 => x"52",
          2070 => x"b9",
          2071 => x"33",
          2072 => x"70",
          2073 => x"ff",
          2074 => x"f3",
          2075 => x"f3",
          2076 => x"b0",
          2077 => x"eb",
          2078 => x"02",
          2079 => x"80",
          2080 => x"26",
          2081 => x"8b",
          2082 => x"72",
          2083 => x"a0",
          2084 => x"5e",
          2085 => x"76",
          2086 => x"34",
          2087 => x"f8",
          2088 => x"98",
          2089 => x"2b",
          2090 => x"56",
          2091 => x"74",
          2092 => x"70",
          2093 => x"ee",
          2094 => x"f8",
          2095 => x"78",
          2096 => x"e0",
          2097 => x"56",
          2098 => x"90",
          2099 => x"0b",
          2100 => x"11",
          2101 => x"11",
          2102 => x"86",
          2103 => x"33",
          2104 => x"33",
          2105 => x"22",
          2106 => x"29",
          2107 => x"5d",
          2108 => x"31",
          2109 => x"7e",
          2110 => x"7a",
          2111 => x"06",
          2112 => x"57",
          2113 => x"83",
          2114 => x"70",
          2115 => x"06",
          2116 => x"78",
          2117 => x"c1",
          2118 => x"34",
          2119 => x"05",
          2120 => x"80",
          2121 => x"b7",
          2122 => x"b7",
          2123 => x"f8",
          2124 => x"5d",
          2125 => x"27",
          2126 => x"73",
          2127 => x"5a",
          2128 => x"38",
          2129 => x"0b",
          2130 => x"33",
          2131 => x"71",
          2132 => x"56",
          2133 => x"ae",
          2134 => x"38",
          2135 => x"06",
          2136 => x"33",
          2137 => x"80",
          2138 => x"86",
          2139 => x"bc",
          2140 => x"bb",
          2141 => x"f6",
          2142 => x"75",
          2143 => x"58",
          2144 => x"8b",
          2145 => x"29",
          2146 => x"74",
          2147 => x"83",
          2148 => x"70",
          2149 => x"55",
          2150 => x"29",
          2151 => x"06",
          2152 => x"83",
          2153 => x"f2",
          2154 => x"fe",
          2155 => x"80",
          2156 => x"73",
          2157 => x"86",
          2158 => x"34",
          2159 => x"98",
          2160 => x"86",
          2161 => x"80",
          2162 => x"52",
          2163 => x"87",
          2164 => x"56",
          2165 => x"84",
          2166 => x"08",
          2167 => x"51",
          2168 => x"cc",
          2169 => x"53",
          2170 => x"08",
          2171 => x"75",
          2172 => x"34",
          2173 => x"3d",
          2174 => x"b9",
          2175 => x"af",
          2176 => x"33",
          2177 => x"81",
          2178 => x"84",
          2179 => x"83",
          2180 => x"86",
          2181 => x"22",
          2182 => x"05",
          2183 => x"ce",
          2184 => x"2e",
          2185 => x"76",
          2186 => x"83",
          2187 => x"ff",
          2188 => x"55",
          2189 => x"19",
          2190 => x"f8",
          2191 => x"84",
          2192 => x"74",
          2193 => x"33",
          2194 => x"72",
          2195 => x"9a",
          2196 => x"33",
          2197 => x"05",
          2198 => x"34",
          2199 => x"27",
          2200 => x"38",
          2201 => x"15",
          2202 => x"34",
          2203 => x"81",
          2204 => x"38",
          2205 => x"75",
          2206 => x"81",
          2207 => x"54",
          2208 => x"72",
          2209 => x"33",
          2210 => x"55",
          2211 => x"b0",
          2212 => x"ff",
          2213 => x"54",
          2214 => x"98",
          2215 => x"53",
          2216 => x"81",
          2217 => x"55",
          2218 => x"81",
          2219 => x"bb",
          2220 => x"5a",
          2221 => x"53",
          2222 => x"0d",
          2223 => x"f8",
          2224 => x"84",
          2225 => x"7a",
          2226 => x"fe",
          2227 => x"05",
          2228 => x"75",
          2229 => x"73",
          2230 => x"33",
          2231 => x"56",
          2232 => x"ae",
          2233 => x"9a",
          2234 => x"a0",
          2235 => x"70",
          2236 => x"72",
          2237 => x"e0",
          2238 => x"05",
          2239 => x"38",
          2240 => x"bc",
          2241 => x"f8",
          2242 => x"19",
          2243 => x"59",
          2244 => x"02",
          2245 => x"70",
          2246 => x"83",
          2247 => x"84",
          2248 => x"86",
          2249 => x"0b",
          2250 => x"04",
          2251 => x"f8",
          2252 => x"52",
          2253 => x"51",
          2254 => x"84",
          2255 => x"83",
          2256 => x"09",
          2257 => x"53",
          2258 => x"39",
          2259 => x"b7",
          2260 => x"70",
          2261 => x"83",
          2262 => x"c8",
          2263 => x"f9",
          2264 => x"9f",
          2265 => x"70",
          2266 => x"b9",
          2267 => x"f8",
          2268 => x"33",
          2269 => x"25",
          2270 => x"f9",
          2271 => x"86",
          2272 => x"f9",
          2273 => x"bb",
          2274 => x"25",
          2275 => x"83",
          2276 => x"3d",
          2277 => x"b1",
          2278 => x"c4",
          2279 => x"f8",
          2280 => x"84",
          2281 => x"2a",
          2282 => x"f0",
          2283 => x"f2",
          2284 => x"84",
          2285 => x"83",
          2286 => x"07",
          2287 => x"0b",
          2288 => x"04",
          2289 => x"51",
          2290 => x"83",
          2291 => x"07",
          2292 => x"39",
          2293 => x"80",
          2294 => x"0d",
          2295 => x"06",
          2296 => x"34",
          2297 => x"87",
          2298 => x"ff",
          2299 => x"fd",
          2300 => x"f4",
          2301 => x"33",
          2302 => x"83",
          2303 => x"f8",
          2304 => x"51",
          2305 => x"39",
          2306 => x"51",
          2307 => x"39",
          2308 => x"80",
          2309 => x"34",
          2310 => x"81",
          2311 => x"f8",
          2312 => x"f4",
          2313 => x"51",
          2314 => x"39",
          2315 => x"80",
          2316 => x"34",
          2317 => x"81",
          2318 => x"f8",
          2319 => x"f4",
          2320 => x"f8",
          2321 => x"f4",
          2322 => x"70",
          2323 => x"f3",
          2324 => x"84",
          2325 => x"f8",
          2326 => x"f9",
          2327 => x"5f",
          2328 => x"a1",
          2329 => x"81",
          2330 => x"be",
          2331 => x"7a",
          2332 => x"f6",
          2333 => x"3d",
          2334 => x"06",
          2335 => x"34",
          2336 => x"0b",
          2337 => x"f8",
          2338 => x"23",
          2339 => x"84",
          2340 => x"33",
          2341 => x"83",
          2342 => x"7d",
          2343 => x"b7",
          2344 => x"7b",
          2345 => x"f9",
          2346 => x"84",
          2347 => x"c0",
          2348 => x"a8",
          2349 => x"83",
          2350 => x"58",
          2351 => x"c9",
          2352 => x"53",
          2353 => x"80",
          2354 => x"33",
          2355 => x"79",
          2356 => x"53",
          2357 => x"db",
          2358 => x"84",
          2359 => x"7a",
          2360 => x"ff",
          2361 => x"34",
          2362 => x"83",
          2363 => x"23",
          2364 => x"0d",
          2365 => x"81",
          2366 => x"83",
          2367 => x"f9",
          2368 => x"83",
          2369 => x"84",
          2370 => x"51",
          2371 => x"f7",
          2372 => x"84",
          2373 => x"83",
          2374 => x"fc",
          2375 => x"70",
          2376 => x"f9",
          2377 => x"05",
          2378 => x"f9",
          2379 => x"29",
          2380 => x"f8",
          2381 => x"7c",
          2382 => x"83",
          2383 => x"57",
          2384 => x"75",
          2385 => x"24",
          2386 => x"85",
          2387 => x"84",
          2388 => x"83",
          2389 => x"55",
          2390 => x"86",
          2391 => x"bc",
          2392 => x"f6",
          2393 => x"56",
          2394 => x"83",
          2395 => x"58",
          2396 => x"b0",
          2397 => x"70",
          2398 => x"83",
          2399 => x"57",
          2400 => x"33",
          2401 => x"70",
          2402 => x"26",
          2403 => x"58",
          2404 => x"72",
          2405 => x"33",
          2406 => x"b7",
          2407 => x"fb",
          2408 => x"89",
          2409 => x"38",
          2410 => x"8a",
          2411 => x"81",
          2412 => x"0b",
          2413 => x"83",
          2414 => x"c4",
          2415 => x"09",
          2416 => x"76",
          2417 => x"13",
          2418 => x"83",
          2419 => x"51",
          2420 => x"ff",
          2421 => x"38",
          2422 => x"34",
          2423 => x"f9",
          2424 => x"0c",
          2425 => x"2e",
          2426 => x"f8",
          2427 => x"ff",
          2428 => x"72",
          2429 => x"51",
          2430 => x"70",
          2431 => x"73",
          2432 => x"f8",
          2433 => x"83",
          2434 => x"ef",
          2435 => x"75",
          2436 => x"e6",
          2437 => x"84",
          2438 => x"2e",
          2439 => x"82",
          2440 => x"78",
          2441 => x"2e",
          2442 => x"8f",
          2443 => x"f8",
          2444 => x"29",
          2445 => x"19",
          2446 => x"84",
          2447 => x"83",
          2448 => x"5a",
          2449 => x"18",
          2450 => x"29",
          2451 => x"33",
          2452 => x"84",
          2453 => x"83",
          2454 => x"72",
          2455 => x"59",
          2456 => x"1f",
          2457 => x"42",
          2458 => x"84",
          2459 => x"38",
          2460 => x"34",
          2461 => x"3d",
          2462 => x"38",
          2463 => x"b8",
          2464 => x"2e",
          2465 => x"c4",
          2466 => x"f8",
          2467 => x"29",
          2468 => x"19",
          2469 => x"84",
          2470 => x"83",
          2471 => x"41",
          2472 => x"1f",
          2473 => x"29",
          2474 => x"86",
          2475 => x"bc",
          2476 => x"f6",
          2477 => x"29",
          2478 => x"f8",
          2479 => x"34",
          2480 => x"41",
          2481 => x"83",
          2482 => x"c8",
          2483 => x"2e",
          2484 => x"81",
          2485 => x"fd",
          2486 => x"34",
          2487 => x"3d",
          2488 => x"38",
          2489 => x"d0",
          2490 => x"59",
          2491 => x"84",
          2492 => x"06",
          2493 => x"34",
          2494 => x"3d",
          2495 => x"38",
          2496 => x"b7",
          2497 => x"f8",
          2498 => x"40",
          2499 => x"a7",
          2500 => x"33",
          2501 => x"22",
          2502 => x"56",
          2503 => x"f8",
          2504 => x"57",
          2505 => x"80",
          2506 => x"81",
          2507 => x"f8",
          2508 => x"42",
          2509 => x"60",
          2510 => x"58",
          2511 => x"ea",
          2512 => x"34",
          2513 => x"83",
          2514 => x"83",
          2515 => x"86",
          2516 => x"22",
          2517 => x"70",
          2518 => x"33",
          2519 => x"2e",
          2520 => x"ff",
          2521 => x"76",
          2522 => x"90",
          2523 => x"80",
          2524 => x"84",
          2525 => x"cb",
          2526 => x"80",
          2527 => x"0d",
          2528 => x"b0",
          2529 => x"b1",
          2530 => x"b2",
          2531 => x"80",
          2532 => x"0d",
          2533 => x"06",
          2534 => x"84",
          2535 => x"83",
          2536 => x"72",
          2537 => x"05",
          2538 => x"7b",
          2539 => x"83",
          2540 => x"42",
          2541 => x"38",
          2542 => x"56",
          2543 => x"f8",
          2544 => x"81",
          2545 => x"72",
          2546 => x"e4",
          2547 => x"84",
          2548 => x"83",
          2549 => x"5a",
          2550 => x"fa",
          2551 => x"71",
          2552 => x"f4",
          2553 => x"84",
          2554 => x"83",
          2555 => x"72",
          2556 => x"59",
          2557 => x"9a",
          2558 => x"06",
          2559 => x"38",
          2560 => x"d0",
          2561 => x"f9",
          2562 => x"ff",
          2563 => x"39",
          2564 => x"bd",
          2565 => x"95",
          2566 => x"7e",
          2567 => x"75",
          2568 => x"10",
          2569 => x"04",
          2570 => x"52",
          2571 => x"84",
          2572 => x"83",
          2573 => x"70",
          2574 => x"70",
          2575 => x"86",
          2576 => x"22",
          2577 => x"83",
          2578 => x"46",
          2579 => x"81",
          2580 => x"81",
          2581 => x"81",
          2582 => x"58",
          2583 => x"a0",
          2584 => x"83",
          2585 => x"72",
          2586 => x"a0",
          2587 => x"f8",
          2588 => x"5e",
          2589 => x"80",
          2590 => x"81",
          2591 => x"f8",
          2592 => x"44",
          2593 => x"84",
          2594 => x"70",
          2595 => x"26",
          2596 => x"58",
          2597 => x"75",
          2598 => x"81",
          2599 => x"f7",
          2600 => x"b7",
          2601 => x"81",
          2602 => x"81",
          2603 => x"5b",
          2604 => x"33",
          2605 => x"b7",
          2606 => x"f8",
          2607 => x"41",
          2608 => x"1c",
          2609 => x"29",
          2610 => x"86",
          2611 => x"bc",
          2612 => x"f6",
          2613 => x"29",
          2614 => x"f8",
          2615 => x"60",
          2616 => x"58",
          2617 => x"83",
          2618 => x"0b",
          2619 => x"b9",
          2620 => x"f8",
          2621 => x"19",
          2622 => x"70",
          2623 => x"f9",
          2624 => x"34",
          2625 => x"3d",
          2626 => x"5b",
          2627 => x"83",
          2628 => x"83",
          2629 => x"5c",
          2630 => x"9c",
          2631 => x"ff",
          2632 => x"80",
          2633 => x"33",
          2634 => x"c9",
          2635 => x"02",
          2636 => x"9c",
          2637 => x"fa",
          2638 => x"33",
          2639 => x"b7",
          2640 => x"5b",
          2641 => x"33",
          2642 => x"33",
          2643 => x"84",
          2644 => x"a0",
          2645 => x"83",
          2646 => x"72",
          2647 => x"78",
          2648 => x"f8",
          2649 => x"83",
          2650 => x"80",
          2651 => x"81",
          2652 => x"f8",
          2653 => x"5f",
          2654 => x"84",
          2655 => x"81",
          2656 => x"90",
          2657 => x"77",
          2658 => x"83",
          2659 => x"c4",
          2660 => x"80",
          2661 => x"33",
          2662 => x"81",
          2663 => x"b9",
          2664 => x"b9",
          2665 => x"b9",
          2666 => x"b9",
          2667 => x"23",
          2668 => x"84",
          2669 => x"84",
          2670 => x"84",
          2671 => x"b8",
          2672 => x"93",
          2673 => x"86",
          2674 => x"83",
          2675 => x"f8",
          2676 => x"83",
          2677 => x"57",
          2678 => x"fe",
          2679 => x"ff",
          2680 => x"05",
          2681 => x"76",
          2682 => x"bd",
          2683 => x"b8",
          2684 => x"06",
          2685 => x"77",
          2686 => x"33",
          2687 => x"38",
          2688 => x"5f",
          2689 => x"5e",
          2690 => x"f8",
          2691 => x"71",
          2692 => x"06",
          2693 => x"f8",
          2694 => x"c9",
          2695 => x"38",
          2696 => x"81",
          2697 => x"57",
          2698 => x"75",
          2699 => x"80",
          2700 => x"f8",
          2701 => x"7b",
          2702 => x"56",
          2703 => x"39",
          2704 => x"f8",
          2705 => x"05",
          2706 => x"38",
          2707 => x"34",
          2708 => x"40",
          2709 => x"f8",
          2710 => x"71",
          2711 => x"06",
          2712 => x"f8",
          2713 => x"c9",
          2714 => x"38",
          2715 => x"2e",
          2716 => x"b7",
          2717 => x"f8",
          2718 => x"a7",
          2719 => x"43",
          2720 => x"70",
          2721 => x"08",
          2722 => x"5d",
          2723 => x"bf",
          2724 => x"fb",
          2725 => x"79",
          2726 => x"9c",
          2727 => x"06",
          2728 => x"cd",
          2729 => x"33",
          2730 => x"84",
          2731 => x"5d",
          2732 => x"11",
          2733 => x"38",
          2734 => x"fb",
          2735 => x"76",
          2736 => x"9d",
          2737 => x"05",
          2738 => x"41",
          2739 => x"57",
          2740 => x"39",
          2741 => x"3f",
          2742 => x"57",
          2743 => x"10",
          2744 => x"5a",
          2745 => x"3f",
          2746 => x"b8",
          2747 => x"82",
          2748 => x"7d",
          2749 => x"22",
          2750 => x"57",
          2751 => x"d5",
          2752 => x"c9",
          2753 => x"38",
          2754 => x"81",
          2755 => x"05",
          2756 => x"33",
          2757 => x"43",
          2758 => x"27",
          2759 => x"f6",
          2760 => x"58",
          2761 => x"57",
          2762 => x"bc",
          2763 => x"27",
          2764 => x"f8",
          2765 => x"c9",
          2766 => x"38",
          2767 => x"33",
          2768 => x"38",
          2769 => x"33",
          2770 => x"33",
          2771 => x"80",
          2772 => x"71",
          2773 => x"06",
          2774 => x"59",
          2775 => x"38",
          2776 => x"31",
          2777 => x"38",
          2778 => x"27",
          2779 => x"83",
          2780 => x"70",
          2781 => x"8e",
          2782 => x"76",
          2783 => x"56",
          2784 => x"ff",
          2785 => x"80",
          2786 => x"77",
          2787 => x"71",
          2788 => x"86",
          2789 => x"80",
          2790 => x"06",
          2791 => x"5c",
          2792 => x"98",
          2793 => x"5f",
          2794 => x"81",
          2795 => x"58",
          2796 => x"81",
          2797 => x"bb",
          2798 => x"5e",
          2799 => x"e0",
          2800 => x"1f",
          2801 => x"76",
          2802 => x"81",
          2803 => x"bc",
          2804 => x"29",
          2805 => x"26",
          2806 => x"b8",
          2807 => x"e0",
          2808 => x"51",
          2809 => x"0b",
          2810 => x"b8",
          2811 => x"78",
          2812 => x"56",
          2813 => x"be",
          2814 => x"81",
          2815 => x"43",
          2816 => x"38",
          2817 => x"26",
          2818 => x"56",
          2819 => x"76",
          2820 => x"f5",
          2821 => x"90",
          2822 => x"11",
          2823 => x"80",
          2824 => x"75",
          2825 => x"76",
          2826 => x"70",
          2827 => x"88",
          2828 => x"52",
          2829 => x"80",
          2830 => x"76",
          2831 => x"26",
          2832 => x"b7",
          2833 => x"06",
          2834 => x"22",
          2835 => x"59",
          2836 => x"78",
          2837 => x"57",
          2838 => x"76",
          2839 => x"33",
          2840 => x"0b",
          2841 => x"81",
          2842 => x"76",
          2843 => x"e0",
          2844 => x"5a",
          2845 => x"d6",
          2846 => x"81",
          2847 => x"83",
          2848 => x"71",
          2849 => x"2a",
          2850 => x"2e",
          2851 => x"0b",
          2852 => x"81",
          2853 => x"83",
          2854 => x"c4",
          2855 => x"33",
          2856 => x"22",
          2857 => x"5d",
          2858 => x"87",
          2859 => x"81",
          2860 => x"f4",
          2861 => x"fd",
          2862 => x"f4",
          2863 => x"81",
          2864 => x"f8",
          2865 => x"33",
          2866 => x"83",
          2867 => x"f4",
          2868 => x"75",
          2869 => x"80",
          2870 => x"18",
          2871 => x"a4",
          2872 => x"06",
          2873 => x"8f",
          2874 => x"06",
          2875 => x"34",
          2876 => x"81",
          2877 => x"83",
          2878 => x"f8",
          2879 => x"07",
          2880 => x"d7",
          2881 => x"06",
          2882 => x"34",
          2883 => x"81",
          2884 => x"f8",
          2885 => x"f4",
          2886 => x"75",
          2887 => x"83",
          2888 => x"07",
          2889 => x"8f",
          2890 => x"06",
          2891 => x"ff",
          2892 => x"07",
          2893 => x"ef",
          2894 => x"07",
          2895 => x"df",
          2896 => x"06",
          2897 => x"f4",
          2898 => x"33",
          2899 => x"83",
          2900 => x"0b",
          2901 => x"51",
          2902 => x"b9",
          2903 => x"b9",
          2904 => x"b9",
          2905 => x"23",
          2906 => x"c7",
          2907 => x"80",
          2908 => x"0d",
          2909 => x"f8",
          2910 => x"ff",
          2911 => x"cc",
          2912 => x"05",
          2913 => x"c8",
          2914 => x"84",
          2915 => x"c8",
          2916 => x"9c",
          2917 => x"34",
          2918 => x"81",
          2919 => x"34",
          2920 => x"80",
          2921 => x"23",
          2922 => x"39",
          2923 => x"52",
          2924 => x"f9",
          2925 => x"05",
          2926 => x"f8",
          2927 => x"fb",
          2928 => x"eb",
          2929 => x"f9",
          2930 => x"2c",
          2931 => x"39",
          2932 => x"b7",
          2933 => x"eb",
          2934 => x"e3",
          2935 => x"70",
          2936 => x"40",
          2937 => x"33",
          2938 => x"11",
          2939 => x"c0",
          2940 => x"b7",
          2941 => x"5c",
          2942 => x"f8",
          2943 => x"81",
          2944 => x"74",
          2945 => x"83",
          2946 => x"29",
          2947 => x"f7",
          2948 => x"5d",
          2949 => x"83",
          2950 => x"80",
          2951 => x"bb",
          2952 => x"38",
          2953 => x"23",
          2954 => x"57",
          2955 => x"b7",
          2956 => x"ec",
          2957 => x"f8",
          2958 => x"f6",
          2959 => x"26",
          2960 => x"7e",
          2961 => x"5e",
          2962 => x"5b",
          2963 => x"06",
          2964 => x"1d",
          2965 => x"ec",
          2966 => x"e0",
          2967 => x"1e",
          2968 => x"76",
          2969 => x"81",
          2970 => x"bc",
          2971 => x"29",
          2972 => x"27",
          2973 => x"5e",
          2974 => x"81",
          2975 => x"58",
          2976 => x"81",
          2977 => x"bb",
          2978 => x"5d",
          2979 => x"eb",
          2980 => x"5c",
          2981 => x"83",
          2982 => x"83",
          2983 => x"5f",
          2984 => x"eb",
          2985 => x"81",
          2986 => x"76",
          2987 => x"83",
          2988 => x"ff",
          2989 => x"38",
          2990 => x"84",
          2991 => x"ff",
          2992 => x"eb",
          2993 => x"f9",
          2994 => x"33",
          2995 => x"11",
          2996 => x"ca",
          2997 => x"81",
          2998 => x"83",
          2999 => x"83",
          3000 => x"57",
          3001 => x"b8",
          3002 => x"75",
          3003 => x"ff",
          3004 => x"fc",
          3005 => x"83",
          3006 => x"7d",
          3007 => x"38",
          3008 => x"83",
          3009 => x"59",
          3010 => x"80",
          3011 => x"f8",
          3012 => x"34",
          3013 => x"39",
          3014 => x"f6",
          3015 => x"f8",
          3016 => x"f8",
          3017 => x"83",
          3018 => x"0b",
          3019 => x"83",
          3020 => x"c4",
          3021 => x"f7",
          3022 => x"0d",
          3023 => x"33",
          3024 => x"73",
          3025 => x"b9",
          3026 => x"52",
          3027 => x"84",
          3028 => x"f3",
          3029 => x"ff",
          3030 => x"ff",
          3031 => x"55",
          3032 => x"38",
          3033 => x"34",
          3034 => x"8f",
          3035 => x"54",
          3036 => x"73",
          3037 => x"09",
          3038 => x"72",
          3039 => x"54",
          3040 => x"38",
          3041 => x"70",
          3042 => x"79",
          3043 => x"bc",
          3044 => x"f8",
          3045 => x"a0",
          3046 => x"59",
          3047 => x"ff",
          3048 => x"59",
          3049 => x"38",
          3050 => x"80",
          3051 => x"0c",
          3052 => x"80",
          3053 => x"08",
          3054 => x"81",
          3055 => x"81",
          3056 => x"83",
          3057 => x"06",
          3058 => x"55",
          3059 => x"81",
          3060 => x"f6",
          3061 => x"5a",
          3062 => x"75",
          3063 => x"e8",
          3064 => x"81",
          3065 => x"89",
          3066 => x"f0",
          3067 => x"58",
          3068 => x"73",
          3069 => x"32",
          3070 => x"80",
          3071 => x"f7",
          3072 => x"72",
          3073 => x"83",
          3074 => x"a1",
          3075 => x"a2",
          3076 => x"f7",
          3077 => x"5e",
          3078 => x"74",
          3079 => x"90",
          3080 => x"82",
          3081 => x"72",
          3082 => x"90",
          3083 => x"74",
          3084 => x"2e",
          3085 => x"53",
          3086 => x"81",
          3087 => x"84",
          3088 => x"54",
          3089 => x"f7",
          3090 => x"98",
          3091 => x"83",
          3092 => x"9c",
          3093 => x"16",
          3094 => x"76",
          3095 => x"a3",
          3096 => x"9e",
          3097 => x"38",
          3098 => x"5a",
          3099 => x"54",
          3100 => x"14",
          3101 => x"7d",
          3102 => x"83",
          3103 => x"2e",
          3104 => x"ce",
          3105 => x"f7",
          3106 => x"77",
          3107 => x"17",
          3108 => x"76",
          3109 => x"83",
          3110 => x"82",
          3111 => x"38",
          3112 => x"fc",
          3113 => x"80",
          3114 => x"2e",
          3115 => x"06",
          3116 => x"ed",
          3117 => x"79",
          3118 => x"75",
          3119 => x"a1",
          3120 => x"17",
          3121 => x"fe",
          3122 => x"57",
          3123 => x"e1",
          3124 => x"05",
          3125 => x"f3",
          3126 => x"78",
          3127 => x"9c",
          3128 => x"7d",
          3129 => x"ff",
          3130 => x"ff",
          3131 => x"38",
          3132 => x"54",
          3133 => x"82",
          3134 => x"07",
          3135 => x"83",
          3136 => x"78",
          3137 => x"72",
          3138 => x"70",
          3139 => x"ba",
          3140 => x"54",
          3141 => x"b7",
          3142 => x"9a",
          3143 => x"f9",
          3144 => x"82",
          3145 => x"c8",
          3146 => x"34",
          3147 => x"81",
          3148 => x"14",
          3149 => x"90",
          3150 => x"83",
          3151 => x"f6",
          3152 => x"86",
          3153 => x"ff",
          3154 => x"96",
          3155 => x"81",
          3156 => x"ff",
          3157 => x"06",
          3158 => x"81",
          3159 => x"54",
          3160 => x"87",
          3161 => x"0c",
          3162 => x"39",
          3163 => x"f9",
          3164 => x"73",
          3165 => x"38",
          3166 => x"83",
          3167 => x"83",
          3168 => x"33",
          3169 => x"5e",
          3170 => x"82",
          3171 => x"7a",
          3172 => x"79",
          3173 => x"38",
          3174 => x"f0",
          3175 => x"b7",
          3176 => x"81",
          3177 => x"59",
          3178 => x"be",
          3179 => x"54",
          3180 => x"f7",
          3181 => x"08",
          3182 => x"83",
          3183 => x"b7",
          3184 => x"11",
          3185 => x"38",
          3186 => x"73",
          3187 => x"80",
          3188 => x"83",
          3189 => x"70",
          3190 => x"80",
          3191 => x"83",
          3192 => x"39",
          3193 => x"3f",
          3194 => x"fc",
          3195 => x"f7",
          3196 => x"0b",
          3197 => x"33",
          3198 => x"81",
          3199 => x"04",
          3200 => x"d4",
          3201 => x"82",
          3202 => x"80",
          3203 => x"d4",
          3204 => x"34",
          3205 => x"87",
          3206 => x"08",
          3207 => x"c0",
          3208 => x"9c",
          3209 => x"81",
          3210 => x"56",
          3211 => x"81",
          3212 => x"a4",
          3213 => x"80",
          3214 => x"80",
          3215 => x"80",
          3216 => x"9c",
          3217 => x"55",
          3218 => x"33",
          3219 => x"70",
          3220 => x"2e",
          3221 => x"55",
          3222 => x"71",
          3223 => x"57",
          3224 => x"81",
          3225 => x"74",
          3226 => x"c8",
          3227 => x"84",
          3228 => x"fa",
          3229 => x"05",
          3230 => x"d4",
          3231 => x"80",
          3232 => x"55",
          3233 => x"90",
          3234 => x"90",
          3235 => x"86",
          3236 => x"74",
          3237 => x"51",
          3238 => x"f3",
          3239 => x"15",
          3240 => x"34",
          3241 => x"d4",
          3242 => x"87",
          3243 => x"98",
          3244 => x"38",
          3245 => x"08",
          3246 => x"71",
          3247 => x"98",
          3248 => x"27",
          3249 => x"2e",
          3250 => x"08",
          3251 => x"98",
          3252 => x"08",
          3253 => x"14",
          3254 => x"52",
          3255 => x"ff",
          3256 => x"08",
          3257 => x"52",
          3258 => x"06",
          3259 => x"38",
          3260 => x"d4",
          3261 => x"56",
          3262 => x"84",
          3263 => x"27",
          3264 => x"33",
          3265 => x"71",
          3266 => x"0c",
          3267 => x"b9",
          3268 => x"51",
          3269 => x"84",
          3270 => x"0b",
          3271 => x"87",
          3272 => x"2a",
          3273 => x"15",
          3274 => x"15",
          3275 => x"15",
          3276 => x"f3",
          3277 => x"13",
          3278 => x"97",
          3279 => x"72",
          3280 => x"26",
          3281 => x"74",
          3282 => x"55",
          3283 => x"f3",
          3284 => x"15",
          3285 => x"34",
          3286 => x"d4",
          3287 => x"87",
          3288 => x"98",
          3289 => x"38",
          3290 => x"08",
          3291 => x"71",
          3292 => x"98",
          3293 => x"27",
          3294 => x"2e",
          3295 => x"08",
          3296 => x"98",
          3297 => x"08",
          3298 => x"14",
          3299 => x"52",
          3300 => x"ff",
          3301 => x"08",
          3302 => x"52",
          3303 => x"06",
          3304 => x"74",
          3305 => x"38",
          3306 => x"73",
          3307 => x"84",
          3308 => x"ff",
          3309 => x"f3",
          3310 => x"85",
          3311 => x"fe",
          3312 => x"f0",
          3313 => x"08",
          3314 => x"90",
          3315 => x"52",
          3316 => x"72",
          3317 => x"c0",
          3318 => x"27",
          3319 => x"38",
          3320 => x"53",
          3321 => x"53",
          3322 => x"c0",
          3323 => x"53",
          3324 => x"c0",
          3325 => x"f6",
          3326 => x"9c",
          3327 => x"38",
          3328 => x"c0",
          3329 => x"83",
          3330 => x"70",
          3331 => x"2e",
          3332 => x"73",
          3333 => x"0d",
          3334 => x"3f",
          3335 => x"84",
          3336 => x"2a",
          3337 => x"2b",
          3338 => x"71",
          3339 => x"11",
          3340 => x"2b",
          3341 => x"53",
          3342 => x"53",
          3343 => x"16",
          3344 => x"8b",
          3345 => x"70",
          3346 => x"71",
          3347 => x"59",
          3348 => x"38",
          3349 => x"8b",
          3350 => x"76",
          3351 => x"86",
          3352 => x"73",
          3353 => x"70",
          3354 => x"71",
          3355 => x"55",
          3356 => x"71",
          3357 => x"16",
          3358 => x"0b",
          3359 => x"53",
          3360 => x"34",
          3361 => x"81",
          3362 => x"80",
          3363 => x"52",
          3364 => x"34",
          3365 => x"87",
          3366 => x"2b",
          3367 => x"17",
          3368 => x"2a",
          3369 => x"71",
          3370 => x"84",
          3371 => x"33",
          3372 => x"83",
          3373 => x"05",
          3374 => x"88",
          3375 => x"59",
          3376 => x"13",
          3377 => x"33",
          3378 => x"81",
          3379 => x"5a",
          3380 => x"13",
          3381 => x"70",
          3382 => x"71",
          3383 => x"81",
          3384 => x"83",
          3385 => x"7b",
          3386 => x"5a",
          3387 => x"73",
          3388 => x"70",
          3389 => x"8b",
          3390 => x"70",
          3391 => x"07",
          3392 => x"5f",
          3393 => x"77",
          3394 => x"b9",
          3395 => x"83",
          3396 => x"2b",
          3397 => x"33",
          3398 => x"58",
          3399 => x"70",
          3400 => x"81",
          3401 => x"80",
          3402 => x"54",
          3403 => x"84",
          3404 => x"81",
          3405 => x"2b",
          3406 => x"15",
          3407 => x"2a",
          3408 => x"53",
          3409 => x"34",
          3410 => x"79",
          3411 => x"80",
          3412 => x"38",
          3413 => x"0d",
          3414 => x"b8",
          3415 => x"23",
          3416 => x"ff",
          3417 => x"b9",
          3418 => x"0b",
          3419 => x"54",
          3420 => x"15",
          3421 => x"86",
          3422 => x"84",
          3423 => x"ff",
          3424 => x"ff",
          3425 => x"55",
          3426 => x"17",
          3427 => x"10",
          3428 => x"05",
          3429 => x"0b",
          3430 => x"3d",
          3431 => x"84",
          3432 => x"2a",
          3433 => x"51",
          3434 => x"b9",
          3435 => x"33",
          3436 => x"5a",
          3437 => x"80",
          3438 => x"10",
          3439 => x"88",
          3440 => x"79",
          3441 => x"7a",
          3442 => x"72",
          3443 => x"85",
          3444 => x"33",
          3445 => x"57",
          3446 => x"ff",
          3447 => x"80",
          3448 => x"81",
          3449 => x"81",
          3450 => x"59",
          3451 => x"59",
          3452 => x"38",
          3453 => x"38",
          3454 => x"16",
          3455 => x"80",
          3456 => x"56",
          3457 => x"15",
          3458 => x"88",
          3459 => x"75",
          3460 => x"70",
          3461 => x"88",
          3462 => x"f8",
          3463 => x"06",
          3464 => x"59",
          3465 => x"81",
          3466 => x"84",
          3467 => x"34",
          3468 => x"08",
          3469 => x"33",
          3470 => x"74",
          3471 => x"84",
          3472 => x"b9",
          3473 => x"86",
          3474 => x"2b",
          3475 => x"59",
          3476 => x"34",
          3477 => x"11",
          3478 => x"71",
          3479 => x"5c",
          3480 => x"87",
          3481 => x"16",
          3482 => x"12",
          3483 => x"2a",
          3484 => x"34",
          3485 => x"08",
          3486 => x"c8",
          3487 => x"33",
          3488 => x"83",
          3489 => x"85",
          3490 => x"88",
          3491 => x"74",
          3492 => x"84",
          3493 => x"33",
          3494 => x"83",
          3495 => x"87",
          3496 => x"88",
          3497 => x"57",
          3498 => x"1a",
          3499 => x"33",
          3500 => x"81",
          3501 => x"57",
          3502 => x"18",
          3503 => x"05",
          3504 => x"79",
          3505 => x"80",
          3506 => x"38",
          3507 => x"0d",
          3508 => x"b9",
          3509 => x"3d",
          3510 => x"b9",
          3511 => x"b4",
          3512 => x"84",
          3513 => x"84",
          3514 => x"81",
          3515 => x"08",
          3516 => x"85",
          3517 => x"76",
          3518 => x"34",
          3519 => x"22",
          3520 => x"83",
          3521 => x"51",
          3522 => x"89",
          3523 => x"10",
          3524 => x"f8",
          3525 => x"81",
          3526 => x"80",
          3527 => x"ed",
          3528 => x"70",
          3529 => x"76",
          3530 => x"2e",
          3531 => x"d7",
          3532 => x"38",
          3533 => x"70",
          3534 => x"83",
          3535 => x"2a",
          3536 => x"2b",
          3537 => x"71",
          3538 => x"83",
          3539 => x"fc",
          3540 => x"33",
          3541 => x"70",
          3542 => x"45",
          3543 => x"48",
          3544 => x"24",
          3545 => x"16",
          3546 => x"10",
          3547 => x"71",
          3548 => x"5c",
          3549 => x"85",
          3550 => x"38",
          3551 => x"a2",
          3552 => x"60",
          3553 => x"38",
          3554 => x"f7",
          3555 => x"33",
          3556 => x"7a",
          3557 => x"98",
          3558 => x"59",
          3559 => x"24",
          3560 => x"33",
          3561 => x"83",
          3562 => x"87",
          3563 => x"2b",
          3564 => x"15",
          3565 => x"2a",
          3566 => x"53",
          3567 => x"79",
          3568 => x"70",
          3569 => x"71",
          3570 => x"05",
          3571 => x"88",
          3572 => x"5e",
          3573 => x"16",
          3574 => x"b8",
          3575 => x"71",
          3576 => x"70",
          3577 => x"79",
          3578 => x"b8",
          3579 => x"12",
          3580 => x"07",
          3581 => x"71",
          3582 => x"5c",
          3583 => x"79",
          3584 => x"b8",
          3585 => x"33",
          3586 => x"74",
          3587 => x"71",
          3588 => x"5c",
          3589 => x"82",
          3590 => x"b9",
          3591 => x"83",
          3592 => x"57",
          3593 => x"5a",
          3594 => x"c4",
          3595 => x"84",
          3596 => x"ff",
          3597 => x"26",
          3598 => x"b9",
          3599 => x"ff",
          3600 => x"80",
          3601 => x"80",
          3602 => x"fe",
          3603 => x"5e",
          3604 => x"34",
          3605 => x"1e",
          3606 => x"b9",
          3607 => x"81",
          3608 => x"08",
          3609 => x"80",
          3610 => x"70",
          3611 => x"88",
          3612 => x"b9",
          3613 => x"b9",
          3614 => x"60",
          3615 => x"34",
          3616 => x"d3",
          3617 => x"7e",
          3618 => x"7f",
          3619 => x"08",
          3620 => x"04",
          3621 => x"83",
          3622 => x"70",
          3623 => x"07",
          3624 => x"48",
          3625 => x"60",
          3626 => x"08",
          3627 => x"82",
          3628 => x"b9",
          3629 => x"12",
          3630 => x"2b",
          3631 => x"83",
          3632 => x"5c",
          3633 => x"82",
          3634 => x"60",
          3635 => x"08",
          3636 => x"1c",
          3637 => x"84",
          3638 => x"fd",
          3639 => x"ff",
          3640 => x"77",
          3641 => x"83",
          3642 => x"18",
          3643 => x"10",
          3644 => x"71",
          3645 => x"5e",
          3646 => x"80",
          3647 => x"61",
          3648 => x"24",
          3649 => x"06",
          3650 => x"fe",
          3651 => x"b9",
          3652 => x"b4",
          3653 => x"84",
          3654 => x"84",
          3655 => x"81",
          3656 => x"08",
          3657 => x"85",
          3658 => x"7e",
          3659 => x"34",
          3660 => x"22",
          3661 => x"83",
          3662 => x"56",
          3663 => x"73",
          3664 => x"22",
          3665 => x"08",
          3666 => x"82",
          3667 => x"fc",
          3668 => x"38",
          3669 => x"7b",
          3670 => x"76",
          3671 => x"ea",
          3672 => x"c8",
          3673 => x"82",
          3674 => x"2b",
          3675 => x"11",
          3676 => x"71",
          3677 => x"33",
          3678 => x"70",
          3679 => x"46",
          3680 => x"84",
          3681 => x"84",
          3682 => x"33",
          3683 => x"83",
          3684 => x"87",
          3685 => x"88",
          3686 => x"5d",
          3687 => x"64",
          3688 => x"16",
          3689 => x"2b",
          3690 => x"2a",
          3691 => x"79",
          3692 => x"70",
          3693 => x"71",
          3694 => x"05",
          3695 => x"2b",
          3696 => x"40",
          3697 => x"75",
          3698 => x"70",
          3699 => x"8b",
          3700 => x"82",
          3701 => x"2b",
          3702 => x"5b",
          3703 => x"34",
          3704 => x"08",
          3705 => x"33",
          3706 => x"56",
          3707 => x"7e",
          3708 => x"3f",
          3709 => x"78",
          3710 => x"99",
          3711 => x"b8",
          3712 => x"23",
          3713 => x"ff",
          3714 => x"b9",
          3715 => x"0b",
          3716 => x"55",
          3717 => x"16",
          3718 => x"86",
          3719 => x"84",
          3720 => x"ff",
          3721 => x"ff",
          3722 => x"44",
          3723 => x"1f",
          3724 => x"10",
          3725 => x"05",
          3726 => x"0b",
          3727 => x"3f",
          3728 => x"33",
          3729 => x"83",
          3730 => x"85",
          3731 => x"88",
          3732 => x"76",
          3733 => x"05",
          3734 => x"84",
          3735 => x"2b",
          3736 => x"14",
          3737 => x"07",
          3738 => x"59",
          3739 => x"34",
          3740 => x"b8",
          3741 => x"71",
          3742 => x"70",
          3743 => x"78",
          3744 => x"b8",
          3745 => x"33",
          3746 => x"74",
          3747 => x"88",
          3748 => x"f8",
          3749 => x"5d",
          3750 => x"7f",
          3751 => x"84",
          3752 => x"81",
          3753 => x"2b",
          3754 => x"33",
          3755 => x"06",
          3756 => x"46",
          3757 => x"60",
          3758 => x"06",
          3759 => x"87",
          3760 => x"2b",
          3761 => x"19",
          3762 => x"2a",
          3763 => x"84",
          3764 => x"b9",
          3765 => x"85",
          3766 => x"2b",
          3767 => x"15",
          3768 => x"2a",
          3769 => x"56",
          3770 => x"87",
          3771 => x"70",
          3772 => x"07",
          3773 => x"5b",
          3774 => x"81",
          3775 => x"1f",
          3776 => x"2b",
          3777 => x"33",
          3778 => x"70",
          3779 => x"05",
          3780 => x"58",
          3781 => x"34",
          3782 => x"08",
          3783 => x"71",
          3784 => x"05",
          3785 => x"2b",
          3786 => x"2a",
          3787 => x"55",
          3788 => x"84",
          3789 => x"33",
          3790 => x"83",
          3791 => x"87",
          3792 => x"2b",
          3793 => x"15",
          3794 => x"2a",
          3795 => x"53",
          3796 => x"34",
          3797 => x"08",
          3798 => x"33",
          3799 => x"74",
          3800 => x"71",
          3801 => x"42",
          3802 => x"86",
          3803 => x"b9",
          3804 => x"33",
          3805 => x"06",
          3806 => x"76",
          3807 => x"b9",
          3808 => x"83",
          3809 => x"2b",
          3810 => x"33",
          3811 => x"41",
          3812 => x"79",
          3813 => x"b9",
          3814 => x"12",
          3815 => x"07",
          3816 => x"33",
          3817 => x"41",
          3818 => x"79",
          3819 => x"84",
          3820 => x"33",
          3821 => x"66",
          3822 => x"52",
          3823 => x"fe",
          3824 => x"1e",
          3825 => x"83",
          3826 => x"d5",
          3827 => x"71",
          3828 => x"05",
          3829 => x"88",
          3830 => x"5d",
          3831 => x"34",
          3832 => x"b8",
          3833 => x"12",
          3834 => x"07",
          3835 => x"33",
          3836 => x"5b",
          3837 => x"73",
          3838 => x"05",
          3839 => x"33",
          3840 => x"81",
          3841 => x"5f",
          3842 => x"16",
          3843 => x"70",
          3844 => x"71",
          3845 => x"81",
          3846 => x"83",
          3847 => x"63",
          3848 => x"5e",
          3849 => x"7b",
          3850 => x"70",
          3851 => x"8b",
          3852 => x"70",
          3853 => x"07",
          3854 => x"47",
          3855 => x"7f",
          3856 => x"83",
          3857 => x"7e",
          3858 => x"b9",
          3859 => x"80",
          3860 => x"84",
          3861 => x"3f",
          3862 => x"61",
          3863 => x"39",
          3864 => x"b9",
          3865 => x"b7",
          3866 => x"84",
          3867 => x"77",
          3868 => x"08",
          3869 => x"e6",
          3870 => x"c8",
          3871 => x"84",
          3872 => x"84",
          3873 => x"a0",
          3874 => x"80",
          3875 => x"51",
          3876 => x"08",
          3877 => x"16",
          3878 => x"84",
          3879 => x"84",
          3880 => x"34",
          3881 => x"b8",
          3882 => x"fe",
          3883 => x"06",
          3884 => x"74",
          3885 => x"84",
          3886 => x"84",
          3887 => x"55",
          3888 => x"15",
          3889 => x"c6",
          3890 => x"02",
          3891 => x"72",
          3892 => x"33",
          3893 => x"3d",
          3894 => x"05",
          3895 => x"9d",
          3896 => x"b9",
          3897 => x"87",
          3898 => x"84",
          3899 => x"b9",
          3900 => x"3d",
          3901 => x"af",
          3902 => x"54",
          3903 => x"c4",
          3904 => x"83",
          3905 => x"0b",
          3906 => x"75",
          3907 => x"b9",
          3908 => x"80",
          3909 => x"08",
          3910 => x"d6",
          3911 => x"73",
          3912 => x"55",
          3913 => x"0d",
          3914 => x"81",
          3915 => x"26",
          3916 => x"0d",
          3917 => x"05",
          3918 => x"76",
          3919 => x"17",
          3920 => x"55",
          3921 => x"87",
          3922 => x"52",
          3923 => x"c8",
          3924 => x"2e",
          3925 => x"54",
          3926 => x"38",
          3927 => x"80",
          3928 => x"74",
          3929 => x"04",
          3930 => x"ff",
          3931 => x"ff",
          3932 => x"78",
          3933 => x"88",
          3934 => x"81",
          3935 => x"b9",
          3936 => x"54",
          3937 => x"87",
          3938 => x"73",
          3939 => x"38",
          3940 => x"72",
          3941 => x"04",
          3942 => x"b9",
          3943 => x"80",
          3944 => x"0c",
          3945 => x"87",
          3946 => x"cd",
          3947 => x"06",
          3948 => x"87",
          3949 => x"38",
          3950 => x"ca",
          3951 => x"8c",
          3952 => x"73",
          3953 => x"82",
          3954 => x"39",
          3955 => x"83",
          3956 => x"77",
          3957 => x"33",
          3958 => x"80",
          3959 => x"fe",
          3960 => x"2e",
          3961 => x"c8",
          3962 => x"b4",
          3963 => x"81",
          3964 => x"81",
          3965 => x"09",
          3966 => x"08",
          3967 => x"a8",
          3968 => x"b9",
          3969 => x"76",
          3970 => x"55",
          3971 => x"8e",
          3972 => x"52",
          3973 => x"76",
          3974 => x"09",
          3975 => x"33",
          3976 => x"fe",
          3977 => x"7a",
          3978 => x"57",
          3979 => x"80",
          3980 => x"aa",
          3981 => x"7a",
          3982 => x"80",
          3983 => x"0b",
          3984 => x"9c",
          3985 => x"19",
          3986 => x"34",
          3987 => x"94",
          3988 => x"34",
          3989 => x"19",
          3990 => x"a2",
          3991 => x"84",
          3992 => x"7a",
          3993 => x"55",
          3994 => x"2a",
          3995 => x"98",
          3996 => x"a4",
          3997 => x"0c",
          3998 => x"81",
          3999 => x"84",
          4000 => x"18",
          4001 => x"c8",
          4002 => x"b2",
          4003 => x"08",
          4004 => x"38",
          4005 => x"81",
          4006 => x"3d",
          4007 => x"74",
          4008 => x"24",
          4009 => x"81",
          4010 => x"70",
          4011 => x"5a",
          4012 => x"b0",
          4013 => x"2e",
          4014 => x"54",
          4015 => x"33",
          4016 => x"08",
          4017 => x"5b",
          4018 => x"38",
          4019 => x"33",
          4020 => x"08",
          4021 => x"08",
          4022 => x"18",
          4023 => x"2e",
          4024 => x"54",
          4025 => x"33",
          4026 => x"08",
          4027 => x"5a",
          4028 => x"38",
          4029 => x"33",
          4030 => x"06",
          4031 => x"5d",
          4032 => x"06",
          4033 => x"04",
          4034 => x"59",
          4035 => x"80",
          4036 => x"5b",
          4037 => x"c2",
          4038 => x"52",
          4039 => x"84",
          4040 => x"ff",
          4041 => x"79",
          4042 => x"06",
          4043 => x"71",
          4044 => x"c8",
          4045 => x"74",
          4046 => x"38",
          4047 => x"59",
          4048 => x"80",
          4049 => x"5b",
          4050 => x"81",
          4051 => x"52",
          4052 => x"84",
          4053 => x"ff",
          4054 => x"79",
          4055 => x"fc",
          4056 => x"33",
          4057 => x"88",
          4058 => x"07",
          4059 => x"ff",
          4060 => x"0c",
          4061 => x"3d",
          4062 => x"53",
          4063 => x"52",
          4064 => x"b9",
          4065 => x"fe",
          4066 => x"18",
          4067 => x"31",
          4068 => x"a0",
          4069 => x"17",
          4070 => x"06",
          4071 => x"08",
          4072 => x"81",
          4073 => x"5a",
          4074 => x"08",
          4075 => x"33",
          4076 => x"c8",
          4077 => x"81",
          4078 => x"34",
          4079 => x"5d",
          4080 => x"82",
          4081 => x"cb",
          4082 => x"de",
          4083 => x"b8",
          4084 => x"5c",
          4085 => x"c8",
          4086 => x"ff",
          4087 => x"34",
          4088 => x"84",
          4089 => x"18",
          4090 => x"33",
          4091 => x"fd",
          4092 => x"a0",
          4093 => x"17",
          4094 => x"fd",
          4095 => x"53",
          4096 => x"52",
          4097 => x"b9",
          4098 => x"fb",
          4099 => x"18",
          4100 => x"31",
          4101 => x"a0",
          4102 => x"17",
          4103 => x"06",
          4104 => x"08",
          4105 => x"81",
          4106 => x"5a",
          4107 => x"08",
          4108 => x"81",
          4109 => x"86",
          4110 => x"fa",
          4111 => x"64",
          4112 => x"27",
          4113 => x"95",
          4114 => x"96",
          4115 => x"74",
          4116 => x"b9",
          4117 => x"88",
          4118 => x"0b",
          4119 => x"2e",
          4120 => x"5b",
          4121 => x"83",
          4122 => x"19",
          4123 => x"3f",
          4124 => x"38",
          4125 => x"0c",
          4126 => x"10",
          4127 => x"ff",
          4128 => x"34",
          4129 => x"34",
          4130 => x"b9",
          4131 => x"83",
          4132 => x"75",
          4133 => x"80",
          4134 => x"78",
          4135 => x"7c",
          4136 => x"06",
          4137 => x"b8",
          4138 => x"8e",
          4139 => x"85",
          4140 => x"1a",
          4141 => x"75",
          4142 => x"b8",
          4143 => x"8f",
          4144 => x"41",
          4145 => x"88",
          4146 => x"90",
          4147 => x"98",
          4148 => x"0b",
          4149 => x"81",
          4150 => x"08",
          4151 => x"76",
          4152 => x"1a",
          4153 => x"2e",
          4154 => x"54",
          4155 => x"33",
          4156 => x"08",
          4157 => x"5c",
          4158 => x"fd",
          4159 => x"b8",
          4160 => x"5f",
          4161 => x"38",
          4162 => x"33",
          4163 => x"77",
          4164 => x"89",
          4165 => x"0b",
          4166 => x"2e",
          4167 => x"b8",
          4168 => x"57",
          4169 => x"c8",
          4170 => x"c7",
          4171 => x"34",
          4172 => x"31",
          4173 => x"5b",
          4174 => x"38",
          4175 => x"82",
          4176 => x"52",
          4177 => x"84",
          4178 => x"ff",
          4179 => x"77",
          4180 => x"19",
          4181 => x"7c",
          4182 => x"81",
          4183 => x"5c",
          4184 => x"34",
          4185 => x"b8",
          4186 => x"5d",
          4187 => x"c8",
          4188 => x"88",
          4189 => x"34",
          4190 => x"31",
          4191 => x"5d",
          4192 => x"ca",
          4193 => x"2e",
          4194 => x"54",
          4195 => x"33",
          4196 => x"aa",
          4197 => x"70",
          4198 => x"ad",
          4199 => x"7d",
          4200 => x"84",
          4201 => x"19",
          4202 => x"1b",
          4203 => x"56",
          4204 => x"82",
          4205 => x"81",
          4206 => x"1f",
          4207 => x"ed",
          4208 => x"81",
          4209 => x"81",
          4210 => x"81",
          4211 => x"09",
          4212 => x"c8",
          4213 => x"70",
          4214 => x"84",
          4215 => x"7e",
          4216 => x"33",
          4217 => x"fa",
          4218 => x"76",
          4219 => x"3f",
          4220 => x"79",
          4221 => x"51",
          4222 => x"39",
          4223 => x"05",
          4224 => x"58",
          4225 => x"5a",
          4226 => x"7e",
          4227 => x"2b",
          4228 => x"83",
          4229 => x"06",
          4230 => x"5f",
          4231 => x"2a",
          4232 => x"2a",
          4233 => x"2a",
          4234 => x"39",
          4235 => x"5b",
          4236 => x"19",
          4237 => x"38",
          4238 => x"38",
          4239 => x"80",
          4240 => x"81",
          4241 => x"9c",
          4242 => x"56",
          4243 => x"52",
          4244 => x"c8",
          4245 => x"58",
          4246 => x"38",
          4247 => x"70",
          4248 => x"51",
          4249 => x"75",
          4250 => x"38",
          4251 => x"8c",
          4252 => x"39",
          4253 => x"7a",
          4254 => x"55",
          4255 => x"38",
          4256 => x"c8",
          4257 => x"08",
          4258 => x"7a",
          4259 => x"9c",
          4260 => x"56",
          4261 => x"80",
          4262 => x"81",
          4263 => x"70",
          4264 => x"7b",
          4265 => x"51",
          4266 => x"b9",
          4267 => x"19",
          4268 => x"38",
          4269 => x"38",
          4270 => x"75",
          4271 => x"75",
          4272 => x"b9",
          4273 => x"70",
          4274 => x"56",
          4275 => x"80",
          4276 => x"19",
          4277 => x"58",
          4278 => x"94",
          4279 => x"5a",
          4280 => x"84",
          4281 => x"80",
          4282 => x"0d",
          4283 => x"da",
          4284 => x"75",
          4285 => x"3f",
          4286 => x"39",
          4287 => x"0c",
          4288 => x"81",
          4289 => x"b6",
          4290 => x"08",
          4291 => x"26",
          4292 => x"72",
          4293 => x"88",
          4294 => x"76",
          4295 => x"38",
          4296 => x"18",
          4297 => x"38",
          4298 => x"94",
          4299 => x"56",
          4300 => x"2a",
          4301 => x"06",
          4302 => x"56",
          4303 => x"0d",
          4304 => x"8a",
          4305 => x"74",
          4306 => x"22",
          4307 => x"27",
          4308 => x"15",
          4309 => x"73",
          4310 => x"71",
          4311 => x"78",
          4312 => x"52",
          4313 => x"c8",
          4314 => x"2e",
          4315 => x"08",
          4316 => x"53",
          4317 => x"91",
          4318 => x"27",
          4319 => x"84",
          4320 => x"f3",
          4321 => x"08",
          4322 => x"0a",
          4323 => x"18",
          4324 => x"74",
          4325 => x"06",
          4326 => x"18",
          4327 => x"85",
          4328 => x"76",
          4329 => x"0c",
          4330 => x"05",
          4331 => x"b9",
          4332 => x"98",
          4333 => x"7a",
          4334 => x"75",
          4335 => x"b9",
          4336 => x"84",
          4337 => x"56",
          4338 => x"38",
          4339 => x"26",
          4340 => x"98",
          4341 => x"f9",
          4342 => x"87",
          4343 => x"ff",
          4344 => x"08",
          4345 => x"84",
          4346 => x"38",
          4347 => x"5f",
          4348 => x"9c",
          4349 => x"5c",
          4350 => x"22",
          4351 => x"5d",
          4352 => x"58",
          4353 => x"70",
          4354 => x"74",
          4355 => x"55",
          4356 => x"54",
          4357 => x"33",
          4358 => x"08",
          4359 => x"39",
          4360 => x"b9",
          4361 => x"54",
          4362 => x"53",
          4363 => x"3f",
          4364 => x"84",
          4365 => x"19",
          4366 => x"a0",
          4367 => x"19",
          4368 => x"06",
          4369 => x"08",
          4370 => x"81",
          4371 => x"c5",
          4372 => x"ff",
          4373 => x"81",
          4374 => x"fe",
          4375 => x"56",
          4376 => x"38",
          4377 => x"1b",
          4378 => x"f8",
          4379 => x"8f",
          4380 => x"66",
          4381 => x"81",
          4382 => x"5e",
          4383 => x"19",
          4384 => x"08",
          4385 => x"33",
          4386 => x"81",
          4387 => x"53",
          4388 => x"e1",
          4389 => x"2e",
          4390 => x"b4",
          4391 => x"38",
          4392 => x"76",
          4393 => x"33",
          4394 => x"41",
          4395 => x"32",
          4396 => x"72",
          4397 => x"45",
          4398 => x"7a",
          4399 => x"81",
          4400 => x"38",
          4401 => x"fa",
          4402 => x"84",
          4403 => x"1c",
          4404 => x"84",
          4405 => x"81",
          4406 => x"81",
          4407 => x"57",
          4408 => x"81",
          4409 => x"08",
          4410 => x"1a",
          4411 => x"5b",
          4412 => x"38",
          4413 => x"09",
          4414 => x"b4",
          4415 => x"7e",
          4416 => x"3f",
          4417 => x"2e",
          4418 => x"86",
          4419 => x"93",
          4420 => x"06",
          4421 => x"0c",
          4422 => x"38",
          4423 => x"39",
          4424 => x"06",
          4425 => x"80",
          4426 => x"c8",
          4427 => x"fd",
          4428 => x"77",
          4429 => x"19",
          4430 => x"71",
          4431 => x"ff",
          4432 => x"06",
          4433 => x"76",
          4434 => x"78",
          4435 => x"88",
          4436 => x"2e",
          4437 => x"ff",
          4438 => x"5c",
          4439 => x"81",
          4440 => x"77",
          4441 => x"57",
          4442 => x"fe",
          4443 => x"05",
          4444 => x"81",
          4445 => x"75",
          4446 => x"ff",
          4447 => x"7c",
          4448 => x"81",
          4449 => x"5a",
          4450 => x"06",
          4451 => x"38",
          4452 => x"0b",
          4453 => x"0c",
          4454 => x"63",
          4455 => x"51",
          4456 => x"5a",
          4457 => x"81",
          4458 => x"1d",
          4459 => x"56",
          4460 => x"82",
          4461 => x"55",
          4462 => x"df",
          4463 => x"52",
          4464 => x"84",
          4465 => x"ff",
          4466 => x"76",
          4467 => x"08",
          4468 => x"84",
          4469 => x"70",
          4470 => x"1d",
          4471 => x"38",
          4472 => x"8f",
          4473 => x"38",
          4474 => x"aa",
          4475 => x"74",
          4476 => x"78",
          4477 => x"05",
          4478 => x"56",
          4479 => x"80",
          4480 => x"57",
          4481 => x"59",
          4482 => x"78",
          4483 => x"31",
          4484 => x"80",
          4485 => x"e1",
          4486 => x"1d",
          4487 => x"3f",
          4488 => x"c8",
          4489 => x"84",
          4490 => x"81",
          4491 => x"81",
          4492 => x"57",
          4493 => x"81",
          4494 => x"08",
          4495 => x"1c",
          4496 => x"59",
          4497 => x"38",
          4498 => x"09",
          4499 => x"b4",
          4500 => x"7d",
          4501 => x"3f",
          4502 => x"fd",
          4503 => x"2a",
          4504 => x"38",
          4505 => x"80",
          4506 => x"81",
          4507 => x"ac",
          4508 => x"2e",
          4509 => x"80",
          4510 => x"b9",
          4511 => x"80",
          4512 => x"75",
          4513 => x"5d",
          4514 => x"39",
          4515 => x"09",
          4516 => x"9b",
          4517 => x"2b",
          4518 => x"38",
          4519 => x"f3",
          4520 => x"83",
          4521 => x"11",
          4522 => x"52",
          4523 => x"38",
          4524 => x"76",
          4525 => x"c8",
          4526 => x"53",
          4527 => x"f6",
          4528 => x"09",
          4529 => x"81",
          4530 => x"38",
          4531 => x"56",
          4532 => x"80",
          4533 => x"70",
          4534 => x"ff",
          4535 => x"fe",
          4536 => x"0c",
          4537 => x"ff",
          4538 => x"fe",
          4539 => x"08",
          4540 => x"58",
          4541 => x"b5",
          4542 => x"57",
          4543 => x"81",
          4544 => x"56",
          4545 => x"1f",
          4546 => x"55",
          4547 => x"70",
          4548 => x"74",
          4549 => x"70",
          4550 => x"82",
          4551 => x"34",
          4552 => x"1c",
          4553 => x"5a",
          4554 => x"33",
          4555 => x"15",
          4556 => x"80",
          4557 => x"74",
          4558 => x"5a",
          4559 => x"10",
          4560 => x"ff",
          4561 => x"58",
          4562 => x"76",
          4563 => x"58",
          4564 => x"55",
          4565 => x"80",
          4566 => x"bf",
          4567 => x"87",
          4568 => x"ff",
          4569 => x"76",
          4570 => x"79",
          4571 => x"27",
          4572 => x"2e",
          4573 => x"27",
          4574 => x"56",
          4575 => x"ea",
          4576 => x"87",
          4577 => x"ec",
          4578 => x"41",
          4579 => x"f4",
          4580 => x"b9",
          4581 => x"80",
          4582 => x"56",
          4583 => x"84",
          4584 => x"08",
          4585 => x"38",
          4586 => x"34",
          4587 => x"05",
          4588 => x"06",
          4589 => x"38",
          4590 => x"b0",
          4591 => x"80",
          4592 => x"b9",
          4593 => x"81",
          4594 => x"19",
          4595 => x"57",
          4596 => x"38",
          4597 => x"09",
          4598 => x"75",
          4599 => x"51",
          4600 => x"80",
          4601 => x"75",
          4602 => x"38",
          4603 => x"74",
          4604 => x"30",
          4605 => x"74",
          4606 => x"59",
          4607 => x"52",
          4608 => x"c8",
          4609 => x"2e",
          4610 => x"2e",
          4611 => x"83",
          4612 => x"38",
          4613 => x"77",
          4614 => x"57",
          4615 => x"76",
          4616 => x"51",
          4617 => x"80",
          4618 => x"76",
          4619 => x"c3",
          4620 => x"55",
          4621 => x"ff",
          4622 => x"9c",
          4623 => x"70",
          4624 => x"05",
          4625 => x"38",
          4626 => x"06",
          4627 => x"0b",
          4628 => x"b9",
          4629 => x"75",
          4630 => x"40",
          4631 => x"81",
          4632 => x"b9",
          4633 => x"80",
          4634 => x"81",
          4635 => x"81",
          4636 => x"b9",
          4637 => x"83",
          4638 => x"19",
          4639 => x"31",
          4640 => x"38",
          4641 => x"84",
          4642 => x"fd",
          4643 => x"08",
          4644 => x"e9",
          4645 => x"b9",
          4646 => x"b9",
          4647 => x"81",
          4648 => x"70",
          4649 => x"70",
          4650 => x"5d",
          4651 => x"b8",
          4652 => x"80",
          4653 => x"38",
          4654 => x"09",
          4655 => x"76",
          4656 => x"51",
          4657 => x"80",
          4658 => x"76",
          4659 => x"83",
          4660 => x"61",
          4661 => x"8d",
          4662 => x"75",
          4663 => x"75",
          4664 => x"05",
          4665 => x"ff",
          4666 => x"70",
          4667 => x"e5",
          4668 => x"75",
          4669 => x"2a",
          4670 => x"83",
          4671 => x"78",
          4672 => x"2e",
          4673 => x"22",
          4674 => x"38",
          4675 => x"34",
          4676 => x"84",
          4677 => x"08",
          4678 => x"7f",
          4679 => x"54",
          4680 => x"53",
          4681 => x"3f",
          4682 => x"83",
          4683 => x"34",
          4684 => x"84",
          4685 => x"1d",
          4686 => x"33",
          4687 => x"fb",
          4688 => x"a0",
          4689 => x"1c",
          4690 => x"fb",
          4691 => x"33",
          4692 => x"09",
          4693 => x"39",
          4694 => x"fa",
          4695 => x"c0",
          4696 => x"b4",
          4697 => x"33",
          4698 => x"08",
          4699 => x"84",
          4700 => x"1c",
          4701 => x"a0",
          4702 => x"33",
          4703 => x"b9",
          4704 => x"ff",
          4705 => x"98",
          4706 => x"f7",
          4707 => x"80",
          4708 => x"81",
          4709 => x"05",
          4710 => x"ce",
          4711 => x"b4",
          4712 => x"7c",
          4713 => x"3f",
          4714 => x"61",
          4715 => x"96",
          4716 => x"82",
          4717 => x"80",
          4718 => x"05",
          4719 => x"58",
          4720 => x"74",
          4721 => x"56",
          4722 => x"14",
          4723 => x"76",
          4724 => x"79",
          4725 => x"55",
          4726 => x"80",
          4727 => x"5e",
          4728 => x"82",
          4729 => x"57",
          4730 => x"81",
          4731 => x"b2",
          4732 => x"75",
          4733 => x"80",
          4734 => x"90",
          4735 => x"77",
          4736 => x"58",
          4737 => x"81",
          4738 => x"38",
          4739 => x"81",
          4740 => x"a5",
          4741 => x"96",
          4742 => x"05",
          4743 => x"1c",
          4744 => x"89",
          4745 => x"08",
          4746 => x"9c",
          4747 => x"82",
          4748 => x"2b",
          4749 => x"88",
          4750 => x"59",
          4751 => x"88",
          4752 => x"56",
          4753 => x"15",
          4754 => x"07",
          4755 => x"3d",
          4756 => x"39",
          4757 => x"31",
          4758 => x"90",
          4759 => x"3f",
          4760 => x"06",
          4761 => x"81",
          4762 => x"2a",
          4763 => x"34",
          4764 => x"1f",
          4765 => x"70",
          4766 => x"38",
          4767 => x"70",
          4768 => x"07",
          4769 => x"74",
          4770 => x"0b",
          4771 => x"72",
          4772 => x"77",
          4773 => x"1e",
          4774 => x"ff",
          4775 => x"a4",
          4776 => x"54",
          4777 => x"84",
          4778 => x"80",
          4779 => x"ff",
          4780 => x"81",
          4781 => x"81",
          4782 => x"59",
          4783 => x"b4",
          4784 => x"80",
          4785 => x"73",
          4786 => x"39",
          4787 => x"42",
          4788 => x"55",
          4789 => x"53",
          4790 => x"72",
          4791 => x"08",
          4792 => x"94",
          4793 => x"82",
          4794 => x"58",
          4795 => x"52",
          4796 => x"72",
          4797 => x"38",
          4798 => x"76",
          4799 => x"17",
          4800 => x"af",
          4801 => x"80",
          4802 => x"82",
          4803 => x"89",
          4804 => x"83",
          4805 => x"70",
          4806 => x"80",
          4807 => x"8f",
          4808 => x"ff",
          4809 => x"72",
          4810 => x"38",
          4811 => x"76",
          4812 => x"17",
          4813 => x"56",
          4814 => x"38",
          4815 => x"32",
          4816 => x"51",
          4817 => x"38",
          4818 => x"33",
          4819 => x"72",
          4820 => x"25",
          4821 => x"38",
          4822 => x"3d",
          4823 => x"26",
          4824 => x"52",
          4825 => x"b9",
          4826 => x"73",
          4827 => x"b9",
          4828 => x"e4",
          4829 => x"53",
          4830 => x"39",
          4831 => x"52",
          4832 => x"c8",
          4833 => x"0d",
          4834 => x"30",
          4835 => x"5a",
          4836 => x"14",
          4837 => x"56",
          4838 => x"dc",
          4839 => x"07",
          4840 => x"61",
          4841 => x"76",
          4842 => x"2e",
          4843 => x"80",
          4844 => x"fe",
          4845 => x"30",
          4846 => x"56",
          4847 => x"89",
          4848 => x"76",
          4849 => x"76",
          4850 => x"22",
          4851 => x"5d",
          4852 => x"38",
          4853 => x"ae",
          4854 => x"aa",
          4855 => x"5a",
          4856 => x"10",
          4857 => x"76",
          4858 => x"22",
          4859 => x"06",
          4860 => x"53",
          4861 => x"ff",
          4862 => x"5c",
          4863 => x"19",
          4864 => x"80",
          4865 => x"38",
          4866 => x"25",
          4867 => x"ce",
          4868 => x"7c",
          4869 => x"77",
          4870 => x"25",
          4871 => x"72",
          4872 => x"2e",
          4873 => x"38",
          4874 => x"9e",
          4875 => x"82",
          4876 => x"5f",
          4877 => x"58",
          4878 => x"1c",
          4879 => x"84",
          4880 => x"7d",
          4881 => x"ed",
          4882 => x"2e",
          4883 => x"06",
          4884 => x"5d",
          4885 => x"07",
          4886 => x"7d",
          4887 => x"5a",
          4888 => x"ec",
          4889 => x"33",
          4890 => x"2e",
          4891 => x"84",
          4892 => x"74",
          4893 => x"2e",
          4894 => x"06",
          4895 => x"65",
          4896 => x"58",
          4897 => x"70",
          4898 => x"56",
          4899 => x"80",
          4900 => x"5a",
          4901 => x"75",
          4902 => x"38",
          4903 => x"81",
          4904 => x"5b",
          4905 => x"56",
          4906 => x"38",
          4907 => x"57",
          4908 => x"e9",
          4909 => x"1d",
          4910 => x"b9",
          4911 => x"84",
          4912 => x"82",
          4913 => x"38",
          4914 => x"06",
          4915 => x"38",
          4916 => x"05",
          4917 => x"33",
          4918 => x"57",
          4919 => x"38",
          4920 => x"55",
          4921 => x"74",
          4922 => x"59",
          4923 => x"79",
          4924 => x"81",
          4925 => x"70",
          4926 => x"09",
          4927 => x"07",
          4928 => x"1d",
          4929 => x"fc",
          4930 => x"ab",
          4931 => x"0c",
          4932 => x"26",
          4933 => x"c9",
          4934 => x"81",
          4935 => x"18",
          4936 => x"82",
          4937 => x"81",
          4938 => x"83",
          4939 => x"06",
          4940 => x"74",
          4941 => x"33",
          4942 => x"b9",
          4943 => x"83",
          4944 => x"70",
          4945 => x"80",
          4946 => x"8f",
          4947 => x"ff",
          4948 => x"72",
          4949 => x"38",
          4950 => x"8a",
          4951 => x"06",
          4952 => x"99",
          4953 => x"81",
          4954 => x"ff",
          4955 => x"a0",
          4956 => x"5b",
          4957 => x"53",
          4958 => x"70",
          4959 => x"2e",
          4960 => x"07",
          4961 => x"74",
          4962 => x"80",
          4963 => x"71",
          4964 => x"07",
          4965 => x"39",
          4966 => x"54",
          4967 => x"11",
          4968 => x"81",
          4969 => x"07",
          4970 => x"e5",
          4971 => x"fd",
          4972 => x"5c",
          4973 => x"b9",
          4974 => x"3d",
          4975 => x"e7",
          4976 => x"0c",
          4977 => x"79",
          4978 => x"81",
          4979 => x"56",
          4980 => x"ed",
          4981 => x"84",
          4982 => x"85",
          4983 => x"90",
          4984 => x"76",
          4985 => x"0c",
          4986 => x"59",
          4987 => x"33",
          4988 => x"c8",
          4989 => x"5e",
          4990 => x"80",
          4991 => x"bc",
          4992 => x"81",
          4993 => x"84",
          4994 => x"81",
          4995 => x"c2",
          4996 => x"82",
          4997 => x"84",
          4998 => x"34",
          4999 => x"5a",
          5000 => x"70",
          5001 => x"bb",
          5002 => x"2e",
          5003 => x"b4",
          5004 => x"84",
          5005 => x"71",
          5006 => x"74",
          5007 => x"75",
          5008 => x"1d",
          5009 => x"58",
          5010 => x"58",
          5011 => x"c4",
          5012 => x"88",
          5013 => x"2e",
          5014 => x"cf",
          5015 => x"88",
          5016 => x"80",
          5017 => x"33",
          5018 => x"81",
          5019 => x"75",
          5020 => x"5e",
          5021 => x"c8",
          5022 => x"17",
          5023 => x"5f",
          5024 => x"82",
          5025 => x"71",
          5026 => x"5a",
          5027 => x"80",
          5028 => x"06",
          5029 => x"17",
          5030 => x"2b",
          5031 => x"74",
          5032 => x"7c",
          5033 => x"80",
          5034 => x"56",
          5035 => x"83",
          5036 => x"2b",
          5037 => x"70",
          5038 => x"07",
          5039 => x"80",
          5040 => x"71",
          5041 => x"7b",
          5042 => x"7a",
          5043 => x"81",
          5044 => x"51",
          5045 => x"08",
          5046 => x"81",
          5047 => x"ff",
          5048 => x"5d",
          5049 => x"82",
          5050 => x"38",
          5051 => x"0c",
          5052 => x"a8",
          5053 => x"57",
          5054 => x"88",
          5055 => x"2e",
          5056 => x"0c",
          5057 => x"38",
          5058 => x"81",
          5059 => x"89",
          5060 => x"08",
          5061 => x"0c",
          5062 => x"0b",
          5063 => x"96",
          5064 => x"22",
          5065 => x"23",
          5066 => x"0b",
          5067 => x"0c",
          5068 => x"97",
          5069 => x"c8",
          5070 => x"d0",
          5071 => x"58",
          5072 => x"78",
          5073 => x"78",
          5074 => x"08",
          5075 => x"08",
          5076 => x"5c",
          5077 => x"ff",
          5078 => x"26",
          5079 => x"06",
          5080 => x"99",
          5081 => x"ff",
          5082 => x"2a",
          5083 => x"06",
          5084 => x"7a",
          5085 => x"2a",
          5086 => x"2e",
          5087 => x"5e",
          5088 => x"61",
          5089 => x"fe",
          5090 => x"5e",
          5091 => x"58",
          5092 => x"59",
          5093 => x"83",
          5094 => x"70",
          5095 => x"5b",
          5096 => x"e8",
          5097 => x"57",
          5098 => x"70",
          5099 => x"84",
          5100 => x"71",
          5101 => x"ff",
          5102 => x"83",
          5103 => x"5b",
          5104 => x"05",
          5105 => x"59",
          5106 => x"b9",
          5107 => x"2a",
          5108 => x"10",
          5109 => x"5d",
          5110 => x"83",
          5111 => x"80",
          5112 => x"18",
          5113 => x"2e",
          5114 => x"17",
          5115 => x"86",
          5116 => x"85",
          5117 => x"18",
          5118 => x"1f",
          5119 => x"5d",
          5120 => x"2e",
          5121 => x"b8",
          5122 => x"2e",
          5123 => x"70",
          5124 => x"42",
          5125 => x"2e",
          5126 => x"06",
          5127 => x"33",
          5128 => x"06",
          5129 => x"f8",
          5130 => x"38",
          5131 => x"7a",
          5132 => x"83",
          5133 => x"40",
          5134 => x"33",
          5135 => x"71",
          5136 => x"77",
          5137 => x"2e",
          5138 => x"83",
          5139 => x"81",
          5140 => x"40",
          5141 => x"58",
          5142 => x"38",
          5143 => x"fe",
          5144 => x"38",
          5145 => x"0d",
          5146 => x"dc",
          5147 => x"e4",
          5148 => x"8d",
          5149 => x"0d",
          5150 => x"e4",
          5151 => x"05",
          5152 => x"33",
          5153 => x"5f",
          5154 => x"74",
          5155 => x"8a",
          5156 => x"78",
          5157 => x"81",
          5158 => x"1b",
          5159 => x"84",
          5160 => x"93",
          5161 => x"83",
          5162 => x"e9",
          5163 => x"88",
          5164 => x"09",
          5165 => x"58",
          5166 => x"b1",
          5167 => x"2e",
          5168 => x"54",
          5169 => x"33",
          5170 => x"c8",
          5171 => x"81",
          5172 => x"99",
          5173 => x"17",
          5174 => x"2b",
          5175 => x"2e",
          5176 => x"17",
          5177 => x"90",
          5178 => x"33",
          5179 => x"71",
          5180 => x"59",
          5181 => x"09",
          5182 => x"17",
          5183 => x"90",
          5184 => x"33",
          5185 => x"71",
          5186 => x"5e",
          5187 => x"09",
          5188 => x"17",
          5189 => x"90",
          5190 => x"33",
          5191 => x"71",
          5192 => x"1c",
          5193 => x"90",
          5194 => x"33",
          5195 => x"71",
          5196 => x"49",
          5197 => x"5a",
          5198 => x"81",
          5199 => x"7c",
          5200 => x"8c",
          5201 => x"f7",
          5202 => x"38",
          5203 => x"39",
          5204 => x"17",
          5205 => x"ff",
          5206 => x"7a",
          5207 => x"84",
          5208 => x"17",
          5209 => x"a0",
          5210 => x"33",
          5211 => x"84",
          5212 => x"74",
          5213 => x"85",
          5214 => x"5c",
          5215 => x"17",
          5216 => x"2b",
          5217 => x"d2",
          5218 => x"ca",
          5219 => x"82",
          5220 => x"2b",
          5221 => x"88",
          5222 => x"0c",
          5223 => x"40",
          5224 => x"75",
          5225 => x"f9",
          5226 => x"38",
          5227 => x"f7",
          5228 => x"38",
          5229 => x"08",
          5230 => x"81",
          5231 => x"fc",
          5232 => x"d3",
          5233 => x"41",
          5234 => x"80",
          5235 => x"05",
          5236 => x"74",
          5237 => x"38",
          5238 => x"d1",
          5239 => x"c4",
          5240 => x"05",
          5241 => x"84",
          5242 => x"80",
          5243 => x"54",
          5244 => x"2e",
          5245 => x"53",
          5246 => x"b9",
          5247 => x"0c",
          5248 => x"b9",
          5249 => x"33",
          5250 => x"56",
          5251 => x"16",
          5252 => x"58",
          5253 => x"7f",
          5254 => x"7b",
          5255 => x"05",
          5256 => x"33",
          5257 => x"99",
          5258 => x"ff",
          5259 => x"76",
          5260 => x"81",
          5261 => x"9f",
          5262 => x"81",
          5263 => x"77",
          5264 => x"9f",
          5265 => x"80",
          5266 => x"5d",
          5267 => x"7f",
          5268 => x"f7",
          5269 => x"8b",
          5270 => x"05",
          5271 => x"56",
          5272 => x"06",
          5273 => x"9e",
          5274 => x"3f",
          5275 => x"c8",
          5276 => x"0c",
          5277 => x"9c",
          5278 => x"90",
          5279 => x"84",
          5280 => x"08",
          5281 => x"06",
          5282 => x"76",
          5283 => x"2e",
          5284 => x"76",
          5285 => x"06",
          5286 => x"66",
          5287 => x"88",
          5288 => x"5e",
          5289 => x"38",
          5290 => x"8f",
          5291 => x"80",
          5292 => x"a0",
          5293 => x"5e",
          5294 => x"9b",
          5295 => x"2e",
          5296 => x"9c",
          5297 => x"80",
          5298 => x"1c",
          5299 => x"34",
          5300 => x"b4",
          5301 => x"5f",
          5302 => x"17",
          5303 => x"57",
          5304 => x"80",
          5305 => x"5b",
          5306 => x"78",
          5307 => x"38",
          5308 => x"05",
          5309 => x"56",
          5310 => x"81",
          5311 => x"75",
          5312 => x"77",
          5313 => x"2e",
          5314 => x"7e",
          5315 => x"a4",
          5316 => x"12",
          5317 => x"40",
          5318 => x"81",
          5319 => x"16",
          5320 => x"90",
          5321 => x"33",
          5322 => x"71",
          5323 => x"60",
          5324 => x"5e",
          5325 => x"90",
          5326 => x"80",
          5327 => x"81",
          5328 => x"38",
          5329 => x"94",
          5330 => x"2b",
          5331 => x"78",
          5332 => x"27",
          5333 => x"5f",
          5334 => x"77",
          5335 => x"84",
          5336 => x"08",
          5337 => x"b9",
          5338 => x"75",
          5339 => x"c2",
          5340 => x"38",
          5341 => x"80",
          5342 => x"79",
          5343 => x"79",
          5344 => x"79",
          5345 => x"ca",
          5346 => x"07",
          5347 => x"8b",
          5348 => x"fe",
          5349 => x"33",
          5350 => x"7d",
          5351 => x"7c",
          5352 => x"74",
          5353 => x"84",
          5354 => x"08",
          5355 => x"c8",
          5356 => x"b9",
          5357 => x"80",
          5358 => x"82",
          5359 => x"38",
          5360 => x"08",
          5361 => x"af",
          5362 => x"17",
          5363 => x"34",
          5364 => x"38",
          5365 => x"34",
          5366 => x"39",
          5367 => x"98",
          5368 => x"5e",
          5369 => x"80",
          5370 => x"17",
          5371 => x"66",
          5372 => x"67",
          5373 => x"80",
          5374 => x"7c",
          5375 => x"38",
          5376 => x"5e",
          5377 => x"2e",
          5378 => x"7d",
          5379 => x"54",
          5380 => x"33",
          5381 => x"c8",
          5382 => x"81",
          5383 => x"7a",
          5384 => x"80",
          5385 => x"f9",
          5386 => x"53",
          5387 => x"52",
          5388 => x"c8",
          5389 => x"aa",
          5390 => x"34",
          5391 => x"84",
          5392 => x"17",
          5393 => x"33",
          5394 => x"ff",
          5395 => x"a0",
          5396 => x"16",
          5397 => x"5b",
          5398 => x"76",
          5399 => x"0c",
          5400 => x"06",
          5401 => x"7e",
          5402 => x"5f",
          5403 => x"38",
          5404 => x"1c",
          5405 => x"f9",
          5406 => x"1a",
          5407 => x"94",
          5408 => x"81",
          5409 => x"84",
          5410 => x"f7",
          5411 => x"9f",
          5412 => x"66",
          5413 => x"89",
          5414 => x"08",
          5415 => x"33",
          5416 => x"16",
          5417 => x"78",
          5418 => x"41",
          5419 => x"1a",
          5420 => x"1a",
          5421 => x"80",
          5422 => x"8c",
          5423 => x"75",
          5424 => x"81",
          5425 => x"06",
          5426 => x"22",
          5427 => x"7a",
          5428 => x"1a",
          5429 => x"38",
          5430 => x"98",
          5431 => x"fe",
          5432 => x"57",
          5433 => x"19",
          5434 => x"05",
          5435 => x"38",
          5436 => x"77",
          5437 => x"55",
          5438 => x"31",
          5439 => x"81",
          5440 => x"84",
          5441 => x"83",
          5442 => x"a9",
          5443 => x"75",
          5444 => x"71",
          5445 => x"75",
          5446 => x"81",
          5447 => x"ef",
          5448 => x"31",
          5449 => x"94",
          5450 => x"0c",
          5451 => x"56",
          5452 => x"0d",
          5453 => x"3d",
          5454 => x"9c",
          5455 => x"84",
          5456 => x"27",
          5457 => x"19",
          5458 => x"83",
          5459 => x"7f",
          5460 => x"81",
          5461 => x"19",
          5462 => x"b9",
          5463 => x"56",
          5464 => x"81",
          5465 => x"ff",
          5466 => x"05",
          5467 => x"38",
          5468 => x"70",
          5469 => x"75",
          5470 => x"81",
          5471 => x"59",
          5472 => x"fe",
          5473 => x"53",
          5474 => x"52",
          5475 => x"84",
          5476 => x"06",
          5477 => x"83",
          5478 => x"08",
          5479 => x"74",
          5480 => x"82",
          5481 => x"81",
          5482 => x"19",
          5483 => x"52",
          5484 => x"3f",
          5485 => x"1b",
          5486 => x"39",
          5487 => x"a3",
          5488 => x"fc",
          5489 => x"9c",
          5490 => x"06",
          5491 => x"08",
          5492 => x"91",
          5493 => x"0c",
          5494 => x"1b",
          5495 => x"92",
          5496 => x"65",
          5497 => x"7e",
          5498 => x"38",
          5499 => x"38",
          5500 => x"38",
          5501 => x"59",
          5502 => x"55",
          5503 => x"38",
          5504 => x"38",
          5505 => x"06",
          5506 => x"82",
          5507 => x"5d",
          5508 => x"09",
          5509 => x"76",
          5510 => x"38",
          5511 => x"89",
          5512 => x"76",
          5513 => x"74",
          5514 => x"2e",
          5515 => x"8c",
          5516 => x"08",
          5517 => x"56",
          5518 => x"81",
          5519 => x"9c",
          5520 => x"77",
          5521 => x"70",
          5522 => x"57",
          5523 => x"15",
          5524 => x"2e",
          5525 => x"7f",
          5526 => x"77",
          5527 => x"33",
          5528 => x"c8",
          5529 => x"08",
          5530 => x"a5",
          5531 => x"72",
          5532 => x"81",
          5533 => x"59",
          5534 => x"60",
          5535 => x"2b",
          5536 => x"7f",
          5537 => x"70",
          5538 => x"5a",
          5539 => x"83",
          5540 => x"7a",
          5541 => x"77",
          5542 => x"34",
          5543 => x"92",
          5544 => x"0c",
          5545 => x"55",
          5546 => x"a2",
          5547 => x"76",
          5548 => x"5a",
          5549 => x"59",
          5550 => x"b6",
          5551 => x"5e",
          5552 => x"06",
          5553 => x"b8",
          5554 => x"98",
          5555 => x"2e",
          5556 => x"b4",
          5557 => x"94",
          5558 => x"58",
          5559 => x"80",
          5560 => x"58",
          5561 => x"ff",
          5562 => x"81",
          5563 => x"81",
          5564 => x"70",
          5565 => x"98",
          5566 => x"08",
          5567 => x"38",
          5568 => x"b4",
          5569 => x"b9",
          5570 => x"08",
          5571 => x"55",
          5572 => x"e3",
          5573 => x"17",
          5574 => x"33",
          5575 => x"fe",
          5576 => x"1a",
          5577 => x"33",
          5578 => x"b4",
          5579 => x"7b",
          5580 => x"39",
          5581 => x"ab",
          5582 => x"84",
          5583 => x"1a",
          5584 => x"79",
          5585 => x"c8",
          5586 => x"bd",
          5587 => x"08",
          5588 => x"33",
          5589 => x"b9",
          5590 => x"c8",
          5591 => x"a8",
          5592 => x"08",
          5593 => x"5c",
          5594 => x"fc",
          5595 => x"17",
          5596 => x"33",
          5597 => x"fb",
          5598 => x"95",
          5599 => x"06",
          5600 => x"08",
          5601 => x"b4",
          5602 => x"81",
          5603 => x"3f",
          5604 => x"84",
          5605 => x"16",
          5606 => x"a0",
          5607 => x"16",
          5608 => x"06",
          5609 => x"08",
          5610 => x"81",
          5611 => x"60",
          5612 => x"58",
          5613 => x"1b",
          5614 => x"92",
          5615 => x"34",
          5616 => x"3d",
          5617 => x"89",
          5618 => x"08",
          5619 => x"33",
          5620 => x"16",
          5621 => x"77",
          5622 => x"5c",
          5623 => x"18",
          5624 => x"57",
          5625 => x"a0",
          5626 => x"79",
          5627 => x"7a",
          5628 => x"b8",
          5629 => x"93",
          5630 => x"2e",
          5631 => x"b4",
          5632 => x"18",
          5633 => x"57",
          5634 => x"19",
          5635 => x"5a",
          5636 => x"2a",
          5637 => x"76",
          5638 => x"83",
          5639 => x"55",
          5640 => x"7a",
          5641 => x"75",
          5642 => x"78",
          5643 => x"0b",
          5644 => x"34",
          5645 => x"0b",
          5646 => x"34",
          5647 => x"7b",
          5648 => x"c8",
          5649 => x"5b",
          5650 => x"b9",
          5651 => x"54",
          5652 => x"53",
          5653 => x"b5",
          5654 => x"fe",
          5655 => x"18",
          5656 => x"31",
          5657 => x"a0",
          5658 => x"17",
          5659 => x"06",
          5660 => x"08",
          5661 => x"81",
          5662 => x"79",
          5663 => x"55",
          5664 => x"56",
          5665 => x"55",
          5666 => x"7a",
          5667 => x"75",
          5668 => x"78",
          5669 => x"0b",
          5670 => x"34",
          5671 => x"0b",
          5672 => x"34",
          5673 => x"7b",
          5674 => x"c8",
          5675 => x"5b",
          5676 => x"39",
          5677 => x"3f",
          5678 => x"74",
          5679 => x"5a",
          5680 => x"70",
          5681 => x"c8",
          5682 => x"38",
          5683 => x"74",
          5684 => x"72",
          5685 => x"86",
          5686 => x"71",
          5687 => x"58",
          5688 => x"0c",
          5689 => x"0d",
          5690 => x"bc",
          5691 => x"53",
          5692 => x"56",
          5693 => x"70",
          5694 => x"38",
          5695 => x"9f",
          5696 => x"38",
          5697 => x"38",
          5698 => x"24",
          5699 => x"80",
          5700 => x"0d",
          5701 => x"8c",
          5702 => x"70",
          5703 => x"89",
          5704 => x"ff",
          5705 => x"2e",
          5706 => x"b8",
          5707 => x"76",
          5708 => x"81",
          5709 => x"54",
          5710 => x"12",
          5711 => x"9f",
          5712 => x"e0",
          5713 => x"71",
          5714 => x"73",
          5715 => x"ff",
          5716 => x"70",
          5717 => x"52",
          5718 => x"18",
          5719 => x"ff",
          5720 => x"77",
          5721 => x"51",
          5722 => x"53",
          5723 => x"51",
          5724 => x"55",
          5725 => x"38",
          5726 => x"0d",
          5727 => x"d0",
          5728 => x"c8",
          5729 => x"c6",
          5730 => x"98",
          5731 => x"e2",
          5732 => x"2a",
          5733 => x"b2",
          5734 => x"12",
          5735 => x"5e",
          5736 => x"a4",
          5737 => x"b9",
          5738 => x"b9",
          5739 => x"ff",
          5740 => x"0c",
          5741 => x"94",
          5742 => x"2b",
          5743 => x"54",
          5744 => x"58",
          5745 => x"0d",
          5746 => x"3d",
          5747 => x"80",
          5748 => x"fd",
          5749 => x"cf",
          5750 => x"84",
          5751 => x"80",
          5752 => x"08",
          5753 => x"3d",
          5754 => x"cc",
          5755 => x"5b",
          5756 => x"3f",
          5757 => x"c8",
          5758 => x"3d",
          5759 => x"2e",
          5760 => x"17",
          5761 => x"81",
          5762 => x"16",
          5763 => x"b9",
          5764 => x"57",
          5765 => x"82",
          5766 => x"11",
          5767 => x"07",
          5768 => x"56",
          5769 => x"80",
          5770 => x"ff",
          5771 => x"59",
          5772 => x"80",
          5773 => x"84",
          5774 => x"08",
          5775 => x"11",
          5776 => x"07",
          5777 => x"56",
          5778 => x"7a",
          5779 => x"52",
          5780 => x"b9",
          5781 => x"80",
          5782 => x"83",
          5783 => x"e4",
          5784 => x"ff",
          5785 => x"33",
          5786 => x"82",
          5787 => x"33",
          5788 => x"17",
          5789 => x"76",
          5790 => x"05",
          5791 => x"11",
          5792 => x"58",
          5793 => x"ff",
          5794 => x"58",
          5795 => x"5a",
          5796 => x"82",
          5797 => x"33",
          5798 => x"70",
          5799 => x"5a",
          5800 => x"70",
          5801 => x"f5",
          5802 => x"ab",
          5803 => x"38",
          5804 => x"81",
          5805 => x"77",
          5806 => x"05",
          5807 => x"06",
          5808 => x"34",
          5809 => x"3d",
          5810 => x"33",
          5811 => x"79",
          5812 => x"95",
          5813 => x"2b",
          5814 => x"dd",
          5815 => x"51",
          5816 => x"08",
          5817 => x"fd",
          5818 => x"b4",
          5819 => x"81",
          5820 => x"3f",
          5821 => x"be",
          5822 => x"34",
          5823 => x"84",
          5824 => x"17",
          5825 => x"33",
          5826 => x"fb",
          5827 => x"a0",
          5828 => x"16",
          5829 => x"59",
          5830 => x"3d",
          5831 => x"80",
          5832 => x"10",
          5833 => x"33",
          5834 => x"2e",
          5835 => x"f1",
          5836 => x"19",
          5837 => x"05",
          5838 => x"38",
          5839 => x"59",
          5840 => x"5e",
          5841 => x"f5",
          5842 => x"84",
          5843 => x"04",
          5844 => x"89",
          5845 => x"08",
          5846 => x"33",
          5847 => x"14",
          5848 => x"78",
          5849 => x"5a",
          5850 => x"15",
          5851 => x"15",
          5852 => x"38",
          5853 => x"78",
          5854 => x"22",
          5855 => x"78",
          5856 => x"17",
          5857 => x"c8",
          5858 => x"55",
          5859 => x"c8",
          5860 => x"30",
          5861 => x"71",
          5862 => x"73",
          5863 => x"27",
          5864 => x"16",
          5865 => x"33",
          5866 => x"57",
          5867 => x"52",
          5868 => x"b9",
          5869 => x"80",
          5870 => x"98",
          5871 => x"79",
          5872 => x"aa",
          5873 => x"39",
          5874 => x"72",
          5875 => x"04",
          5876 => x"06",
          5877 => x"94",
          5878 => x"78",
          5879 => x"77",
          5880 => x"75",
          5881 => x"0c",
          5882 => x"76",
          5883 => x"59",
          5884 => x"08",
          5885 => x"0c",
          5886 => x"3d",
          5887 => x"88",
          5888 => x"fe",
          5889 => x"2e",
          5890 => x"b9",
          5891 => x"94",
          5892 => x"75",
          5893 => x"9c",
          5894 => x"73",
          5895 => x"22",
          5896 => x"78",
          5897 => x"80",
          5898 => x"56",
          5899 => x"ff",
          5900 => x"54",
          5901 => x"ff",
          5902 => x"81",
          5903 => x"75",
          5904 => x"52",
          5905 => x"b9",
          5906 => x"81",
          5907 => x"ff",
          5908 => x"08",
          5909 => x"fe",
          5910 => x"82",
          5911 => x"0d",
          5912 => x"54",
          5913 => x"8c",
          5914 => x"05",
          5915 => x"08",
          5916 => x"8f",
          5917 => x"84",
          5918 => x"7a",
          5919 => x"b9",
          5920 => x"84",
          5921 => x"16",
          5922 => x"78",
          5923 => x"84",
          5924 => x"2e",
          5925 => x"11",
          5926 => x"07",
          5927 => x"57",
          5928 => x"17",
          5929 => x"17",
          5930 => x"b9",
          5931 => x"84",
          5932 => x"84",
          5933 => x"85",
          5934 => x"95",
          5935 => x"2b",
          5936 => x"19",
          5937 => x"3d",
          5938 => x"2e",
          5939 => x"2e",
          5940 => x"2e",
          5941 => x"22",
          5942 => x"80",
          5943 => x"75",
          5944 => x"3d",
          5945 => x"ff",
          5946 => x"06",
          5947 => x"53",
          5948 => x"7c",
          5949 => x"9f",
          5950 => x"97",
          5951 => x"8f",
          5952 => x"59",
          5953 => x"80",
          5954 => x"c7",
          5955 => x"75",
          5956 => x"84",
          5957 => x"08",
          5958 => x"08",
          5959 => x"b2",
          5960 => x"99",
          5961 => x"32",
          5962 => x"84",
          5963 => x"72",
          5964 => x"04",
          5965 => x"b1",
          5966 => x"99",
          5967 => x"32",
          5968 => x"84",
          5969 => x"cf",
          5970 => x"f9",
          5971 => x"c8",
          5972 => x"33",
          5973 => x"c8",
          5974 => x"38",
          5975 => x"39",
          5976 => x"89",
          5977 => x"c1",
          5978 => x"84",
          5979 => x"74",
          5980 => x"04",
          5981 => x"3f",
          5982 => x"c8",
          5983 => x"33",
          5984 => x"24",
          5985 => x"76",
          5986 => x"74",
          5987 => x"04",
          5988 => x"3d",
          5989 => x"56",
          5990 => x"52",
          5991 => x"b9",
          5992 => x"9a",
          5993 => x"11",
          5994 => x"57",
          5995 => x"75",
          5996 => x"95",
          5997 => x"77",
          5998 => x"93",
          5999 => x"c8",
          6000 => x"38",
          6001 => x"b4",
          6002 => x"83",
          6003 => x"8d",
          6004 => x"52",
          6005 => x"3f",
          6006 => x"38",
          6007 => x"0c",
          6008 => x"38",
          6009 => x"8d",
          6010 => x"33",
          6011 => x"88",
          6012 => x"07",
          6013 => x"ff",
          6014 => x"80",
          6015 => x"ff",
          6016 => x"53",
          6017 => x"78",
          6018 => x"94",
          6019 => x"58",
          6020 => x"c8",
          6021 => x"b4",
          6022 => x"81",
          6023 => x"3f",
          6024 => x"f8",
          6025 => x"34",
          6026 => x"84",
          6027 => x"18",
          6028 => x"33",
          6029 => x"fe",
          6030 => x"a0",
          6031 => x"17",
          6032 => x"5e",
          6033 => x"3d",
          6034 => x"81",
          6035 => x"2e",
          6036 => x"81",
          6037 => x"08",
          6038 => x"80",
          6039 => x"58",
          6040 => x"ca",
          6041 => x"0c",
          6042 => x"84",
          6043 => x"b8",
          6044 => x"88",
          6045 => x"1f",
          6046 => x"5f",
          6047 => x"fd",
          6048 => x"fd",
          6049 => x"7f",
          6050 => x"33",
          6051 => x"fe",
          6052 => x"39",
          6053 => x"76",
          6054 => x"74",
          6055 => x"73",
          6056 => x"84",
          6057 => x"81",
          6058 => x"80",
          6059 => x"80",
          6060 => x"2a",
          6061 => x"80",
          6062 => x"54",
          6063 => x"73",
          6064 => x"08",
          6065 => x"9c",
          6066 => x"56",
          6067 => x"08",
          6068 => x"59",
          6069 => x"85",
          6070 => x"74",
          6071 => x"04",
          6072 => x"38",
          6073 => x"3f",
          6074 => x"c8",
          6075 => x"b9",
          6076 => x"84",
          6077 => x"38",
          6078 => x"85",
          6079 => x"c8",
          6080 => x"18",
          6081 => x"ff",
          6082 => x"84",
          6083 => x"17",
          6084 => x"a0",
          6085 => x"fe",
          6086 => x"81",
          6087 => x"77",
          6088 => x"0b",
          6089 => x"80",
          6090 => x"98",
          6091 => x"b9",
          6092 => x"81",
          6093 => x"2e",
          6094 => x"79",
          6095 => x"08",
          6096 => x"08",
          6097 => x"54",
          6098 => x"81",
          6099 => x"17",
          6100 => x"2e",
          6101 => x"51",
          6102 => x"08",
          6103 => x"38",
          6104 => x"3f",
          6105 => x"c8",
          6106 => x"b9",
          6107 => x"84",
          6108 => x"38",
          6109 => x"83",
          6110 => x"e6",
          6111 => x"18",
          6112 => x"90",
          6113 => x"16",
          6114 => x"34",
          6115 => x"38",
          6116 => x"58",
          6117 => x"39",
          6118 => x"fc",
          6119 => x"0b",
          6120 => x"39",
          6121 => x"59",
          6122 => x"18",
          6123 => x"b9",
          6124 => x"ff",
          6125 => x"a7",
          6126 => x"51",
          6127 => x"08",
          6128 => x"8a",
          6129 => x"3d",
          6130 => x"52",
          6131 => x"f8",
          6132 => x"b9",
          6133 => x"05",
          6134 => x"57",
          6135 => x"2b",
          6136 => x"80",
          6137 => x"57",
          6138 => x"a3",
          6139 => x"33",
          6140 => x"5e",
          6141 => x"d5",
          6142 => x"76",
          6143 => x"98",
          6144 => x"77",
          6145 => x"52",
          6146 => x"f9",
          6147 => x"b9",
          6148 => x"c8",
          6149 => x"3f",
          6150 => x"c8",
          6151 => x"c8",
          6152 => x"33",
          6153 => x"90",
          6154 => x"ff",
          6155 => x"2e",
          6156 => x"a1",
          6157 => x"57",
          6158 => x"38",
          6159 => x"3f",
          6160 => x"c8",
          6161 => x"70",
          6162 => x"80",
          6163 => x"38",
          6164 => x"27",
          6165 => x"81",
          6166 => x"38",
          6167 => x"b9",
          6168 => x"3d",
          6169 => x"08",
          6170 => x"2e",
          6171 => x"59",
          6172 => x"80",
          6173 => x"17",
          6174 => x"ee",
          6175 => x"85",
          6176 => x"18",
          6177 => x"19",
          6178 => x"83",
          6179 => x"fe",
          6180 => x"8b",
          6181 => x"84",
          6182 => x"38",
          6183 => x"cd",
          6184 => x"54",
          6185 => x"17",
          6186 => x"58",
          6187 => x"81",
          6188 => x"08",
          6189 => x"18",
          6190 => x"55",
          6191 => x"38",
          6192 => x"09",
          6193 => x"b4",
          6194 => x"7c",
          6195 => x"c5",
          6196 => x"55",
          6197 => x"52",
          6198 => x"b9",
          6199 => x"80",
          6200 => x"08",
          6201 => x"c8",
          6202 => x"53",
          6203 => x"3f",
          6204 => x"17",
          6205 => x"5c",
          6206 => x"81",
          6207 => x"81",
          6208 => x"55",
          6209 => x"56",
          6210 => x"39",
          6211 => x"39",
          6212 => x"0d",
          6213 => x"52",
          6214 => x"84",
          6215 => x"08",
          6216 => x"c8",
          6217 => x"6f",
          6218 => x"a6",
          6219 => x"84",
          6220 => x"84",
          6221 => x"84",
          6222 => x"06",
          6223 => x"70",
          6224 => x"56",
          6225 => x"52",
          6226 => x"c0",
          6227 => x"5c",
          6228 => x"56",
          6229 => x"f9",
          6230 => x"81",
          6231 => x"84",
          6232 => x"5a",
          6233 => x"9c",
          6234 => x"5b",
          6235 => x"22",
          6236 => x"5c",
          6237 => x"59",
          6238 => x"70",
          6239 => x"74",
          6240 => x"55",
          6241 => x"54",
          6242 => x"33",
          6243 => x"c8",
          6244 => x"dc",
          6245 => x"54",
          6246 => x"53",
          6247 => x"a5",
          6248 => x"be",
          6249 => x"34",
          6250 => x"55",
          6251 => x"38",
          6252 => x"09",
          6253 => x"b4",
          6254 => x"77",
          6255 => x"e5",
          6256 => x"7d",
          6257 => x"b4",
          6258 => x"ac",
          6259 => x"f9",
          6260 => x"b9",
          6261 => x"84",
          6262 => x"38",
          6263 => x"84",
          6264 => x"fe",
          6265 => x"fc",
          6266 => x"94",
          6267 => x"27",
          6268 => x"84",
          6269 => x"18",
          6270 => x"a1",
          6271 => x"3d",
          6272 => x"83",
          6273 => x"78",
          6274 => x"8b",
          6275 => x"70",
          6276 => x"75",
          6277 => x"18",
          6278 => x"19",
          6279 => x"34",
          6280 => x"80",
          6281 => x"d1",
          6282 => x"06",
          6283 => x"77",
          6284 => x"34",
          6285 => x"cc",
          6286 => x"1a",
          6287 => x"81",
          6288 => x"59",
          6289 => x"7d",
          6290 => x"64",
          6291 => x"57",
          6292 => x"88",
          6293 => x"75",
          6294 => x"38",
          6295 => x"79",
          6296 => x"c8",
          6297 => x"b6",
          6298 => x"96",
          6299 => x"17",
          6300 => x"cc",
          6301 => x"5d",
          6302 => x"59",
          6303 => x"79",
          6304 => x"90",
          6305 => x"0b",
          6306 => x"80",
          6307 => x"84",
          6308 => x"76",
          6309 => x"34",
          6310 => x"17",
          6311 => x"5b",
          6312 => x"2a",
          6313 => x"59",
          6314 => x"57",
          6315 => x"2a",
          6316 => x"2a",
          6317 => x"90",
          6318 => x"0b",
          6319 => x"98",
          6320 => x"96",
          6321 => x"3d",
          6322 => x"2e",
          6323 => x"33",
          6324 => x"2e",
          6325 => x"ba",
          6326 => x"3d",
          6327 => x"ff",
          6328 => x"56",
          6329 => x"38",
          6330 => x"0d",
          6331 => x"08",
          6332 => x"9f",
          6333 => x"84",
          6334 => x"bb",
          6335 => x"56",
          6336 => x"ae",
          6337 => x"81",
          6338 => x"59",
          6339 => x"99",
          6340 => x"55",
          6341 => x"70",
          6342 => x"74",
          6343 => x"51",
          6344 => x"08",
          6345 => x"38",
          6346 => x"38",
          6347 => x"3d",
          6348 => x"81",
          6349 => x"26",
          6350 => x"06",
          6351 => x"80",
          6352 => x"b8",
          6353 => x"5c",
          6354 => x"70",
          6355 => x"5a",
          6356 => x"e0",
          6357 => x"ff",
          6358 => x"38",
          6359 => x"55",
          6360 => x"75",
          6361 => x"77",
          6362 => x"30",
          6363 => x"5d",
          6364 => x"81",
          6365 => x"24",
          6366 => x"5b",
          6367 => x"b4",
          6368 => x"3d",
          6369 => x"ff",
          6370 => x"56",
          6371 => x"fd",
          6372 => x"09",
          6373 => x"ff",
          6374 => x"56",
          6375 => x"6f",
          6376 => x"05",
          6377 => x"70",
          6378 => x"05",
          6379 => x"38",
          6380 => x"34",
          6381 => x"06",
          6382 => x"07",
          6383 => x"81",
          6384 => x"70",
          6385 => x"80",
          6386 => x"6b",
          6387 => x"33",
          6388 => x"72",
          6389 => x"2e",
          6390 => x"08",
          6391 => x"82",
          6392 => x"29",
          6393 => x"80",
          6394 => x"58",
          6395 => x"83",
          6396 => x"81",
          6397 => x"17",
          6398 => x"b9",
          6399 => x"58",
          6400 => x"57",
          6401 => x"fb",
          6402 => x"ae",
          6403 => x"70",
          6404 => x"80",
          6405 => x"77",
          6406 => x"7a",
          6407 => x"75",
          6408 => x"34",
          6409 => x"18",
          6410 => x"34",
          6411 => x"08",
          6412 => x"38",
          6413 => x"3f",
          6414 => x"c8",
          6415 => x"98",
          6416 => x"08",
          6417 => x"7a",
          6418 => x"06",
          6419 => x"b8",
          6420 => x"e2",
          6421 => x"2e",
          6422 => x"b4",
          6423 => x"9c",
          6424 => x"0b",
          6425 => x"27",
          6426 => x"fc",
          6427 => x"84",
          6428 => x"38",
          6429 => x"38",
          6430 => x"51",
          6431 => x"08",
          6432 => x"04",
          6433 => x"3d",
          6434 => x"33",
          6435 => x"78",
          6436 => x"84",
          6437 => x"38",
          6438 => x"a0",
          6439 => x"3d",
          6440 => x"53",
          6441 => x"e2",
          6442 => x"08",
          6443 => x"38",
          6444 => x"b4",
          6445 => x"b9",
          6446 => x"08",
          6447 => x"5d",
          6448 => x"93",
          6449 => x"17",
          6450 => x"33",
          6451 => x"fd",
          6452 => x"53",
          6453 => x"52",
          6454 => x"84",
          6455 => x"b9",
          6456 => x"08",
          6457 => x"08",
          6458 => x"fc",
          6459 => x"82",
          6460 => x"81",
          6461 => x"05",
          6462 => x"fe",
          6463 => x"39",
          6464 => x"33",
          6465 => x"56",
          6466 => x"52",
          6467 => x"84",
          6468 => x"08",
          6469 => x"c8",
          6470 => x"66",
          6471 => x"96",
          6472 => x"84",
          6473 => x"cf",
          6474 => x"56",
          6475 => x"71",
          6476 => x"74",
          6477 => x"8b",
          6478 => x"16",
          6479 => x"84",
          6480 => x"96",
          6481 => x"57",
          6482 => x"97",
          6483 => x"b9",
          6484 => x"80",
          6485 => x"0c",
          6486 => x"52",
          6487 => x"d8",
          6488 => x"b9",
          6489 => x"05",
          6490 => x"75",
          6491 => x"19",
          6492 => x"56",
          6493 => x"55",
          6494 => x"58",
          6495 => x"54",
          6496 => x"0b",
          6497 => x"88",
          6498 => x"c8",
          6499 => x"0d",
          6500 => x"3d",
          6501 => x"a0",
          6502 => x"b9",
          6503 => x"08",
          6504 => x"80",
          6505 => x"5a",
          6506 => x"70",
          6507 => x"80",
          6508 => x"06",
          6509 => x"38",
          6510 => x"5a",
          6511 => x"38",
          6512 => x"7a",
          6513 => x"81",
          6514 => x"16",
          6515 => x"b9",
          6516 => x"57",
          6517 => x"57",
          6518 => x"58",
          6519 => x"38",
          6520 => x"38",
          6521 => x"11",
          6522 => x"71",
          6523 => x"72",
          6524 => x"62",
          6525 => x"76",
          6526 => x"04",
          6527 => x"3d",
          6528 => x"84",
          6529 => x"08",
          6530 => x"2e",
          6531 => x"7b",
          6532 => x"54",
          6533 => x"53",
          6534 => x"ad",
          6535 => x"7a",
          6536 => x"84",
          6537 => x"16",
          6538 => x"c8",
          6539 => x"27",
          6540 => x"74",
          6541 => x"38",
          6542 => x"08",
          6543 => x"51",
          6544 => x"54",
          6545 => x"33",
          6546 => x"c8",
          6547 => x"86",
          6548 => x"bb",
          6549 => x"b9",
          6550 => x"c8",
          6551 => x"59",
          6552 => x"57",
          6553 => x"19",
          6554 => x"70",
          6555 => x"80",
          6556 => x"11",
          6557 => x"2e",
          6558 => x"fd",
          6559 => x"a1",
          6560 => x"51",
          6561 => x"08",
          6562 => x"38",
          6563 => x"a0",
          6564 => x"15",
          6565 => x"08",
          6566 => x"58",
          6567 => x"38",
          6568 => x"81",
          6569 => x"81",
          6570 => x"ff",
          6571 => x"a1",
          6572 => x"c8",
          6573 => x"c8",
          6574 => x"80",
          6575 => x"0b",
          6576 => x"06",
          6577 => x"d6",
          6578 => x"38",
          6579 => x"06",
          6580 => x"38",
          6581 => x"38",
          6582 => x"a3",
          6583 => x"38",
          6584 => x"ff",
          6585 => x"55",
          6586 => x"81",
          6587 => x"5d",
          6588 => x"33",
          6589 => x"5a",
          6590 => x"3d",
          6591 => x"2e",
          6592 => x"02",
          6593 => x"5c",
          6594 => x"87",
          6595 => x"7d",
          6596 => x"70",
          6597 => x"b9",
          6598 => x"80",
          6599 => x"b9",
          6600 => x"b5",
          6601 => x"b9",
          6602 => x"74",
          6603 => x"b9",
          6604 => x"e6",
          6605 => x"52",
          6606 => x"b9",
          6607 => x"80",
          6608 => x"38",
          6609 => x"70",
          6610 => x"05",
          6611 => x"38",
          6612 => x"7d",
          6613 => x"c8",
          6614 => x"8a",
          6615 => x"ff",
          6616 => x"2e",
          6617 => x"55",
          6618 => x"08",
          6619 => x"b1",
          6620 => x"b9",
          6621 => x"81",
          6622 => x"19",
          6623 => x"59",
          6624 => x"83",
          6625 => x"81",
          6626 => x"53",
          6627 => x"fe",
          6628 => x"80",
          6629 => x"76",
          6630 => x"38",
          6631 => x"5a",
          6632 => x"38",
          6633 => x"56",
          6634 => x"81",
          6635 => x"81",
          6636 => x"84",
          6637 => x"08",
          6638 => x"76",
          6639 => x"76",
          6640 => x"80",
          6641 => x"15",
          6642 => x"0b",
          6643 => x"57",
          6644 => x"76",
          6645 => x"55",
          6646 => x"70",
          6647 => x"05",
          6648 => x"38",
          6649 => x"34",
          6650 => x"7d",
          6651 => x"c8",
          6652 => x"fe",
          6653 => x"53",
          6654 => x"d4",
          6655 => x"2e",
          6656 => x"b9",
          6657 => x"08",
          6658 => x"19",
          6659 => x"55",
          6660 => x"c8",
          6661 => x"81",
          6662 => x"84",
          6663 => x"08",
          6664 => x"39",
          6665 => x"fd",
          6666 => x"b4",
          6667 => x"7a",
          6668 => x"fd",
          6669 => x"60",
          6670 => x"33",
          6671 => x"2e",
          6672 => x"2e",
          6673 => x"2e",
          6674 => x"22",
          6675 => x"38",
          6676 => x"38",
          6677 => x"38",
          6678 => x"17",
          6679 => x"70",
          6680 => x"80",
          6681 => x"22",
          6682 => x"57",
          6683 => x"15",
          6684 => x"9f",
          6685 => x"1c",
          6686 => x"81",
          6687 => x"78",
          6688 => x"56",
          6689 => x"fe",
          6690 => x"55",
          6691 => x"82",
          6692 => x"81",
          6693 => x"2e",
          6694 => x"81",
          6695 => x"2e",
          6696 => x"06",
          6697 => x"84",
          6698 => x"87",
          6699 => x"0d",
          6700 => x"ac",
          6701 => x"54",
          6702 => x"55",
          6703 => x"81",
          6704 => x"80",
          6705 => x"81",
          6706 => x"52",
          6707 => x"b9",
          6708 => x"ff",
          6709 => x"57",
          6710 => x"90",
          6711 => x"8c",
          6712 => x"18",
          6713 => x"5c",
          6714 => x"fe",
          6715 => x"7a",
          6716 => x"94",
          6717 => x"5d",
          6718 => x"d6",
          6719 => x"5b",
          6720 => x"fe",
          6721 => x"ff",
          6722 => x"d4",
          6723 => x"a5",
          6724 => x"05",
          6725 => x"3d",
          6726 => x"2e",
          6727 => x"5b",
          6728 => x"ba",
          6729 => x"75",
          6730 => x"a4",
          6731 => x"38",
          6732 => x"70",
          6733 => x"38",
          6734 => x"bc",
          6735 => x"40",
          6736 => x"ce",
          6737 => x"ff",
          6738 => x"57",
          6739 => x"81",
          6740 => x"38",
          6741 => x"79",
          6742 => x"c8",
          6743 => x"80",
          6744 => x"80",
          6745 => x"06",
          6746 => x"2e",
          6747 => x"f8",
          6748 => x"f0",
          6749 => x"83",
          6750 => x"08",
          6751 => x"4c",
          6752 => x"38",
          6753 => x"56",
          6754 => x"7d",
          6755 => x"74",
          6756 => x"be",
          6757 => x"83",
          6758 => x"61",
          6759 => x"07",
          6760 => x"d5",
          6761 => x"7d",
          6762 => x"33",
          6763 => x"38",
          6764 => x"12",
          6765 => x"07",
          6766 => x"2b",
          6767 => x"83",
          6768 => x"2b",
          6769 => x"70",
          6770 => x"07",
          6771 => x"0c",
          6772 => x"59",
          6773 => x"57",
          6774 => x"93",
          6775 => x"38",
          6776 => x"49",
          6777 => x"87",
          6778 => x"61",
          6779 => x"83",
          6780 => x"58",
          6781 => x"ae",
          6782 => x"83",
          6783 => x"2e",
          6784 => x"83",
          6785 => x"70",
          6786 => x"86",
          6787 => x"52",
          6788 => x"b9",
          6789 => x"b9",
          6790 => x"81",
          6791 => x"b9",
          6792 => x"83",
          6793 => x"89",
          6794 => x"1f",
          6795 => x"05",
          6796 => x"57",
          6797 => x"74",
          6798 => x"60",
          6799 => x"f2",
          6800 => x"53",
          6801 => x"98",
          6802 => x"83",
          6803 => x"09",
          6804 => x"f5",
          6805 => x"ac",
          6806 => x"55",
          6807 => x"74",
          6808 => x"84",
          6809 => x"b9",
          6810 => x"39",
          6811 => x"3d",
          6812 => x"33",
          6813 => x"57",
          6814 => x"1d",
          6815 => x"58",
          6816 => x"0b",
          6817 => x"7d",
          6818 => x"33",
          6819 => x"9f",
          6820 => x"89",
          6821 => x"58",
          6822 => x"26",
          6823 => x"06",
          6824 => x"5a",
          6825 => x"85",
          6826 => x"32",
          6827 => x"7b",
          6828 => x"80",
          6829 => x"5c",
          6830 => x"56",
          6831 => x"53",
          6832 => x"3f",
          6833 => x"b6",
          6834 => x"b9",
          6835 => x"bf",
          6836 => x"26",
          6837 => x"fb",
          6838 => x"7b",
          6839 => x"a3",
          6840 => x"81",
          6841 => x"fd",
          6842 => x"46",
          6843 => x"08",
          6844 => x"38",
          6845 => x"fb",
          6846 => x"c8",
          6847 => x"0c",
          6848 => x"99",
          6849 => x"74",
          6850 => x"ae",
          6851 => x"76",
          6852 => x"55",
          6853 => x"84",
          6854 => x"58",
          6855 => x"ff",
          6856 => x"05",
          6857 => x"05",
          6858 => x"83",
          6859 => x"05",
          6860 => x"8f",
          6861 => x"62",
          6862 => x"61",
          6863 => x"06",
          6864 => x"56",
          6865 => x"38",
          6866 => x"61",
          6867 => x"6b",
          6868 => x"05",
          6869 => x"61",
          6870 => x"34",
          6871 => x"9c",
          6872 => x"61",
          6873 => x"6b",
          6874 => x"84",
          6875 => x"61",
          6876 => x"f7",
          6877 => x"61",
          6878 => x"34",
          6879 => x"83",
          6880 => x"05",
          6881 => x"97",
          6882 => x"34",
          6883 => x"ab",
          6884 => x"76",
          6885 => x"81",
          6886 => x"ef",
          6887 => x"d5",
          6888 => x"ff",
          6889 => x"60",
          6890 => x"81",
          6891 => x"38",
          6892 => x"9c",
          6893 => x"70",
          6894 => x"74",
          6895 => x"83",
          6896 => x"f8",
          6897 => x"57",
          6898 => x"45",
          6899 => x"34",
          6900 => x"81",
          6901 => x"75",
          6902 => x"66",
          6903 => x"7a",
          6904 => x"9d",
          6905 => x"38",
          6906 => x"70",
          6907 => x"74",
          6908 => x"58",
          6909 => x"40",
          6910 => x"56",
          6911 => x"65",
          6912 => x"55",
          6913 => x"51",
          6914 => x"08",
          6915 => x"31",
          6916 => x"62",
          6917 => x"83",
          6918 => x"62",
          6919 => x"84",
          6920 => x"5e",
          6921 => x"56",
          6922 => x"34",
          6923 => x"d5",
          6924 => x"83",
          6925 => x"67",
          6926 => x"34",
          6927 => x"84",
          6928 => x"52",
          6929 => x"fe",
          6930 => x"08",
          6931 => x"86",
          6932 => x"87",
          6933 => x"34",
          6934 => x"61",
          6935 => x"08",
          6936 => x"83",
          6937 => x"64",
          6938 => x"2a",
          6939 => x"62",
          6940 => x"05",
          6941 => x"79",
          6942 => x"84",
          6943 => x"53",
          6944 => x"3f",
          6945 => x"b6",
          6946 => x"c8",
          6947 => x"0c",
          6948 => x"1c",
          6949 => x"7a",
          6950 => x"0b",
          6951 => x"80",
          6952 => x"38",
          6953 => x"17",
          6954 => x"2e",
          6955 => x"77",
          6956 => x"84",
          6957 => x"05",
          6958 => x"80",
          6959 => x"8a",
          6960 => x"77",
          6961 => x"e4",
          6962 => x"f5",
          6963 => x"38",
          6964 => x"38",
          6965 => x"06",
          6966 => x"83",
          6967 => x"05",
          6968 => x"a1",
          6969 => x"61",
          6970 => x"76",
          6971 => x"80",
          6972 => x"80",
          6973 => x"05",
          6974 => x"34",
          6975 => x"2a",
          6976 => x"90",
          6977 => x"7c",
          6978 => x"34",
          6979 => x"ad",
          6980 => x"80",
          6981 => x"05",
          6982 => x"61",
          6983 => x"34",
          6984 => x"a9",
          6985 => x"80",
          6986 => x"55",
          6987 => x"70",
          6988 => x"74",
          6989 => x"81",
          6990 => x"58",
          6991 => x"f9",
          6992 => x"52",
          6993 => x"57",
          6994 => x"7d",
          6995 => x"83",
          6996 => x"c8",
          6997 => x"bf",
          6998 => x"84",
          6999 => x"b9",
          7000 => x"4a",
          7001 => x"ff",
          7002 => x"6a",
          7003 => x"61",
          7004 => x"34",
          7005 => x"88",
          7006 => x"ff",
          7007 => x"7c",
          7008 => x"1f",
          7009 => x"d5",
          7010 => x"75",
          7011 => x"57",
          7012 => x"7c",
          7013 => x"80",
          7014 => x"80",
          7015 => x"80",
          7016 => x"e4",
          7017 => x"05",
          7018 => x"34",
          7019 => x"7f",
          7020 => x"05",
          7021 => x"83",
          7022 => x"75",
          7023 => x"2a",
          7024 => x"82",
          7025 => x"83",
          7026 => x"05",
          7027 => x"80",
          7028 => x"81",
          7029 => x"51",
          7030 => x"1f",
          7031 => x"a5",
          7032 => x"39",
          7033 => x"80",
          7034 => x"76",
          7035 => x"8e",
          7036 => x"52",
          7037 => x"81",
          7038 => x"3d",
          7039 => x"74",
          7040 => x"17",
          7041 => x"77",
          7042 => x"55",
          7043 => x"b9",
          7044 => x"3d",
          7045 => x"33",
          7046 => x"38",
          7047 => x"9e",
          7048 => x"05",
          7049 => x"55",
          7050 => x"18",
          7051 => x"3d",
          7052 => x"74",
          7053 => x"ff",
          7054 => x"30",
          7055 => x"84",
          7056 => x"5a",
          7057 => x"51",
          7058 => x"3d",
          7059 => x"3d",
          7060 => x"80",
          7061 => x"15",
          7062 => x"77",
          7063 => x"7c",
          7064 => x"7d",
          7065 => x"75",
          7066 => x"b8",
          7067 => x"88",
          7068 => x"9e",
          7069 => x"75",
          7070 => x"ff",
          7071 => x"86",
          7072 => x"0b",
          7073 => x"04",
          7074 => x"54",
          7075 => x"9d",
          7076 => x"70",
          7077 => x"5a",
          7078 => x"76",
          7079 => x"7d",
          7080 => x"04",
          7081 => x"9a",
          7082 => x"80",
          7083 => x"ff",
          7084 => x"85",
          7085 => x"27",
          7086 => x"06",
          7087 => x"83",
          7088 => x"9c",
          7089 => x"06",
          7090 => x"38",
          7091 => x"22",
          7092 => x"70",
          7093 => x"53",
          7094 => x"02",
          7095 => x"05",
          7096 => x"ff",
          7097 => x"b9",
          7098 => x"83",
          7099 => x"70",
          7100 => x"83",
          7101 => x"c8",
          7102 => x"3d",
          7103 => x"26",
          7104 => x"06",
          7105 => x"ff",
          7106 => x"05",
          7107 => x"25",
          7108 => x"53",
          7109 => x"53",
          7110 => x"81",
          7111 => x"76",
          7112 => x"10",
          7113 => x"54",
          7114 => x"26",
          7115 => x"cb",
          7116 => x"0c",
          7117 => x"55",
          7118 => x"38",
          7119 => x"54",
          7120 => x"83",
          7121 => x"d3",
          7122 => x"ff",
          7123 => x"70",
          7124 => x"39",
          7125 => x"57",
          7126 => x"ff",
          7127 => x"16",
          7128 => x"c5",
          7129 => x"06",
          7130 => x"31",
          7131 => x"ff",
          7132 => x"39",
          7133 => x"22",
          7134 => x"00",
          7135 => x"ff",
          7136 => x"00",
          7137 => x"00",
          7138 => x"00",
          7139 => x"00",
          7140 => x"00",
          7141 => x"00",
          7142 => x"00",
          7143 => x"00",
          7144 => x"00",
          7145 => x"00",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"74",
          7374 => x"74",
          7375 => x"74",
          7376 => x"64",
          7377 => x"63",
          7378 => x"61",
          7379 => x"79",
          7380 => x"66",
          7381 => x"70",
          7382 => x"6d",
          7383 => x"68",
          7384 => x"68",
          7385 => x"63",
          7386 => x"6a",
          7387 => x"61",
          7388 => x"74",
          7389 => x"00",
          7390 => x"00",
          7391 => x"7a",
          7392 => x"69",
          7393 => x"69",
          7394 => x"00",
          7395 => x"55",
          7396 => x"65",
          7397 => x"50",
          7398 => x"72",
          7399 => x"72",
          7400 => x"54",
          7401 => x"20",
          7402 => x"6c",
          7403 => x"49",
          7404 => x"69",
          7405 => x"6f",
          7406 => x"46",
          7407 => x"6c",
          7408 => x"54",
          7409 => x"20",
          7410 => x"6f",
          7411 => x"6c",
          7412 => x"46",
          7413 => x"62",
          7414 => x"4e",
          7415 => x"74",
          7416 => x"6c",
          7417 => x"20",
          7418 => x"6e",
          7419 => x"44",
          7420 => x"20",
          7421 => x"2e",
          7422 => x"65",
          7423 => x"20",
          7424 => x"6c",
          7425 => x"53",
          7426 => x"69",
          7427 => x"65",
          7428 => x"46",
          7429 => x"64",
          7430 => x"6c",
          7431 => x"46",
          7432 => x"65",
          7433 => x"73",
          7434 => x"41",
          7435 => x"65",
          7436 => x"49",
          7437 => x"66",
          7438 => x"2e",
          7439 => x"61",
          7440 => x"64",
          7441 => x"69",
          7442 => x"64",
          7443 => x"20",
          7444 => x"64",
          7445 => x"72",
          7446 => x"6f",
          7447 => x"20",
          7448 => x"53",
          7449 => x"00",
          7450 => x"20",
          7451 => x"73",
          7452 => x"20",
          7453 => x"65",
          7454 => x"72",
          7455 => x"25",
          7456 => x"3a",
          7457 => x"00",
          7458 => x"7c",
          7459 => x"25",
          7460 => x"20",
          7461 => x"00",
          7462 => x"2a",
          7463 => x"31",
          7464 => x"32",
          7465 => x"61",
          7466 => x"2c",
          7467 => x"32",
          7468 => x"73",
          7469 => x"4f",
          7470 => x"42",
          7471 => x"72",
          7472 => x"20",
          7473 => x"20",
          7474 => x"0a",
          7475 => x"41",
          7476 => x"65",
          7477 => x"20",
          7478 => x"20",
          7479 => x"0a",
          7480 => x"49",
          7481 => x"74",
          7482 => x"72",
          7483 => x"31",
          7484 => x"65",
          7485 => x"55",
          7486 => x"20",
          7487 => x"70",
          7488 => x"30",
          7489 => x"65",
          7490 => x"55",
          7491 => x"20",
          7492 => x"70",
          7493 => x"4c",
          7494 => x"65",
          7495 => x"49",
          7496 => x"20",
          7497 => x"70",
          7498 => x"69",
          7499 => x"74",
          7500 => x"72",
          7501 => x"75",
          7502 => x"69",
          7503 => x"69",
          7504 => x"45",
          7505 => x"20",
          7506 => x"2e",
          7507 => x"65",
          7508 => x"00",
          7509 => x"7a",
          7510 => x"46",
          7511 => x"6f",
          7512 => x"6c",
          7513 => x"63",
          7514 => x"70",
          7515 => x"6e",
          7516 => x"61",
          7517 => x"2a",
          7518 => x"25",
          7519 => x"42",
          7520 => x"61",
          7521 => x"5a",
          7522 => x"25",
          7523 => x"73",
          7524 => x"43",
          7525 => x"6f",
          7526 => x"2e",
          7527 => x"61",
          7528 => x"70",
          7529 => x"6f",
          7530 => x"43",
          7531 => x"63",
          7532 => x"30",
          7533 => x"0a",
          7534 => x"20",
          7535 => x"64",
          7536 => x"25",
          7537 => x"45",
          7538 => x"67",
          7539 => x"20",
          7540 => x"2e",
          7541 => x"58",
          7542 => x"00",
          7543 => x"58",
          7544 => x"43",
          7545 => x"67",
          7546 => x"25",
          7547 => x"38",
          7548 => x"6c",
          7549 => x"0a",
          7550 => x"69",
          7551 => x"25",
          7552 => x"32",
          7553 => x"72",
          7554 => x"00",
          7555 => x"20",
          7556 => x"0a",
          7557 => x"65",
          7558 => x"25",
          7559 => x"4d",
          7560 => x"78",
          7561 => x"2c",
          7562 => x"20",
          7563 => x"20",
          7564 => x"2e",
          7565 => x"25",
          7566 => x"20",
          7567 => x"64",
          7568 => x"53",
          7569 => x"69",
          7570 => x"6e",
          7571 => x"76",
          7572 => x"70",
          7573 => x"64",
          7574 => x"65",
          7575 => x"20",
          7576 => x"52",
          7577 => x"63",
          7578 => x"72",
          7579 => x"30",
          7580 => x"20",
          7581 => x"4d",
          7582 => x"74",
          7583 => x"72",
          7584 => x"30",
          7585 => x"20",
          7586 => x"6b",
          7587 => x"41",
          7588 => x"20",
          7589 => x"30",
          7590 => x"4d",
          7591 => x"20",
          7592 => x"49",
          7593 => x"20",
          7594 => x"20",
          7595 => x"30",
          7596 => x"20",
          7597 => x"65",
          7598 => x"20",
          7599 => x"20",
          7600 => x"64",
          7601 => x"7a",
          7602 => x"57",
          7603 => x"20",
          7604 => x"6c",
          7605 => x"71",
          7606 => x"34",
          7607 => x"20",
          7608 => x"4d",
          7609 => x"46",
          7610 => x"20",
          7611 => x"64",
          7612 => x"7a",
          7613 => x"53",
          7614 => x"50",
          7615 => x"49",
          7616 => x"20",
          7617 => x"32",
          7618 => x"57",
          7619 => x"20",
          7620 => x"20",
          7621 => x"20",
          7622 => x"68",
          7623 => x"25",
          7624 => x"20",
          7625 => x"52",
          7626 => x"69",
          7627 => x"25",
          7628 => x"20",
          7629 => x"41",
          7630 => x"65",
          7631 => x"25",
          7632 => x"20",
          7633 => x"20",
          7634 => x"30",
          7635 => x"29",
          7636 => x"42",
          7637 => x"20",
          7638 => x"25",
          7639 => x"20",
          7640 => x"20",
          7641 => x"30",
          7642 => x"29",
          7643 => x"53",
          7644 => x"20",
          7645 => x"25",
          7646 => x"20",
          7647 => x"44",
          7648 => x"30",
          7649 => x"29",
          7650 => x"6f",
          7651 => x"6f",
          7652 => x"55",
          7653 => x"45",
          7654 => x"53",
          7655 => x"4d",
          7656 => x"46",
          7657 => x"45",
          7658 => x"01",
          7659 => x"00",
          7660 => x"00",
          7661 => x"01",
          7662 => x"00",
          7663 => x"00",
          7664 => x"01",
          7665 => x"00",
          7666 => x"00",
          7667 => x"01",
          7668 => x"00",
          7669 => x"00",
          7670 => x"01",
          7671 => x"00",
          7672 => x"00",
          7673 => x"01",
          7674 => x"00",
          7675 => x"00",
          7676 => x"04",
          7677 => x"00",
          7678 => x"00",
          7679 => x"03",
          7680 => x"00",
          7681 => x"00",
          7682 => x"04",
          7683 => x"00",
          7684 => x"00",
          7685 => x"03",
          7686 => x"00",
          7687 => x"00",
          7688 => x"03",
          7689 => x"00",
          7690 => x"00",
          7691 => x"1b",
          7692 => x"1b",
          7693 => x"1b",
          7694 => x"1b",
          7695 => x"1b",
          7696 => x"10",
          7697 => x"0d",
          7698 => x"08",
          7699 => x"05",
          7700 => x"03",
          7701 => x"01",
          7702 => x"6f",
          7703 => x"63",
          7704 => x"69",
          7705 => x"69",
          7706 => x"61",
          7707 => x"68",
          7708 => x"68",
          7709 => x"21",
          7710 => x"75",
          7711 => x"46",
          7712 => x"6f",
          7713 => x"74",
          7714 => x"6f",
          7715 => x"20",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"1b",
          7720 => x"1b",
          7721 => x"7e",
          7722 => x"7e",
          7723 => x"7e",
          7724 => x"7e",
          7725 => x"7e",
          7726 => x"7e",
          7727 => x"7e",
          7728 => x"7e",
          7729 => x"7e",
          7730 => x"7e",
          7731 => x"00",
          7732 => x"00",
          7733 => x"1b",
          7734 => x"1b",
          7735 => x"58",
          7736 => x"25",
          7737 => x"2c",
          7738 => x"00",
          7739 => x"2d",
          7740 => x"63",
          7741 => x"25",
          7742 => x"4b",
          7743 => x"25",
          7744 => x"25",
          7745 => x"52",
          7746 => x"72",
          7747 => x"72",
          7748 => x"30",
          7749 => x"00",
          7750 => x"30",
          7751 => x"00",
          7752 => x"30",
          7753 => x"4e",
          7754 => x"64",
          7755 => x"00",
          7756 => x"22",
          7757 => x"00",
          7758 => x"5b",
          7759 => x"46",
          7760 => x"eb",
          7761 => x"35",
          7762 => x"41",
          7763 => x"41",
          7764 => x"4e",
          7765 => x"20",
          7766 => x"20",
          7767 => x"00",
          7768 => x"00",
          7769 => x"09",
          7770 => x"1e",
          7771 => x"8e",
          7772 => x"49",
          7773 => x"99",
          7774 => x"9c",
          7775 => x"a5",
          7776 => x"ac",
          7777 => x"b4",
          7778 => x"bc",
          7779 => x"c4",
          7780 => x"cc",
          7781 => x"d4",
          7782 => x"dc",
          7783 => x"e4",
          7784 => x"ec",
          7785 => x"f4",
          7786 => x"fc",
          7787 => x"3d",
          7788 => x"3c",
          7789 => x"00",
          7790 => x"01",
          7791 => x"00",
          7792 => x"00",
          7793 => x"00",
          7794 => x"00",
          7795 => x"00",
          7796 => x"00",
          7797 => x"00",
          7798 => x"00",
          7799 => x"00",
          7800 => x"00",
          7801 => x"00",
          7802 => x"00",
          7803 => x"00",
          7804 => x"00",
          7805 => x"25",
          7806 => x"25",
          7807 => x"25",
          7808 => x"25",
          7809 => x"25",
          7810 => x"25",
          7811 => x"25",
          7812 => x"25",
          7813 => x"25",
          7814 => x"25",
          7815 => x"25",
          7816 => x"25",
          7817 => x"03",
          7818 => x"03",
          7819 => x"03",
          7820 => x"22",
          7821 => x"22",
          7822 => x"23",
          7823 => x"00",
          7824 => x"20",
          7825 => x"00",
          7826 => x"00",
          7827 => x"01",
          7828 => x"01",
          7829 => x"01",
          7830 => x"00",
          7831 => x"01",
          7832 => x"01",
          7833 => x"01",
          7834 => x"01",
          7835 => x"01",
          7836 => x"01",
          7837 => x"01",
          7838 => x"01",
          7839 => x"01",
          7840 => x"01",
          7841 => x"01",
          7842 => x"01",
          7843 => x"01",
          7844 => x"01",
          7845 => x"01",
          7846 => x"01",
          7847 => x"01",
          7848 => x"01",
          7849 => x"01",
          7850 => x"01",
          7851 => x"01",
          7852 => x"01",
          7853 => x"02",
          7854 => x"2c",
          7855 => x"2c",
          7856 => x"02",
          7857 => x"00",
          7858 => x"01",
          7859 => x"02",
          7860 => x"02",
          7861 => x"02",
          7862 => x"02",
          7863 => x"02",
          7864 => x"02",
          7865 => x"01",
          7866 => x"02",
          7867 => x"02",
          7868 => x"02",
          7869 => x"02",
          7870 => x"02",
          7871 => x"01",
          7872 => x"02",
          7873 => x"01",
          7874 => x"03",
          7875 => x"03",
          7876 => x"03",
          7877 => x"03",
          7878 => x"03",
          7879 => x"03",
          7880 => x"00",
          7881 => x"03",
          7882 => x"03",
          7883 => x"03",
          7884 => x"01",
          7885 => x"01",
          7886 => x"04",
          7887 => x"00",
          7888 => x"2c",
          7889 => x"01",
          7890 => x"06",
          7891 => x"06",
          7892 => x"00",
          7893 => x"1f",
          7894 => x"1f",
          7895 => x"1f",
          7896 => x"1f",
          7897 => x"1f",
          7898 => x"1f",
          7899 => x"1f",
          7900 => x"1f",
          7901 => x"1f",
          7902 => x"1f",
          7903 => x"06",
          7904 => x"1f",
          7905 => x"00",
          7906 => x"21",
          7907 => x"05",
          7908 => x"01",
          7909 => x"01",
          7910 => x"08",
          7911 => x"00",
          7912 => x"01",
          7913 => x"00",
          7914 => x"01",
          7915 => x"00",
          7916 => x"01",
          7917 => x"00",
          7918 => x"01",
          7919 => x"00",
          7920 => x"01",
          7921 => x"00",
          7922 => x"01",
          7923 => x"00",
          7924 => x"01",
          7925 => x"00",
          7926 => x"01",
          7927 => x"00",
          7928 => x"01",
          7929 => x"00",
          7930 => x"01",
          7931 => x"00",
          7932 => x"01",
          7933 => x"00",
          7934 => x"01",
          7935 => x"00",
          7936 => x"01",
          7937 => x"00",
          7938 => x"01",
          7939 => x"00",
          7940 => x"01",
          7941 => x"00",
          7942 => x"01",
          7943 => x"00",
          7944 => x"01",
          7945 => x"00",
          7946 => x"01",
          7947 => x"00",
          7948 => x"01",
          7949 => x"00",
          7950 => x"01",
          7951 => x"00",
          7952 => x"01",
          7953 => x"00",
          7954 => x"01",
          7955 => x"00",
          7956 => x"01",
          7957 => x"00",
          7958 => x"01",
          7959 => x"00",
          7960 => x"01",
          7961 => x"00",
          7962 => x"01",
          7963 => x"00",
          7964 => x"01",
          7965 => x"00",
          7966 => x"01",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"01",
          7973 => x"00",
          7974 => x"00",
          7975 => x"05",
          7976 => x"05",
          7977 => x"01",
          7978 => x"01",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"00",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"f0",
          7996 => x"5d",
          7997 => x"75",
          7998 => x"6d",
          7999 => x"65",
          8000 => x"35",
          8001 => x"30",
          8002 => x"f1",
          8003 => x"f0",
          8004 => x"84",
          8005 => x"f0",
          8006 => x"5d",
          8007 => x"55",
          8008 => x"4d",
          8009 => x"45",
          8010 => x"35",
          8011 => x"30",
          8012 => x"f1",
          8013 => x"f0",
          8014 => x"84",
          8015 => x"f0",
          8016 => x"7d",
          8017 => x"55",
          8018 => x"4d",
          8019 => x"45",
          8020 => x"25",
          8021 => x"20",
          8022 => x"f9",
          8023 => x"f0",
          8024 => x"89",
          8025 => x"f0",
          8026 => x"1d",
          8027 => x"15",
          8028 => x"0d",
          8029 => x"05",
          8030 => x"f0",
          8031 => x"f0",
          8032 => x"f0",
          8033 => x"f0",
          8034 => x"84",
          8035 => x"f0",
          8036 => x"b7",
          8037 => x"39",
          8038 => x"1d",
          8039 => x"74",
          8040 => x"7a",
          8041 => x"9d",
          8042 => x"c3",
          8043 => x"f0",
          8044 => x"84",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"f8",
          8059 => x"f3",
          8060 => x"f4",
          8061 => x"f1",
          8062 => x"f2",
          8063 => x"80",
          8064 => x"81",
          8065 => x"82",
          8066 => x"83",
          8067 => x"84",
          8068 => x"85",
          8069 => x"86",
          8070 => x"87",
          8071 => x"88",
          8072 => x"89",
          8073 => x"f6",
          8074 => x"7f",
          8075 => x"f9",
          8076 => x"e0",
          8077 => x"e1",
          8078 => x"71",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"50",
          9080 => x"cc",
          9081 => x"f8",
          9082 => x"e1",
          9083 => x"e3",
          9084 => x"00",
          9085 => x"68",
          9086 => x"20",
          9087 => x"28",
          9088 => x"55",
          9089 => x"08",
          9090 => x"10",
          9091 => x"18",
          9092 => x"c7",
          9093 => x"88",
          9094 => x"90",
          9095 => x"98",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"01",
        others => X"00"
    );

    signal RAM0_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM1_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM2_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM3_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM4_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM5_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM6_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM7_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM0_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM1_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM2_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM3_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM4_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM5_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM6_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM7_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal lowDataA          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataA         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.
    signal lowDataB          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataB         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.

begin

    -- Correctly assign the Little Endian value to the correct array, byte writes the data is in '7 downto 0', h-word writes
    -- the data is in '15 downto 0', word writes the data is in '31 downto 0'. Long words (64bits) are treated as two words for Endianness,
    -- and not as one continuous long word, this is because the ZPU is 32bit even when accessing a 64bit chunk.
    --
    RAM0_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '0'
                 else (others => '0');
    RAM1_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '0' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM4_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '1'
                 else (others => '0');
    RAM5_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM6_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM7_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '1' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "011") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "010") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "001") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "000") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM4_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "111") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM5_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "110") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM6_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "101") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';
    RAM7_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "100") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';

    memARead  <= lowDataA  when memAAddr(2) = '0'
                 else
                 highDataA;
    memBRead  <= lowDataB & highDataB;

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM0_DATA;
            else
                lowDataA(7 downto 0)    <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM1_DATA;
            else
                lowDataA(15 downto 8)   <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM2_DATA;
            else
                lowDataA(23 downto 16)  <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM3_DATA;
            else
                lowDataA(31 downto 24)  <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 4 - Port A - bits 39 to 32 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM4_WREN = '1' then
                RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM4_DATA;
            else
                highDataA(7 downto 0)   <= RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 5 - Port A - bits 47 to 40 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM5_WREN = '1' then
                RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM5_DATA;
            else
                highDataA(15 downto 8)  <= RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 6 - Port A - bits 56 to 48
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM6_WREN = '1' then
                RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM6_DATA;
            else
                highDataA(23 downto 16) <= RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 7 - Port A - bits 63 to 57 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM7_WREN = '1' then
                RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM7_DATA;
            else
                highDataA(31 downto 24) <= RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;


    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(7 downto 0);
                lowDataB(7 downto 0)    <= memBWrite(7 downto 0);
            else
                lowDataB(7 downto 0)    <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(15 downto 8);
                lowDataB(15 downto 8)    <= memBWrite(15 downto 8);
            else
                lowDataB(15 downto 8)    <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(23 downto 16);
                lowDataB(23 downto 16)  <= memBWrite(23 downto 16);
            else
                lowDataB(23 downto 16)  <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(31 downto 24);
                lowDataB(31 downto 24)  <= memBWrite(31 downto 24);
            else
                lowDataB(31 downto 24)  <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 4 - Port B - bits 39 downto 32
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(39 downto 32);
                highDataB(7 downto 0)   <= memBWrite(39 downto 32);
            else
                highDataB(7 downto 0)   <= RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 5 - Port B - bits 47 downto 40
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(47 downto 40);
                highDataB(15 downto 8)  <= memBWrite(47 downto 40);
            else
                highDataB(15 downto 8)  <= RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 6 - Port B - bits 55 downto 48
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(55 downto 48);
                highDataB(23 downto 16)  <= memBWrite(55 downto 48);
            else
                highDataB(23 downto 16)  <= RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 7 - Port B - bits 63 downto 56 
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(63 downto 56);
                highDataB(31 downto 24)  <= memBWrite(63 downto 56);
            else
                highDataB(31 downto 24)  <= RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

end arch;
