-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b93",
             1 => x"8c040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b92",
            73 => x"f0040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b92d3",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b81e1",
           162 => x"b0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"92d80400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b94",
           171 => x"912d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b95",
           179 => x"fd2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"94040b0b",
           269 => x"0b8ca304",
           270 => x"0b0b0b8c",
           271 => x"b2040b0b",
           272 => x"0b8cc104",
           273 => x"0b0b0b8c",
           274 => x"d0040b0b",
           275 => x"0b8cdf04",
           276 => x"0b0b0b8c",
           277 => x"ee040b0b",
           278 => x"0b8cfd04",
           279 => x"0b0b0b8d",
           280 => x"8c040b0b",
           281 => x"0b8d9b04",
           282 => x"0b0b0b8d",
           283 => x"aa040b0b",
           284 => x"0b8db904",
           285 => x"0b0b0b8d",
           286 => x"c8040b0b",
           287 => x"0b8dd704",
           288 => x"0b0b0b8d",
           289 => x"e6040b0b",
           290 => x"0b8df504",
           291 => x"0b0b0b8e",
           292 => x"84040b0b",
           293 => x"0b8e9304",
           294 => x"0b0b0b8e",
           295 => x"a3040b0b",
           296 => x"0b8eb304",
           297 => x"0b0b0b8e",
           298 => x"c3040b0b",
           299 => x"0b8ed304",
           300 => x"0b0b0b8e",
           301 => x"e3040b0b",
           302 => x"0b8ef304",
           303 => x"0b0b0b8f",
           304 => x"83040b0b",
           305 => x"0b8f9304",
           306 => x"0b0b0b8f",
           307 => x"a3040b0b",
           308 => x"0b8fb304",
           309 => x"0b0b0b8f",
           310 => x"c3040b0b",
           311 => x"0b8fd304",
           312 => x"0b0b0b8f",
           313 => x"e3040b0b",
           314 => x"0b8ff304",
           315 => x"0b0b0b90",
           316 => x"83040b0b",
           317 => x"0b909304",
           318 => x"0b0b0b90",
           319 => x"a3040b0b",
           320 => x"0b90b304",
           321 => x"0b0b0b90",
           322 => x"c3040b0b",
           323 => x"0b90d304",
           324 => x"0b0b0b90",
           325 => x"e3040b0b",
           326 => x"0b90f304",
           327 => x"0b0b0b91",
           328 => x"83040b0b",
           329 => x"0b919304",
           330 => x"0b0b0b91",
           331 => x"a3040b0b",
           332 => x"0b91b304",
           333 => x"0b0b0b91",
           334 => x"c3040b0b",
           335 => x"0b91d304",
           336 => x"0b0b0b91",
           337 => x"e3040b0b",
           338 => x"0b91f304",
           339 => x"0b0b0b92",
           340 => x"82040b0b",
           341 => x"0b929104",
           342 => x"0b0b0b92",
           343 => x"a004ffff",
           344 => x"ffffffff",
           345 => x"ffffffff",
           346 => x"ffffffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0481fefc",
           386 => x"0ca3ff2d",
           387 => x"81fefc08",
           388 => x"83809004",
           389 => x"81fefc0c",
           390 => x"b5c82d81",
           391 => x"fefc0883",
           392 => x"80900481",
           393 => x"fefc0cb6",
           394 => x"872d81fe",
           395 => x"fc088380",
           396 => x"900481fe",
           397 => x"fc0cb6a5",
           398 => x"2d81fefc",
           399 => x"08838090",
           400 => x"0481fefc",
           401 => x"0cbce32d",
           402 => x"81fefc08",
           403 => x"83809004",
           404 => x"81fefc0c",
           405 => x"bde12d81",
           406 => x"fefc0883",
           407 => x"80900481",
           408 => x"fefc0cb6",
           409 => x"c82d81fe",
           410 => x"fc088380",
           411 => x"900481fe",
           412 => x"fc0cbdfe",
           413 => x"2d81fefc",
           414 => x"08838090",
           415 => x"0481fefc",
           416 => x"0cbff02d",
           417 => x"81fefc08",
           418 => x"83809004",
           419 => x"81fefc0c",
           420 => x"bc892d81",
           421 => x"fefc0883",
           422 => x"80900481",
           423 => x"fefc0cb6",
           424 => x"fa2d81fe",
           425 => x"fc088380",
           426 => x"900481fe",
           427 => x"fc0cbc9f",
           428 => x"2d81fefc",
           429 => x"08838090",
           430 => x"0481fefc",
           431 => x"0cbcc32d",
           432 => x"81fefc08",
           433 => x"83809004",
           434 => x"81fefc0c",
           435 => x"a68c2d81",
           436 => x"fefc0883",
           437 => x"80900481",
           438 => x"fefc0ca6",
           439 => x"dd2d81fe",
           440 => x"fc088380",
           441 => x"900481fe",
           442 => x"fc0c9ef9",
           443 => x"2d81fefc",
           444 => x"08838090",
           445 => x"0481fefc",
           446 => x"0ca0ae2d",
           447 => x"81fefc08",
           448 => x"83809004",
           449 => x"81fefc0c",
           450 => x"a1e12d81",
           451 => x"fefc0883",
           452 => x"80900481",
           453 => x"fefc0c81",
           454 => x"84c32d81",
           455 => x"fefc0883",
           456 => x"80900481",
           457 => x"fefc0c81",
           458 => x"91b42d81",
           459 => x"fefc0883",
           460 => x"80900481",
           461 => x"fefc0c81",
           462 => x"89a82d81",
           463 => x"fefc0883",
           464 => x"80900481",
           465 => x"fefc0c81",
           466 => x"8ca52d81",
           467 => x"fefc0883",
           468 => x"80900481",
           469 => x"fefc0c81",
           470 => x"96c32d81",
           471 => x"fefc0883",
           472 => x"80900481",
           473 => x"fefc0c81",
           474 => x"9fa32d81",
           475 => x"fefc0883",
           476 => x"80900481",
           477 => x"fefc0c81",
           478 => x"90962d81",
           479 => x"fefc0883",
           480 => x"80900481",
           481 => x"fefc0c81",
           482 => x"99e22d81",
           483 => x"fefc0883",
           484 => x"80900481",
           485 => x"fefc0c81",
           486 => x"9b812d81",
           487 => x"fefc0883",
           488 => x"80900481",
           489 => x"fefc0c81",
           490 => x"9ba02d81",
           491 => x"fefc0883",
           492 => x"80900481",
           493 => x"fefc0c81",
           494 => x"a38a2d81",
           495 => x"fefc0883",
           496 => x"80900481",
           497 => x"fefc0c81",
           498 => x"a0f02d81",
           499 => x"fefc0883",
           500 => x"80900481",
           501 => x"fefc0c81",
           502 => x"a5de2d81",
           503 => x"fefc0883",
           504 => x"80900481",
           505 => x"fefc0c81",
           506 => x"9ca42d81",
           507 => x"fefc0883",
           508 => x"80900481",
           509 => x"fefc0c81",
           510 => x"a8de2d81",
           511 => x"fefc0883",
           512 => x"80900481",
           513 => x"fefc0c81",
           514 => x"a9df2d81",
           515 => x"fefc0883",
           516 => x"80900481",
           517 => x"fefc0c81",
           518 => x"92942d81",
           519 => x"fefc0883",
           520 => x"80900481",
           521 => x"fefc0c81",
           522 => x"91ed2d81",
           523 => x"fefc0883",
           524 => x"80900481",
           525 => x"fefc0c81",
           526 => x"93982d81",
           527 => x"fefc0883",
           528 => x"80900481",
           529 => x"fefc0c81",
           530 => x"9cfb2d81",
           531 => x"fefc0883",
           532 => x"80900481",
           533 => x"fefc0c81",
           534 => x"aad02d81",
           535 => x"fefc0883",
           536 => x"80900481",
           537 => x"fefc0c81",
           538 => x"acda2d81",
           539 => x"fefc0883",
           540 => x"80900481",
           541 => x"fefc0c81",
           542 => x"b09c2d81",
           543 => x"fefc0883",
           544 => x"80900481",
           545 => x"fefc0c81",
           546 => x"83e22d81",
           547 => x"fefc0883",
           548 => x"80900481",
           549 => x"fefc0c81",
           550 => x"b3882d81",
           551 => x"fefc0883",
           552 => x"80900481",
           553 => x"fefc0c81",
           554 => x"c1bd2d81",
           555 => x"fefc0883",
           556 => x"80900481",
           557 => x"fefc0c81",
           558 => x"bfa92d81",
           559 => x"fefc0883",
           560 => x"80900481",
           561 => x"fefc0c80",
           562 => x"d59d2d81",
           563 => x"fefc0883",
           564 => x"80900481",
           565 => x"fefc0c80",
           566 => x"d7872d81",
           567 => x"fefc0883",
           568 => x"80900481",
           569 => x"fefc0c80",
           570 => x"d8eb2d81",
           571 => x"fefc0883",
           572 => x"80900481",
           573 => x"fefc0c9f",
           574 => x"a22d81fe",
           575 => x"fc088380",
           576 => x"900481fe",
           577 => x"fc0ca084",
           578 => x"2d81fefc",
           579 => x"08838090",
           580 => x"0481fefc",
           581 => x"0ca2f12d",
           582 => x"81fefc08",
           583 => x"83809004",
           584 => x"81fefc0c",
           585 => x"81c2d82d",
           586 => x"81fefc08",
           587 => x"83809004",
           588 => x"3c040000",
           589 => x"10101010",
           590 => x"10101010",
           591 => x"10101010",
           592 => x"10101010",
           593 => x"10101010",
           594 => x"10101010",
           595 => x"10101010",
           596 => x"10101053",
           597 => x"51040000",
           598 => x"7381ff06",
           599 => x"73830609",
           600 => x"81058305",
           601 => x"1010102b",
           602 => x"0772fc06",
           603 => x"0c515104",
           604 => x"72728072",
           605 => x"8106ff05",
           606 => x"09720605",
           607 => x"71105272",
           608 => x"0a100a53",
           609 => x"72ed3851",
           610 => x"51535104",
           611 => x"81fef070",
           612 => x"8296b027",
           613 => x"8e388071",
           614 => x"70840553",
           615 => x"0c0b0b0b",
           616 => x"938f048c",
           617 => x"815181e0",
           618 => x"80040081",
           619 => x"fefc0802",
           620 => x"81fefc0c",
           621 => x"fd3d0d80",
           622 => x"5381fefc",
           623 => x"088c0508",
           624 => x"5281fefc",
           625 => x"08880508",
           626 => x"5183d43f",
           627 => x"81fef008",
           628 => x"7081fef0",
           629 => x"0c54853d",
           630 => x"0d81fefc",
           631 => x"0c0481fe",
           632 => x"fc080281",
           633 => x"fefc0cfd",
           634 => x"3d0d8153",
           635 => x"81fefc08",
           636 => x"8c050852",
           637 => x"81fefc08",
           638 => x"88050851",
           639 => x"83a13f81",
           640 => x"fef00870",
           641 => x"81fef00c",
           642 => x"54853d0d",
           643 => x"81fefc0c",
           644 => x"0481fefc",
           645 => x"080281fe",
           646 => x"fc0cf93d",
           647 => x"0d800b81",
           648 => x"fefc08fc",
           649 => x"050c81fe",
           650 => x"fc088805",
           651 => x"088025b9",
           652 => x"3881fefc",
           653 => x"08880508",
           654 => x"3081fefc",
           655 => x"0888050c",
           656 => x"800b81fe",
           657 => x"fc08f405",
           658 => x"0c81fefc",
           659 => x"08fc0508",
           660 => x"8a38810b",
           661 => x"81fefc08",
           662 => x"f4050c81",
           663 => x"fefc08f4",
           664 => x"050881fe",
           665 => x"fc08fc05",
           666 => x"0c81fefc",
           667 => x"088c0508",
           668 => x"8025b938",
           669 => x"81fefc08",
           670 => x"8c050830",
           671 => x"81fefc08",
           672 => x"8c050c80",
           673 => x"0b81fefc",
           674 => x"08f0050c",
           675 => x"81fefc08",
           676 => x"fc05088a",
           677 => x"38810b81",
           678 => x"fefc08f0",
           679 => x"050c81fe",
           680 => x"fc08f005",
           681 => x"0881fefc",
           682 => x"08fc050c",
           683 => x"805381fe",
           684 => x"fc088c05",
           685 => x"085281fe",
           686 => x"fc088805",
           687 => x"085181df",
           688 => x"3f81fef0",
           689 => x"087081fe",
           690 => x"fc08f805",
           691 => x"0c5481fe",
           692 => x"fc08fc05",
           693 => x"08802e90",
           694 => x"3881fefc",
           695 => x"08f80508",
           696 => x"3081fefc",
           697 => x"08f8050c",
           698 => x"81fefc08",
           699 => x"f8050870",
           700 => x"81fef00c",
           701 => x"54893d0d",
           702 => x"81fefc0c",
           703 => x"0481fefc",
           704 => x"080281fe",
           705 => x"fc0cfb3d",
           706 => x"0d800b81",
           707 => x"fefc08fc",
           708 => x"050c81fe",
           709 => x"fc088805",
           710 => x"08802599",
           711 => x"3881fefc",
           712 => x"08880508",
           713 => x"3081fefc",
           714 => x"0888050c",
           715 => x"810b81fe",
           716 => x"fc08fc05",
           717 => x"0c81fefc",
           718 => x"088c0508",
           719 => x"80259038",
           720 => x"81fefc08",
           721 => x"8c050830",
           722 => x"81fefc08",
           723 => x"8c050c81",
           724 => x"5381fefc",
           725 => x"088c0508",
           726 => x"5281fefc",
           727 => x"08880508",
           728 => x"51bd3f81",
           729 => x"fef00870",
           730 => x"81fefc08",
           731 => x"f8050c54",
           732 => x"81fefc08",
           733 => x"fc050880",
           734 => x"2e903881",
           735 => x"fefc08f8",
           736 => x"05083081",
           737 => x"fefc08f8",
           738 => x"050c81fe",
           739 => x"fc08f805",
           740 => x"087081fe",
           741 => x"f00c5487",
           742 => x"3d0d81fe",
           743 => x"fc0c0481",
           744 => x"fefc0802",
           745 => x"81fefc0c",
           746 => x"fd3d0d81",
           747 => x"0b81fefc",
           748 => x"08fc050c",
           749 => x"800b81fe",
           750 => x"fc08f805",
           751 => x"0c81fefc",
           752 => x"088c0508",
           753 => x"81fefc08",
           754 => x"88050827",
           755 => x"b93881fe",
           756 => x"fc08fc05",
           757 => x"08802eae",
           758 => x"38800b81",
           759 => x"fefc088c",
           760 => x"050824a2",
           761 => x"3881fefc",
           762 => x"088c0508",
           763 => x"1081fefc",
           764 => x"088c050c",
           765 => x"81fefc08",
           766 => x"fc050810",
           767 => x"81fefc08",
           768 => x"fc050cff",
           769 => x"b83981fe",
           770 => x"fc08fc05",
           771 => x"08802e80",
           772 => x"e13881fe",
           773 => x"fc088c05",
           774 => x"0881fefc",
           775 => x"08880508",
           776 => x"26ad3881",
           777 => x"fefc0888",
           778 => x"050881fe",
           779 => x"fc088c05",
           780 => x"083181fe",
           781 => x"fc088805",
           782 => x"0c81fefc",
           783 => x"08f80508",
           784 => x"81fefc08",
           785 => x"fc050807",
           786 => x"81fefc08",
           787 => x"f8050c81",
           788 => x"fefc08fc",
           789 => x"0508812a",
           790 => x"81fefc08",
           791 => x"fc050c81",
           792 => x"fefc088c",
           793 => x"0508812a",
           794 => x"81fefc08",
           795 => x"8c050cff",
           796 => x"953981fe",
           797 => x"fc089005",
           798 => x"08802e93",
           799 => x"3881fefc",
           800 => x"08880508",
           801 => x"7081fefc",
           802 => x"08f4050c",
           803 => x"51913981",
           804 => x"fefc08f8",
           805 => x"05087081",
           806 => x"fefc08f4",
           807 => x"050c5181",
           808 => x"fefc08f4",
           809 => x"050881fe",
           810 => x"f00c853d",
           811 => x"0d81fefc",
           812 => x"0c04fc3d",
           813 => x"0d767079",
           814 => x"7b555555",
           815 => x"558f7227",
           816 => x"8c387275",
           817 => x"07830651",
           818 => x"70802ea9",
           819 => x"38ff1252",
           820 => x"71ff2e98",
           821 => x"38727081",
           822 => x"05543374",
           823 => x"70810556",
           824 => x"34ff1252",
           825 => x"71ff2e09",
           826 => x"8106ea38",
           827 => x"7481fef0",
           828 => x"0c863d0d",
           829 => x"04745172",
           830 => x"70840554",
           831 => x"08717084",
           832 => x"05530c72",
           833 => x"70840554",
           834 => x"08717084",
           835 => x"05530c72",
           836 => x"70840554",
           837 => x"08717084",
           838 => x"05530c72",
           839 => x"70840554",
           840 => x"08717084",
           841 => x"05530cf0",
           842 => x"1252718f",
           843 => x"26c93883",
           844 => x"72279538",
           845 => x"72708405",
           846 => x"54087170",
           847 => x"8405530c",
           848 => x"fc125271",
           849 => x"8326ed38",
           850 => x"7054ff81",
           851 => x"39fc3d0d",
           852 => x"76797102",
           853 => x"8c059f05",
           854 => x"33575553",
           855 => x"55837227",
           856 => x"8a387483",
           857 => x"06517080",
           858 => x"2ea438ff",
           859 => x"125271ff",
           860 => x"2e933873",
           861 => x"73708105",
           862 => x"5534ff12",
           863 => x"5271ff2e",
           864 => x"098106ef",
           865 => x"387481fe",
           866 => x"f00c863d",
           867 => x"0d047474",
           868 => x"882b7507",
           869 => x"7071902b",
           870 => x"07515451",
           871 => x"8f7227a5",
           872 => x"38727170",
           873 => x"8405530c",
           874 => x"72717084",
           875 => x"05530c72",
           876 => x"71708405",
           877 => x"530c7271",
           878 => x"70840553",
           879 => x"0cf01252",
           880 => x"718f26dd",
           881 => x"38837227",
           882 => x"90387271",
           883 => x"70840553",
           884 => x"0cfc1252",
           885 => x"718326f2",
           886 => x"387053ff",
           887 => x"8e39fc3d",
           888 => x"0d767079",
           889 => x"70730783",
           890 => x"06545454",
           891 => x"557080c3",
           892 => x"38717008",
           893 => x"700970f7",
           894 => x"fbfdff13",
           895 => x"0670f884",
           896 => x"82818006",
           897 => x"51515353",
           898 => x"5470a638",
           899 => x"84147274",
           900 => x"70840556",
           901 => x"0c700870",
           902 => x"0970f7fb",
           903 => x"fdff1306",
           904 => x"70f88482",
           905 => x"81800651",
           906 => x"51535354",
           907 => x"70802edc",
           908 => x"38735271",
           909 => x"70810553",
           910 => x"33517073",
           911 => x"70810555",
           912 => x"3470f038",
           913 => x"7481fef0",
           914 => x"0c863d0d",
           915 => x"04fd3d0d",
           916 => x"75707183",
           917 => x"06535552",
           918 => x"70b83871",
           919 => x"70087009",
           920 => x"f7fbfdff",
           921 => x"120670f8",
           922 => x"84828180",
           923 => x"06515152",
           924 => x"53709d38",
           925 => x"84137008",
           926 => x"7009f7fb",
           927 => x"fdff1206",
           928 => x"70f88482",
           929 => x"81800651",
           930 => x"51525370",
           931 => x"802ee538",
           932 => x"72527133",
           933 => x"5170802e",
           934 => x"8a388112",
           935 => x"70335252",
           936 => x"70f83871",
           937 => x"743181fe",
           938 => x"f00c853d",
           939 => x"0d04fa3d",
           940 => x"0d787a7c",
           941 => x"70545555",
           942 => x"5272802e",
           943 => x"80d93871",
           944 => x"74078306",
           945 => x"5170802e",
           946 => x"80d638ff",
           947 => x"135372ff",
           948 => x"2eb13871",
           949 => x"33743356",
           950 => x"5174712e",
           951 => x"098106a9",
           952 => x"3872802e",
           953 => x"81893870",
           954 => x"81ff0651",
           955 => x"70802e80",
           956 => x"fe388112",
           957 => x"8115ff15",
           958 => x"55555272",
           959 => x"ff2e0981",
           960 => x"06d13871",
           961 => x"33743356",
           962 => x"517081ff",
           963 => x"067581ff",
           964 => x"06717131",
           965 => x"51525270",
           966 => x"81fef00c",
           967 => x"883d0d04",
           968 => x"71745755",
           969 => x"83732788",
           970 => x"38710874",
           971 => x"082e8838",
           972 => x"74765552",
           973 => x"ff9539fc",
           974 => x"13537280",
           975 => x"2eb13874",
           976 => x"087009f7",
           977 => x"fbfdff12",
           978 => x"0670f884",
           979 => x"82818006",
           980 => x"51515170",
           981 => x"9a388415",
           982 => x"84175755",
           983 => x"837327d0",
           984 => x"38740876",
           985 => x"082ed038",
           986 => x"74765552",
           987 => x"fedd3980",
           988 => x"0b81fef0",
           989 => x"0c883d0d",
           990 => x"04fe3d0d",
           991 => x"80528353",
           992 => x"71882b52",
           993 => x"87863f81",
           994 => x"fef00881",
           995 => x"ff067207",
           996 => x"ff145452",
           997 => x"728025e8",
           998 => x"387181fe",
           999 => x"f00c843d",
          1000 => x"0d04fb3d",
          1001 => x"0d777008",
          1002 => x"70535356",
          1003 => x"71802e80",
          1004 => x"ca387133",
          1005 => x"5170a02e",
          1006 => x"09810686",
          1007 => x"38811252",
          1008 => x"f1397153",
          1009 => x"84398113",
          1010 => x"53807333",
          1011 => x"7081ff06",
          1012 => x"53555570",
          1013 => x"a02e8338",
          1014 => x"81557080",
          1015 => x"2e843874",
          1016 => x"e5387381",
          1017 => x"ff065170",
          1018 => x"a02e0981",
          1019 => x"06883880",
          1020 => x"73708105",
          1021 => x"55347276",
          1022 => x"0c715170",
          1023 => x"81fef00c",
          1024 => x"873d0d04",
          1025 => x"fc3d0d76",
          1026 => x"53720880",
          1027 => x"2e913886",
          1028 => x"3dfc0552",
          1029 => x"72519fd8",
          1030 => x"3f81fef0",
          1031 => x"08853880",
          1032 => x"53833974",
          1033 => x"537281fe",
          1034 => x"f00c863d",
          1035 => x"0d04fc3d",
          1036 => x"0d768211",
          1037 => x"33ff0552",
          1038 => x"53815270",
          1039 => x"8b268198",
          1040 => x"38831333",
          1041 => x"ff055182",
          1042 => x"52709e26",
          1043 => x"818a3884",
          1044 => x"13335183",
          1045 => x"52709726",
          1046 => x"80fe3885",
          1047 => x"13335184",
          1048 => x"5270bb26",
          1049 => x"80f23886",
          1050 => x"13335185",
          1051 => x"5270bb26",
          1052 => x"80e63888",
          1053 => x"13225586",
          1054 => x"527487e7",
          1055 => x"2680d938",
          1056 => x"8a132254",
          1057 => x"87527387",
          1058 => x"e72680cc",
          1059 => x"38810b87",
          1060 => x"c0989c0c",
          1061 => x"722287c0",
          1062 => x"98bc0c82",
          1063 => x"133387c0",
          1064 => x"98b80c83",
          1065 => x"133387c0",
          1066 => x"98b40c84",
          1067 => x"133387c0",
          1068 => x"98b00c85",
          1069 => x"133387c0",
          1070 => x"98ac0c86",
          1071 => x"133387c0",
          1072 => x"98a80c74",
          1073 => x"87c098a4",
          1074 => x"0c7387c0",
          1075 => x"98a00c80",
          1076 => x"0b87c098",
          1077 => x"9c0c8052",
          1078 => x"7181fef0",
          1079 => x"0c863d0d",
          1080 => x"04f33d0d",
          1081 => x"7f5b87c0",
          1082 => x"989c5d81",
          1083 => x"7d0c87c0",
          1084 => x"98bc085e",
          1085 => x"7d7b2387",
          1086 => x"c098b808",
          1087 => x"5a79821c",
          1088 => x"3487c098",
          1089 => x"b4085a79",
          1090 => x"831c3487",
          1091 => x"c098b008",
          1092 => x"5a79841c",
          1093 => x"3487c098",
          1094 => x"ac085a79",
          1095 => x"851c3487",
          1096 => x"c098a808",
          1097 => x"5a79861c",
          1098 => x"3487c098",
          1099 => x"a4085c7b",
          1100 => x"881c2387",
          1101 => x"c098a008",
          1102 => x"5a798a1c",
          1103 => x"23807d0c",
          1104 => x"7983ffff",
          1105 => x"06597b83",
          1106 => x"ffff0658",
          1107 => x"861b3357",
          1108 => x"851b3356",
          1109 => x"841b3355",
          1110 => x"831b3354",
          1111 => x"821b3353",
          1112 => x"7d83ffff",
          1113 => x"065281e2",
          1114 => x"d451999d",
          1115 => x"3f8f3d0d",
          1116 => x"04ff3d0d",
          1117 => x"028f0533",
          1118 => x"7030709f",
          1119 => x"2a515252",
          1120 => x"700b0b81",
          1121 => x"f9e83483",
          1122 => x"3d0d04fb",
          1123 => x"3d0d770b",
          1124 => x"0b81f9e8",
          1125 => x"337081ff",
          1126 => x"06575556",
          1127 => x"87c09484",
          1128 => x"5174802e",
          1129 => x"863887c0",
          1130 => x"94945170",
          1131 => x"0870962a",
          1132 => x"70810653",
          1133 => x"54527080",
          1134 => x"2e8c3871",
          1135 => x"912a7081",
          1136 => x"06515170",
          1137 => x"d7387281",
          1138 => x"32708106",
          1139 => x"51517080",
          1140 => x"2e8d3871",
          1141 => x"932a7081",
          1142 => x"06515170",
          1143 => x"ffbe3873",
          1144 => x"81ff0651",
          1145 => x"87c09480",
          1146 => x"5270802e",
          1147 => x"863887c0",
          1148 => x"94905275",
          1149 => x"720c7581",
          1150 => x"fef00c87",
          1151 => x"3d0d04fb",
          1152 => x"3d0d029f",
          1153 => x"05330b0b",
          1154 => x"81f9e833",
          1155 => x"7081ff06",
          1156 => x"57555687",
          1157 => x"c0948451",
          1158 => x"74802e86",
          1159 => x"3887c094",
          1160 => x"94517008",
          1161 => x"70962a70",
          1162 => x"81065354",
          1163 => x"5270802e",
          1164 => x"8c387191",
          1165 => x"2a708106",
          1166 => x"515170d7",
          1167 => x"38728132",
          1168 => x"70810651",
          1169 => x"5170802e",
          1170 => x"8d387193",
          1171 => x"2a708106",
          1172 => x"515170ff",
          1173 => x"be387381",
          1174 => x"ff065187",
          1175 => x"c0948052",
          1176 => x"70802e86",
          1177 => x"3887c094",
          1178 => x"90527572",
          1179 => x"0c873d0d",
          1180 => x"04f93d0d",
          1181 => x"79548074",
          1182 => x"337081ff",
          1183 => x"06535357",
          1184 => x"70772e80",
          1185 => x"fe387181",
          1186 => x"ff068115",
          1187 => x"0b0b81f9",
          1188 => x"e8337081",
          1189 => x"ff065957",
          1190 => x"555887c0",
          1191 => x"94845175",
          1192 => x"802e8638",
          1193 => x"87c09494",
          1194 => x"51700870",
          1195 => x"962a7081",
          1196 => x"06535452",
          1197 => x"70802e8c",
          1198 => x"3871912a",
          1199 => x"70810651",
          1200 => x"5170d738",
          1201 => x"72813270",
          1202 => x"81065151",
          1203 => x"70802e8d",
          1204 => x"3871932a",
          1205 => x"70810651",
          1206 => x"5170ffbe",
          1207 => x"387481ff",
          1208 => x"065187c0",
          1209 => x"94805270",
          1210 => x"802e8638",
          1211 => x"87c09490",
          1212 => x"5277720c",
          1213 => x"81177433",
          1214 => x"7081ff06",
          1215 => x"53535770",
          1216 => x"ff843876",
          1217 => x"81fef00c",
          1218 => x"893d0d04",
          1219 => x"fe3d0d0b",
          1220 => x"0b81f9e8",
          1221 => x"337081ff",
          1222 => x"06545287",
          1223 => x"c0948451",
          1224 => x"72802e86",
          1225 => x"3887c094",
          1226 => x"94517008",
          1227 => x"70822a70",
          1228 => x"81065151",
          1229 => x"5170802e",
          1230 => x"e2387181",
          1231 => x"ff065187",
          1232 => x"c0948052",
          1233 => x"70802e86",
          1234 => x"3887c094",
          1235 => x"90527108",
          1236 => x"7081ff06",
          1237 => x"81fef00c",
          1238 => x"51843d0d",
          1239 => x"04fe3d0d",
          1240 => x"0b0b81f9",
          1241 => x"e8337081",
          1242 => x"ff065253",
          1243 => x"87c09484",
          1244 => x"5270802e",
          1245 => x"863887c0",
          1246 => x"94945271",
          1247 => x"0870822a",
          1248 => x"70810651",
          1249 => x"5151ff52",
          1250 => x"70802ea0",
          1251 => x"387281ff",
          1252 => x"065187c0",
          1253 => x"94805270",
          1254 => x"802e8638",
          1255 => x"87c09490",
          1256 => x"52710870",
          1257 => x"982b7098",
          1258 => x"2c515351",
          1259 => x"7181fef0",
          1260 => x"0c843d0d",
          1261 => x"04ff3d0d",
          1262 => x"87c09e80",
          1263 => x"08709c2a",
          1264 => x"8a065151",
          1265 => x"70802e84",
          1266 => x"b43887c0",
          1267 => x"9ea40881",
          1268 => x"f9ec0c87",
          1269 => x"c09ea808",
          1270 => x"81f9f00c",
          1271 => x"87c09e94",
          1272 => x"0881f9f4",
          1273 => x"0c87c09e",
          1274 => x"980881f9",
          1275 => x"f80c87c0",
          1276 => x"9e9c0881",
          1277 => x"f9fc0c87",
          1278 => x"c09ea008",
          1279 => x"81fa800c",
          1280 => x"87c09eac",
          1281 => x"0881fa84",
          1282 => x"0c87c09e",
          1283 => x"b00881fa",
          1284 => x"880c87c0",
          1285 => x"9eb40881",
          1286 => x"fa8c0c87",
          1287 => x"c09eb808",
          1288 => x"81fa900c",
          1289 => x"87c09ebc",
          1290 => x"0881fa94",
          1291 => x"0c87c09e",
          1292 => x"c00881fa",
          1293 => x"980c87c0",
          1294 => x"9ec40881",
          1295 => x"fa9c0c87",
          1296 => x"c09e8008",
          1297 => x"517081fa",
          1298 => x"a02387c0",
          1299 => x"9e840881",
          1300 => x"faa40c87",
          1301 => x"c09e8808",
          1302 => x"81faa80c",
          1303 => x"87c09e8c",
          1304 => x"0881faac",
          1305 => x"0c810b81",
          1306 => x"fab03480",
          1307 => x"0b87c09e",
          1308 => x"90087084",
          1309 => x"800a0651",
          1310 => x"52527080",
          1311 => x"2e833881",
          1312 => x"527181fa",
          1313 => x"b134800b",
          1314 => x"87c09e90",
          1315 => x"08708880",
          1316 => x"0a065152",
          1317 => x"5270802e",
          1318 => x"83388152",
          1319 => x"7181fab2",
          1320 => x"34800b87",
          1321 => x"c09e9008",
          1322 => x"7090800a",
          1323 => x"06515252",
          1324 => x"70802e83",
          1325 => x"38815271",
          1326 => x"81fab334",
          1327 => x"800b87c0",
          1328 => x"9e900870",
          1329 => x"88808006",
          1330 => x"51525270",
          1331 => x"802e8338",
          1332 => x"81527181",
          1333 => x"fab43480",
          1334 => x"0b87c09e",
          1335 => x"900870a0",
          1336 => x"80800651",
          1337 => x"52527080",
          1338 => x"2e833881",
          1339 => x"527181fa",
          1340 => x"b534800b",
          1341 => x"87c09e90",
          1342 => x"08709080",
          1343 => x"80065152",
          1344 => x"5270802e",
          1345 => x"83388152",
          1346 => x"7181fab6",
          1347 => x"34800b87",
          1348 => x"c09e9008",
          1349 => x"70848080",
          1350 => x"06515252",
          1351 => x"70802e83",
          1352 => x"38815271",
          1353 => x"81fab734",
          1354 => x"800b87c0",
          1355 => x"9e900870",
          1356 => x"82808006",
          1357 => x"51525270",
          1358 => x"802e8338",
          1359 => x"81527181",
          1360 => x"fab83480",
          1361 => x"0b87c09e",
          1362 => x"90087081",
          1363 => x"80800651",
          1364 => x"52527080",
          1365 => x"2e833881",
          1366 => x"527181fa",
          1367 => x"b934800b",
          1368 => x"87c09e90",
          1369 => x"087080c0",
          1370 => x"80065152",
          1371 => x"5270802e",
          1372 => x"83388152",
          1373 => x"7181faba",
          1374 => x"34800b87",
          1375 => x"c09e9008",
          1376 => x"70a08006",
          1377 => x"51525270",
          1378 => x"802e8338",
          1379 => x"81527181",
          1380 => x"fabb3487",
          1381 => x"c09e9008",
          1382 => x"70988006",
          1383 => x"708a2a51",
          1384 => x"51517081",
          1385 => x"fabc3480",
          1386 => x"0b87c09e",
          1387 => x"90087084",
          1388 => x"80065152",
          1389 => x"5270802e",
          1390 => x"83388152",
          1391 => x"7181fabd",
          1392 => x"3487c09e",
          1393 => x"90087083",
          1394 => x"f0067084",
          1395 => x"2a515151",
          1396 => x"7081fabe",
          1397 => x"34800b87",
          1398 => x"c09e9008",
          1399 => x"70880651",
          1400 => x"52527080",
          1401 => x"2e833881",
          1402 => x"527181fa",
          1403 => x"bf3487c0",
          1404 => x"9e900870",
          1405 => x"87065151",
          1406 => x"7081fac0",
          1407 => x"34833d0d",
          1408 => x"04fb3d0d",
          1409 => x"81e2ec51",
          1410 => x"8a9b3f81",
          1411 => x"fab03354",
          1412 => x"73802e88",
          1413 => x"3881e380",
          1414 => x"518a8a3f",
          1415 => x"81e39451",
          1416 => x"8a833f81",
          1417 => x"fab23354",
          1418 => x"73802e93",
          1419 => x"3881fa8c",
          1420 => x"0881fa90",
          1421 => x"08115452",
          1422 => x"81e3ac51",
          1423 => x"8fcb3f81",
          1424 => x"fab73354",
          1425 => x"73802e93",
          1426 => x"3881fa84",
          1427 => x"0881fa88",
          1428 => x"08115452",
          1429 => x"81e3c851",
          1430 => x"8faf3f81",
          1431 => x"fab43354",
          1432 => x"73802e93",
          1433 => x"3881f9ec",
          1434 => x"0881f9f0",
          1435 => x"08115452",
          1436 => x"81e3e451",
          1437 => x"8f933f81",
          1438 => x"fab53354",
          1439 => x"73802e93",
          1440 => x"3881f9f4",
          1441 => x"0881f9f8",
          1442 => x"08115452",
          1443 => x"81e48051",
          1444 => x"8ef73f81",
          1445 => x"fab63354",
          1446 => x"73802e93",
          1447 => x"3881f9fc",
          1448 => x"0881fa80",
          1449 => x"08115452",
          1450 => x"81e49c51",
          1451 => x"8edb3f81",
          1452 => x"fabb3354",
          1453 => x"73802e8d",
          1454 => x"3881fabc",
          1455 => x"335281e4",
          1456 => x"b8518ec5",
          1457 => x"3f81fabf",
          1458 => x"33547380",
          1459 => x"2e8d3881",
          1460 => x"fac03352",
          1461 => x"81e4d851",
          1462 => x"8eaf3f81",
          1463 => x"fabd3354",
          1464 => x"73802e8d",
          1465 => x"3881fabe",
          1466 => x"335281e4",
          1467 => x"f8518e99",
          1468 => x"3f81fab1",
          1469 => x"33547380",
          1470 => x"2e883881",
          1471 => x"e5985188",
          1472 => x"a43f81fa",
          1473 => x"b3335473",
          1474 => x"802e8838",
          1475 => x"81e5ac51",
          1476 => x"88933f81",
          1477 => x"fab83354",
          1478 => x"73802e88",
          1479 => x"3881e5b8",
          1480 => x"5188823f",
          1481 => x"81fab933",
          1482 => x"5473802e",
          1483 => x"883881e5",
          1484 => x"c45187f1",
          1485 => x"3f81faba",
          1486 => x"33547380",
          1487 => x"2e883881",
          1488 => x"e5d05187",
          1489 => x"e03f81e5",
          1490 => x"dc5187d9",
          1491 => x"3f81fa94",
          1492 => x"085281e5",
          1493 => x"e8518db1",
          1494 => x"3f81fa98",
          1495 => x"085281e6",
          1496 => x"90518da5",
          1497 => x"3f81fa9c",
          1498 => x"085281e6",
          1499 => x"b8518d99",
          1500 => x"3f81e6e0",
          1501 => x"5187ae3f",
          1502 => x"81faa022",
          1503 => x"5281e6e8",
          1504 => x"518d863f",
          1505 => x"81faa408",
          1506 => x"56bd84c0",
          1507 => x"527551e4",
          1508 => x"9a3f81fe",
          1509 => x"f008bd84",
          1510 => x"c0297671",
          1511 => x"31545481",
          1512 => x"fef00852",
          1513 => x"81e79051",
          1514 => x"8cdf3f81",
          1515 => x"fab73354",
          1516 => x"73802ea8",
          1517 => x"3881faa8",
          1518 => x"0856bd84",
          1519 => x"c0527551",
          1520 => x"e3e93f81",
          1521 => x"fef008bd",
          1522 => x"84c02976",
          1523 => x"71315454",
          1524 => x"81fef008",
          1525 => x"5281e7bc",
          1526 => x"518cae3f",
          1527 => x"81fab233",
          1528 => x"5473802e",
          1529 => x"a83881fa",
          1530 => x"ac0856bd",
          1531 => x"84c05275",
          1532 => x"51e3b83f",
          1533 => x"81fef008",
          1534 => x"bd84c029",
          1535 => x"76713154",
          1536 => x"5481fef0",
          1537 => x"085281e7",
          1538 => x"e8518bfd",
          1539 => x"3f81f5e4",
          1540 => x"5186923f",
          1541 => x"873d0d04",
          1542 => x"fe3d0d02",
          1543 => x"920533ff",
          1544 => x"05527184",
          1545 => x"26aa3871",
          1546 => x"842981e1",
          1547 => x"c0055271",
          1548 => x"080481e8",
          1549 => x"94519d39",
          1550 => x"81e89c51",
          1551 => x"973981e8",
          1552 => x"a4519139",
          1553 => x"81e8ac51",
          1554 => x"8b3981e8",
          1555 => x"b0518539",
          1556 => x"81e8b851",
          1557 => x"85cf3f84",
          1558 => x"3d0d0471",
          1559 => x"88800c04",
          1560 => x"ff3d0d87",
          1561 => x"c0968470",
          1562 => x"08525280",
          1563 => x"720c7074",
          1564 => x"077081fa",
          1565 => x"c40c720c",
          1566 => x"833d0d04",
          1567 => x"ff3d0d87",
          1568 => x"c0968470",
          1569 => x"0881fac4",
          1570 => x"0c528072",
          1571 => x"0c730970",
          1572 => x"81fac408",
          1573 => x"067081fa",
          1574 => x"c40c730c",
          1575 => x"51833d0d",
          1576 => x"04800b87",
          1577 => x"c096840c",
          1578 => x"0481fac4",
          1579 => x"0887c096",
          1580 => x"840c04fe",
          1581 => x"3d0d81ff",
          1582 => x"80088938",
          1583 => x"8296b00b",
          1584 => x"81ff800c",
          1585 => x"81ff8008",
          1586 => x"75115252",
          1587 => x"ff537083",
          1588 => x"b7f82688",
          1589 => x"387081ff",
          1590 => x"800c7153",
          1591 => x"7281fef0",
          1592 => x"0c843d0d",
          1593 => x"04f93d0d",
          1594 => x"797b8412",
          1595 => x"08a01290",
          1596 => x"14089415",
          1597 => x"0890165e",
          1598 => x"5a585459",
          1599 => x"57537077",
          1600 => x"26ba3875",
          1601 => x"13881408",
          1602 => x"53518171",
          1603 => x"0c767631",
          1604 => x"84120c80",
          1605 => x"730c7584",
          1606 => x"140c728c",
          1607 => x"120c7188",
          1608 => x"120c708c",
          1609 => x"130c7088",
          1610 => x"140c7390",
          1611 => x"120c7494",
          1612 => x"120c7094",
          1613 => x"150c7090",
          1614 => x"160c8c39",
          1615 => x"80730c73",
          1616 => x"90160c74",
          1617 => x"94150c77",
          1618 => x"81fef00c",
          1619 => x"893d0d04",
          1620 => x"fc3d0d76",
          1621 => x"8c110888",
          1622 => x"12085653",
          1623 => x"53710881",
          1624 => x"2e098106",
          1625 => x"a3388412",
          1626 => x"08701352",
          1627 => x"5570732e",
          1628 => x"09810694",
          1629 => x"38841308",
          1630 => x"1584130c",
          1631 => x"7388130c",
          1632 => x"718c150c",
          1633 => x"71539f39",
          1634 => x"81730c81",
          1635 => x"fad80890",
          1636 => x"140c81fa",
          1637 => x"c80b9414",
          1638 => x"0c7281fa",
          1639 => x"d80c9013",
          1640 => x"08739412",
          1641 => x"0c517308",
          1642 => x"812e0981",
          1643 => x"06b33884",
          1644 => x"13087014",
          1645 => x"52527074",
          1646 => x"2e098106",
          1647 => x"a4388414",
          1648 => x"08128414",
          1649 => x"0c941408",
          1650 => x"90150870",
          1651 => x"90130c52",
          1652 => x"94120c8c",
          1653 => x"14088815",
          1654 => x"08708813",
          1655 => x"0c528c12",
          1656 => x"0c7281fe",
          1657 => x"f00c863d",
          1658 => x"0d04f93d",
          1659 => x"0d797055",
          1660 => x"5776802e",
          1661 => x"81b5389f",
          1662 => x"17f00681",
          1663 => x"fad80857",
          1664 => x"57750882",
          1665 => x"2e8f3884",
          1666 => x"16087727",
          1667 => x"80c73890",
          1668 => x"160856ed",
          1669 => x"3983ffff",
          1670 => x"17fc8080",
          1671 => x"06705258",
          1672 => x"fd913f81",
          1673 => x"fef00881",
          1674 => x"fef00830",
          1675 => x"7081fef0",
          1676 => x"08078025",
          1677 => x"81fef008",
          1678 => x"09703070",
          1679 => x"72078025",
          1680 => x"73075358",
          1681 => x"58515456",
          1682 => x"80547274",
          1683 => x"2e098106",
          1684 => x"80d93888",
          1685 => x"39765275",
          1686 => x"5180c839",
          1687 => x"810b81fe",
          1688 => x"f0080c77",
          1689 => x"81fef008",
          1690 => x"84050c81",
          1691 => x"fad40853",
          1692 => x"7208822e",
          1693 => x"8c387573",
          1694 => x"2687388c",
          1695 => x"130853f0",
          1696 => x"39881308",
          1697 => x"88170c72",
          1698 => x"8c170c75",
          1699 => x"88140c88",
          1700 => x"1608768c",
          1701 => x"120c5375",
          1702 => x"51fdb53f",
          1703 => x"765281fe",
          1704 => x"f00851fc",
          1705 => x"c03f81fe",
          1706 => x"f0085473",
          1707 => x"81fef00c",
          1708 => x"893d0d04",
          1709 => x"ff3d0d73",
          1710 => x"5271802e",
          1711 => x"8738f012",
          1712 => x"51fd8d3f",
          1713 => x"833d0d04",
          1714 => x"fe3d0d02",
          1715 => x"93053353",
          1716 => x"728a2e09",
          1717 => x"81068538",
          1718 => x"8d51ed3f",
          1719 => x"81ff8c08",
          1720 => x"5271802e",
          1721 => x"90387272",
          1722 => x"3481ff8c",
          1723 => x"08810581",
          1724 => x"ff8c0c8f",
          1725 => x"3981ff84",
          1726 => x"08527180",
          1727 => x"2e853872",
          1728 => x"51712d84",
          1729 => x"3d0d04fe",
          1730 => x"3d0d0297",
          1731 => x"053381ff",
          1732 => x"84087681",
          1733 => x"ff840c54",
          1734 => x"51ffad3f",
          1735 => x"7281ff84",
          1736 => x"0c843d0d",
          1737 => x"04fd3d0d",
          1738 => x"75547333",
          1739 => x"7081ff06",
          1740 => x"53537180",
          1741 => x"2e8e3872",
          1742 => x"81ff0651",
          1743 => x"811454ff",
          1744 => x"873fe739",
          1745 => x"853d0d04",
          1746 => x"fc3d0d77",
          1747 => x"81ff8408",
          1748 => x"7881ff84",
          1749 => x"0c565473",
          1750 => x"337081ff",
          1751 => x"06535371",
          1752 => x"802e8e38",
          1753 => x"7281ff06",
          1754 => x"51811454",
          1755 => x"feda3fe7",
          1756 => x"397481ff",
          1757 => x"840c863d",
          1758 => x"0d04ec3d",
          1759 => x"0d666859",
          1760 => x"59787081",
          1761 => x"055a3356",
          1762 => x"75802e84",
          1763 => x"f83875a5",
          1764 => x"2e098106",
          1765 => x"82de3880",
          1766 => x"707a7081",
          1767 => x"055c3358",
          1768 => x"5b5b75b0",
          1769 => x"2e098106",
          1770 => x"8538815a",
          1771 => x"8b3975ad",
          1772 => x"2e098106",
          1773 => x"8a38825a",
          1774 => x"78708105",
          1775 => x"5a335675",
          1776 => x"aa2e0981",
          1777 => x"06923877",
          1778 => x"84197108",
          1779 => x"7b708105",
          1780 => x"5d33595d",
          1781 => x"59539d39",
          1782 => x"d0165372",
          1783 => x"89269538",
          1784 => x"7a88297b",
          1785 => x"10057605",
          1786 => x"d0057970",
          1787 => x"81055b33",
          1788 => x"575be539",
          1789 => x"7580ec32",
          1790 => x"70307072",
          1791 => x"07802578",
          1792 => x"80cc3270",
          1793 => x"30707207",
          1794 => x"80257307",
          1795 => x"53545851",
          1796 => x"55537380",
          1797 => x"2e8c3879",
          1798 => x"84077970",
          1799 => x"81055b33",
          1800 => x"575a7580",
          1801 => x"2e83de38",
          1802 => x"755480e0",
          1803 => x"76278938",
          1804 => x"e0167081",
          1805 => x"ff065553",
          1806 => x"7380cf2e",
          1807 => x"81aa3873",
          1808 => x"80cf24a2",
          1809 => x"387380c3",
          1810 => x"2e818e38",
          1811 => x"7380c324",
          1812 => x"8b387380",
          1813 => x"c22e818c",
          1814 => x"38819939",
          1815 => x"7380c42e",
          1816 => x"818a3881",
          1817 => x"8f397380",
          1818 => x"d52e8180",
          1819 => x"387380d5",
          1820 => x"248a3873",
          1821 => x"80d32e8e",
          1822 => x"3880f939",
          1823 => x"7380d82e",
          1824 => x"80ee3880",
          1825 => x"ef397784",
          1826 => x"19710856",
          1827 => x"59538074",
          1828 => x"33545572",
          1829 => x"752e8d38",
          1830 => x"81157015",
          1831 => x"70335154",
          1832 => x"5572f538",
          1833 => x"79812a56",
          1834 => x"90397481",
          1835 => x"16565372",
          1836 => x"7b278f38",
          1837 => x"a051fc90",
          1838 => x"3f758106",
          1839 => x"5372802e",
          1840 => x"e9387351",
          1841 => x"fcdf3f74",
          1842 => x"81165653",
          1843 => x"727b27fd",
          1844 => x"b038a051",
          1845 => x"fbf23fef",
          1846 => x"39778419",
          1847 => x"83123353",
          1848 => x"59539339",
          1849 => x"825c9539",
          1850 => x"885c9139",
          1851 => x"8a5c8d39",
          1852 => x"905c8939",
          1853 => x"7551fbd0",
          1854 => x"3ffd8639",
          1855 => x"79822a70",
          1856 => x"81065153",
          1857 => x"72802e88",
          1858 => x"38778419",
          1859 => x"59538639",
          1860 => x"84187854",
          1861 => x"58720874",
          1862 => x"80c43270",
          1863 => x"30707207",
          1864 => x"80255155",
          1865 => x"55557480",
          1866 => x"258d3872",
          1867 => x"802e8838",
          1868 => x"74307a90",
          1869 => x"075b5580",
          1870 => x"0b8f3d5e",
          1871 => x"577b5274",
          1872 => x"51d99b3f",
          1873 => x"81fef008",
          1874 => x"81ff067c",
          1875 => x"53755254",
          1876 => x"d8d93f81",
          1877 => x"fef00855",
          1878 => x"89742792",
          1879 => x"38a71453",
          1880 => x"7580f82e",
          1881 => x"84388714",
          1882 => x"537281ff",
          1883 => x"0654b014",
          1884 => x"53727d70",
          1885 => x"81055f34",
          1886 => x"81177530",
          1887 => x"7077079f",
          1888 => x"2a515457",
          1889 => x"769f2685",
          1890 => x"3872ffb1",
          1891 => x"3879842a",
          1892 => x"70810651",
          1893 => x"5372802e",
          1894 => x"8e38963d",
          1895 => x"7705e005",
          1896 => x"53ad7334",
          1897 => x"81175776",
          1898 => x"7a810654",
          1899 => x"55b05472",
          1900 => x"8338a054",
          1901 => x"79812a70",
          1902 => x"81065456",
          1903 => x"729f3881",
          1904 => x"1755767b",
          1905 => x"27973873",
          1906 => x"51f9fd3f",
          1907 => x"75810653",
          1908 => x"728b3874",
          1909 => x"81165653",
          1910 => x"7a7326eb",
          1911 => x"38963d77",
          1912 => x"05e00553",
          1913 => x"ff17ff14",
          1914 => x"70335354",
          1915 => x"57f9d93f",
          1916 => x"76f23874",
          1917 => x"81165653",
          1918 => x"727b27fb",
          1919 => x"8438a051",
          1920 => x"f9c63fef",
          1921 => x"39963d0d",
          1922 => x"04fd3d0d",
          1923 => x"863d7070",
          1924 => x"84055208",
          1925 => x"55527351",
          1926 => x"fae03f85",
          1927 => x"3d0d04fe",
          1928 => x"3d0d7481",
          1929 => x"ff8c0c85",
          1930 => x"3d880552",
          1931 => x"7551faca",
          1932 => x"3f81ff8c",
          1933 => x"08538073",
          1934 => x"34800b81",
          1935 => x"ff8c0c84",
          1936 => x"3d0d04fd",
          1937 => x"3d0d81ff",
          1938 => x"84087681",
          1939 => x"ff840c87",
          1940 => x"3d880553",
          1941 => x"775253fa",
          1942 => x"a13f7281",
          1943 => x"ff840c85",
          1944 => x"3d0d04fb",
          1945 => x"3d0d7779",
          1946 => x"81ff8808",
          1947 => x"70565457",
          1948 => x"55805471",
          1949 => x"802e80e0",
          1950 => x"3881ff88",
          1951 => x"0852712d",
          1952 => x"81fef008",
          1953 => x"81ff0653",
          1954 => x"72802e80",
          1955 => x"cb38728d",
          1956 => x"2eb93872",
          1957 => x"88327030",
          1958 => x"70802551",
          1959 => x"51527380",
          1960 => x"2e8b3871",
          1961 => x"802e8638",
          1962 => x"ff145497",
          1963 => x"399f7325",
          1964 => x"c838ff16",
          1965 => x"52737225",
          1966 => x"c0387414",
          1967 => x"52727234",
          1968 => x"81145472",
          1969 => x"51f8813f",
          1970 => x"ffaf3973",
          1971 => x"15528072",
          1972 => x"348a51f7",
          1973 => x"f33f8153",
          1974 => x"7281fef0",
          1975 => x"0c873d0d",
          1976 => x"04fe3d0d",
          1977 => x"81ff8808",
          1978 => x"7581ff88",
          1979 => x"0c775376",
          1980 => x"5253feef",
          1981 => x"3f7281ff",
          1982 => x"880c843d",
          1983 => x"0d04f83d",
          1984 => x"0d7a7c5a",
          1985 => x"5680707a",
          1986 => x"0c587508",
          1987 => x"70335553",
          1988 => x"73a02e09",
          1989 => x"81068738",
          1990 => x"8113760c",
          1991 => x"ed3973ad",
          1992 => x"2e098106",
          1993 => x"8e388176",
          1994 => x"0811770c",
          1995 => x"76087033",
          1996 => x"56545873",
          1997 => x"b02e0981",
          1998 => x"0680c238",
          1999 => x"75088105",
          2000 => x"760c7508",
          2001 => x"70335553",
          2002 => x"7380e22e",
          2003 => x"8b389057",
          2004 => x"7380f82e",
          2005 => x"85388f39",
          2006 => x"82578113",
          2007 => x"760c7508",
          2008 => x"70335553",
          2009 => x"ac398155",
          2010 => x"a0742780",
          2011 => x"fa38d014",
          2012 => x"53805588",
          2013 => x"57897327",
          2014 => x"983880eb",
          2015 => x"39d01453",
          2016 => x"80557289",
          2017 => x"2680e038",
          2018 => x"86398055",
          2019 => x"80d9398a",
          2020 => x"578055a0",
          2021 => x"742780c2",
          2022 => x"3880e074",
          2023 => x"278938e0",
          2024 => x"147081ff",
          2025 => x"065553d0",
          2026 => x"147081ff",
          2027 => x"06555390",
          2028 => x"74278e38",
          2029 => x"f9147081",
          2030 => x"ff065553",
          2031 => x"897427ca",
          2032 => x"38737727",
          2033 => x"c5387477",
          2034 => x"29147608",
          2035 => x"8105770c",
          2036 => x"76087033",
          2037 => x"565455ff",
          2038 => x"ba397780",
          2039 => x"2e843874",
          2040 => x"30557479",
          2041 => x"0c815574",
          2042 => x"81fef00c",
          2043 => x"8a3d0d04",
          2044 => x"f83d0d7a",
          2045 => x"7c5a5680",
          2046 => x"707a0c58",
          2047 => x"75087033",
          2048 => x"555373a0",
          2049 => x"2e098106",
          2050 => x"87388113",
          2051 => x"760ced39",
          2052 => x"73ad2e09",
          2053 => x"81068e38",
          2054 => x"81760811",
          2055 => x"770c7608",
          2056 => x"70335654",
          2057 => x"5873b02e",
          2058 => x"09810680",
          2059 => x"c2387508",
          2060 => x"8105760c",
          2061 => x"75087033",
          2062 => x"55537380",
          2063 => x"e22e8b38",
          2064 => x"90577380",
          2065 => x"f82e8538",
          2066 => x"8f398257",
          2067 => x"8113760c",
          2068 => x"75087033",
          2069 => x"5553ac39",
          2070 => x"8155a074",
          2071 => x"2780fa38",
          2072 => x"d0145380",
          2073 => x"55885789",
          2074 => x"73279838",
          2075 => x"80eb39d0",
          2076 => x"14538055",
          2077 => x"72892680",
          2078 => x"e0388639",
          2079 => x"805580d9",
          2080 => x"398a5780",
          2081 => x"55a07427",
          2082 => x"80c23880",
          2083 => x"e0742789",
          2084 => x"38e01470",
          2085 => x"81ff0655",
          2086 => x"53d01470",
          2087 => x"81ff0655",
          2088 => x"53907427",
          2089 => x"8e38f914",
          2090 => x"7081ff06",
          2091 => x"55538974",
          2092 => x"27ca3873",
          2093 => x"7727c538",
          2094 => x"74772914",
          2095 => x"76088105",
          2096 => x"770c7608",
          2097 => x"70335654",
          2098 => x"55ffba39",
          2099 => x"77802e84",
          2100 => x"38743055",
          2101 => x"74790c81",
          2102 => x"557481fe",
          2103 => x"f00c8a3d",
          2104 => x"0d04fd3d",
          2105 => x"0d76982b",
          2106 => x"70982c79",
          2107 => x"982b7098",
          2108 => x"2c721013",
          2109 => x"70822b51",
          2110 => x"53515451",
          2111 => x"51800b81",
          2112 => x"e9cc1233",
          2113 => x"55537174",
          2114 => x"259c3881",
          2115 => x"e9c81108",
          2116 => x"12028405",
          2117 => x"97053371",
          2118 => x"33525252",
          2119 => x"70722e09",
          2120 => x"81068338",
          2121 => x"81537281",
          2122 => x"fef00c85",
          2123 => x"3d0d04fc",
          2124 => x"3d0d7802",
          2125 => x"84059f05",
          2126 => x"33713354",
          2127 => x"55537180",
          2128 => x"2e9f3888",
          2129 => x"51f3813f",
          2130 => x"a051f2fc",
          2131 => x"3f8851f2",
          2132 => x"f73f7233",
          2133 => x"ff055271",
          2134 => x"73347181",
          2135 => x"ff0652de",
          2136 => x"397651f3",
          2137 => x"c03f7373",
          2138 => x"34863d0d",
          2139 => x"04f63d0d",
          2140 => x"7c028405",
          2141 => x"b7053302",
          2142 => x"8805bb05",
          2143 => x"3381fbbc",
          2144 => x"33708429",
          2145 => x"81fae405",
          2146 => x"70085159",
          2147 => x"595a5859",
          2148 => x"74802e86",
          2149 => x"387451f2",
          2150 => x"9b3f81fb",
          2151 => x"bc337084",
          2152 => x"2981fae4",
          2153 => x"05811970",
          2154 => x"5458565a",
          2155 => x"f0bc3f81",
          2156 => x"fef00875",
          2157 => x"0c81fbbc",
          2158 => x"33708429",
          2159 => x"81fae405",
          2160 => x"70085156",
          2161 => x"5a74802e",
          2162 => x"a6387553",
          2163 => x"78527451",
          2164 => x"d5e03f81",
          2165 => x"fbbc3381",
          2166 => x"05557481",
          2167 => x"fbbc3474",
          2168 => x"81ff0655",
          2169 => x"93752787",
          2170 => x"38800b81",
          2171 => x"fbbc3477",
          2172 => x"802eb638",
          2173 => x"81fbb808",
          2174 => x"5675802e",
          2175 => x"ac3881fb",
          2176 => x"b4335574",
          2177 => x"a4388c3d",
          2178 => x"fc055476",
          2179 => x"53785275",
          2180 => x"5180c891",
          2181 => x"3f81fbb8",
          2182 => x"08528a51",
          2183 => x"80fd9e3f",
          2184 => x"81fbb808",
          2185 => x"5180cbee",
          2186 => x"3f8c3d0d",
          2187 => x"04dc3d0d",
          2188 => x"81578052",
          2189 => x"81fbb808",
          2190 => x"5180d287",
          2191 => x"3f81fef0",
          2192 => x"0880d138",
          2193 => x"81fbb808",
          2194 => x"5380f852",
          2195 => x"883d7052",
          2196 => x"5680fad5",
          2197 => x"3f81fef0",
          2198 => x"08802eb8",
          2199 => x"387551d7",
          2200 => x"ec3f81fe",
          2201 => x"f0085580",
          2202 => x"0b81fef0",
          2203 => x"08259c38",
          2204 => x"81fef008",
          2205 => x"ff057017",
          2206 => x"55558074",
          2207 => x"34755376",
          2208 => x"52811781",
          2209 => x"e8e05257",
          2210 => x"f6ff3f74",
          2211 => x"ff2e0981",
          2212 => x"06ffb138",
          2213 => x"a63d0d04",
          2214 => x"d93d0daa",
          2215 => x"3d08ad3d",
          2216 => x"085a5a81",
          2217 => x"70585880",
          2218 => x"5281fbb8",
          2219 => x"085180d1",
          2220 => x"923f81fe",
          2221 => x"f0088191",
          2222 => x"38ff0b81",
          2223 => x"fbb80854",
          2224 => x"5580f852",
          2225 => x"8b3d7052",
          2226 => x"5680f9dd",
          2227 => x"3f81fef0",
          2228 => x"08802ea4",
          2229 => x"387551d6",
          2230 => x"f43f81fe",
          2231 => x"f0088118",
          2232 => x"5855800b",
          2233 => x"81fef008",
          2234 => x"258e3881",
          2235 => x"fef008ff",
          2236 => x"05701755",
          2237 => x"55807434",
          2238 => x"74097030",
          2239 => x"7072079f",
          2240 => x"2a515555",
          2241 => x"78772e85",
          2242 => x"3873ffad",
          2243 => x"3881fbb8",
          2244 => x"088c1108",
          2245 => x"535180d0",
          2246 => x"aa3f81fe",
          2247 => x"f008802e",
          2248 => x"883881e8",
          2249 => x"ec51effd",
          2250 => x"3f78772e",
          2251 => x"09810699",
          2252 => x"38755279",
          2253 => x"51d5a73f",
          2254 => x"7951d691",
          2255 => x"3fab3d08",
          2256 => x"5481fef0",
          2257 => x"08743480",
          2258 => x"587781fe",
          2259 => x"f00ca93d",
          2260 => x"0d04f63d",
          2261 => x"0d7c7e71",
          2262 => x"5c717233",
          2263 => x"57595a58",
          2264 => x"73a02e09",
          2265 => x"8106a238",
          2266 => x"78337805",
          2267 => x"56777627",
          2268 => x"98388117",
          2269 => x"705b7071",
          2270 => x"33565855",
          2271 => x"73a02e09",
          2272 => x"81068638",
          2273 => x"757526ea",
          2274 => x"38805473",
          2275 => x"882981fb",
          2276 => x"c0057008",
          2277 => x"5255d5b5",
          2278 => x"3f81fef0",
          2279 => x"08537952",
          2280 => x"740851d6",
          2281 => x"893f81fe",
          2282 => x"f00880c4",
          2283 => x"38841533",
          2284 => x"5574812e",
          2285 => x"88387482",
          2286 => x"2e8838b4",
          2287 => x"39fcee3f",
          2288 => x"ab39811a",
          2289 => x"5a8c3dfc",
          2290 => x"1153f805",
          2291 => x"51f6af3f",
          2292 => x"81fef008",
          2293 => x"802e9938",
          2294 => x"7a537852",
          2295 => x"7751fdb8",
          2296 => x"3f81fef0",
          2297 => x"0881ff06",
          2298 => x"55748538",
          2299 => x"74549139",
          2300 => x"81147081",
          2301 => x"ff065154",
          2302 => x"827427ff",
          2303 => x"8e388054",
          2304 => x"7381fef0",
          2305 => x"0c8c3d0d",
          2306 => x"04d33d0d",
          2307 => x"b03d0802",
          2308 => x"840581c3",
          2309 => x"05335f5a",
          2310 => x"800baf3d",
          2311 => x"3481fbbc",
          2312 => x"335b81fb",
          2313 => x"b80881a3",
          2314 => x"3881fbb4",
          2315 => x"33547381",
          2316 => x"9a38a851",
          2317 => x"ebb43f81",
          2318 => x"fef00881",
          2319 => x"fbb80c81",
          2320 => x"fef00880",
          2321 => x"2e80fe38",
          2322 => x"935381fa",
          2323 => x"e0085281",
          2324 => x"fef00851",
          2325 => x"bbed3f81",
          2326 => x"fef00880",
          2327 => x"2e8b3881",
          2328 => x"e99851f3",
          2329 => x"a43f80e3",
          2330 => x"3981fbb8",
          2331 => x"085380f8",
          2332 => x"52903d70",
          2333 => x"525480f6",
          2334 => x"b03f81fe",
          2335 => x"f0085681",
          2336 => x"fef00874",
          2337 => x"2e098106",
          2338 => x"80c13881",
          2339 => x"fef00851",
          2340 => x"d3bb3f81",
          2341 => x"fef00855",
          2342 => x"800b81fe",
          2343 => x"f008259a",
          2344 => x"3881fef0",
          2345 => x"08ff0570",
          2346 => x"17555580",
          2347 => x"74348053",
          2348 => x"7481ff06",
          2349 => x"527551f9",
          2350 => x"b43f74ff",
          2351 => x"2e098106",
          2352 => x"ffa73887",
          2353 => x"39810b81",
          2354 => x"fbb4348f",
          2355 => x"3d5ddd8d",
          2356 => x"3f81fef0",
          2357 => x"08982b70",
          2358 => x"982c5159",
          2359 => x"78ff2eee",
          2360 => x"387881ff",
          2361 => x"0681ff94",
          2362 => x"3370982b",
          2363 => x"70982c81",
          2364 => x"ff903370",
          2365 => x"982b7097",
          2366 => x"2c71982c",
          2367 => x"05708429",
          2368 => x"81e9c805",
          2369 => x"70081570",
          2370 => x"33515151",
          2371 => x"51595951",
          2372 => x"595d5881",
          2373 => x"5673782e",
          2374 => x"80e93877",
          2375 => x"7427b438",
          2376 => x"7481800a",
          2377 => x"2981ff0a",
          2378 => x"0570982c",
          2379 => x"51558075",
          2380 => x"2480ce38",
          2381 => x"76537452",
          2382 => x"7751f7a6",
          2383 => x"3f81fef0",
          2384 => x"0881ff06",
          2385 => x"5473802e",
          2386 => x"d7387481",
          2387 => x"ff903481",
          2388 => x"56b13974",
          2389 => x"81800a29",
          2390 => x"81800a05",
          2391 => x"70982c70",
          2392 => x"81ff0656",
          2393 => x"5155738a",
          2394 => x"26973876",
          2395 => x"53745277",
          2396 => x"51f6ef3f",
          2397 => x"81fef008",
          2398 => x"81ff0654",
          2399 => x"73cc38d3",
          2400 => x"39805675",
          2401 => x"802e80ca",
          2402 => x"38811c55",
          2403 => x"7481ff94",
          2404 => x"3474982b",
          2405 => x"70982c81",
          2406 => x"ff903370",
          2407 => x"982b7098",
          2408 => x"2c701011",
          2409 => x"70822b81",
          2410 => x"e9cc1133",
          2411 => x"5e515151",
          2412 => x"57585155",
          2413 => x"74772e09",
          2414 => x"8106fe92",
          2415 => x"3881e9d0",
          2416 => x"14087d0c",
          2417 => x"800b81ff",
          2418 => x"9434800b",
          2419 => x"81ff9034",
          2420 => x"92397581",
          2421 => x"ff943475",
          2422 => x"81ff9034",
          2423 => x"78af3d34",
          2424 => x"757d0c7e",
          2425 => x"54738b26",
          2426 => x"fde13873",
          2427 => x"842981e1",
          2428 => x"d4055473",
          2429 => x"080481ff",
          2430 => x"9c335473",
          2431 => x"7e2efdcb",
          2432 => x"3881ff98",
          2433 => x"33557375",
          2434 => x"27ab3874",
          2435 => x"982b7098",
          2436 => x"2c515573",
          2437 => x"75249e38",
          2438 => x"741a5473",
          2439 => x"33811534",
          2440 => x"7481800a",
          2441 => x"2981ff0a",
          2442 => x"0570982c",
          2443 => x"81ff9c33",
          2444 => x"565155df",
          2445 => x"3981ff9c",
          2446 => x"33811156",
          2447 => x"547481ff",
          2448 => x"9c34731a",
          2449 => x"54ae3d33",
          2450 => x"743481ff",
          2451 => x"98335473",
          2452 => x"7e278938",
          2453 => x"81145473",
          2454 => x"81ff9834",
          2455 => x"81ff9c33",
          2456 => x"7081800a",
          2457 => x"2981ff0a",
          2458 => x"0570982c",
          2459 => x"81ff9833",
          2460 => x"5a515656",
          2461 => x"747725a2",
          2462 => x"38741a70",
          2463 => x"335254e8",
          2464 => x"c73f7481",
          2465 => x"800a2981",
          2466 => x"800a0570",
          2467 => x"982c81ff",
          2468 => x"98335651",
          2469 => x"55737524",
          2470 => x"e03881ff",
          2471 => x"9c337098",
          2472 => x"2b70982c",
          2473 => x"81ff9833",
          2474 => x"5a515656",
          2475 => x"747725fc",
          2476 => x"9a388851",
          2477 => x"e8923f74",
          2478 => x"81800a29",
          2479 => x"81800a05",
          2480 => x"70982c81",
          2481 => x"ff983356",
          2482 => x"51557375",
          2483 => x"24e438fb",
          2484 => x"fa3981ff",
          2485 => x"9c337081",
          2486 => x"ff065555",
          2487 => x"73802efb",
          2488 => x"ea3881ff",
          2489 => x"9833ff05",
          2490 => x"547381ff",
          2491 => x"9834ff15",
          2492 => x"547381ff",
          2493 => x"9c348851",
          2494 => x"e7ce3f81",
          2495 => x"ff9c3370",
          2496 => x"982b7098",
          2497 => x"2c81ff98",
          2498 => x"33575156",
          2499 => x"57747425",
          2500 => x"a738741a",
          2501 => x"54811433",
          2502 => x"74347333",
          2503 => x"51e7a93f",
          2504 => x"7481800a",
          2505 => x"2981800a",
          2506 => x"0570982c",
          2507 => x"81ff9833",
          2508 => x"58515575",
          2509 => x"7524db38",
          2510 => x"a051e78c",
          2511 => x"3f81ff9c",
          2512 => x"3370982b",
          2513 => x"70982c81",
          2514 => x"ff983357",
          2515 => x"51565774",
          2516 => x"7424faf7",
          2517 => x"388851e6",
          2518 => x"ef3f7481",
          2519 => x"800a2981",
          2520 => x"800a0570",
          2521 => x"982c81ff",
          2522 => x"98335851",
          2523 => x"55757525",
          2524 => x"e438fad7",
          2525 => x"3981ff98",
          2526 => x"337a0554",
          2527 => x"8074348a",
          2528 => x"51e6c53f",
          2529 => x"81ff9852",
          2530 => x"7951f7c6",
          2531 => x"3f81fef0",
          2532 => x"0881ff06",
          2533 => x"54739838",
          2534 => x"81ff9833",
          2535 => x"5473802e",
          2536 => x"84c93881",
          2537 => x"53735279",
          2538 => x"51f3c23f",
          2539 => x"84bd3980",
          2540 => x"7a3484b7",
          2541 => x"3981ff9c",
          2542 => x"33547380",
          2543 => x"2efa8c38",
          2544 => x"8851e684",
          2545 => x"3f81ff9c",
          2546 => x"33ff0554",
          2547 => x"7381ff9c",
          2548 => x"347381ff",
          2549 => x"0654e339",
          2550 => x"81ff9c33",
          2551 => x"81ff9833",
          2552 => x"55557375",
          2553 => x"2ef9e438",
          2554 => x"ff145473",
          2555 => x"81ff9834",
          2556 => x"74982b70",
          2557 => x"982c7581",
          2558 => x"ff065651",
          2559 => x"55747425",
          2560 => x"a738741a",
          2561 => x"54811433",
          2562 => x"74347333",
          2563 => x"51e5b93f",
          2564 => x"7481800a",
          2565 => x"2981800a",
          2566 => x"0570982c",
          2567 => x"81ff9833",
          2568 => x"58515575",
          2569 => x"7524db38",
          2570 => x"a051e59c",
          2571 => x"3f81ff9c",
          2572 => x"3370982b",
          2573 => x"70982c81",
          2574 => x"ff983357",
          2575 => x"51565774",
          2576 => x"7424f987",
          2577 => x"388851e4",
          2578 => x"ff3f7481",
          2579 => x"800a2981",
          2580 => x"800a0570",
          2581 => x"982c81ff",
          2582 => x"98335851",
          2583 => x"55757525",
          2584 => x"e438f8e7",
          2585 => x"3981ff9c",
          2586 => x"337081ff",
          2587 => x"0681ff98",
          2588 => x"33595654",
          2589 => x"747727f8",
          2590 => x"d2388114",
          2591 => x"547381ff",
          2592 => x"9c34741a",
          2593 => x"70335254",
          2594 => x"e4be3f81",
          2595 => x"ff9c3370",
          2596 => x"81ff0681",
          2597 => x"ff983358",
          2598 => x"56547575",
          2599 => x"26dc38f8",
          2600 => x"aa397aae",
          2601 => x"3881fbb0",
          2602 => x"08557480",
          2603 => x"2ea43874",
          2604 => x"51cb9a3f",
          2605 => x"81fef008",
          2606 => x"81ff9834",
          2607 => x"81fef008",
          2608 => x"81ff0681",
          2609 => x"05537452",
          2610 => x"7951c7e6",
          2611 => x"3f935b81",
          2612 => x"c1397a84",
          2613 => x"2981fae4",
          2614 => x"05fc1108",
          2615 => x"56547480",
          2616 => x"2ea53874",
          2617 => x"51cae63f",
          2618 => x"81fef008",
          2619 => x"81ff9834",
          2620 => x"81fef008",
          2621 => x"81ff0681",
          2622 => x"05537452",
          2623 => x"7951c7b2",
          2624 => x"3fff1b54",
          2625 => x"80de3973",
          2626 => x"08557480",
          2627 => x"2ef7bc38",
          2628 => x"7451cab9",
          2629 => x"3f80e239",
          2630 => x"7a932e09",
          2631 => x"81069338",
          2632 => x"81fae408",
          2633 => x"5574802e",
          2634 => x"89387451",
          2635 => x"ca9f3f80",
          2636 => x"c8397a84",
          2637 => x"2981fae4",
          2638 => x"05841108",
          2639 => x"56547480",
          2640 => x"2ea93874",
          2641 => x"51ca863f",
          2642 => x"81fef008",
          2643 => x"81ff9834",
          2644 => x"81fef008",
          2645 => x"81ff0681",
          2646 => x"05537452",
          2647 => x"7951c6d2",
          2648 => x"3f811b54",
          2649 => x"7381ff06",
          2650 => x"5ba83973",
          2651 => x"08557480",
          2652 => x"2ef6d838",
          2653 => x"7451c9d5",
          2654 => x"3f81fef0",
          2655 => x"0881ff98",
          2656 => x"3481fef0",
          2657 => x"0881ff06",
          2658 => x"81055374",
          2659 => x"527951c6",
          2660 => x"a13f81ff",
          2661 => x"9c5381ff",
          2662 => x"98335279",
          2663 => x"51ef903f",
          2664 => x"f6a93981",
          2665 => x"ff9c3370",
          2666 => x"81ff0681",
          2667 => x"ff983359",
          2668 => x"56547477",
          2669 => x"27f69438",
          2670 => x"81145473",
          2671 => x"81ff9c34",
          2672 => x"741a7033",
          2673 => x"5254e280",
          2674 => x"3ff68039",
          2675 => x"81ff9c33",
          2676 => x"5473802e",
          2677 => x"f5f53888",
          2678 => x"51e1ed3f",
          2679 => x"81ff9c33",
          2680 => x"ff055473",
          2681 => x"81ff9c34",
          2682 => x"f5e13980",
          2683 => x"0b81ff9c",
          2684 => x"34800b81",
          2685 => x"ff983479",
          2686 => x"81fef00c",
          2687 => x"af3d0d04",
          2688 => x"ff3d0d02",
          2689 => x"8f053351",
          2690 => x"81527072",
          2691 => x"26873881",
          2692 => x"fbd81133",
          2693 => x"527181fe",
          2694 => x"f00c833d",
          2695 => x"0d04fc3d",
          2696 => x"0d029b05",
          2697 => x"33028405",
          2698 => x"9f053356",
          2699 => x"53835172",
          2700 => x"812680e0",
          2701 => x"3872842b",
          2702 => x"87c0928c",
          2703 => x"11535188",
          2704 => x"5474802e",
          2705 => x"84388188",
          2706 => x"5473720c",
          2707 => x"87c0928c",
          2708 => x"11518171",
          2709 => x"0c850b87",
          2710 => x"c0988c0c",
          2711 => x"70527108",
          2712 => x"70820651",
          2713 => x"5170802e",
          2714 => x"8a3887c0",
          2715 => x"988c0851",
          2716 => x"70ec3871",
          2717 => x"08fc8080",
          2718 => x"06527192",
          2719 => x"3887c098",
          2720 => x"8c085170",
          2721 => x"802e8738",
          2722 => x"7181fbd8",
          2723 => x"143481fb",
          2724 => x"d8133351",
          2725 => x"7081fef0",
          2726 => x"0c863d0d",
          2727 => x"04f33d0d",
          2728 => x"60626402",
          2729 => x"8c05bf05",
          2730 => x"33574058",
          2731 => x"5b837452",
          2732 => x"5afecd3f",
          2733 => x"81fef008",
          2734 => x"81067a54",
          2735 => x"527181be",
          2736 => x"38717275",
          2737 => x"842b87c0",
          2738 => x"92801187",
          2739 => x"c0928c12",
          2740 => x"87c09284",
          2741 => x"13415a40",
          2742 => x"575a5885",
          2743 => x"0b87c098",
          2744 => x"8c0c767d",
          2745 => x"0c84760c",
          2746 => x"75087085",
          2747 => x"2a708106",
          2748 => x"51535471",
          2749 => x"802e8e38",
          2750 => x"7b085271",
          2751 => x"7b708105",
          2752 => x"5d348119",
          2753 => x"598074a2",
          2754 => x"06535371",
          2755 => x"732e8338",
          2756 => x"81537883",
          2757 => x"ff268f38",
          2758 => x"72802e8a",
          2759 => x"3887c098",
          2760 => x"8c085271",
          2761 => x"c33887c0",
          2762 => x"988c0852",
          2763 => x"71802e87",
          2764 => x"38788480",
          2765 => x"2e993881",
          2766 => x"760c87c0",
          2767 => x"928c1553",
          2768 => x"72087082",
          2769 => x"06515271",
          2770 => x"f738ff1a",
          2771 => x"5a8d3984",
          2772 => x"80178119",
          2773 => x"7081ff06",
          2774 => x"5a535779",
          2775 => x"802e9038",
          2776 => x"73fc8080",
          2777 => x"06527187",
          2778 => x"387d7826",
          2779 => x"feed3873",
          2780 => x"fc808006",
          2781 => x"5271802e",
          2782 => x"83388152",
          2783 => x"71537281",
          2784 => x"fef00c8f",
          2785 => x"3d0d04f3",
          2786 => x"3d0d6062",
          2787 => x"64028c05",
          2788 => x"bf053357",
          2789 => x"40585b83",
          2790 => x"59807452",
          2791 => x"58fce13f",
          2792 => x"81fef008",
          2793 => x"81067954",
          2794 => x"5271782e",
          2795 => x"09810681",
          2796 => x"b1387774",
          2797 => x"842b87c0",
          2798 => x"92801187",
          2799 => x"c0928c12",
          2800 => x"87c09284",
          2801 => x"1340595f",
          2802 => x"565a850b",
          2803 => x"87c0988c",
          2804 => x"0c767d0c",
          2805 => x"82760c80",
          2806 => x"58750870",
          2807 => x"842a7081",
          2808 => x"06515354",
          2809 => x"71802e8c",
          2810 => x"387a7081",
          2811 => x"055c337c",
          2812 => x"0c811858",
          2813 => x"73812a70",
          2814 => x"81065152",
          2815 => x"71802e8a",
          2816 => x"3887c098",
          2817 => x"8c085271",
          2818 => x"d03887c0",
          2819 => x"988c0852",
          2820 => x"71802e87",
          2821 => x"38778480",
          2822 => x"2e993881",
          2823 => x"760c87c0",
          2824 => x"928c1553",
          2825 => x"72087082",
          2826 => x"06515271",
          2827 => x"f738ff19",
          2828 => x"598d3981",
          2829 => x"1a7081ff",
          2830 => x"06848019",
          2831 => x"595b5278",
          2832 => x"802e9038",
          2833 => x"73fc8080",
          2834 => x"06527187",
          2835 => x"387d7a26",
          2836 => x"fef83873",
          2837 => x"fc808006",
          2838 => x"5271802e",
          2839 => x"83388152",
          2840 => x"71537281",
          2841 => x"fef00c8f",
          2842 => x"3d0d04fa",
          2843 => x"3d0d7a02",
          2844 => x"8405a305",
          2845 => x"33028805",
          2846 => x"a7053371",
          2847 => x"54545657",
          2848 => x"fafe3f81",
          2849 => x"fef00881",
          2850 => x"06538354",
          2851 => x"7280fe38",
          2852 => x"850b87c0",
          2853 => x"988c0c81",
          2854 => x"5671762e",
          2855 => x"80dc3871",
          2856 => x"76249338",
          2857 => x"74842b87",
          2858 => x"c0928c11",
          2859 => x"54547180",
          2860 => x"2e8d3880",
          2861 => x"d4397183",
          2862 => x"2e80c638",
          2863 => x"80cb3972",
          2864 => x"0870812a",
          2865 => x"70810651",
          2866 => x"51527180",
          2867 => x"2e8a3887",
          2868 => x"c0988c08",
          2869 => x"5271e838",
          2870 => x"87c0988c",
          2871 => x"08527196",
          2872 => x"3881730c",
          2873 => x"87c0928c",
          2874 => x"14537208",
          2875 => x"70820651",
          2876 => x"5271f738",
          2877 => x"96398056",
          2878 => x"92398880",
          2879 => x"0a770c85",
          2880 => x"39818077",
          2881 => x"0c725683",
          2882 => x"39845675",
          2883 => x"547381fe",
          2884 => x"f00c883d",
          2885 => x"0d04fe3d",
          2886 => x"0d748111",
          2887 => x"33713371",
          2888 => x"882b0781",
          2889 => x"fef00c53",
          2890 => x"51843d0d",
          2891 => x"04fd3d0d",
          2892 => x"75831133",
          2893 => x"82123371",
          2894 => x"902b7188",
          2895 => x"2b078114",
          2896 => x"33707207",
          2897 => x"882b7533",
          2898 => x"710781fe",
          2899 => x"f00c5253",
          2900 => x"54565452",
          2901 => x"853d0d04",
          2902 => x"ff3d0d73",
          2903 => x"02840592",
          2904 => x"05225252",
          2905 => x"70727081",
          2906 => x"05543470",
          2907 => x"882a5170",
          2908 => x"7234833d",
          2909 => x"0d04ff3d",
          2910 => x"0d737552",
          2911 => x"52707270",
          2912 => x"81055434",
          2913 => x"70882a51",
          2914 => x"70727081",
          2915 => x"05543470",
          2916 => x"882a5170",
          2917 => x"72708105",
          2918 => x"54347088",
          2919 => x"2a517072",
          2920 => x"34833d0d",
          2921 => x"04fe3d0d",
          2922 => x"76757754",
          2923 => x"54517080",
          2924 => x"2e923871",
          2925 => x"70810553",
          2926 => x"33737081",
          2927 => x"055534ff",
          2928 => x"1151eb39",
          2929 => x"843d0d04",
          2930 => x"fe3d0d75",
          2931 => x"77765452",
          2932 => x"53727270",
          2933 => x"81055434",
          2934 => x"ff115170",
          2935 => x"f438843d",
          2936 => x"0d04fc3d",
          2937 => x"0d787779",
          2938 => x"56565374",
          2939 => x"70810556",
          2940 => x"33747081",
          2941 => x"05563371",
          2942 => x"7131ff16",
          2943 => x"56525252",
          2944 => x"72802e86",
          2945 => x"3871802e",
          2946 => x"e2387181",
          2947 => x"fef00c86",
          2948 => x"3d0d04fe",
          2949 => x"3d0d7476",
          2950 => x"54518939",
          2951 => x"71732e8a",
          2952 => x"38811151",
          2953 => x"70335271",
          2954 => x"f3387033",
          2955 => x"81fef00c",
          2956 => x"843d0d04",
          2957 => x"800b81fe",
          2958 => x"f00c0480",
          2959 => x"0b81fef0",
          2960 => x"0c04f73d",
          2961 => x"0d7b5680",
          2962 => x"0b831733",
          2963 => x"565a747a",
          2964 => x"2e80d638",
          2965 => x"8154b016",
          2966 => x"0853b416",
          2967 => x"70538117",
          2968 => x"335259fa",
          2969 => x"a23f81fe",
          2970 => x"f0087a2e",
          2971 => x"098106b7",
          2972 => x"3881fef0",
          2973 => x"08831734",
          2974 => x"b0160870",
          2975 => x"a4180831",
          2976 => x"9c180859",
          2977 => x"56587477",
          2978 => x"279f3882",
          2979 => x"16335574",
          2980 => x"822e0981",
          2981 => x"06933881",
          2982 => x"54761853",
          2983 => x"78528116",
          2984 => x"3351f9e3",
          2985 => x"3f833981",
          2986 => x"5a7981fe",
          2987 => x"f00c8b3d",
          2988 => x"0d04fa3d",
          2989 => x"0d787a56",
          2990 => x"56805774",
          2991 => x"b017082e",
          2992 => x"af387551",
          2993 => x"fefc3f81",
          2994 => x"fef00857",
          2995 => x"81fef008",
          2996 => x"9f388154",
          2997 => x"7453b416",
          2998 => x"52811633",
          2999 => x"51f7be3f",
          3000 => x"81fef008",
          3001 => x"802e8538",
          3002 => x"ff558157",
          3003 => x"74b0170c",
          3004 => x"7681fef0",
          3005 => x"0c883d0d",
          3006 => x"04f83d0d",
          3007 => x"7a705257",
          3008 => x"fec03f81",
          3009 => x"fef00858",
          3010 => x"81fef008",
          3011 => x"81913876",
          3012 => x"33557483",
          3013 => x"2e098106",
          3014 => x"80f03884",
          3015 => x"17335978",
          3016 => x"812e0981",
          3017 => x"0680e338",
          3018 => x"84805381",
          3019 => x"fef00852",
          3020 => x"b4177052",
          3021 => x"56fd913f",
          3022 => x"82d4d552",
          3023 => x"84b21751",
          3024 => x"fc963f84",
          3025 => x"8b85a4d2",
          3026 => x"527551fc",
          3027 => x"a93f868a",
          3028 => x"85e4f252",
          3029 => x"84981751",
          3030 => x"fc9c3f90",
          3031 => x"17085284",
          3032 => x"9c1751fc",
          3033 => x"913f8c17",
          3034 => x"085284a0",
          3035 => x"1751fc86",
          3036 => x"3fa01708",
          3037 => x"810570b0",
          3038 => x"190c7955",
          3039 => x"53755281",
          3040 => x"173351f8",
          3041 => x"823f7784",
          3042 => x"18348053",
          3043 => x"80528117",
          3044 => x"3351f9d7",
          3045 => x"3f81fef0",
          3046 => x"08802e83",
          3047 => x"38815877",
          3048 => x"81fef00c",
          3049 => x"8a3d0d04",
          3050 => x"fb3d0d77",
          3051 => x"fe1a9812",
          3052 => x"08fe0555",
          3053 => x"56548056",
          3054 => x"7473278d",
          3055 => x"388a1422",
          3056 => x"757129ac",
          3057 => x"16080557",
          3058 => x"537581fe",
          3059 => x"f00c873d",
          3060 => x"0d04f93d",
          3061 => x"0d7a7a70",
          3062 => x"08565457",
          3063 => x"81772781",
          3064 => x"df387698",
          3065 => x"15082781",
          3066 => x"d738ff74",
          3067 => x"33545872",
          3068 => x"822e80f5",
          3069 => x"38728224",
          3070 => x"89387281",
          3071 => x"2e8d3881",
          3072 => x"bf397283",
          3073 => x"2e818e38",
          3074 => x"81b63976",
          3075 => x"812a1770",
          3076 => x"892aa416",
          3077 => x"08055374",
          3078 => x"5255fd96",
          3079 => x"3f81fef0",
          3080 => x"08819f38",
          3081 => x"7483ff06",
          3082 => x"14b41133",
          3083 => x"81177089",
          3084 => x"2aa41808",
          3085 => x"05557654",
          3086 => x"575753fc",
          3087 => x"f53f81fe",
          3088 => x"f00880fe",
          3089 => x"387483ff",
          3090 => x"0614b411",
          3091 => x"3370882b",
          3092 => x"78077981",
          3093 => x"0671842a",
          3094 => x"5c525851",
          3095 => x"537280e2",
          3096 => x"38759fff",
          3097 => x"065880da",
          3098 => x"3976882a",
          3099 => x"a4150805",
          3100 => x"527351fc",
          3101 => x"bd3f81fe",
          3102 => x"f00880c6",
          3103 => x"38761083",
          3104 => x"fe067405",
          3105 => x"b40551f9",
          3106 => x"8d3f81fe",
          3107 => x"f00883ff",
          3108 => x"ff0658ae",
          3109 => x"3976872a",
          3110 => x"a4150805",
          3111 => x"527351fc",
          3112 => x"913f81fe",
          3113 => x"f0089b38",
          3114 => x"76822b83",
          3115 => x"fc067405",
          3116 => x"b40551f8",
          3117 => x"f83f81fe",
          3118 => x"f008f00a",
          3119 => x"06588339",
          3120 => x"81587781",
          3121 => x"fef00c89",
          3122 => x"3d0d04f8",
          3123 => x"3d0d7a7c",
          3124 => x"7e5a5856",
          3125 => x"82598177",
          3126 => x"27829e38",
          3127 => x"76981708",
          3128 => x"27829638",
          3129 => x"75335372",
          3130 => x"792e819d",
          3131 => x"38727924",
          3132 => x"89387281",
          3133 => x"2e8d3882",
          3134 => x"80397283",
          3135 => x"2e81b838",
          3136 => x"81f73976",
          3137 => x"812a1770",
          3138 => x"892aa418",
          3139 => x"08055376",
          3140 => x"5255fb9e",
          3141 => x"3f81fef0",
          3142 => x"085981fe",
          3143 => x"f00881d9",
          3144 => x"387483ff",
          3145 => x"0616b405",
          3146 => x"81167881",
          3147 => x"06595654",
          3148 => x"77537680",
          3149 => x"2e8f3877",
          3150 => x"842b9ff0",
          3151 => x"0674338f",
          3152 => x"06710751",
          3153 => x"53727434",
          3154 => x"810b8317",
          3155 => x"3474892a",
          3156 => x"a4170805",
          3157 => x"527551fa",
          3158 => x"d93f81fe",
          3159 => x"f0085981",
          3160 => x"fef00881",
          3161 => x"94387483",
          3162 => x"ff0616b4",
          3163 => x"0578842a",
          3164 => x"5454768f",
          3165 => x"3877882a",
          3166 => x"743381f0",
          3167 => x"06718f06",
          3168 => x"07515372",
          3169 => x"743480ec",
          3170 => x"3976882a",
          3171 => x"a4170805",
          3172 => x"527551fa",
          3173 => x"9d3f81fe",
          3174 => x"f0085981",
          3175 => x"fef00880",
          3176 => x"d8387783",
          3177 => x"ffff0652",
          3178 => x"761083fe",
          3179 => x"067605b4",
          3180 => x"0551f7a4",
          3181 => x"3fbe3976",
          3182 => x"872aa417",
          3183 => x"08055275",
          3184 => x"51f9ef3f",
          3185 => x"81fef008",
          3186 => x"5981fef0",
          3187 => x"08ab3877",
          3188 => x"f00a0677",
          3189 => x"822b83fc",
          3190 => x"067018b4",
          3191 => x"05705451",
          3192 => x"5454f6c9",
          3193 => x"3f81fef0",
          3194 => x"088f0a06",
          3195 => x"74075272",
          3196 => x"51f7833f",
          3197 => x"810b8317",
          3198 => x"347881fe",
          3199 => x"f00c8a3d",
          3200 => x"0d04f83d",
          3201 => x"0d7a7c7e",
          3202 => x"72085956",
          3203 => x"56598175",
          3204 => x"27a43874",
          3205 => x"98170827",
          3206 => x"9d387380",
          3207 => x"2eaa38ff",
          3208 => x"53735275",
          3209 => x"51fda43f",
          3210 => x"81fef008",
          3211 => x"5481fef0",
          3212 => x"0880f238",
          3213 => x"93398254",
          3214 => x"80eb3981",
          3215 => x"5480e639",
          3216 => x"81fef008",
          3217 => x"5480de39",
          3218 => x"74527851",
          3219 => x"fb843f81",
          3220 => x"fef00858",
          3221 => x"81fef008",
          3222 => x"802e80c7",
          3223 => x"3881fef0",
          3224 => x"08812ed2",
          3225 => x"3881fef0",
          3226 => x"08ff2ecf",
          3227 => x"38805374",
          3228 => x"527551fc",
          3229 => x"d63f81fe",
          3230 => x"f008c538",
          3231 => x"981608fe",
          3232 => x"11901808",
          3233 => x"57555774",
          3234 => x"74279038",
          3235 => x"81159017",
          3236 => x"0c841633",
          3237 => x"81075473",
          3238 => x"84173477",
          3239 => x"55767826",
          3240 => x"ffa63880",
          3241 => x"547381fe",
          3242 => x"f00c8a3d",
          3243 => x"0d04f63d",
          3244 => x"0d7c7e71",
          3245 => x"08595b5b",
          3246 => x"7995388c",
          3247 => x"17085877",
          3248 => x"802e8838",
          3249 => x"98170878",
          3250 => x"26b23881",
          3251 => x"58ae3979",
          3252 => x"527a51f9",
          3253 => x"fd3f8155",
          3254 => x"7481fef0",
          3255 => x"082782e0",
          3256 => x"3881fef0",
          3257 => x"085581fe",
          3258 => x"f008ff2e",
          3259 => x"82d23898",
          3260 => x"170881fe",
          3261 => x"f0082682",
          3262 => x"c7387958",
          3263 => x"90170870",
          3264 => x"56547380",
          3265 => x"2e82b938",
          3266 => x"777a2e09",
          3267 => x"810680e2",
          3268 => x"38811a56",
          3269 => x"98170876",
          3270 => x"26833882",
          3271 => x"5675527a",
          3272 => x"51f9af3f",
          3273 => x"805981fe",
          3274 => x"f008812e",
          3275 => x"09810686",
          3276 => x"3881fef0",
          3277 => x"085981fe",
          3278 => x"f0080970",
          3279 => x"30707207",
          3280 => x"8025707c",
          3281 => x"0781fef0",
          3282 => x"08545151",
          3283 => x"55557381",
          3284 => x"ef3881fe",
          3285 => x"f008802e",
          3286 => x"95388c17",
          3287 => x"08548174",
          3288 => x"27903873",
          3289 => x"98180827",
          3290 => x"89387358",
          3291 => x"85397580",
          3292 => x"db387756",
          3293 => x"81165698",
          3294 => x"17087626",
          3295 => x"89388256",
          3296 => x"75782681",
          3297 => x"ac387552",
          3298 => x"7a51f8c6",
          3299 => x"3f81fef0",
          3300 => x"08802eb8",
          3301 => x"38805981",
          3302 => x"fef00881",
          3303 => x"2e098106",
          3304 => x"863881fe",
          3305 => x"f0085981",
          3306 => x"fef00809",
          3307 => x"70307072",
          3308 => x"07802570",
          3309 => x"7c075151",
          3310 => x"55557380",
          3311 => x"f8387578",
          3312 => x"2e098106",
          3313 => x"ffae3873",
          3314 => x"5580f539",
          3315 => x"ff537552",
          3316 => x"7651f9f7",
          3317 => x"3f81fef0",
          3318 => x"0881fef0",
          3319 => x"08307081",
          3320 => x"fef00807",
          3321 => x"80255155",
          3322 => x"5579802e",
          3323 => x"94387380",
          3324 => x"2e8f3875",
          3325 => x"53795276",
          3326 => x"51f9d03f",
          3327 => x"81fef008",
          3328 => x"5574a538",
          3329 => x"758c180c",
          3330 => x"981708fe",
          3331 => x"05901808",
          3332 => x"56547474",
          3333 => x"268638ff",
          3334 => x"1590180c",
          3335 => x"84173381",
          3336 => x"07547384",
          3337 => x"18349739",
          3338 => x"ff567481",
          3339 => x"2e90388c",
          3340 => x"3980558c",
          3341 => x"3981fef0",
          3342 => x"08558539",
          3343 => x"81567555",
          3344 => x"7481fef0",
          3345 => x"0c8c3d0d",
          3346 => x"04f83d0d",
          3347 => x"7a705255",
          3348 => x"f3f03f81",
          3349 => x"fef00858",
          3350 => x"815681fe",
          3351 => x"f00880d8",
          3352 => x"387b5274",
          3353 => x"51f6c13f",
          3354 => x"81fef008",
          3355 => x"81fef008",
          3356 => x"b0170c59",
          3357 => x"84805377",
          3358 => x"52b41570",
          3359 => x"5257f2c8",
          3360 => x"3f775684",
          3361 => x"39811656",
          3362 => x"8a152258",
          3363 => x"75782797",
          3364 => x"38815475",
          3365 => x"19537652",
          3366 => x"81153351",
          3367 => x"ede93f81",
          3368 => x"fef00880",
          3369 => x"2edf388a",
          3370 => x"15227632",
          3371 => x"70307072",
          3372 => x"07709f2a",
          3373 => x"53515656",
          3374 => x"7581fef0",
          3375 => x"0c8a3d0d",
          3376 => x"04f83d0d",
          3377 => x"7a7c7108",
          3378 => x"58565774",
          3379 => x"f0800a26",
          3380 => x"80f13874",
          3381 => x"9f065372",
          3382 => x"80e93874",
          3383 => x"90180c88",
          3384 => x"17085473",
          3385 => x"aa387533",
          3386 => x"53827327",
          3387 => x"8838a816",
          3388 => x"0854739b",
          3389 => x"3874852a",
          3390 => x"53820b88",
          3391 => x"17225a58",
          3392 => x"72792780",
          3393 => x"fe38a816",
          3394 => x"0898180c",
          3395 => x"80cd398a",
          3396 => x"16227089",
          3397 => x"2b545872",
          3398 => x"7526b238",
          3399 => x"73527651",
          3400 => x"f5b03f81",
          3401 => x"fef00854",
          3402 => x"81fef008",
          3403 => x"ff2ebd38",
          3404 => x"810b81fe",
          3405 => x"f008278b",
          3406 => x"38981608",
          3407 => x"81fef008",
          3408 => x"26853882",
          3409 => x"58bd3974",
          3410 => x"733155cb",
          3411 => x"39735275",
          3412 => x"51f4d53f",
          3413 => x"81fef008",
          3414 => x"98180c73",
          3415 => x"94180c98",
          3416 => x"17085382",
          3417 => x"5872802e",
          3418 => x"9a388539",
          3419 => x"81589439",
          3420 => x"74892a13",
          3421 => x"98180c74",
          3422 => x"83ff0616",
          3423 => x"b4059c18",
          3424 => x"0c805877",
          3425 => x"81fef00c",
          3426 => x"8a3d0d04",
          3427 => x"f83d0d7a",
          3428 => x"70089012",
          3429 => x"08a00559",
          3430 => x"5754f080",
          3431 => x"0a772786",
          3432 => x"38800b98",
          3433 => x"150c9814",
          3434 => x"08538455",
          3435 => x"72802e81",
          3436 => x"cb387683",
          3437 => x"ff065877",
          3438 => x"81b53881",
          3439 => x"1398150c",
          3440 => x"94140855",
          3441 => x"74923876",
          3442 => x"852a8817",
          3443 => x"22565374",
          3444 => x"7326819b",
          3445 => x"3880c039",
          3446 => x"8a1622ff",
          3447 => x"0577892a",
          3448 => x"06537281",
          3449 => x"8a387452",
          3450 => x"7351f3e6",
          3451 => x"3f81fef0",
          3452 => x"08538255",
          3453 => x"810b81fe",
          3454 => x"f0082780",
          3455 => x"ff388155",
          3456 => x"81fef008",
          3457 => x"ff2e80f4",
          3458 => x"38981608",
          3459 => x"81fef008",
          3460 => x"2680ca38",
          3461 => x"7b8a3877",
          3462 => x"98150c84",
          3463 => x"5580dd39",
          3464 => x"94140852",
          3465 => x"7351f986",
          3466 => x"3f81fef0",
          3467 => x"08538755",
          3468 => x"81fef008",
          3469 => x"802e80c4",
          3470 => x"38825581",
          3471 => x"fef00881",
          3472 => x"2eba3881",
          3473 => x"5581fef0",
          3474 => x"08ff2eb0",
          3475 => x"3881fef0",
          3476 => x"08527551",
          3477 => x"fbf33f81",
          3478 => x"fef008a0",
          3479 => x"38729415",
          3480 => x"0c725275",
          3481 => x"51f2c13f",
          3482 => x"81fef008",
          3483 => x"98150c76",
          3484 => x"90150c77",
          3485 => x"16b4059c",
          3486 => x"150c8055",
          3487 => x"7481fef0",
          3488 => x"0c8a3d0d",
          3489 => x"04f73d0d",
          3490 => x"7b7d7108",
          3491 => x"5b5b5780",
          3492 => x"527651fc",
          3493 => x"ac3f81fe",
          3494 => x"f0085481",
          3495 => x"fef00880",
          3496 => x"ec3881fe",
          3497 => x"f0085698",
          3498 => x"17085278",
          3499 => x"51f0833f",
          3500 => x"81fef008",
          3501 => x"5481fef0",
          3502 => x"0880d238",
          3503 => x"81fef008",
          3504 => x"9c180870",
          3505 => x"33515458",
          3506 => x"7281e52e",
          3507 => x"09810683",
          3508 => x"38815881",
          3509 => x"fef00855",
          3510 => x"72833881",
          3511 => x"55777507",
          3512 => x"5372802e",
          3513 => x"8e388116",
          3514 => x"56757a2e",
          3515 => x"09810688",
          3516 => x"38a53981",
          3517 => x"fef00856",
          3518 => x"81527651",
          3519 => x"fd8e3f81",
          3520 => x"fef00854",
          3521 => x"81fef008",
          3522 => x"802eff9b",
          3523 => x"3873842e",
          3524 => x"09810683",
          3525 => x"38875473",
          3526 => x"81fef00c",
          3527 => x"8b3d0d04",
          3528 => x"fd3d0d76",
          3529 => x"9a115254",
          3530 => x"ebec3f81",
          3531 => x"fef00883",
          3532 => x"ffff0676",
          3533 => x"70335153",
          3534 => x"5371832e",
          3535 => x"09810690",
          3536 => x"38941451",
          3537 => x"ebd03f81",
          3538 => x"fef00890",
          3539 => x"2b730753",
          3540 => x"7281fef0",
          3541 => x"0c853d0d",
          3542 => x"04fc3d0d",
          3543 => x"77797083",
          3544 => x"ffff0654",
          3545 => x"9a125355",
          3546 => x"55ebed3f",
          3547 => x"76703351",
          3548 => x"5372832e",
          3549 => x"0981068b",
          3550 => x"3873902a",
          3551 => x"52941551",
          3552 => x"ebd63f86",
          3553 => x"3d0d04f7",
          3554 => x"3d0d7b7d",
          3555 => x"5b558475",
          3556 => x"085a5898",
          3557 => x"1508802e",
          3558 => x"818a3898",
          3559 => x"15085278",
          3560 => x"51ee8f3f",
          3561 => x"81fef008",
          3562 => x"5881fef0",
          3563 => x"0880f538",
          3564 => x"9c150870",
          3565 => x"33555373",
          3566 => x"86388458",
          3567 => x"80e6398b",
          3568 => x"133370bf",
          3569 => x"067081ff",
          3570 => x"06585153",
          3571 => x"72861634",
          3572 => x"81fef008",
          3573 => x"537381e5",
          3574 => x"2e833881",
          3575 => x"5373ae2e",
          3576 => x"a9388170",
          3577 => x"74065457",
          3578 => x"72802e9e",
          3579 => x"38758f2e",
          3580 => x"993881fe",
          3581 => x"f00876df",
          3582 => x"06545472",
          3583 => x"882e0981",
          3584 => x"06833876",
          3585 => x"54737a2e",
          3586 => x"a0388052",
          3587 => x"7451fafc",
          3588 => x"3f81fef0",
          3589 => x"085881fe",
          3590 => x"f0088938",
          3591 => x"981508fe",
          3592 => x"fa388639",
          3593 => x"800b9816",
          3594 => x"0c7781fe",
          3595 => x"f00c8b3d",
          3596 => x"0d04fb3d",
          3597 => x"0d777008",
          3598 => x"57548152",
          3599 => x"7351fcc5",
          3600 => x"3f81fef0",
          3601 => x"085581fe",
          3602 => x"f008b438",
          3603 => x"98140852",
          3604 => x"7551ecde",
          3605 => x"3f81fef0",
          3606 => x"085581fe",
          3607 => x"f008a038",
          3608 => x"a05381fe",
          3609 => x"f008529c",
          3610 => x"140851ea",
          3611 => x"db3f8b53",
          3612 => x"a014529c",
          3613 => x"140851ea",
          3614 => x"ac3f810b",
          3615 => x"83173474",
          3616 => x"81fef00c",
          3617 => x"873d0d04",
          3618 => x"fd3d0d75",
          3619 => x"70089812",
          3620 => x"08547053",
          3621 => x"5553ec9a",
          3622 => x"3f81fef0",
          3623 => x"088d389c",
          3624 => x"130853e5",
          3625 => x"7334810b",
          3626 => x"83153485",
          3627 => x"3d0d04fa",
          3628 => x"3d0d787a",
          3629 => x"5757800b",
          3630 => x"89173498",
          3631 => x"1708802e",
          3632 => x"81823880",
          3633 => x"70891855",
          3634 => x"55559c17",
          3635 => x"08147033",
          3636 => x"81165651",
          3637 => x"5271a02e",
          3638 => x"a8387185",
          3639 => x"2e098106",
          3640 => x"843881e5",
          3641 => x"5273892e",
          3642 => x"0981068b",
          3643 => x"38ae7370",
          3644 => x"81055534",
          3645 => x"81155571",
          3646 => x"73708105",
          3647 => x"55348115",
          3648 => x"558a7427",
          3649 => x"c5387515",
          3650 => x"88055280",
          3651 => x"0b811334",
          3652 => x"9c170852",
          3653 => x"8b123388",
          3654 => x"17349c17",
          3655 => x"089c1152",
          3656 => x"52e88a3f",
          3657 => x"81fef008",
          3658 => x"760c9612",
          3659 => x"51e7e73f",
          3660 => x"81fef008",
          3661 => x"86172398",
          3662 => x"1251e7da",
          3663 => x"3f81fef0",
          3664 => x"08841723",
          3665 => x"883d0d04",
          3666 => x"f33d0d7f",
          3667 => x"70085e5b",
          3668 => x"80617033",
          3669 => x"51555573",
          3670 => x"af2e8338",
          3671 => x"81557380",
          3672 => x"dc2e9138",
          3673 => x"74802e8c",
          3674 => x"38941d08",
          3675 => x"881c0caa",
          3676 => x"39811541",
          3677 => x"80617033",
          3678 => x"56565673",
          3679 => x"af2e0981",
          3680 => x"06833881",
          3681 => x"567380dc",
          3682 => x"32703070",
          3683 => x"80257807",
          3684 => x"51515473",
          3685 => x"dc387388",
          3686 => x"1c0c6070",
          3687 => x"33515473",
          3688 => x"9f269638",
          3689 => x"ff800bab",
          3690 => x"1c348052",
          3691 => x"7a51f691",
          3692 => x"3f81fef0",
          3693 => x"08558598",
          3694 => x"39913d61",
          3695 => x"a01d5c5a",
          3696 => x"5e8b53a0",
          3697 => x"527951e7",
          3698 => x"ff3f8070",
          3699 => x"59578879",
          3700 => x"33555c73",
          3701 => x"ae2e0981",
          3702 => x"0680d438",
          3703 => x"78187033",
          3704 => x"811a71ae",
          3705 => x"32703070",
          3706 => x"9f2a7382",
          3707 => x"26075151",
          3708 => x"535a5754",
          3709 => x"738c3879",
          3710 => x"17547574",
          3711 => x"34811757",
          3712 => x"db3975af",
          3713 => x"32703070",
          3714 => x"9f2a5151",
          3715 => x"547580dc",
          3716 => x"2e8c3873",
          3717 => x"802e8738",
          3718 => x"75a02682",
          3719 => x"bd387719",
          3720 => x"7e0ca454",
          3721 => x"a0762782",
          3722 => x"bd38a054",
          3723 => x"82b83978",
          3724 => x"18703381",
          3725 => x"1a5a5754",
          3726 => x"a0762781",
          3727 => x"fc3875af",
          3728 => x"32703077",
          3729 => x"80dc3270",
          3730 => x"30728025",
          3731 => x"71802507",
          3732 => x"51515651",
          3733 => x"5573802e",
          3734 => x"ac388439",
          3735 => x"81185880",
          3736 => x"781a7033",
          3737 => x"51555573",
          3738 => x"af2e0981",
          3739 => x"06833881",
          3740 => x"557380dc",
          3741 => x"32703070",
          3742 => x"80257707",
          3743 => x"51515473",
          3744 => x"db3881b5",
          3745 => x"3975ae2e",
          3746 => x"09810683",
          3747 => x"38815476",
          3748 => x"7c277407",
          3749 => x"5473802e",
          3750 => x"a2387b8b",
          3751 => x"32703077",
          3752 => x"ae327030",
          3753 => x"72802571",
          3754 => x"9f2a0753",
          3755 => x"51565155",
          3756 => x"7481a738",
          3757 => x"88578b5c",
          3758 => x"fef53975",
          3759 => x"982b5473",
          3760 => x"80258c38",
          3761 => x"7580ff06",
          3762 => x"81ebdc11",
          3763 => x"33575475",
          3764 => x"51e6e13f",
          3765 => x"81fef008",
          3766 => x"802eb238",
          3767 => x"78187033",
          3768 => x"811a7154",
          3769 => x"5a5654e6",
          3770 => x"d23f81fe",
          3771 => x"f008802e",
          3772 => x"80e838ff",
          3773 => x"1c547674",
          3774 => x"2780df38",
          3775 => x"79175475",
          3776 => x"74348117",
          3777 => x"7a115557",
          3778 => x"747434a7",
          3779 => x"39755281",
          3780 => x"eafc51e5",
          3781 => x"fe3f81fe",
          3782 => x"f008bf38",
          3783 => x"ff9f1654",
          3784 => x"73992689",
          3785 => x"38e01670",
          3786 => x"81ff0657",
          3787 => x"54791754",
          3788 => x"75743481",
          3789 => x"1757fdf7",
          3790 => x"3977197e",
          3791 => x"0c76802e",
          3792 => x"99387933",
          3793 => x"547381e5",
          3794 => x"2e098106",
          3795 => x"8438857a",
          3796 => x"348454a0",
          3797 => x"76278f38",
          3798 => x"8b398655",
          3799 => x"81f23984",
          3800 => x"5680f339",
          3801 => x"8054738b",
          3802 => x"1b34807b",
          3803 => x"0858527a",
          3804 => x"51f2ce3f",
          3805 => x"81fef008",
          3806 => x"5681fef0",
          3807 => x"0880d738",
          3808 => x"981b0852",
          3809 => x"7651e6aa",
          3810 => x"3f81fef0",
          3811 => x"085681fe",
          3812 => x"f00880c2",
          3813 => x"389c1b08",
          3814 => x"70335555",
          3815 => x"73802eff",
          3816 => x"be388b15",
          3817 => x"33bf0654",
          3818 => x"73861c34",
          3819 => x"8b153370",
          3820 => x"832a7081",
          3821 => x"06515558",
          3822 => x"7392388b",
          3823 => x"53795274",
          3824 => x"51e49f3f",
          3825 => x"81fef008",
          3826 => x"802e8b38",
          3827 => x"75527a51",
          3828 => x"f3ba3fff",
          3829 => x"9f3975ab",
          3830 => x"1c335755",
          3831 => x"74802ebb",
          3832 => x"3874842e",
          3833 => x"09810680",
          3834 => x"e7387585",
          3835 => x"2a708106",
          3836 => x"77822a58",
          3837 => x"51547380",
          3838 => x"2e963875",
          3839 => x"81065473",
          3840 => x"802efbb5",
          3841 => x"38ff800b",
          3842 => x"ab1c3480",
          3843 => x"5580c139",
          3844 => x"75810654",
          3845 => x"73ba3885",
          3846 => x"55b63975",
          3847 => x"822a7081",
          3848 => x"06515473",
          3849 => x"ab38861b",
          3850 => x"3370842a",
          3851 => x"70810651",
          3852 => x"55557380",
          3853 => x"2ee13890",
          3854 => x"1b0883ff",
          3855 => x"061db405",
          3856 => x"527c51f5",
          3857 => x"db3f81fe",
          3858 => x"f008881c",
          3859 => x"0cfaea39",
          3860 => x"7481fef0",
          3861 => x"0c8f3d0d",
          3862 => x"04f63d0d",
          3863 => x"7c5bff7b",
          3864 => x"08707173",
          3865 => x"55595c55",
          3866 => x"5973802e",
          3867 => x"81c63875",
          3868 => x"70810557",
          3869 => x"3370a026",
          3870 => x"525271ba",
          3871 => x"2e8d3870",
          3872 => x"ee3871ba",
          3873 => x"2e098106",
          3874 => x"81a53873",
          3875 => x"33d01170",
          3876 => x"81ff0651",
          3877 => x"52537089",
          3878 => x"26913882",
          3879 => x"147381ff",
          3880 => x"06d00556",
          3881 => x"5271762e",
          3882 => x"80f73880",
          3883 => x"0b81ebcc",
          3884 => x"59557708",
          3885 => x"7a555776",
          3886 => x"70810558",
          3887 => x"33747081",
          3888 => x"055633ff",
          3889 => x"9f125353",
          3890 => x"53709926",
          3891 => x"8938e013",
          3892 => x"7081ff06",
          3893 => x"5451ff9f",
          3894 => x"12517099",
          3895 => x"268938e0",
          3896 => x"127081ff",
          3897 => x"06535172",
          3898 => x"30709f2a",
          3899 => x"51517272",
          3900 => x"2e098106",
          3901 => x"853870ff",
          3902 => x"be387230",
          3903 => x"74773270",
          3904 => x"30707207",
          3905 => x"9f2a739f",
          3906 => x"2a075354",
          3907 => x"54517080",
          3908 => x"2e8f3881",
          3909 => x"15841959",
          3910 => x"55837525",
          3911 => x"ff94388b",
          3912 => x"39748324",
          3913 => x"86387476",
          3914 => x"7c0c5978",
          3915 => x"51863981",
          3916 => x"ffb43351",
          3917 => x"7081fef0",
          3918 => x"0c8c3d0d",
          3919 => x"04fa3d0d",
          3920 => x"7856800b",
          3921 => x"831734ff",
          3922 => x"0bb0170c",
          3923 => x"79527551",
          3924 => x"e2e03f84",
          3925 => x"5581fef0",
          3926 => x"08818038",
          3927 => x"84b21651",
          3928 => x"dfb43f81",
          3929 => x"fef00883",
          3930 => x"ffff0654",
          3931 => x"83557382",
          3932 => x"d4d52e09",
          3933 => x"810680e3",
          3934 => x"38800bb4",
          3935 => x"17335657",
          3936 => x"7481e92e",
          3937 => x"09810683",
          3938 => x"38815774",
          3939 => x"81eb3270",
          3940 => x"30708025",
          3941 => x"79075151",
          3942 => x"54738a38",
          3943 => x"7481e82e",
          3944 => x"098106b5",
          3945 => x"38835381",
          3946 => x"eb8c5280",
          3947 => x"ea1651e0",
          3948 => x"b13f81fe",
          3949 => x"f0085581",
          3950 => x"fef00880",
          3951 => x"2e9d3885",
          3952 => x"5381eb90",
          3953 => x"52818616",
          3954 => x"51e0973f",
          3955 => x"81fef008",
          3956 => x"5581fef0",
          3957 => x"08802e83",
          3958 => x"38825574",
          3959 => x"81fef00c",
          3960 => x"883d0d04",
          3961 => x"f23d0d61",
          3962 => x"02840580",
          3963 => x"cb053358",
          3964 => x"5580750c",
          3965 => x"6051fce1",
          3966 => x"3f81fef0",
          3967 => x"08588b56",
          3968 => x"800b81fe",
          3969 => x"f0082486",
          3970 => x"fc3881fe",
          3971 => x"f0088429",
          3972 => x"81ffa005",
          3973 => x"70085553",
          3974 => x"8c567380",
          3975 => x"2e86e638",
          3976 => x"73750c76",
          3977 => x"81fe0674",
          3978 => x"33545772",
          3979 => x"802eae38",
          3980 => x"81143351",
          3981 => x"d7ca3f81",
          3982 => x"fef00881",
          3983 => x"ff067081",
          3984 => x"06545572",
          3985 => x"98387680",
          3986 => x"2e86b838",
          3987 => x"74822a70",
          3988 => x"81065153",
          3989 => x"8a567286",
          3990 => x"ac3886a7",
          3991 => x"39807434",
          3992 => x"77811534",
          3993 => x"81528114",
          3994 => x"3351d7b2",
          3995 => x"3f81fef0",
          3996 => x"0881ff06",
          3997 => x"70810654",
          3998 => x"55835672",
          3999 => x"86873876",
          4000 => x"802e8f38",
          4001 => x"74822a70",
          4002 => x"81065153",
          4003 => x"8a567285",
          4004 => x"f4388070",
          4005 => x"5374525b",
          4006 => x"fda33f81",
          4007 => x"fef00881",
          4008 => x"ff065776",
          4009 => x"822e0981",
          4010 => x"0680e238",
          4011 => x"8c3d7456",
          4012 => x"58835683",
          4013 => x"f6153370",
          4014 => x"58537280",
          4015 => x"2e8d3883",
          4016 => x"fa1551dc",
          4017 => x"e83f81fe",
          4018 => x"f0085776",
          4019 => x"78708405",
          4020 => x"5a0cff16",
          4021 => x"90165656",
          4022 => x"758025d7",
          4023 => x"38800b8d",
          4024 => x"3d545672",
          4025 => x"70840554",
          4026 => x"085b8357",
          4027 => x"7a802e95",
          4028 => x"387a5273",
          4029 => x"51fcc63f",
          4030 => x"81fef008",
          4031 => x"81ff0657",
          4032 => x"81772789",
          4033 => x"38811656",
          4034 => x"837627d7",
          4035 => x"38815676",
          4036 => x"842e84f1",
          4037 => x"388d5676",
          4038 => x"812684e9",
          4039 => x"38bf1451",
          4040 => x"dbf43f81",
          4041 => x"fef00883",
          4042 => x"ffff0653",
          4043 => x"7284802e",
          4044 => x"09810684",
          4045 => x"d03880ca",
          4046 => x"1451dbda",
          4047 => x"3f81fef0",
          4048 => x"0883ffff",
          4049 => x"0658778d",
          4050 => x"3880d814",
          4051 => x"51dbde3f",
          4052 => x"81fef008",
          4053 => x"58779c15",
          4054 => x"0c80c414",
          4055 => x"33821534",
          4056 => x"80c41433",
          4057 => x"ff117081",
          4058 => x"ff065154",
          4059 => x"558d5672",
          4060 => x"81268491",
          4061 => x"387481ff",
          4062 => x"06787129",
          4063 => x"80c11633",
          4064 => x"52595372",
          4065 => x"8a152372",
          4066 => x"802e8b38",
          4067 => x"ff137306",
          4068 => x"5372802e",
          4069 => x"86388d56",
          4070 => x"83eb3980",
          4071 => x"c51451da",
          4072 => x"f53f81fe",
          4073 => x"f0085381",
          4074 => x"fef00888",
          4075 => x"1523728f",
          4076 => x"06578d56",
          4077 => x"7683ce38",
          4078 => x"80c71451",
          4079 => x"dad83f81",
          4080 => x"fef00883",
          4081 => x"ffff0655",
          4082 => x"748d3880",
          4083 => x"d41451da",
          4084 => x"dc3f81fe",
          4085 => x"f0085580",
          4086 => x"c21451da",
          4087 => x"b93f81fe",
          4088 => x"f00883ff",
          4089 => x"ff06538d",
          4090 => x"5672802e",
          4091 => x"83973888",
          4092 => x"14227814",
          4093 => x"71842a05",
          4094 => x"5a5a7875",
          4095 => x"26838638",
          4096 => x"8a142252",
          4097 => x"74793151",
          4098 => x"ff93a03f",
          4099 => x"81fef008",
          4100 => x"5581fef0",
          4101 => x"08802e82",
          4102 => x"ec3881fe",
          4103 => x"f00880ff",
          4104 => x"fffff526",
          4105 => x"83388357",
          4106 => x"7483fff5",
          4107 => x"26833882",
          4108 => x"57749ff5",
          4109 => x"26853881",
          4110 => x"5789398d",
          4111 => x"5676802e",
          4112 => x"82c33882",
          4113 => x"15709816",
          4114 => x"0c7ba016",
          4115 => x"0c731c70",
          4116 => x"a4170c7a",
          4117 => x"1dac170c",
          4118 => x"54557683",
          4119 => x"2e098106",
          4120 => x"af3880de",
          4121 => x"1451d9ae",
          4122 => x"3f81fef0",
          4123 => x"0883ffff",
          4124 => x"06538d56",
          4125 => x"72828e38",
          4126 => x"79828a38",
          4127 => x"80e01451",
          4128 => x"d9ab3f81",
          4129 => x"fef008a8",
          4130 => x"150c7482",
          4131 => x"2b53a239",
          4132 => x"8d567980",
          4133 => x"2e81ee38",
          4134 => x"7713a815",
          4135 => x"0c741553",
          4136 => x"76822e8d",
          4137 => x"38741015",
          4138 => x"70812a76",
          4139 => x"81060551",
          4140 => x"5383ff13",
          4141 => x"892a538d",
          4142 => x"56729c15",
          4143 => x"082681c5",
          4144 => x"38ff0b90",
          4145 => x"150cff0b",
          4146 => x"8c150cff",
          4147 => x"800b8415",
          4148 => x"3476832e",
          4149 => x"09810681",
          4150 => x"923880e4",
          4151 => x"1451d8b6",
          4152 => x"3f81fef0",
          4153 => x"0883ffff",
          4154 => x"06537281",
          4155 => x"2e098106",
          4156 => x"80f93881",
          4157 => x"1b527351",
          4158 => x"dbb83f81",
          4159 => x"fef00880",
          4160 => x"ea3881fe",
          4161 => x"f0088415",
          4162 => x"3484b214",
          4163 => x"51d8873f",
          4164 => x"81fef008",
          4165 => x"83ffff06",
          4166 => x"537282d4",
          4167 => x"d52e0981",
          4168 => x"0680c838",
          4169 => x"b41451d8",
          4170 => x"843f81fe",
          4171 => x"f008848b",
          4172 => x"85a4d22e",
          4173 => x"098106b3",
          4174 => x"38849814",
          4175 => x"51d7ee3f",
          4176 => x"81fef008",
          4177 => x"868a85e4",
          4178 => x"f22e0981",
          4179 => x"069d3884",
          4180 => x"9c1451d7",
          4181 => x"d83f81fe",
          4182 => x"f0089015",
          4183 => x"0c84a014",
          4184 => x"51d7ca3f",
          4185 => x"81fef008",
          4186 => x"8c150c76",
          4187 => x"743481ff",
          4188 => x"b0228105",
          4189 => x"537281ff",
          4190 => x"b0237286",
          4191 => x"1523800b",
          4192 => x"94150c80",
          4193 => x"567581fe",
          4194 => x"f00c903d",
          4195 => x"0d04fb3d",
          4196 => x"0d775489",
          4197 => x"5573802e",
          4198 => x"b9387308",
          4199 => x"5372802e",
          4200 => x"b1387233",
          4201 => x"5271802e",
          4202 => x"a9388613",
          4203 => x"22841522",
          4204 => x"57527176",
          4205 => x"2e098106",
          4206 => x"99388113",
          4207 => x"3351d0c0",
          4208 => x"3f81fef0",
          4209 => x"08810652",
          4210 => x"71883871",
          4211 => x"74085455",
          4212 => x"83398053",
          4213 => x"7873710c",
          4214 => x"527481fe",
          4215 => x"f00c873d",
          4216 => x"0d04fa3d",
          4217 => x"0d02ab05",
          4218 => x"337a5889",
          4219 => x"3dfc0552",
          4220 => x"56f4e63f",
          4221 => x"8b54800b",
          4222 => x"81fef008",
          4223 => x"24bc3881",
          4224 => x"fef00884",
          4225 => x"2981ffa0",
          4226 => x"05700855",
          4227 => x"5573802e",
          4228 => x"84388074",
          4229 => x"34785473",
          4230 => x"802e8438",
          4231 => x"80743478",
          4232 => x"750c7554",
          4233 => x"75802e92",
          4234 => x"38805389",
          4235 => x"3d705384",
          4236 => x"0551f7b0",
          4237 => x"3f81fef0",
          4238 => x"08547381",
          4239 => x"fef00c88",
          4240 => x"3d0d04eb",
          4241 => x"3d0d6702",
          4242 => x"840580e7",
          4243 => x"05335959",
          4244 => x"89547880",
          4245 => x"2e84c838",
          4246 => x"77bf0670",
          4247 => x"54983dd0",
          4248 => x"0553993d",
          4249 => x"84055258",
          4250 => x"f6fa3f81",
          4251 => x"fef00855",
          4252 => x"81fef008",
          4253 => x"84a4387a",
          4254 => x"5c68528c",
          4255 => x"3d705256",
          4256 => x"edc63f81",
          4257 => x"fef00855",
          4258 => x"81fef008",
          4259 => x"92380280",
          4260 => x"d7053370",
          4261 => x"982b5557",
          4262 => x"73802583",
          4263 => x"38865577",
          4264 => x"9c065473",
          4265 => x"802e81ab",
          4266 => x"3874802e",
          4267 => x"95387484",
          4268 => x"2e098106",
          4269 => x"aa387551",
          4270 => x"eaf83f81",
          4271 => x"fef00855",
          4272 => x"9e3902b2",
          4273 => x"05339106",
          4274 => x"547381b8",
          4275 => x"3877822a",
          4276 => x"70810651",
          4277 => x"5473802e",
          4278 => x"8e388855",
          4279 => x"83bc3977",
          4280 => x"88075874",
          4281 => x"83b43877",
          4282 => x"832a7081",
          4283 => x"06515473",
          4284 => x"802e81af",
          4285 => x"3862527a",
          4286 => x"51e8a53f",
          4287 => x"81fef008",
          4288 => x"568288b2",
          4289 => x"0a52628e",
          4290 => x"0551d4ea",
          4291 => x"3f6254a0",
          4292 => x"0b8b1534",
          4293 => x"80536252",
          4294 => x"7a51e8bd",
          4295 => x"3f805262",
          4296 => x"9c0551d4",
          4297 => x"d13f7a54",
          4298 => x"810b8315",
          4299 => x"3475802e",
          4300 => x"80f1387a",
          4301 => x"b0110851",
          4302 => x"54805375",
          4303 => x"52973dd4",
          4304 => x"0551ddbe",
          4305 => x"3f81fef0",
          4306 => x"085581fe",
          4307 => x"f00882ca",
          4308 => x"38b73974",
          4309 => x"82c43802",
          4310 => x"b2053370",
          4311 => x"842a7081",
          4312 => x"06515556",
          4313 => x"73802e86",
          4314 => x"38845582",
          4315 => x"ad397781",
          4316 => x"2a708106",
          4317 => x"51547380",
          4318 => x"2ea93875",
          4319 => x"81065473",
          4320 => x"802ea038",
          4321 => x"87558292",
          4322 => x"3973527a",
          4323 => x"51d6a33f",
          4324 => x"81fef008",
          4325 => x"7bff188c",
          4326 => x"120c5555",
          4327 => x"81fef008",
          4328 => x"81f83877",
          4329 => x"832a7081",
          4330 => x"06515473",
          4331 => x"802e8638",
          4332 => x"7780c007",
          4333 => x"587ab011",
          4334 => x"08a01b0c",
          4335 => x"63a41b0c",
          4336 => x"63537052",
          4337 => x"57e6d93f",
          4338 => x"81fef008",
          4339 => x"81fef008",
          4340 => x"881b0c63",
          4341 => x"9c05525a",
          4342 => x"d2d33f81",
          4343 => x"fef00881",
          4344 => x"fef0088c",
          4345 => x"1b0c777a",
          4346 => x"0c568617",
          4347 => x"22841a23",
          4348 => x"77901a34",
          4349 => x"800b911a",
          4350 => x"34800b9c",
          4351 => x"1a0c800b",
          4352 => x"941a0c77",
          4353 => x"852a7081",
          4354 => x"06515473",
          4355 => x"802e818d",
          4356 => x"3881fef0",
          4357 => x"08802e81",
          4358 => x"843881fe",
          4359 => x"f008941a",
          4360 => x"0c8a1722",
          4361 => x"70892b7b",
          4362 => x"525957a8",
          4363 => x"39765278",
          4364 => x"51d79f3f",
          4365 => x"81fef008",
          4366 => x"5781fef0",
          4367 => x"08812683",
          4368 => x"38825581",
          4369 => x"fef008ff",
          4370 => x"2e098106",
          4371 => x"83387955",
          4372 => x"75783156",
          4373 => x"74307076",
          4374 => x"07802551",
          4375 => x"54777627",
          4376 => x"8a388170",
          4377 => x"7506555a",
          4378 => x"73c33876",
          4379 => x"981a0c74",
          4380 => x"a9387583",
          4381 => x"ff065473",
          4382 => x"802ea238",
          4383 => x"76527a51",
          4384 => x"d6a63f81",
          4385 => x"fef00885",
          4386 => x"3882558e",
          4387 => x"3975892a",
          4388 => x"81fef008",
          4389 => x"059c1a0c",
          4390 => x"84398079",
          4391 => x"0c745473",
          4392 => x"81fef00c",
          4393 => x"973d0d04",
          4394 => x"f23d0d60",
          4395 => x"63656440",
          4396 => x"405d5980",
          4397 => x"7e0c903d",
          4398 => x"fc055278",
          4399 => x"51f9cf3f",
          4400 => x"81fef008",
          4401 => x"5581fef0",
          4402 => x"088a3891",
          4403 => x"19335574",
          4404 => x"802e8638",
          4405 => x"745682c4",
          4406 => x"39901933",
          4407 => x"81065587",
          4408 => x"5674802e",
          4409 => x"82b63895",
          4410 => x"39820b91",
          4411 => x"1a348256",
          4412 => x"82aa3981",
          4413 => x"0b911a34",
          4414 => x"815682a0",
          4415 => x"398c1908",
          4416 => x"941a0831",
          4417 => x"55747c27",
          4418 => x"8338745c",
          4419 => x"7b802e82",
          4420 => x"89389419",
          4421 => x"087083ff",
          4422 => x"06565674",
          4423 => x"81b2387e",
          4424 => x"8a1122ff",
          4425 => x"0577892a",
          4426 => x"065b5579",
          4427 => x"a8387587",
          4428 => x"38881908",
          4429 => x"558f3998",
          4430 => x"19085278",
          4431 => x"51d5933f",
          4432 => x"81fef008",
          4433 => x"55817527",
          4434 => x"ff9f3874",
          4435 => x"ff2effa3",
          4436 => x"3874981a",
          4437 => x"0c981908",
          4438 => x"527e51d4",
          4439 => x"cb3f81fe",
          4440 => x"f008802e",
          4441 => x"ff833881",
          4442 => x"fef0081a",
          4443 => x"7c892a59",
          4444 => x"5777802e",
          4445 => x"80d63877",
          4446 => x"1a7f8a11",
          4447 => x"22585c55",
          4448 => x"75752785",
          4449 => x"38757a31",
          4450 => x"58775476",
          4451 => x"537c5281",
          4452 => x"1b3351ca",
          4453 => x"883f81fe",
          4454 => x"f008fed7",
          4455 => x"387e8311",
          4456 => x"33565674",
          4457 => x"802e9f38",
          4458 => x"b0160877",
          4459 => x"31557478",
          4460 => x"27943884",
          4461 => x"8053b416",
          4462 => x"52b01608",
          4463 => x"7731892b",
          4464 => x"7d0551cf",
          4465 => x"e03f7789",
          4466 => x"2b56b939",
          4467 => x"769c1a0c",
          4468 => x"94190883",
          4469 => x"ff068480",
          4470 => x"71315755",
          4471 => x"7b762783",
          4472 => x"387b569c",
          4473 => x"1908527e",
          4474 => x"51d1c73f",
          4475 => x"81fef008",
          4476 => x"fe813875",
          4477 => x"53941908",
          4478 => x"83ff061f",
          4479 => x"b405527c",
          4480 => x"51cfa23f",
          4481 => x"7b76317e",
          4482 => x"08177f0c",
          4483 => x"761e941b",
          4484 => x"0818941c",
          4485 => x"0c5e5cfd",
          4486 => x"f3398056",
          4487 => x"7581fef0",
          4488 => x"0c903d0d",
          4489 => x"04f23d0d",
          4490 => x"60636564",
          4491 => x"40405d58",
          4492 => x"807e0c90",
          4493 => x"3dfc0552",
          4494 => x"7751f6d2",
          4495 => x"3f81fef0",
          4496 => x"085581fe",
          4497 => x"f0088a38",
          4498 => x"91183355",
          4499 => x"74802e86",
          4500 => x"38745683",
          4501 => x"b8399018",
          4502 => x"3370812a",
          4503 => x"70810651",
          4504 => x"56568756",
          4505 => x"74802e83",
          4506 => x"a4389539",
          4507 => x"820b9119",
          4508 => x"34825683",
          4509 => x"9839810b",
          4510 => x"91193481",
          4511 => x"56838e39",
          4512 => x"9418087c",
          4513 => x"11565674",
          4514 => x"76278438",
          4515 => x"75095c7b",
          4516 => x"802e82ec",
          4517 => x"38941808",
          4518 => x"7083ff06",
          4519 => x"56567481",
          4520 => x"fd387e8a",
          4521 => x"1122ff05",
          4522 => x"77892a06",
          4523 => x"5c557abf",
          4524 => x"38758c38",
          4525 => x"88180855",
          4526 => x"749c387a",
          4527 => x"52853998",
          4528 => x"18085277",
          4529 => x"51d7e73f",
          4530 => x"81fef008",
          4531 => x"5581fef0",
          4532 => x"08802e82",
          4533 => x"ab387481",
          4534 => x"2eff9138",
          4535 => x"74ff2eff",
          4536 => x"95387498",
          4537 => x"190c8818",
          4538 => x"08853874",
          4539 => x"88190c7e",
          4540 => x"55b01508",
          4541 => x"9c19082e",
          4542 => x"0981068d",
          4543 => x"387451ce",
          4544 => x"c13f81fe",
          4545 => x"f008feee",
          4546 => x"38981808",
          4547 => x"527e51d1",
          4548 => x"973f81fe",
          4549 => x"f008802e",
          4550 => x"fed23881",
          4551 => x"fef0081b",
          4552 => x"7c892a5a",
          4553 => x"5778802e",
          4554 => x"80d53878",
          4555 => x"1b7f8a11",
          4556 => x"22585b55",
          4557 => x"75752785",
          4558 => x"38757b31",
          4559 => x"59785476",
          4560 => x"537c5281",
          4561 => x"1a3351c8",
          4562 => x"be3f81fe",
          4563 => x"f008fea6",
          4564 => x"387eb011",
          4565 => x"08783156",
          4566 => x"56747927",
          4567 => x"9b388480",
          4568 => x"53b01608",
          4569 => x"7731892b",
          4570 => x"7d0552b4",
          4571 => x"1651ccb5",
          4572 => x"3f7e5580",
          4573 => x"0b831634",
          4574 => x"78892b56",
          4575 => x"80db398c",
          4576 => x"18089419",
          4577 => x"08269338",
          4578 => x"7e51cdb6",
          4579 => x"3f81fef0",
          4580 => x"08fde338",
          4581 => x"7e77b012",
          4582 => x"0c55769c",
          4583 => x"190c9418",
          4584 => x"0883ff06",
          4585 => x"84807131",
          4586 => x"57557b76",
          4587 => x"2783387b",
          4588 => x"569c1808",
          4589 => x"527e51cd",
          4590 => x"f93f81fe",
          4591 => x"f008fdb6",
          4592 => x"3875537c",
          4593 => x"52941808",
          4594 => x"83ff061f",
          4595 => x"b40551cb",
          4596 => x"d43f7e55",
          4597 => x"810b8316",
          4598 => x"347b7631",
          4599 => x"7e08177f",
          4600 => x"0c761e94",
          4601 => x"1a081870",
          4602 => x"941c0c8c",
          4603 => x"1b085858",
          4604 => x"5e5c7476",
          4605 => x"27833875",
          4606 => x"55748c19",
          4607 => x"0cfd9039",
          4608 => x"90183380",
          4609 => x"c0075574",
          4610 => x"90193480",
          4611 => x"567581fe",
          4612 => x"f00c903d",
          4613 => x"0d04f83d",
          4614 => x"0d7a8b3d",
          4615 => x"fc055370",
          4616 => x"5256f2ea",
          4617 => x"3f81fef0",
          4618 => x"085781fe",
          4619 => x"f00880fb",
          4620 => x"38901633",
          4621 => x"70862a70",
          4622 => x"81065155",
          4623 => x"5573802e",
          4624 => x"80e938a0",
          4625 => x"16085278",
          4626 => x"51cce73f",
          4627 => x"81fef008",
          4628 => x"5781fef0",
          4629 => x"0880d438",
          4630 => x"a416088b",
          4631 => x"1133a007",
          4632 => x"5555738b",
          4633 => x"16348816",
          4634 => x"08537452",
          4635 => x"750851dd",
          4636 => x"e83f8c16",
          4637 => x"08529c15",
          4638 => x"51c9fb3f",
          4639 => x"8288b20a",
          4640 => x"52961551",
          4641 => x"c9f03f76",
          4642 => x"52921551",
          4643 => x"c9ca3f78",
          4644 => x"54810b83",
          4645 => x"15347851",
          4646 => x"ccdf3f81",
          4647 => x"fef00890",
          4648 => x"173381bf",
          4649 => x"06555773",
          4650 => x"90173476",
          4651 => x"81fef00c",
          4652 => x"8a3d0d04",
          4653 => x"fc3d0d76",
          4654 => x"705254fe",
          4655 => x"d93f81fe",
          4656 => x"f0085381",
          4657 => x"fef0089c",
          4658 => x"38863dfc",
          4659 => x"05527351",
          4660 => x"f1bc3f81",
          4661 => x"fef00853",
          4662 => x"81fef008",
          4663 => x"873881fe",
          4664 => x"f008740c",
          4665 => x"7281fef0",
          4666 => x"0c863d0d",
          4667 => x"04ff3d0d",
          4668 => x"843d51e6",
          4669 => x"e43f8b52",
          4670 => x"800b81fe",
          4671 => x"f008248b",
          4672 => x"3881fef0",
          4673 => x"0881ffb4",
          4674 => x"34805271",
          4675 => x"81fef00c",
          4676 => x"833d0d04",
          4677 => x"ef3d0d80",
          4678 => x"53933dd0",
          4679 => x"0552943d",
          4680 => x"51e9c13f",
          4681 => x"81fef008",
          4682 => x"5581fef0",
          4683 => x"0880e038",
          4684 => x"76586352",
          4685 => x"933dd405",
          4686 => x"51e08d3f",
          4687 => x"81fef008",
          4688 => x"5581fef0",
          4689 => x"08bc3802",
          4690 => x"80c70533",
          4691 => x"70982b55",
          4692 => x"56738025",
          4693 => x"8938767a",
          4694 => x"94120c54",
          4695 => x"b23902a2",
          4696 => x"05337084",
          4697 => x"2a708106",
          4698 => x"51555673",
          4699 => x"802e9e38",
          4700 => x"767f5370",
          4701 => x"5254dba8",
          4702 => x"3f81fef0",
          4703 => x"0894150c",
          4704 => x"8e3981fe",
          4705 => x"f008842e",
          4706 => x"09810683",
          4707 => x"38855574",
          4708 => x"81fef00c",
          4709 => x"933d0d04",
          4710 => x"e43d0d6f",
          4711 => x"6f5b5b80",
          4712 => x"7a348053",
          4713 => x"9e3dffb8",
          4714 => x"05529f3d",
          4715 => x"51e8b53f",
          4716 => x"81fef008",
          4717 => x"5781fef0",
          4718 => x"0882fc38",
          4719 => x"7b437a7c",
          4720 => x"94110847",
          4721 => x"55586454",
          4722 => x"73802e81",
          4723 => x"ed38a052",
          4724 => x"933d7052",
          4725 => x"55d5ea3f",
          4726 => x"81fef008",
          4727 => x"5781fef0",
          4728 => x"0882d438",
          4729 => x"68527b51",
          4730 => x"c9c83f81",
          4731 => x"fef00857",
          4732 => x"81fef008",
          4733 => x"82c13869",
          4734 => x"527b51da",
          4735 => x"a33f81fe",
          4736 => x"f0084576",
          4737 => x"527451d5",
          4738 => x"b83f81fe",
          4739 => x"f0085781",
          4740 => x"fef00882",
          4741 => x"a2388052",
          4742 => x"7451daeb",
          4743 => x"3f81fef0",
          4744 => x"085781fe",
          4745 => x"f008a438",
          4746 => x"69527b51",
          4747 => x"d9f23f73",
          4748 => x"81fef008",
          4749 => x"2ea63876",
          4750 => x"527451d6",
          4751 => x"cf3f81fe",
          4752 => x"f0085781",
          4753 => x"fef00880",
          4754 => x"2ecc3876",
          4755 => x"842e0981",
          4756 => x"06863882",
          4757 => x"5781e039",
          4758 => x"7681dc38",
          4759 => x"9e3dffbc",
          4760 => x"05527451",
          4761 => x"dcc93f76",
          4762 => x"903d7811",
          4763 => x"81113351",
          4764 => x"565a5673",
          4765 => x"802e9138",
          4766 => x"02b90555",
          4767 => x"81168116",
          4768 => x"70335656",
          4769 => x"5673f538",
          4770 => x"81165473",
          4771 => x"78268190",
          4772 => x"3875802e",
          4773 => x"99387816",
          4774 => x"810555ff",
          4775 => x"186f11ff",
          4776 => x"18ff1858",
          4777 => x"58555874",
          4778 => x"33743475",
          4779 => x"ee38ff18",
          4780 => x"6f115558",
          4781 => x"af7434fe",
          4782 => x"8d39777b",
          4783 => x"2e098106",
          4784 => x"8a38ff18",
          4785 => x"6f115558",
          4786 => x"af743480",
          4787 => x"0b81ffb4",
          4788 => x"33708429",
          4789 => x"81ebcc05",
          4790 => x"70087033",
          4791 => x"525c5656",
          4792 => x"5673762e",
          4793 => x"8d388116",
          4794 => x"701a7033",
          4795 => x"51555673",
          4796 => x"f5388216",
          4797 => x"54737826",
          4798 => x"a7388055",
          4799 => x"74762791",
          4800 => x"38741954",
          4801 => x"73337a70",
          4802 => x"81055c34",
          4803 => x"811555ec",
          4804 => x"39ba7a70",
          4805 => x"81055c34",
          4806 => x"74ff2e09",
          4807 => x"81068538",
          4808 => x"91579439",
          4809 => x"6e188119",
          4810 => x"59547333",
          4811 => x"7a708105",
          4812 => x"5c347a78",
          4813 => x"26ee3880",
          4814 => x"7a347681",
          4815 => x"fef00c9e",
          4816 => x"3d0d04f7",
          4817 => x"3d0d7b7d",
          4818 => x"8d3dfc05",
          4819 => x"54715357",
          4820 => x"55ecbb3f",
          4821 => x"81fef008",
          4822 => x"5381fef0",
          4823 => x"0882fa38",
          4824 => x"91153353",
          4825 => x"7282f238",
          4826 => x"8c150854",
          4827 => x"73762792",
          4828 => x"38901533",
          4829 => x"70812a70",
          4830 => x"81065154",
          4831 => x"57728338",
          4832 => x"73569415",
          4833 => x"08548070",
          4834 => x"94170c58",
          4835 => x"75782e82",
          4836 => x"9738798a",
          4837 => x"11227089",
          4838 => x"2b595153",
          4839 => x"73782eb7",
          4840 => x"387652ff",
          4841 => x"1651fefc",
          4842 => x"823f81fe",
          4843 => x"f008ff15",
          4844 => x"78547053",
          4845 => x"5553fefb",
          4846 => x"f23f81fe",
          4847 => x"f0087326",
          4848 => x"96387630",
          4849 => x"70750670",
          4850 => x"94180c77",
          4851 => x"71319818",
          4852 => x"08575851",
          4853 => x"53b13988",
          4854 => x"15085473",
          4855 => x"a6387352",
          4856 => x"7451cdca",
          4857 => x"3f81fef0",
          4858 => x"085481fe",
          4859 => x"f008812e",
          4860 => x"819a3881",
          4861 => x"fef008ff",
          4862 => x"2e819b38",
          4863 => x"81fef008",
          4864 => x"88160c73",
          4865 => x"98160c73",
          4866 => x"802e819c",
          4867 => x"38767627",
          4868 => x"80dc3875",
          4869 => x"77319416",
          4870 => x"08189417",
          4871 => x"0c901633",
          4872 => x"70812a70",
          4873 => x"81065155",
          4874 => x"5a567280",
          4875 => x"2e9a3873",
          4876 => x"527451cc",
          4877 => x"f93f81fe",
          4878 => x"f0085481",
          4879 => x"fef00894",
          4880 => x"3881fef0",
          4881 => x"0856a739",
          4882 => x"73527451",
          4883 => x"c7843f81",
          4884 => x"fef00854",
          4885 => x"73ff2ebe",
          4886 => x"38817427",
          4887 => x"af387953",
          4888 => x"73981408",
          4889 => x"27a63873",
          4890 => x"98160cff",
          4891 => x"a0399415",
          4892 => x"08169416",
          4893 => x"0c7583ff",
          4894 => x"06537280",
          4895 => x"2eaa3873",
          4896 => x"527951c6",
          4897 => x"a33f81fe",
          4898 => x"f0089438",
          4899 => x"820b9116",
          4900 => x"34825380",
          4901 => x"c439810b",
          4902 => x"91163481",
          4903 => x"53bb3975",
          4904 => x"892a81fe",
          4905 => x"f0080558",
          4906 => x"94150854",
          4907 => x"8c150874",
          4908 => x"27903873",
          4909 => x"8c160c90",
          4910 => x"153380c0",
          4911 => x"07537290",
          4912 => x"16347383",
          4913 => x"ff065372",
          4914 => x"802e8c38",
          4915 => x"779c1608",
          4916 => x"2e853877",
          4917 => x"9c160c80",
          4918 => x"537281fe",
          4919 => x"f00c8b3d",
          4920 => x"0d04f93d",
          4921 => x"0d795689",
          4922 => x"5475802e",
          4923 => x"818a3880",
          4924 => x"53893dfc",
          4925 => x"05528a3d",
          4926 => x"840551e1",
          4927 => x"e73f81fe",
          4928 => x"f0085581",
          4929 => x"fef00880",
          4930 => x"ea387776",
          4931 => x"0c7a5275",
          4932 => x"51d8b53f",
          4933 => x"81fef008",
          4934 => x"5581fef0",
          4935 => x"0880c338",
          4936 => x"ab163370",
          4937 => x"982b5557",
          4938 => x"807424a2",
          4939 => x"38861633",
          4940 => x"70842a70",
          4941 => x"81065155",
          4942 => x"5773802e",
          4943 => x"ad389c16",
          4944 => x"08527751",
          4945 => x"d3da3f81",
          4946 => x"fef00888",
          4947 => x"170c7754",
          4948 => x"86142284",
          4949 => x"17237452",
          4950 => x"7551cee5",
          4951 => x"3f81fef0",
          4952 => x"08557484",
          4953 => x"2e098106",
          4954 => x"85388555",
          4955 => x"86397480",
          4956 => x"2e843880",
          4957 => x"760c7454",
          4958 => x"7381fef0",
          4959 => x"0c893d0d",
          4960 => x"04fc3d0d",
          4961 => x"76873dfc",
          4962 => x"05537052",
          4963 => x"53e7ff3f",
          4964 => x"81fef008",
          4965 => x"873881fe",
          4966 => x"f008730c",
          4967 => x"863d0d04",
          4968 => x"fb3d0d77",
          4969 => x"79893dfc",
          4970 => x"05547153",
          4971 => x"5654e7de",
          4972 => x"3f81fef0",
          4973 => x"085381fe",
          4974 => x"f00880df",
          4975 => x"38749338",
          4976 => x"81fef008",
          4977 => x"527351cd",
          4978 => x"f83f81fe",
          4979 => x"f0085380",
          4980 => x"ca3981fe",
          4981 => x"f0085273",
          4982 => x"51d3ac3f",
          4983 => x"81fef008",
          4984 => x"5381fef0",
          4985 => x"08842e09",
          4986 => x"81068538",
          4987 => x"80538739",
          4988 => x"81fef008",
          4989 => x"a6387452",
          4990 => x"7351d5b3",
          4991 => x"3f725273",
          4992 => x"51cf893f",
          4993 => x"81fef008",
          4994 => x"84327030",
          4995 => x"7072079f",
          4996 => x"2c7081fe",
          4997 => x"f0080651",
          4998 => x"51545472",
          4999 => x"81fef00c",
          5000 => x"873d0d04",
          5001 => x"ee3d0d65",
          5002 => x"57805389",
          5003 => x"3d705396",
          5004 => x"3d5256df",
          5005 => x"af3f81fe",
          5006 => x"f0085581",
          5007 => x"fef008b2",
          5008 => x"38645275",
          5009 => x"51d6813f",
          5010 => x"81fef008",
          5011 => x"5581fef0",
          5012 => x"08a03802",
          5013 => x"80cb0533",
          5014 => x"70982b55",
          5015 => x"58738025",
          5016 => x"85388655",
          5017 => x"8d397680",
          5018 => x"2e883876",
          5019 => x"527551d4",
          5020 => x"be3f7481",
          5021 => x"fef00c94",
          5022 => x"3d0d04f0",
          5023 => x"3d0d6365",
          5024 => x"555c8053",
          5025 => x"923dec05",
          5026 => x"52933d51",
          5027 => x"ded63f81",
          5028 => x"fef0085b",
          5029 => x"81fef008",
          5030 => x"8280387c",
          5031 => x"740c7308",
          5032 => x"981108fe",
          5033 => x"11901308",
          5034 => x"59565855",
          5035 => x"75742691",
          5036 => x"38757c0c",
          5037 => x"81e43981",
          5038 => x"5b81cc39",
          5039 => x"825b81c7",
          5040 => x"3981fef0",
          5041 => x"08753355",
          5042 => x"5973812e",
          5043 => x"098106bf",
          5044 => x"3882755f",
          5045 => x"57765292",
          5046 => x"3df00551",
          5047 => x"c1f43f81",
          5048 => x"fef008ff",
          5049 => x"2ed13881",
          5050 => x"fef00881",
          5051 => x"2ece3881",
          5052 => x"fef00830",
          5053 => x"7081fef0",
          5054 => x"08078025",
          5055 => x"7a058119",
          5056 => x"7f53595a",
          5057 => x"54981408",
          5058 => x"7726ca38",
          5059 => x"80f939a4",
          5060 => x"150881fe",
          5061 => x"f0085758",
          5062 => x"75983877",
          5063 => x"5281187d",
          5064 => x"5258ffbf",
          5065 => x"8d3f81fe",
          5066 => x"f0085b81",
          5067 => x"fef00880",
          5068 => x"d6387c70",
          5069 => x"337712ff",
          5070 => x"1a5d5256",
          5071 => x"5474822e",
          5072 => x"0981069e",
          5073 => x"38b41451",
          5074 => x"ffbbcb3f",
          5075 => x"81fef008",
          5076 => x"83ffff06",
          5077 => x"70307080",
          5078 => x"251b8219",
          5079 => x"595b5154",
          5080 => x"9b39b414",
          5081 => x"51ffbbc5",
          5082 => x"3f81fef0",
          5083 => x"08f00a06",
          5084 => x"70307080",
          5085 => x"251b8419",
          5086 => x"595b5154",
          5087 => x"7583ff06",
          5088 => x"7a585679",
          5089 => x"ff923878",
          5090 => x"7c0c7c79",
          5091 => x"90120c84",
          5092 => x"11338107",
          5093 => x"56547484",
          5094 => x"15347a81",
          5095 => x"fef00c92",
          5096 => x"3d0d04f9",
          5097 => x"3d0d798a",
          5098 => x"3dfc0553",
          5099 => x"705257e3",
          5100 => x"dd3f81fe",
          5101 => x"f0085681",
          5102 => x"fef00881",
          5103 => x"a8389117",
          5104 => x"33567581",
          5105 => x"a0389017",
          5106 => x"3370812a",
          5107 => x"70810651",
          5108 => x"55558755",
          5109 => x"73802e81",
          5110 => x"8e389417",
          5111 => x"0854738c",
          5112 => x"18082781",
          5113 => x"8038739b",
          5114 => x"3881fef0",
          5115 => x"08538817",
          5116 => x"08527651",
          5117 => x"c48c3f81",
          5118 => x"fef00874",
          5119 => x"88190c56",
          5120 => x"80c93998",
          5121 => x"17085276",
          5122 => x"51ffbfc6",
          5123 => x"3f81fef0",
          5124 => x"08ff2e09",
          5125 => x"81068338",
          5126 => x"815681fe",
          5127 => x"f008812e",
          5128 => x"09810685",
          5129 => x"388256a3",
          5130 => x"3975a038",
          5131 => x"775481fe",
          5132 => x"f0089815",
          5133 => x"08279438",
          5134 => x"98170853",
          5135 => x"81fef008",
          5136 => x"527651c3",
          5137 => x"bd3f81fe",
          5138 => x"f0085694",
          5139 => x"17088c18",
          5140 => x"0c901733",
          5141 => x"80c00754",
          5142 => x"73901834",
          5143 => x"75802e85",
          5144 => x"38759118",
          5145 => x"34755574",
          5146 => x"81fef00c",
          5147 => x"893d0d04",
          5148 => x"e23d0d82",
          5149 => x"53a03dff",
          5150 => x"a40552a1",
          5151 => x"3d51dae4",
          5152 => x"3f81fef0",
          5153 => x"085581fe",
          5154 => x"f00881f5",
          5155 => x"387845a1",
          5156 => x"3d085295",
          5157 => x"3d705258",
          5158 => x"d1ae3f81",
          5159 => x"fef00855",
          5160 => x"81fef008",
          5161 => x"81db3802",
          5162 => x"80fb0533",
          5163 => x"70852a70",
          5164 => x"81065155",
          5165 => x"56865573",
          5166 => x"81c73875",
          5167 => x"982b5480",
          5168 => x"742481bd",
          5169 => x"380280d6",
          5170 => x"05337081",
          5171 => x"06585487",
          5172 => x"557681ad",
          5173 => x"386b5278",
          5174 => x"51ccc53f",
          5175 => x"81fef008",
          5176 => x"74842a70",
          5177 => x"81065155",
          5178 => x"5673802e",
          5179 => x"80d43878",
          5180 => x"5481fef0",
          5181 => x"08941508",
          5182 => x"2e818638",
          5183 => x"735a81fe",
          5184 => x"f0085c76",
          5185 => x"528a3d70",
          5186 => x"5254c7b5",
          5187 => x"3f81fef0",
          5188 => x"085581fe",
          5189 => x"f00880e9",
          5190 => x"3881fef0",
          5191 => x"08527351",
          5192 => x"cce53f81",
          5193 => x"fef00855",
          5194 => x"81fef008",
          5195 => x"86388755",
          5196 => x"80cf3981",
          5197 => x"fef00884",
          5198 => x"2e883881",
          5199 => x"fef00880",
          5200 => x"c0387751",
          5201 => x"cec23f81",
          5202 => x"fef00881",
          5203 => x"fef00830",
          5204 => x"7081fef0",
          5205 => x"08078025",
          5206 => x"51555575",
          5207 => x"802e9438",
          5208 => x"73802e8f",
          5209 => x"38805375",
          5210 => x"527751c1",
          5211 => x"953f81fe",
          5212 => x"f0085574",
          5213 => x"8c387851",
          5214 => x"ffbafe3f",
          5215 => x"81fef008",
          5216 => x"557481fe",
          5217 => x"f00ca03d",
          5218 => x"0d04e93d",
          5219 => x"0d825399",
          5220 => x"3dc00552",
          5221 => x"9a3d51d8",
          5222 => x"cb3f81fe",
          5223 => x"f0085481",
          5224 => x"fef00882",
          5225 => x"b038785e",
          5226 => x"69528e3d",
          5227 => x"705258cf",
          5228 => x"973f81fe",
          5229 => x"f0085481",
          5230 => x"fef00886",
          5231 => x"38885482",
          5232 => x"943981fe",
          5233 => x"f008842e",
          5234 => x"09810682",
          5235 => x"88380280",
          5236 => x"df053370",
          5237 => x"852a8106",
          5238 => x"51558654",
          5239 => x"7481f638",
          5240 => x"785a7452",
          5241 => x"8a3d7052",
          5242 => x"57c1c33f",
          5243 => x"81fef008",
          5244 => x"75555681",
          5245 => x"fef00883",
          5246 => x"38875481",
          5247 => x"fef00881",
          5248 => x"2e098106",
          5249 => x"83388254",
          5250 => x"81fef008",
          5251 => x"ff2e0981",
          5252 => x"06863881",
          5253 => x"5481b439",
          5254 => x"7381b038",
          5255 => x"81fef008",
          5256 => x"527851c4",
          5257 => x"a43f81fe",
          5258 => x"f0085481",
          5259 => x"fef00881",
          5260 => x"9a388b53",
          5261 => x"a052b419",
          5262 => x"51ffb78c",
          5263 => x"3f7854ae",
          5264 => x"0bb41534",
          5265 => x"7854900b",
          5266 => x"bf153482",
          5267 => x"88b20a52",
          5268 => x"80ca1951",
          5269 => x"ffb69f3f",
          5270 => x"755378b4",
          5271 => x"115351c9",
          5272 => x"f83fa053",
          5273 => x"78b41153",
          5274 => x"80d40551",
          5275 => x"ffb6b63f",
          5276 => x"7854ae0b",
          5277 => x"80d51534",
          5278 => x"7f537880",
          5279 => x"d4115351",
          5280 => x"c9d73f78",
          5281 => x"54810b83",
          5282 => x"15347751",
          5283 => x"cba43f81",
          5284 => x"fef00854",
          5285 => x"81fef008",
          5286 => x"b2388288",
          5287 => x"b20a5264",
          5288 => x"960551ff",
          5289 => x"b5d03f75",
          5290 => x"53645278",
          5291 => x"51c9aa3f",
          5292 => x"6454900b",
          5293 => x"8b153478",
          5294 => x"54810b83",
          5295 => x"15347851",
          5296 => x"ffb8b63f",
          5297 => x"81fef008",
          5298 => x"548b3980",
          5299 => x"53755276",
          5300 => x"51ffbeae",
          5301 => x"3f7381fe",
          5302 => x"f00c993d",
          5303 => x"0d04da3d",
          5304 => x"0da93d84",
          5305 => x"0551d2f1",
          5306 => x"3f8253a8",
          5307 => x"3dff8405",
          5308 => x"52a93d51",
          5309 => x"d5ee3f81",
          5310 => x"fef00855",
          5311 => x"81fef008",
          5312 => x"82d33878",
          5313 => x"4da93d08",
          5314 => x"529d3d70",
          5315 => x"5258ccb8",
          5316 => x"3f81fef0",
          5317 => x"085581fe",
          5318 => x"f00882b9",
          5319 => x"3802819b",
          5320 => x"053381a0",
          5321 => x"06548655",
          5322 => x"7382aa38",
          5323 => x"a053a43d",
          5324 => x"0852a83d",
          5325 => x"ff880551",
          5326 => x"ffb4ea3f",
          5327 => x"ac537752",
          5328 => x"923d7052",
          5329 => x"54ffb4dd",
          5330 => x"3faa3d08",
          5331 => x"527351cb",
          5332 => x"f73f81fe",
          5333 => x"f0085581",
          5334 => x"fef00895",
          5335 => x"38636f2e",
          5336 => x"09810688",
          5337 => x"3865a23d",
          5338 => x"082e9238",
          5339 => x"885581e5",
          5340 => x"3981fef0",
          5341 => x"08842e09",
          5342 => x"810681b8",
          5343 => x"387351c9",
          5344 => x"b13f81fe",
          5345 => x"f0085581",
          5346 => x"fef00881",
          5347 => x"c8386856",
          5348 => x"9353a83d",
          5349 => x"ff950552",
          5350 => x"8d1651ff",
          5351 => x"b4873f02",
          5352 => x"af05338b",
          5353 => x"17348b16",
          5354 => x"3370842a",
          5355 => x"70810651",
          5356 => x"55557389",
          5357 => x"3874a007",
          5358 => x"54738b17",
          5359 => x"34785481",
          5360 => x"0b831534",
          5361 => x"8b163370",
          5362 => x"842a7081",
          5363 => x"06515555",
          5364 => x"73802e80",
          5365 => x"e5386e64",
          5366 => x"2e80df38",
          5367 => x"75527851",
          5368 => x"c6be3f81",
          5369 => x"fef00852",
          5370 => x"7851ffb7",
          5371 => x"bb3f8255",
          5372 => x"81fef008",
          5373 => x"802e80dd",
          5374 => x"3881fef0",
          5375 => x"08527851",
          5376 => x"ffb5af3f",
          5377 => x"81fef008",
          5378 => x"7980d411",
          5379 => x"58585581",
          5380 => x"fef00880",
          5381 => x"c0388116",
          5382 => x"335473ae",
          5383 => x"2e098106",
          5384 => x"99386353",
          5385 => x"75527651",
          5386 => x"c6af3f78",
          5387 => x"54810b83",
          5388 => x"15348739",
          5389 => x"81fef008",
          5390 => x"9c387751",
          5391 => x"c8ca3f81",
          5392 => x"fef00855",
          5393 => x"81fef008",
          5394 => x"8c387851",
          5395 => x"ffb5aa3f",
          5396 => x"81fef008",
          5397 => x"557481fe",
          5398 => x"f00ca83d",
          5399 => x"0d04ed3d",
          5400 => x"0d0280db",
          5401 => x"05330284",
          5402 => x"0580df05",
          5403 => x"33575782",
          5404 => x"53953dd0",
          5405 => x"0552963d",
          5406 => x"51d2e93f",
          5407 => x"81fef008",
          5408 => x"5581fef0",
          5409 => x"0880cf38",
          5410 => x"785a6552",
          5411 => x"953dd405",
          5412 => x"51c9b53f",
          5413 => x"81fef008",
          5414 => x"5581fef0",
          5415 => x"08b83802",
          5416 => x"80cf0533",
          5417 => x"81a00654",
          5418 => x"865573aa",
          5419 => x"3875a706",
          5420 => x"6171098b",
          5421 => x"12337106",
          5422 => x"7a740607",
          5423 => x"51575556",
          5424 => x"748b1534",
          5425 => x"7854810b",
          5426 => x"83153478",
          5427 => x"51ffb4a9",
          5428 => x"3f81fef0",
          5429 => x"08557481",
          5430 => x"fef00c95",
          5431 => x"3d0d04ef",
          5432 => x"3d0d6456",
          5433 => x"8253933d",
          5434 => x"d0055294",
          5435 => x"3d51d1f4",
          5436 => x"3f81fef0",
          5437 => x"085581fe",
          5438 => x"f00880cb",
          5439 => x"38765863",
          5440 => x"52933dd4",
          5441 => x"0551c8c0",
          5442 => x"3f81fef0",
          5443 => x"085581fe",
          5444 => x"f008b438",
          5445 => x"0280c705",
          5446 => x"3381a006",
          5447 => x"54865573",
          5448 => x"a6388416",
          5449 => x"22861722",
          5450 => x"71902b07",
          5451 => x"5354961f",
          5452 => x"51ffb0c2",
          5453 => x"3f765481",
          5454 => x"0b831534",
          5455 => x"7651ffb3",
          5456 => x"b83f81fe",
          5457 => x"f0085574",
          5458 => x"81fef00c",
          5459 => x"933d0d04",
          5460 => x"ea3d0d69",
          5461 => x"6b5c5a80",
          5462 => x"53983dd0",
          5463 => x"0552993d",
          5464 => x"51d1813f",
          5465 => x"81fef008",
          5466 => x"81fef008",
          5467 => x"307081fe",
          5468 => x"f0080780",
          5469 => x"25515557",
          5470 => x"79802e81",
          5471 => x"85388170",
          5472 => x"75065555",
          5473 => x"73802e80",
          5474 => x"f9387b5d",
          5475 => x"805f8052",
          5476 => x"8d3d7052",
          5477 => x"54ffbea9",
          5478 => x"3f81fef0",
          5479 => x"085781fe",
          5480 => x"f00880d1",
          5481 => x"38745273",
          5482 => x"51c3dc3f",
          5483 => x"81fef008",
          5484 => x"5781fef0",
          5485 => x"08bf3881",
          5486 => x"fef00881",
          5487 => x"fef00865",
          5488 => x"5b595678",
          5489 => x"1881197b",
          5490 => x"18565955",
          5491 => x"74337434",
          5492 => x"8116568a",
          5493 => x"7827ec38",
          5494 => x"8b56751a",
          5495 => x"54807434",
          5496 => x"75802e9e",
          5497 => x"38ff1670",
          5498 => x"1b703351",
          5499 => x"555673a0",
          5500 => x"2ee8388e",
          5501 => x"3976842e",
          5502 => x"09810686",
          5503 => x"38807a34",
          5504 => x"80577630",
          5505 => x"70780780",
          5506 => x"2551547a",
          5507 => x"802e80c1",
          5508 => x"3873802e",
          5509 => x"bc387ba0",
          5510 => x"11085351",
          5511 => x"ffb1933f",
          5512 => x"81fef008",
          5513 => x"5781fef0",
          5514 => x"08a7387b",
          5515 => x"70335555",
          5516 => x"80c35673",
          5517 => x"832e8b38",
          5518 => x"80e45673",
          5519 => x"842e8338",
          5520 => x"a7567515",
          5521 => x"b40551ff",
          5522 => x"ade33f81",
          5523 => x"fef0087b",
          5524 => x"0c7681fe",
          5525 => x"f00c983d",
          5526 => x"0d04e63d",
          5527 => x"0d82539c",
          5528 => x"3dffb805",
          5529 => x"529d3d51",
          5530 => x"cefa3f81",
          5531 => x"fef00881",
          5532 => x"fef00856",
          5533 => x"5481fef0",
          5534 => x"08839838",
          5535 => x"8b53a052",
          5536 => x"8b3d7052",
          5537 => x"59ffaec0",
          5538 => x"3f736d70",
          5539 => x"337081ff",
          5540 => x"06525755",
          5541 => x"579f7427",
          5542 => x"81bc3878",
          5543 => x"587481ff",
          5544 => x"066d8105",
          5545 => x"4e705255",
          5546 => x"ffaf893f",
          5547 => x"81fef008",
          5548 => x"802ea538",
          5549 => x"6c703370",
          5550 => x"535754ff",
          5551 => x"aefd3f81",
          5552 => x"fef00880",
          5553 => x"2e8d3874",
          5554 => x"882b7607",
          5555 => x"6d81054e",
          5556 => x"55863981",
          5557 => x"fef00855",
          5558 => x"ff9f1570",
          5559 => x"83ffff06",
          5560 => x"51547399",
          5561 => x"268a38e0",
          5562 => x"157083ff",
          5563 => x"ff065654",
          5564 => x"80ff7527",
          5565 => x"873881ea",
          5566 => x"dc153355",
          5567 => x"74802ea3",
          5568 => x"38745281",
          5569 => x"ecdc51ff",
          5570 => x"ae893f81",
          5571 => x"fef00893",
          5572 => x"3881ff75",
          5573 => x"27883876",
          5574 => x"89268838",
          5575 => x"8b398a77",
          5576 => x"27863886",
          5577 => x"5581ec39",
          5578 => x"81ff7527",
          5579 => x"8f387488",
          5580 => x"2a547378",
          5581 => x"7081055a",
          5582 => x"34811757",
          5583 => x"74787081",
          5584 => x"055a3481",
          5585 => x"176d7033",
          5586 => x"7081ff06",
          5587 => x"52575557",
          5588 => x"739f26fe",
          5589 => x"c8388b3d",
          5590 => x"33548655",
          5591 => x"7381e52e",
          5592 => x"81b13876",
          5593 => x"802e9938",
          5594 => x"02a70555",
          5595 => x"76157033",
          5596 => x"515473a0",
          5597 => x"2e098106",
          5598 => x"8738ff17",
          5599 => x"5776ed38",
          5600 => x"79418043",
          5601 => x"8052913d",
          5602 => x"705255ff",
          5603 => x"bab33f81",
          5604 => x"fef00854",
          5605 => x"81fef008",
          5606 => x"80f73881",
          5607 => x"527451ff",
          5608 => x"bfe53f81",
          5609 => x"fef00854",
          5610 => x"81fef008",
          5611 => x"8d387680",
          5612 => x"c4386754",
          5613 => x"e5743480",
          5614 => x"c63981fe",
          5615 => x"f008842e",
          5616 => x"09810680",
          5617 => x"cc388054",
          5618 => x"76742e80",
          5619 => x"c4388152",
          5620 => x"7451ffbd",
          5621 => x"b03f81fe",
          5622 => x"f0085481",
          5623 => x"fef008b1",
          5624 => x"38a05381",
          5625 => x"fef00852",
          5626 => x"6751ffab",
          5627 => x"db3f6754",
          5628 => x"880b8b15",
          5629 => x"348b5378",
          5630 => x"526751ff",
          5631 => x"aba73f79",
          5632 => x"54810b83",
          5633 => x"15347951",
          5634 => x"ffadee3f",
          5635 => x"81fef008",
          5636 => x"54735574",
          5637 => x"81fef00c",
          5638 => x"9c3d0d04",
          5639 => x"f23d0d60",
          5640 => x"62028805",
          5641 => x"80cb0533",
          5642 => x"933dfc05",
          5643 => x"55725440",
          5644 => x"5e5ad2da",
          5645 => x"3f81fef0",
          5646 => x"085881fe",
          5647 => x"f00882bd",
          5648 => x"38911a33",
          5649 => x"587782b5",
          5650 => x"387c802e",
          5651 => x"97388c1a",
          5652 => x"08597890",
          5653 => x"38901a33",
          5654 => x"70812a70",
          5655 => x"81065155",
          5656 => x"55739038",
          5657 => x"87548297",
          5658 => x"39825882",
          5659 => x"90398158",
          5660 => x"828b397e",
          5661 => x"8a112270",
          5662 => x"892b7055",
          5663 => x"7f545656",
          5664 => x"56fee2a7",
          5665 => x"3fff147d",
          5666 => x"06703070",
          5667 => x"72079f2a",
          5668 => x"81fef008",
          5669 => x"058c1908",
          5670 => x"7c405a5d",
          5671 => x"55558177",
          5672 => x"27883898",
          5673 => x"16087726",
          5674 => x"83388257",
          5675 => x"76775659",
          5676 => x"80567452",
          5677 => x"7951ffae",
          5678 => x"993f8115",
          5679 => x"7f555598",
          5680 => x"14087526",
          5681 => x"83388255",
          5682 => x"81fef008",
          5683 => x"812eff99",
          5684 => x"3881fef0",
          5685 => x"08ff2eff",
          5686 => x"953881fe",
          5687 => x"f0088e38",
          5688 => x"81165675",
          5689 => x"7b2e0981",
          5690 => x"06873893",
          5691 => x"39745980",
          5692 => x"5674772e",
          5693 => x"098106ff",
          5694 => x"b9388758",
          5695 => x"80ff397d",
          5696 => x"802eba38",
          5697 => x"787b5555",
          5698 => x"7a802eb4",
          5699 => x"38811556",
          5700 => x"73812e09",
          5701 => x"81068338",
          5702 => x"ff567553",
          5703 => x"74527e51",
          5704 => x"ffafa83f",
          5705 => x"81fef008",
          5706 => x"5881fef0",
          5707 => x"0880ce38",
          5708 => x"748116ff",
          5709 => x"1656565c",
          5710 => x"73d33884",
          5711 => x"39ff195c",
          5712 => x"7e7c8c12",
          5713 => x"0c557d80",
          5714 => x"2eb33878",
          5715 => x"881b0c7c",
          5716 => x"8c1b0c90",
          5717 => x"1a3380c0",
          5718 => x"07547390",
          5719 => x"1b349815",
          5720 => x"08fe0590",
          5721 => x"16085754",
          5722 => x"75742691",
          5723 => x"38757b31",
          5724 => x"90160c84",
          5725 => x"15338107",
          5726 => x"54738416",
          5727 => x"34775473",
          5728 => x"81fef00c",
          5729 => x"903d0d04",
          5730 => x"e93d0d6b",
          5731 => x"6d028805",
          5732 => x"80eb0533",
          5733 => x"9d3d545a",
          5734 => x"5c59c5bd",
          5735 => x"3f8b5680",
          5736 => x"0b81fef0",
          5737 => x"08248bf8",
          5738 => x"3881fef0",
          5739 => x"08842981",
          5740 => x"ffa00570",
          5741 => x"08515574",
          5742 => x"802e8438",
          5743 => x"80753481",
          5744 => x"fef00881",
          5745 => x"ff065f81",
          5746 => x"527e51ff",
          5747 => x"a0d03f81",
          5748 => x"fef00881",
          5749 => x"ff067081",
          5750 => x"06565783",
          5751 => x"56748bc0",
          5752 => x"3876822a",
          5753 => x"70810651",
          5754 => x"558a5674",
          5755 => x"8bb23899",
          5756 => x"3dfc0553",
          5757 => x"83527e51",
          5758 => x"ffa4f03f",
          5759 => x"81fef008",
          5760 => x"99386755",
          5761 => x"74802e92",
          5762 => x"38748280",
          5763 => x"80268b38",
          5764 => x"ff157506",
          5765 => x"5574802e",
          5766 => x"83388148",
          5767 => x"78802e87",
          5768 => x"38848079",
          5769 => x"26923878",
          5770 => x"81800a26",
          5771 => x"8b38ff19",
          5772 => x"79065574",
          5773 => x"802e8638",
          5774 => x"93568ae4",
          5775 => x"3978892a",
          5776 => x"6e892a70",
          5777 => x"892b7759",
          5778 => x"4843597a",
          5779 => x"83388156",
          5780 => x"61307080",
          5781 => x"25770751",
          5782 => x"55915674",
          5783 => x"8ac23899",
          5784 => x"3df80553",
          5785 => x"81527e51",
          5786 => x"ffa4803f",
          5787 => x"815681fe",
          5788 => x"f0088aac",
          5789 => x"3877832a",
          5790 => x"70770681",
          5791 => x"fef00843",
          5792 => x"56457483",
          5793 => x"38bf4166",
          5794 => x"558e5660",
          5795 => x"75268a90",
          5796 => x"38746131",
          5797 => x"70485580",
          5798 => x"ff75278a",
          5799 => x"83389356",
          5800 => x"78818026",
          5801 => x"89fa3877",
          5802 => x"812a7081",
          5803 => x"06564374",
          5804 => x"802e9538",
          5805 => x"77870655",
          5806 => x"74822e83",
          5807 => x"8d387781",
          5808 => x"06557480",
          5809 => x"2e838338",
          5810 => x"77810655",
          5811 => x"9356825e",
          5812 => x"74802e89",
          5813 => x"cb38785a",
          5814 => x"7d832e09",
          5815 => x"810680e1",
          5816 => x"3878ae38",
          5817 => x"66912a57",
          5818 => x"810b81ed",
          5819 => x"8022565a",
          5820 => x"74802e9d",
          5821 => x"38747726",
          5822 => x"983881ed",
          5823 => x"80567910",
          5824 => x"82177022",
          5825 => x"57575a74",
          5826 => x"802e8638",
          5827 => x"767527ee",
          5828 => x"38795266",
          5829 => x"51fedd93",
          5830 => x"3f81fef0",
          5831 => x"08842984",
          5832 => x"87057089",
          5833 => x"2a5e55a0",
          5834 => x"5c800b81",
          5835 => x"fef008fc",
          5836 => x"808a0556",
          5837 => x"44fdfff0",
          5838 => x"0a752780",
          5839 => x"ec3888d3",
          5840 => x"3978ae38",
          5841 => x"668c2a57",
          5842 => x"810b81ec",
          5843 => x"f022565a",
          5844 => x"74802e9d",
          5845 => x"38747726",
          5846 => x"983881ec",
          5847 => x"f0567910",
          5848 => x"82177022",
          5849 => x"57575a74",
          5850 => x"802e8638",
          5851 => x"767527ee",
          5852 => x"38795266",
          5853 => x"51fedcb3",
          5854 => x"3f81fef0",
          5855 => x"08108405",
          5856 => x"5781fef0",
          5857 => x"089ff526",
          5858 => x"9638810b",
          5859 => x"81fef008",
          5860 => x"1081fef0",
          5861 => x"08057111",
          5862 => x"722a8305",
          5863 => x"59565e83",
          5864 => x"ff17892a",
          5865 => x"5d815ca0",
          5866 => x"44601c7d",
          5867 => x"11650569",
          5868 => x"7012ff05",
          5869 => x"71307072",
          5870 => x"0674315c",
          5871 => x"52595759",
          5872 => x"407d832e",
          5873 => x"09810689",
          5874 => x"38761c60",
          5875 => x"18415c84",
          5876 => x"39761d5d",
          5877 => x"79902918",
          5878 => x"70623168",
          5879 => x"58515574",
          5880 => x"762687af",
          5881 => x"38757c31",
          5882 => x"7d317a53",
          5883 => x"70653152",
          5884 => x"55fedbb7",
          5885 => x"3f81fef0",
          5886 => x"08587d83",
          5887 => x"2e098106",
          5888 => x"9b3881fe",
          5889 => x"f00883ff",
          5890 => x"f52680dd",
          5891 => x"38788783",
          5892 => x"3879812a",
          5893 => x"5978fdbe",
          5894 => x"3886f839",
          5895 => x"7d822e09",
          5896 => x"810680c5",
          5897 => x"3883fff5",
          5898 => x"0b81fef0",
          5899 => x"0827a038",
          5900 => x"788f3879",
          5901 => x"1a557480",
          5902 => x"c0268638",
          5903 => x"7459fd96",
          5904 => x"39628106",
          5905 => x"5574802e",
          5906 => x"8f38835e",
          5907 => x"fd883981",
          5908 => x"fef0089f",
          5909 => x"f5269238",
          5910 => x"7886b838",
          5911 => x"791a5981",
          5912 => x"807927fc",
          5913 => x"f13886ab",
          5914 => x"3980557d",
          5915 => x"812e0981",
          5916 => x"0683387d",
          5917 => x"559ff578",
          5918 => x"278b3874",
          5919 => x"8106558e",
          5920 => x"5674869c",
          5921 => x"38848053",
          5922 => x"80527a51",
          5923 => x"ffa2b93f",
          5924 => x"8b5381eb",
          5925 => x"98527a51",
          5926 => x"ffa28a3f",
          5927 => x"8480528b",
          5928 => x"1b51ffa1",
          5929 => x"b33f798d",
          5930 => x"1c347b83",
          5931 => x"ffff0652",
          5932 => x"8e1b51ff",
          5933 => x"a1a23f81",
          5934 => x"0b901c34",
          5935 => x"7d833270",
          5936 => x"3070962a",
          5937 => x"84800654",
          5938 => x"5155911b",
          5939 => x"51ffa188",
          5940 => x"3f665574",
          5941 => x"83ffff26",
          5942 => x"90387483",
          5943 => x"ffff0652",
          5944 => x"931b51ff",
          5945 => x"a0f23f8a",
          5946 => x"397452a0",
          5947 => x"1b51ffa1",
          5948 => x"853ff80b",
          5949 => x"951c34bf",
          5950 => x"52981b51",
          5951 => x"ffa0d93f",
          5952 => x"81ff529a",
          5953 => x"1b51ffa0",
          5954 => x"cf3f6052",
          5955 => x"9c1b51ff",
          5956 => x"a0e43f7d",
          5957 => x"832e0981",
          5958 => x"0680cb38",
          5959 => x"8288b20a",
          5960 => x"5280c31b",
          5961 => x"51ffa0ce",
          5962 => x"3f7c52a4",
          5963 => x"1b51ffa0",
          5964 => x"c53f8252",
          5965 => x"ac1b51ff",
          5966 => x"a0bc3f81",
          5967 => x"52b01b51",
          5968 => x"ffa0953f",
          5969 => x"8652b21b",
          5970 => x"51ffa08c",
          5971 => x"3fff800b",
          5972 => x"80c01c34",
          5973 => x"a90b80c2",
          5974 => x"1c349353",
          5975 => x"81eba452",
          5976 => x"80c71b51",
          5977 => x"ae398288",
          5978 => x"b20a52a7",
          5979 => x"1b51ffa0",
          5980 => x"853f7c83",
          5981 => x"ffff0652",
          5982 => x"961b51ff",
          5983 => x"9fda3fff",
          5984 => x"800ba41c",
          5985 => x"34a90ba6",
          5986 => x"1c349353",
          5987 => x"81ebb852",
          5988 => x"ab1b51ff",
          5989 => x"a08f3f82",
          5990 => x"d4d55283",
          5991 => x"fe1b7052",
          5992 => x"59ff9fb4",
          5993 => x"3f815460",
          5994 => x"537a527e",
          5995 => x"51ff9bd7",
          5996 => x"3f815681",
          5997 => x"fef00883",
          5998 => x"e7387d83",
          5999 => x"2e098106",
          6000 => x"80ee3875",
          6001 => x"54608605",
          6002 => x"537a527e",
          6003 => x"51ff9bb7",
          6004 => x"3f848053",
          6005 => x"80527a51",
          6006 => x"ff9fed3f",
          6007 => x"848b85a4",
          6008 => x"d2527a51",
          6009 => x"ff9f8f3f",
          6010 => x"868a85e4",
          6011 => x"f25283e4",
          6012 => x"1b51ff9f",
          6013 => x"813fff18",
          6014 => x"5283e81b",
          6015 => x"51ff9ef6",
          6016 => x"3f825283",
          6017 => x"ec1b51ff",
          6018 => x"9eec3f82",
          6019 => x"d4d55278",
          6020 => x"51ff9ec4",
          6021 => x"3f755460",
          6022 => x"8705537a",
          6023 => x"527e51ff",
          6024 => x"9ae53f75",
          6025 => x"54601653",
          6026 => x"7a527e51",
          6027 => x"ff9ad83f",
          6028 => x"65538052",
          6029 => x"7a51ff9f",
          6030 => x"8f3f7f56",
          6031 => x"80587d83",
          6032 => x"2e098106",
          6033 => x"9a38f852",
          6034 => x"7a51ff9e",
          6035 => x"a93fff52",
          6036 => x"841b51ff",
          6037 => x"9ea03ff0",
          6038 => x"0a52881b",
          6039 => x"51913987",
          6040 => x"fffff855",
          6041 => x"7d812e83",
          6042 => x"38f85574",
          6043 => x"527a51ff",
          6044 => x"9e843f7c",
          6045 => x"55615774",
          6046 => x"62268338",
          6047 => x"74577654",
          6048 => x"75537a52",
          6049 => x"7e51ff99",
          6050 => x"fe3f81fe",
          6051 => x"f0088287",
          6052 => x"38848053",
          6053 => x"81fef008",
          6054 => x"527a51ff",
          6055 => x"9eaa3f76",
          6056 => x"16757831",
          6057 => x"565674cd",
          6058 => x"38811858",
          6059 => x"77802eff",
          6060 => x"8d387955",
          6061 => x"7d832e83",
          6062 => x"38635561",
          6063 => x"57746226",
          6064 => x"83387457",
          6065 => x"76547553",
          6066 => x"7a527e51",
          6067 => x"ff99b83f",
          6068 => x"81fef008",
          6069 => x"81c13876",
          6070 => x"16757831",
          6071 => x"565674db",
          6072 => x"388c567d",
          6073 => x"832e9338",
          6074 => x"86566683",
          6075 => x"ffff268a",
          6076 => x"3884567d",
          6077 => x"822e8338",
          6078 => x"81566481",
          6079 => x"06587780",
          6080 => x"fe388480",
          6081 => x"5377527a",
          6082 => x"51ff9dbc",
          6083 => x"3f82d4d5",
          6084 => x"527851ff",
          6085 => x"9cc23f83",
          6086 => x"be1b5577",
          6087 => x"7534810b",
          6088 => x"81163481",
          6089 => x"0b821634",
          6090 => x"77831634",
          6091 => x"75841634",
          6092 => x"60670556",
          6093 => x"80fdc152",
          6094 => x"7551fed4",
          6095 => x"ee3ffe0b",
          6096 => x"85163481",
          6097 => x"fef00882",
          6098 => x"2abf0756",
          6099 => x"75861634",
          6100 => x"81fef008",
          6101 => x"87163460",
          6102 => x"5283c61b",
          6103 => x"51ff9c96",
          6104 => x"3f665283",
          6105 => x"ca1b51ff",
          6106 => x"9c8c3f81",
          6107 => x"5477537a",
          6108 => x"527e51ff",
          6109 => x"98913f81",
          6110 => x"5681fef0",
          6111 => x"08a23880",
          6112 => x"5380527e",
          6113 => x"51ff99e3",
          6114 => x"3f815681",
          6115 => x"fef00890",
          6116 => x"3889398e",
          6117 => x"568a3981",
          6118 => x"56863981",
          6119 => x"fef00856",
          6120 => x"7581fef0",
          6121 => x"0c993d0d",
          6122 => x"04f53d0d",
          6123 => x"7d605b59",
          6124 => x"807960ff",
          6125 => x"055a5757",
          6126 => x"767825b4",
          6127 => x"388d3df8",
          6128 => x"11555581",
          6129 => x"53fc1552",
          6130 => x"7951c9dc",
          6131 => x"3f7a812e",
          6132 => x"0981069c",
          6133 => x"388c3d33",
          6134 => x"55748d2e",
          6135 => x"db387476",
          6136 => x"70810558",
          6137 => x"34811757",
          6138 => x"748a2e09",
          6139 => x"8106c938",
          6140 => x"80763478",
          6141 => x"55768338",
          6142 => x"76557481",
          6143 => x"fef00c8d",
          6144 => x"3d0d04f7",
          6145 => x"3d0d7b02",
          6146 => x"8405b305",
          6147 => x"33595777",
          6148 => x"8a2e0981",
          6149 => x"0687388d",
          6150 => x"527651e7",
          6151 => x"3f841708",
          6152 => x"56807624",
          6153 => x"be388817",
          6154 => x"0877178c",
          6155 => x"05565977",
          6156 => x"75348116",
          6157 => x"56bb7625",
          6158 => x"a1388b3d",
          6159 => x"fc055475",
          6160 => x"538c1752",
          6161 => x"760851cb",
          6162 => x"dc3f7976",
          6163 => x"32703070",
          6164 => x"72079f2a",
          6165 => x"70305351",
          6166 => x"56567584",
          6167 => x"180c8119",
          6168 => x"88180c8b",
          6169 => x"3d0d04f9",
          6170 => x"3d0d7984",
          6171 => x"11085656",
          6172 => x"807524a7",
          6173 => x"38893dfc",
          6174 => x"05547453",
          6175 => x"8c165275",
          6176 => x"0851cba1",
          6177 => x"3f81fef0",
          6178 => x"08913884",
          6179 => x"1608782e",
          6180 => x"09810687",
          6181 => x"38881608",
          6182 => x"558339ff",
          6183 => x"557481fe",
          6184 => x"f00c893d",
          6185 => x"0d04fd3d",
          6186 => x"0d755480",
          6187 => x"cc538052",
          6188 => x"7351ff9a",
          6189 => x"933f7674",
          6190 => x"0c853d0d",
          6191 => x"04ea3d0d",
          6192 => x"0280e305",
          6193 => x"336a5386",
          6194 => x"3d705354",
          6195 => x"54d83f73",
          6196 => x"527251fe",
          6197 => x"ae3f7251",
          6198 => x"ff8d3f98",
          6199 => x"3d0d04f8",
          6200 => x"3d0d7a70",
          6201 => x"08705656",
          6202 => x"5974802e",
          6203 => x"80e1388c",
          6204 => x"39771579",
          6205 => x"0c851633",
          6206 => x"5480d439",
          6207 => x"74335473",
          6208 => x"a02e0981",
          6209 => x"06863881",
          6210 => x"1555f139",
          6211 => x"80577690",
          6212 => x"2981fbe0",
          6213 => x"05700852",
          6214 => x"56fedab1",
          6215 => x"3f81fef0",
          6216 => x"0881fef0",
          6217 => x"08547553",
          6218 => x"76085258",
          6219 => x"fedaff3f",
          6220 => x"81fef008",
          6221 => x"8b388416",
          6222 => x"33547381",
          6223 => x"2effb238",
          6224 => x"81177081",
          6225 => x"ff065854",
          6226 => x"987727c2",
          6227 => x"38ff5473",
          6228 => x"81fef00c",
          6229 => x"8a3d0d04",
          6230 => x"ff3d0d73",
          6231 => x"52719326",
          6232 => x"818e3871",
          6233 => x"842981e2",
          6234 => x"84055271",
          6235 => x"080481ee",
          6236 => x"b8518180",
          6237 => x"3981eec4",
          6238 => x"5180f939",
          6239 => x"81eed851",
          6240 => x"80f23981",
          6241 => x"eeec5180",
          6242 => x"eb3981ee",
          6243 => x"fc5180e4",
          6244 => x"3981ef8c",
          6245 => x"5180dd39",
          6246 => x"81efa051",
          6247 => x"80d63981",
          6248 => x"efb05180",
          6249 => x"cf3981ef",
          6250 => x"c85180c8",
          6251 => x"3981efe0",
          6252 => x"5180c139",
          6253 => x"81eff851",
          6254 => x"bb3981f0",
          6255 => x"9451b539",
          6256 => x"81f0a851",
          6257 => x"af3981f0",
          6258 => x"d451a939",
          6259 => x"81f0e851",
          6260 => x"a33981f1",
          6261 => x"88519d39",
          6262 => x"81f19c51",
          6263 => x"973981f1",
          6264 => x"b4519139",
          6265 => x"81f1cc51",
          6266 => x"8b3981f1",
          6267 => x"e4518539",
          6268 => x"81f1f051",
          6269 => x"fef2ae3f",
          6270 => x"833d0d04",
          6271 => x"fb3d0d77",
          6272 => x"79565674",
          6273 => x"87e7268a",
          6274 => x"38745275",
          6275 => x"87e82951",
          6276 => x"913987e8",
          6277 => x"527451fe",
          6278 => x"cf913f81",
          6279 => x"fef00852",
          6280 => x"7551fecf",
          6281 => x"863f81fe",
          6282 => x"f0085479",
          6283 => x"53755281",
          6284 => x"f28051fe",
          6285 => x"f7d33f87",
          6286 => x"3d0d04ec",
          6287 => x"3d0d6602",
          6288 => x"840580e3",
          6289 => x"05335b57",
          6290 => x"80687830",
          6291 => x"707a0773",
          6292 => x"25515759",
          6293 => x"59785677",
          6294 => x"87ff2683",
          6295 => x"38815674",
          6296 => x"76077081",
          6297 => x"ff065155",
          6298 => x"93567481",
          6299 => x"80388153",
          6300 => x"76528c3d",
          6301 => x"705256ff",
          6302 => x"bfc93f81",
          6303 => x"fef00857",
          6304 => x"81fef008",
          6305 => x"b83881fe",
          6306 => x"f00887c0",
          6307 => x"98880c81",
          6308 => x"fef00859",
          6309 => x"963dd405",
          6310 => x"54848053",
          6311 => x"77527551",
          6312 => x"c4863f81",
          6313 => x"fef00857",
          6314 => x"81fef008",
          6315 => x"90387a55",
          6316 => x"74802e89",
          6317 => x"38741975",
          6318 => x"195959d8",
          6319 => x"39963dd8",
          6320 => x"0551cbf0",
          6321 => x"3f763070",
          6322 => x"78078025",
          6323 => x"7b30709f",
          6324 => x"2a720651",
          6325 => x"57515674",
          6326 => x"802e9038",
          6327 => x"81f2a453",
          6328 => x"87c09888",
          6329 => x"08527851",
          6330 => x"fe923f76",
          6331 => x"567581fe",
          6332 => x"f00c963d",
          6333 => x"0d04f93d",
          6334 => x"0d7b0284",
          6335 => x"05b30533",
          6336 => x"5758ff57",
          6337 => x"80537a52",
          6338 => x"7951feaf",
          6339 => x"3f81fef0",
          6340 => x"08a43875",
          6341 => x"802e8838",
          6342 => x"75812e98",
          6343 => x"38983960",
          6344 => x"557f5481",
          6345 => x"fef0537e",
          6346 => x"527d5177",
          6347 => x"2d81fef0",
          6348 => x"08578339",
          6349 => x"77047681",
          6350 => x"fef00c89",
          6351 => x"3d0d04f3",
          6352 => x"3d0d7f61",
          6353 => x"63028c05",
          6354 => x"80cf0533",
          6355 => x"73731568",
          6356 => x"415f5c5c",
          6357 => x"5e5e5e7a",
          6358 => x"5281f2ac",
          6359 => x"51fef5a9",
          6360 => x"3f81f2b4",
          6361 => x"51feefbd",
          6362 => x"3f805574",
          6363 => x"792780fc",
          6364 => x"387b902e",
          6365 => x"89387ba0",
          6366 => x"2ea73880",
          6367 => x"c6397418",
          6368 => x"53727a27",
          6369 => x"8e387222",
          6370 => x"5281f2b8",
          6371 => x"51fef4f9",
          6372 => x"3f893981",
          6373 => x"f2c451fe",
          6374 => x"ef8b3f82",
          6375 => x"155580c3",
          6376 => x"39741853",
          6377 => x"727a278e",
          6378 => x"38720852",
          6379 => x"81f2ac51",
          6380 => x"fef4d63f",
          6381 => x"893981f2",
          6382 => x"c051feee",
          6383 => x"e83f8415",
          6384 => x"55a13974",
          6385 => x"1853727a",
          6386 => x"278e3872",
          6387 => x"335281f2",
          6388 => x"cc51fef4",
          6389 => x"b43f8939",
          6390 => x"81f2d451",
          6391 => x"feeec63f",
          6392 => x"811555a0",
          6393 => x"51feede0",
          6394 => x"3fff8039",
          6395 => x"81f2d851",
          6396 => x"feeeb23f",
          6397 => x"80557479",
          6398 => x"27bc3874",
          6399 => x"18703355",
          6400 => x"53805672",
          6401 => x"7a278338",
          6402 => x"81568053",
          6403 => x"9f742783",
          6404 => x"38815375",
          6405 => x"73067081",
          6406 => x"ff065153",
          6407 => x"72802e8b",
          6408 => x"387380fe",
          6409 => x"26853873",
          6410 => x"518339a0",
          6411 => x"51feed98",
          6412 => x"3f811555",
          6413 => x"c13981f2",
          6414 => x"dc51feed",
          6415 => x"e83f7818",
          6416 => x"791c5c58",
          6417 => x"fede963f",
          6418 => x"81fef008",
          6419 => x"982b7098",
          6420 => x"2c515776",
          6421 => x"a02e0981",
          6422 => x"06ab38fe",
          6423 => x"ddff3f81",
          6424 => x"fef00898",
          6425 => x"2b70982c",
          6426 => x"70a03270",
          6427 => x"30729b32",
          6428 => x"70307072",
          6429 => x"07737507",
          6430 => x"06515858",
          6431 => x"59575157",
          6432 => x"807324d7",
          6433 => x"38769b2e",
          6434 => x"09810685",
          6435 => x"3880538c",
          6436 => x"397c1e53",
          6437 => x"727826fd",
          6438 => x"be38ff53",
          6439 => x"7281fef0",
          6440 => x"0c8f3d0d",
          6441 => x"04fc3d0d",
          6442 => x"029b0533",
          6443 => x"81f2e053",
          6444 => x"81f2e852",
          6445 => x"55fef2d1",
          6446 => x"3f81faa0",
          6447 => x"2251fee6",
          6448 => x"d73f81f2",
          6449 => x"f45481f3",
          6450 => x"805381fa",
          6451 => x"a1335281",
          6452 => x"f38851fe",
          6453 => x"f2b33f74",
          6454 => x"802e8538",
          6455 => x"fee2a23f",
          6456 => x"863d0d04",
          6457 => x"fe3d0d87",
          6458 => x"c0968008",
          6459 => x"53fee7b1",
          6460 => x"3f8151fe",
          6461 => x"d8fb3f81",
          6462 => x"f3a451fe",
          6463 => x"daf33f80",
          6464 => x"51fed8ed",
          6465 => x"3f72812a",
          6466 => x"70810651",
          6467 => x"5271802e",
          6468 => x"95388151",
          6469 => x"fed8da3f",
          6470 => x"81f3c051",
          6471 => x"fedad23f",
          6472 => x"8051fed8",
          6473 => x"cc3f7282",
          6474 => x"2a708106",
          6475 => x"51527180",
          6476 => x"2e953881",
          6477 => x"51fed8b9",
          6478 => x"3f81f3d4",
          6479 => x"51fedab1",
          6480 => x"3f8051fe",
          6481 => x"d8ab3f72",
          6482 => x"832a7081",
          6483 => x"06515271",
          6484 => x"802e9538",
          6485 => x"8151fed8",
          6486 => x"983f81f3",
          6487 => x"e451feda",
          6488 => x"903f8051",
          6489 => x"fed88a3f",
          6490 => x"72842a70",
          6491 => x"81065152",
          6492 => x"71802e95",
          6493 => x"388151fe",
          6494 => x"d7f73f81",
          6495 => x"f3f851fe",
          6496 => x"d9ef3f80",
          6497 => x"51fed7e9",
          6498 => x"3f72852a",
          6499 => x"70810651",
          6500 => x"5271802e",
          6501 => x"95388151",
          6502 => x"fed7d63f",
          6503 => x"81f48c51",
          6504 => x"fed9ce3f",
          6505 => x"8051fed7",
          6506 => x"c83f7286",
          6507 => x"2a708106",
          6508 => x"51527180",
          6509 => x"2e953881",
          6510 => x"51fed7b5",
          6511 => x"3f81f4a0",
          6512 => x"51fed9ad",
          6513 => x"3f8051fe",
          6514 => x"d7a73f72",
          6515 => x"872a7081",
          6516 => x"06515271",
          6517 => x"802e9538",
          6518 => x"8151fed7",
          6519 => x"943f81f4",
          6520 => x"b451fed9",
          6521 => x"8c3f8051",
          6522 => x"fed7863f",
          6523 => x"72882a70",
          6524 => x"81065152",
          6525 => x"71802e95",
          6526 => x"388151fe",
          6527 => x"d6f33f81",
          6528 => x"f4c851fe",
          6529 => x"d8eb3f80",
          6530 => x"51fed6e5",
          6531 => x"3ffee599",
          6532 => x"3f843d0d",
          6533 => x"04fb3d0d",
          6534 => x"77028405",
          6535 => x"a3053370",
          6536 => x"55565680",
          6537 => x"527551fe",
          6538 => x"cea33f81",
          6539 => x"fbdc3354",
          6540 => x"73a73881",
          6541 => x"5381f588",
          6542 => x"52829688",
          6543 => x"51ffb883",
          6544 => x"3f81fef0",
          6545 => x"08307081",
          6546 => x"fef00807",
          6547 => x"80258271",
          6548 => x"31515154",
          6549 => x"7381fbdc",
          6550 => x"3481fbdc",
          6551 => x"33547381",
          6552 => x"2e098106",
          6553 => x"ac388296",
          6554 => x"88537452",
          6555 => x"7551f2b9",
          6556 => x"3f81fef0",
          6557 => x"08802e8c",
          6558 => x"3881fef0",
          6559 => x"0851fee9",
          6560 => x"a43f8e39",
          6561 => x"82968851",
          6562 => x"c4aa3f82",
          6563 => x"0b81fbdc",
          6564 => x"3481fbdc",
          6565 => x"33547382",
          6566 => x"2e098106",
          6567 => x"89387452",
          6568 => x"7551fefa",
          6569 => x"e43f800b",
          6570 => x"81fef00c",
          6571 => x"873d0d04",
          6572 => x"ce3d0d80",
          6573 => x"70718296",
          6574 => x"840c5f5d",
          6575 => x"81527c51",
          6576 => x"ff86db3f",
          6577 => x"81fef008",
          6578 => x"81ff0659",
          6579 => x"787d2e09",
          6580 => x"8106a238",
          6581 => x"81f59852",
          6582 => x"963d7052",
          6583 => x"59feeebf",
          6584 => x"3f7c5378",
          6585 => x"528280b4",
          6586 => x"51ffb5f6",
          6587 => x"3f81fef0",
          6588 => x"087d2e88",
          6589 => x"3881f59c",
          6590 => x"5191fe39",
          6591 => x"81705f5d",
          6592 => x"81f5d451",
          6593 => x"fee89e3f",
          6594 => x"963d7046",
          6595 => x"5a80f852",
          6596 => x"7951fe81",
          6597 => x"3fb43dff",
          6598 => x"840551f3",
          6599 => x"c23f81fe",
          6600 => x"f008902b",
          6601 => x"70902c51",
          6602 => x"597880c1",
          6603 => x"2e89f138",
          6604 => x"7880c124",
          6605 => x"80d93878",
          6606 => x"ab2e83c0",
          6607 => x"3878ab24",
          6608 => x"a4387882",
          6609 => x"2e81b338",
          6610 => x"7882248a",
          6611 => x"3878802e",
          6612 => x"ffae388f",
          6613 => x"a5397884",
          6614 => x"2e828638",
          6615 => x"78942e82",
          6616 => x"b1388f96",
          6617 => x"3978bd2e",
          6618 => x"858c3878",
          6619 => x"bd249038",
          6620 => x"78b02e83",
          6621 => x"af3878bc",
          6622 => x"2e849138",
          6623 => x"8efc3978",
          6624 => x"bf2e85d7",
          6625 => x"387880c0",
          6626 => x"2e86d238",
          6627 => x"8eec3978",
          6628 => x"80d52e8d",
          6629 => x"c2387880",
          6630 => x"d524b038",
          6631 => x"7880d02e",
          6632 => x"8cf63878",
          6633 => x"80d02492",
          6634 => x"387880c2",
          6635 => x"2e8a9938",
          6636 => x"7880c32e",
          6637 => x"8bc2388e",
          6638 => x"c1397880",
          6639 => x"d12e8ce9",
          6640 => x"387880d4",
          6641 => x"2e8cf338",
          6642 => x"8eb03978",
          6643 => x"81822e8e",
          6644 => x"86387881",
          6645 => x"82249238",
          6646 => x"7880f82e",
          6647 => x"8d963878",
          6648 => x"80f92e8d",
          6649 => x"b4388e92",
          6650 => x"39788183",
          6651 => x"2e8df738",
          6652 => x"7881852e",
          6653 => x"8dfd388e",
          6654 => x"8139b43d",
          6655 => x"ff801153",
          6656 => x"ff840551",
          6657 => x"feedf73f",
          6658 => x"81fef008",
          6659 => x"883881f5",
          6660 => x"d8518fe5",
          6661 => x"39b43dfe",
          6662 => x"fc1153ff",
          6663 => x"840551fe",
          6664 => x"eddc3f81",
          6665 => x"fef00880",
          6666 => x"2e883881",
          6667 => x"63258338",
          6668 => x"80430280",
          6669 => x"cb053352",
          6670 => x"0280cf05",
          6671 => x"3351ff83",
          6672 => x"dd3f81fe",
          6673 => x"f00881ff",
          6674 => x"0659788e",
          6675 => x"3881f5e8",
          6676 => x"51fee5d1",
          6677 => x"3f815efd",
          6678 => x"a73981f5",
          6679 => x"f85187b9",
          6680 => x"39b43dff",
          6681 => x"801153ff",
          6682 => x"840551fe",
          6683 => x"ed903f81",
          6684 => x"fef00880",
          6685 => x"2efd8938",
          6686 => x"80538052",
          6687 => x"0280cf05",
          6688 => x"3351ff87",
          6689 => x"e63f81fe",
          6690 => x"f0085281",
          6691 => x"f690518c",
          6692 => x"bf39b43d",
          6693 => x"ff801153",
          6694 => x"ff840551",
          6695 => x"feecdf3f",
          6696 => x"81fef008",
          6697 => x"802e8738",
          6698 => x"638926fc",
          6699 => x"d338b43d",
          6700 => x"fefc1153",
          6701 => x"ff840551",
          6702 => x"feecc33f",
          6703 => x"81fef008",
          6704 => x"863881fe",
          6705 => x"f0084363",
          6706 => x"5381f698",
          6707 => x"527951fe",
          6708 => x"eacd3f02",
          6709 => x"80cb0533",
          6710 => x"53795263",
          6711 => x"84b42982",
          6712 => x"80b40551",
          6713 => x"ffb1fb3f",
          6714 => x"81fef008",
          6715 => x"81933881",
          6716 => x"f5e851fe",
          6717 => x"e4af3f81",
          6718 => x"5dfc8539",
          6719 => x"b43dff84",
          6720 => x"0551fecd",
          6721 => x"9d3f81fe",
          6722 => x"f008b53d",
          6723 => x"ff840552",
          6724 => x"5bfecdf0",
          6725 => x"3f815381",
          6726 => x"fef00852",
          6727 => x"7a51f29b",
          6728 => x"3f80d539",
          6729 => x"b43dff84",
          6730 => x"0551fecc",
          6731 => x"f53f81fe",
          6732 => x"f008b53d",
          6733 => x"ff840552",
          6734 => x"5bfecdc8",
          6735 => x"3f81fef0",
          6736 => x"08b53dff",
          6737 => x"8405525a",
          6738 => x"fecdb93f",
          6739 => x"81fef008",
          6740 => x"b53dff84",
          6741 => x"055259fe",
          6742 => x"cdaa3f81",
          6743 => x"f9ec5881",
          6744 => x"ffb85780",
          6745 => x"56805581",
          6746 => x"fef00881",
          6747 => x"ff065478",
          6748 => x"5379527a",
          6749 => x"51f2ff3f",
          6750 => x"81fef008",
          6751 => x"802efb80",
          6752 => x"3881fef0",
          6753 => x"0851efd0",
          6754 => x"3ffaf539",
          6755 => x"b43dff80",
          6756 => x"1153ff84",
          6757 => x"0551feea",
          6758 => x"e53f81fe",
          6759 => x"f008802e",
          6760 => x"fade38b4",
          6761 => x"3dfefc11",
          6762 => x"53ff8405",
          6763 => x"51feeace",
          6764 => x"3f81fef0",
          6765 => x"08802efa",
          6766 => x"c738b43d",
          6767 => x"fef81153",
          6768 => x"ff840551",
          6769 => x"feeab73f",
          6770 => x"81fef008",
          6771 => x"863881fe",
          6772 => x"f0084281",
          6773 => x"f69c51fe",
          6774 => x"e2cb3f63",
          6775 => x"635c5a79",
          6776 => x"7b2781f2",
          6777 => x"38615978",
          6778 => x"7a708405",
          6779 => x"5c0c7a7a",
          6780 => x"26f53881",
          6781 => x"e139b43d",
          6782 => x"ff801153",
          6783 => x"ff840551",
          6784 => x"fee9fb3f",
          6785 => x"81fef008",
          6786 => x"802ef9f4",
          6787 => x"38b43dfe",
          6788 => x"fc1153ff",
          6789 => x"840551fe",
          6790 => x"e9e43f81",
          6791 => x"fef00880",
          6792 => x"2ef9dd38",
          6793 => x"b43dfef8",
          6794 => x"1153ff84",
          6795 => x"0551fee9",
          6796 => x"cd3f81fe",
          6797 => x"f008802e",
          6798 => x"f9c63881",
          6799 => x"f6ac51fe",
          6800 => x"e1e33f63",
          6801 => x"5a796327",
          6802 => x"818c3861",
          6803 => x"59797081",
          6804 => x"055b3379",
          6805 => x"34618105",
          6806 => x"42eb39b4",
          6807 => x"3dff8011",
          6808 => x"53ff8405",
          6809 => x"51fee996",
          6810 => x"3f81fef0",
          6811 => x"08802ef9",
          6812 => x"8f38b43d",
          6813 => x"fefc1153",
          6814 => x"ff840551",
          6815 => x"fee8ff3f",
          6816 => x"81fef008",
          6817 => x"802ef8f8",
          6818 => x"38b43dfe",
          6819 => x"f81153ff",
          6820 => x"840551fe",
          6821 => x"e8e83f81",
          6822 => x"fef00880",
          6823 => x"2ef8e138",
          6824 => x"81f6b851",
          6825 => x"fee0fe3f",
          6826 => x"635a7963",
          6827 => x"27a83861",
          6828 => x"70337b33",
          6829 => x"5e5a5b78",
          6830 => x"7c2e9238",
          6831 => x"78557a54",
          6832 => x"79335379",
          6833 => x"5281f6c8",
          6834 => x"51fee6bd",
          6835 => x"3f811a62",
          6836 => x"8105435a",
          6837 => x"d53981f5",
          6838 => x"e45182bd",
          6839 => x"39b43dff",
          6840 => x"801153ff",
          6841 => x"840551fe",
          6842 => x"e8943f81",
          6843 => x"fef00880",
          6844 => x"df3881fa",
          6845 => x"b4335978",
          6846 => x"802e8938",
          6847 => x"81f9ec08",
          6848 => x"4480cd39",
          6849 => x"81fab533",
          6850 => x"5978802e",
          6851 => x"883881f9",
          6852 => x"f40844bc",
          6853 => x"3981fab6",
          6854 => x"33597880",
          6855 => x"2e883881",
          6856 => x"f9fc0844",
          6857 => x"ab3981fa",
          6858 => x"b7335978",
          6859 => x"802e8838",
          6860 => x"81fa8408",
          6861 => x"449a3981",
          6862 => x"fab23359",
          6863 => x"78802e88",
          6864 => x"3881fa8c",
          6865 => x"08448939",
          6866 => x"81fa9c08",
          6867 => x"fc800544",
          6868 => x"b43dfefc",
          6869 => x"1153ff84",
          6870 => x"0551fee7",
          6871 => x"a13f81fe",
          6872 => x"f00880de",
          6873 => x"3881fab4",
          6874 => x"33597880",
          6875 => x"2e893881",
          6876 => x"f9f00843",
          6877 => x"80cc3981",
          6878 => x"fab53359",
          6879 => x"78802e88",
          6880 => x"3881f9f8",
          6881 => x"0843bb39",
          6882 => x"81fab633",
          6883 => x"5978802e",
          6884 => x"883881fa",
          6885 => x"800843aa",
          6886 => x"3981fab7",
          6887 => x"33597880",
          6888 => x"2e883881",
          6889 => x"fa880843",
          6890 => x"993981fa",
          6891 => x"b2335978",
          6892 => x"802e8838",
          6893 => x"81fa9008",
          6894 => x"43883981",
          6895 => x"fa9c0888",
          6896 => x"0543b43d",
          6897 => x"fef81153",
          6898 => x"ff840551",
          6899 => x"fee6af3f",
          6900 => x"81fef008",
          6901 => x"802ea738",
          6902 => x"80625c5c",
          6903 => x"7a882e83",
          6904 => x"38815c7a",
          6905 => x"90327030",
          6906 => x"7072079f",
          6907 => x"2a707f06",
          6908 => x"51515a5a",
          6909 => x"78802e88",
          6910 => x"387aa02e",
          6911 => x"83388842",
          6912 => x"81f6e451",
          6913 => x"fede9e3f",
          6914 => x"a0556354",
          6915 => x"61536252",
          6916 => x"6351eeab",
          6917 => x"3f81f6f4",
          6918 => x"51fede89",
          6919 => x"3ff5e139",
          6920 => x"b43dff80",
          6921 => x"1153ff84",
          6922 => x"0551fee5",
          6923 => x"d13f81fe",
          6924 => x"f008802e",
          6925 => x"f5ca38b4",
          6926 => x"3dfefc11",
          6927 => x"53ff8405",
          6928 => x"51fee5ba",
          6929 => x"3f81fef0",
          6930 => x"08802ea5",
          6931 => x"38635902",
          6932 => x"80cb0533",
          6933 => x"79346381",
          6934 => x"0544b43d",
          6935 => x"fefc1153",
          6936 => x"ff840551",
          6937 => x"fee5973f",
          6938 => x"81fef008",
          6939 => x"e038f590",
          6940 => x"39637033",
          6941 => x"545281f7",
          6942 => x"8051fee3",
          6943 => x"8c3f80f8",
          6944 => x"527951fe",
          6945 => x"e3dd3f79",
          6946 => x"45793359",
          6947 => x"78ae2ef4",
          6948 => x"ef389f79",
          6949 => x"27a038b4",
          6950 => x"3dfefc11",
          6951 => x"53ff8405",
          6952 => x"51fee4da",
          6953 => x"3f81fef0",
          6954 => x"08802e91",
          6955 => x"38635902",
          6956 => x"80cb0533",
          6957 => x"79346381",
          6958 => x"0544ffb5",
          6959 => x"3981f78c",
          6960 => x"51fedce1",
          6961 => x"3fffaa39",
          6962 => x"b43dfef4",
          6963 => x"1153ff84",
          6964 => x"0551fee6",
          6965 => x"9b3f81fe",
          6966 => x"f008802e",
          6967 => x"f4a238b4",
          6968 => x"3dfef011",
          6969 => x"53ff8405",
          6970 => x"51fee684",
          6971 => x"3f81fef0",
          6972 => x"08802ea6",
          6973 => x"38605902",
          6974 => x"be052279",
          6975 => x"7082055b",
          6976 => x"237841b4",
          6977 => x"3dfef011",
          6978 => x"53ff8405",
          6979 => x"51fee5e0",
          6980 => x"3f81fef0",
          6981 => x"08df38f3",
          6982 => x"e7396070",
          6983 => x"22545281",
          6984 => x"f79451fe",
          6985 => x"e1e33f80",
          6986 => x"f8527951",
          6987 => x"fee2b43f",
          6988 => x"79457933",
          6989 => x"5978ae2e",
          6990 => x"f3c63878",
          6991 => x"9f268738",
          6992 => x"60820541",
          6993 => x"d539b43d",
          6994 => x"fef01153",
          6995 => x"ff840551",
          6996 => x"fee59d3f",
          6997 => x"81fef008",
          6998 => x"802e9238",
          6999 => x"605902be",
          7000 => x"05227970",
          7001 => x"82055b23",
          7002 => x"7841ffae",
          7003 => x"3981f78c",
          7004 => x"51fedbb1",
          7005 => x"3fffa339",
          7006 => x"b43dfef4",
          7007 => x"1153ff84",
          7008 => x"0551fee4",
          7009 => x"eb3f81fe",
          7010 => x"f008802e",
          7011 => x"f2f238b4",
          7012 => x"3dfef011",
          7013 => x"53ff8405",
          7014 => x"51fee4d4",
          7015 => x"3f81fef0",
          7016 => x"08802ea1",
          7017 => x"38606071",
          7018 => x"0c596084",
          7019 => x"0541b43d",
          7020 => x"fef01153",
          7021 => x"ff840551",
          7022 => x"fee4b53f",
          7023 => x"81fef008",
          7024 => x"e438f2bc",
          7025 => x"39607008",
          7026 => x"545281f7",
          7027 => x"a051fee0",
          7028 => x"b83f80f8",
          7029 => x"527951fe",
          7030 => x"e1893f79",
          7031 => x"45793359",
          7032 => x"78ae2ef2",
          7033 => x"9b389f79",
          7034 => x"279c38b4",
          7035 => x"3dfef011",
          7036 => x"53ff8405",
          7037 => x"51fee3f8",
          7038 => x"3f81fef0",
          7039 => x"08802e8d",
          7040 => x"38606071",
          7041 => x"0c596084",
          7042 => x"0541ffb9",
          7043 => x"3981f78c",
          7044 => x"51feda91",
          7045 => x"3fffae39",
          7046 => x"81f7ac51",
          7047 => x"feda863f",
          7048 => x"8251fed4",
          7049 => x"d73ff1d8",
          7050 => x"3981f7c4",
          7051 => x"51fed9f5",
          7052 => x"3fa251fe",
          7053 => x"d4aa3ff1",
          7054 => x"c73981f7",
          7055 => x"dc51fed9",
          7056 => x"e43f8480",
          7057 => x"810b87c0",
          7058 => x"94840c84",
          7059 => x"80810b87",
          7060 => x"c094940c",
          7061 => x"f1aa3981",
          7062 => x"f7f051fe",
          7063 => x"d9c73f8c",
          7064 => x"80830b87",
          7065 => x"c094840c",
          7066 => x"8c80830b",
          7067 => x"87c09494",
          7068 => x"0cf18d39",
          7069 => x"b43dff80",
          7070 => x"1153ff84",
          7071 => x"0551fee0",
          7072 => x"fd3f81fe",
          7073 => x"f008802e",
          7074 => x"f0f63863",
          7075 => x"5281f884",
          7076 => x"51fedef5",
          7077 => x"3f635978",
          7078 => x"04b43dff",
          7079 => x"801153ff",
          7080 => x"840551fe",
          7081 => x"e0d83f81",
          7082 => x"fef00880",
          7083 => x"2ef0d138",
          7084 => x"635281f8",
          7085 => x"a051fede",
          7086 => x"d03f6359",
          7087 => x"782d81fe",
          7088 => x"f008802e",
          7089 => x"f0ba3881",
          7090 => x"fef00852",
          7091 => x"81f8bc51",
          7092 => x"fedeb63f",
          7093 => x"f0aa3981",
          7094 => x"f8d851fe",
          7095 => x"d8c73ffe",
          7096 => x"b5aa3ff0",
          7097 => x"9b3981f8",
          7098 => x"f451fed8",
          7099 => x"b83f8059",
          7100 => x"ffa539fe",
          7101 => x"ce8b3ff0",
          7102 => x"87397945",
          7103 => x"79335978",
          7104 => x"802eeffc",
          7105 => x"387d7d06",
          7106 => x"5978802e",
          7107 => x"81d338b4",
          7108 => x"3dff8405",
          7109 => x"51fec18a",
          7110 => x"3f81fef0",
          7111 => x"085b815c",
          7112 => x"7b822eb2",
          7113 => x"387b8224",
          7114 => x"89387b81",
          7115 => x"2e8c3880",
          7116 => x"cd397b83",
          7117 => x"2eb03880",
          7118 => x"c53981f9",
          7119 => x"88567a55",
          7120 => x"81f98c54",
          7121 => x"805381f9",
          7122 => x"9052b43d",
          7123 => x"ffb00551",
          7124 => x"feddcc3f",
          7125 => x"bb3981f9",
          7126 => x"b052b43d",
          7127 => x"ffb00551",
          7128 => x"feddbc3f",
          7129 => x"ab397a55",
          7130 => x"81f98c54",
          7131 => x"805381f9",
          7132 => x"a052b43d",
          7133 => x"ffb00551",
          7134 => x"fedda43f",
          7135 => x"93397a54",
          7136 => x"805381f9",
          7137 => x"ac52b43d",
          7138 => x"ffb00551",
          7139 => x"fedd903f",
          7140 => x"81f9ec58",
          7141 => x"81ffb857",
          7142 => x"80566455",
          7143 => x"80548380",
          7144 => x"80538380",
          7145 => x"8052b43d",
          7146 => x"ffb00551",
          7147 => x"e6c83f81",
          7148 => x"fef00881",
          7149 => x"fef00809",
          7150 => x"70307072",
          7151 => x"07802551",
          7152 => x"5b5b5f80",
          7153 => x"5a7b8326",
          7154 => x"8338815a",
          7155 => x"787a0659",
          7156 => x"78802e8d",
          7157 => x"38811c70",
          7158 => x"81ff065d",
          7159 => x"597bfec0",
          7160 => x"387d8132",
          7161 => x"7d813207",
          7162 => x"59788a38",
          7163 => x"7eff2e09",
          7164 => x"8106ee8c",
          7165 => x"3881f9b4",
          7166 => x"51fedc8d",
          7167 => x"3fee8139",
          7168 => x"fc3d0d80",
          7169 => x"0b81ffb8",
          7170 => x"3487c094",
          7171 => x"8c700854",
          7172 => x"55878480",
          7173 => x"527251fe",
          7174 => x"b3913f81",
          7175 => x"fef00890",
          7176 => x"2b750855",
          7177 => x"53878480",
          7178 => x"527351fe",
          7179 => x"b2fd3f72",
          7180 => x"81fef008",
          7181 => x"07750c87",
          7182 => x"c0949c70",
          7183 => x"08545587",
          7184 => x"84805272",
          7185 => x"51feb2e3",
          7186 => x"3f81fef0",
          7187 => x"08902b75",
          7188 => x"08555387",
          7189 => x"84805273",
          7190 => x"51feb2cf",
          7191 => x"3f7281fe",
          7192 => x"f0080775",
          7193 => x"0c8c8083",
          7194 => x"0b87c094",
          7195 => x"840c8c80",
          7196 => x"830b87c0",
          7197 => x"94940ca3",
          7198 => x"8b0b81ff",
          7199 => x"840ca68c",
          7200 => x"0b81ff88",
          7201 => x"0cfec6ad",
          7202 => x"3ffed095",
          7203 => x"3f81f9c4",
          7204 => x"51fed591",
          7205 => x"3f81f9d0",
          7206 => x"51fed589",
          7207 => x"3f81c9e4",
          7208 => x"51fecfb7",
          7209 => x"3f8151e7",
          7210 => x"fc3fec84",
          7211 => x"3f800400",
          7212 => x"00ffffff",
          7213 => x"ff00ffff",
          7214 => x"ffff00ff",
          7215 => x"ffffff00",
          7216 => x"00001832",
          7217 => x"00001838",
          7218 => x"0000183e",
          7219 => x"00001844",
          7220 => x"0000184a",
          7221 => x"000025f6",
          7222 => x"000026d2",
          7223 => x"00002775",
          7224 => x"000027b5",
          7225 => x"000027d8",
          7226 => x"00002865",
          7227 => x"000024cb",
          7228 => x"000024cb",
          7229 => x"000028a2",
          7230 => x"00002918",
          7231 => x"000029a3",
          7232 => x"000029cc",
          7233 => x"000061ea",
          7234 => x"0000616e",
          7235 => x"00006175",
          7236 => x"0000617c",
          7237 => x"00006183",
          7238 => x"0000618a",
          7239 => x"00006191",
          7240 => x"00006198",
          7241 => x"0000619f",
          7242 => x"000061a6",
          7243 => x"000061ad",
          7244 => x"000061b4",
          7245 => x"000061ba",
          7246 => x"000061c0",
          7247 => x"000061c6",
          7248 => x"000061cc",
          7249 => x"000061d2",
          7250 => x"000061d8",
          7251 => x"000061de",
          7252 => x"000061e4",
          7253 => x"25642f25",
          7254 => x"642f2564",
          7255 => x"2025643a",
          7256 => x"25643a25",
          7257 => x"642e2564",
          7258 => x"25640a00",
          7259 => x"536f4320",
          7260 => x"436f6e66",
          7261 => x"69677572",
          7262 => x"6174696f",
          7263 => x"6e000000",
          7264 => x"20286672",
          7265 => x"6f6d2053",
          7266 => x"6f432063",
          7267 => x"6f6e6669",
          7268 => x"67290000",
          7269 => x"3a0a4465",
          7270 => x"76696365",
          7271 => x"7320696d",
          7272 => x"706c656d",
          7273 => x"656e7465",
          7274 => x"643a0a00",
          7275 => x"20202020",
          7276 => x"57422053",
          7277 => x"4452414d",
          7278 => x"20202825",
          7279 => x"3038583a",
          7280 => x"25303858",
          7281 => x"292e0a00",
          7282 => x"20202020",
          7283 => x"53445241",
          7284 => x"4d202020",
          7285 => x"20202825",
          7286 => x"3038583a",
          7287 => x"25303858",
          7288 => x"292e0a00",
          7289 => x"20202020",
          7290 => x"494e534e",
          7291 => x"20425241",
          7292 => x"4d202825",
          7293 => x"3038583a",
          7294 => x"25303858",
          7295 => x"292e0a00",
          7296 => x"20202020",
          7297 => x"4252414d",
          7298 => x"20202020",
          7299 => x"20202825",
          7300 => x"3038583a",
          7301 => x"25303858",
          7302 => x"292e0a00",
          7303 => x"20202020",
          7304 => x"52414d20",
          7305 => x"20202020",
          7306 => x"20202825",
          7307 => x"3038583a",
          7308 => x"25303858",
          7309 => x"292e0a00",
          7310 => x"20202020",
          7311 => x"53442043",
          7312 => x"41524420",
          7313 => x"20202844",
          7314 => x"65766963",
          7315 => x"6573203d",
          7316 => x"25303264",
          7317 => x"292e0a00",
          7318 => x"20202020",
          7319 => x"54494d45",
          7320 => x"52312020",
          7321 => x"20202854",
          7322 => x"696d6572",
          7323 => x"7320203d",
          7324 => x"25303264",
          7325 => x"292e0a00",
          7326 => x"20202020",
          7327 => x"494e5452",
          7328 => x"20435452",
          7329 => x"4c202843",
          7330 => x"68616e6e",
          7331 => x"656c733d",
          7332 => x"25303264",
          7333 => x"292e0a00",
          7334 => x"20202020",
          7335 => x"57495348",
          7336 => x"424f4e45",
          7337 => x"20425553",
          7338 => x"0a000000",
          7339 => x"20202020",
          7340 => x"57422049",
          7341 => x"32430a00",
          7342 => x"20202020",
          7343 => x"494f4354",
          7344 => x"4c0a0000",
          7345 => x"20202020",
          7346 => x"5053320a",
          7347 => x"00000000",
          7348 => x"20202020",
          7349 => x"5350490a",
          7350 => x"00000000",
          7351 => x"41646472",
          7352 => x"65737365",
          7353 => x"733a0a00",
          7354 => x"20202020",
          7355 => x"43505520",
          7356 => x"52657365",
          7357 => x"74205665",
          7358 => x"63746f72",
          7359 => x"20416464",
          7360 => x"72657373",
          7361 => x"203d2025",
          7362 => x"3038580a",
          7363 => x"00000000",
          7364 => x"20202020",
          7365 => x"43505520",
          7366 => x"4d656d6f",
          7367 => x"72792053",
          7368 => x"74617274",
          7369 => x"20416464",
          7370 => x"72657373",
          7371 => x"203d2025",
          7372 => x"3038580a",
          7373 => x"00000000",
          7374 => x"20202020",
          7375 => x"53746163",
          7376 => x"6b205374",
          7377 => x"61727420",
          7378 => x"41646472",
          7379 => x"65737320",
          7380 => x"20202020",
          7381 => x"203d2025",
          7382 => x"3038580a",
          7383 => x"00000000",
          7384 => x"4d697363",
          7385 => x"3a0a0000",
          7386 => x"20202020",
          7387 => x"5a505520",
          7388 => x"49642020",
          7389 => x"20202020",
          7390 => x"20202020",
          7391 => x"20202020",
          7392 => x"20202020",
          7393 => x"203d2025",
          7394 => x"3034580a",
          7395 => x"00000000",
          7396 => x"20202020",
          7397 => x"53797374",
          7398 => x"656d2043",
          7399 => x"6c6f636b",
          7400 => x"20467265",
          7401 => x"71202020",
          7402 => x"20202020",
          7403 => x"203d2025",
          7404 => x"642e2530",
          7405 => x"34644d48",
          7406 => x"7a0a0000",
          7407 => x"20202020",
          7408 => x"53445241",
          7409 => x"4d20436c",
          7410 => x"6f636b20",
          7411 => x"46726571",
          7412 => x"20202020",
          7413 => x"20202020",
          7414 => x"203d2025",
          7415 => x"642e2530",
          7416 => x"34644d48",
          7417 => x"7a0a0000",
          7418 => x"20202020",
          7419 => x"57697368",
          7420 => x"626f6e65",
          7421 => x"20534452",
          7422 => x"414d2043",
          7423 => x"6c6f636b",
          7424 => x"20467265",
          7425 => x"713d2025",
          7426 => x"642e2530",
          7427 => x"34644d48",
          7428 => x"7a0a0000",
          7429 => x"536d616c",
          7430 => x"6c000000",
          7431 => x"4d656469",
          7432 => x"756d0000",
          7433 => x"466c6578",
          7434 => x"00000000",
          7435 => x"45564f00",
          7436 => x"45564f6d",
          7437 => x"696e0000",
          7438 => x"556e6b6e",
          7439 => x"6f776e00",
          7440 => x"68697374",
          7441 => x"6f72792e",
          7442 => x"74787400",
          7443 => x"68697374",
          7444 => x"6f727900",
          7445 => x"68697374",
          7446 => x"00000000",
          7447 => x"21000000",
          7448 => x"25303464",
          7449 => x"20202573",
          7450 => x"0a000000",
          7451 => x"4661696c",
          7452 => x"65642074",
          7453 => x"6f207265",
          7454 => x"73657420",
          7455 => x"74686520",
          7456 => x"68697374",
          7457 => x"6f727920",
          7458 => x"66696c65",
          7459 => x"20746f20",
          7460 => x"454f462e",
          7461 => x"0a000000",
          7462 => x"43616e6e",
          7463 => x"6f74206f",
          7464 => x"70656e2f",
          7465 => x"63726561",
          7466 => x"74652068",
          7467 => x"6973746f",
          7468 => x"72792066",
          7469 => x"696c652c",
          7470 => x"20646973",
          7471 => x"61626c69",
          7472 => x"6e672e0a",
          7473 => x"00000000",
          7474 => x"00007574",
          7475 => x"01000000",
          7476 => x"00000001",
          7477 => x"00007570",
          7478 => x"01000000",
          7479 => x"00000002",
          7480 => x"0000756c",
          7481 => x"04000000",
          7482 => x"00000003",
          7483 => x"00007568",
          7484 => x"04000000",
          7485 => x"00000004",
          7486 => x"00007564",
          7487 => x"04000000",
          7488 => x"00000005",
          7489 => x"00007560",
          7490 => x"04000000",
          7491 => x"00000006",
          7492 => x"0000755c",
          7493 => x"04000000",
          7494 => x"00000007",
          7495 => x"00007558",
          7496 => x"03000000",
          7497 => x"00000008",
          7498 => x"00007554",
          7499 => x"03000000",
          7500 => x"00000009",
          7501 => x"00007550",
          7502 => x"03000000",
          7503 => x"0000000a",
          7504 => x"0000754c",
          7505 => x"03000000",
          7506 => x"0000000b",
          7507 => x"1b5b4400",
          7508 => x"1b5b4300",
          7509 => x"1b5b4200",
          7510 => x"1b5b4100",
          7511 => x"1b5b367e",
          7512 => x"1b5b357e",
          7513 => x"1b5b347e",
          7514 => x"1b5b337e",
          7515 => x"1b5b317e",
          7516 => x"0d000000",
          7517 => x"08000000",
          7518 => x"53440000",
          7519 => x"222a2b2c",
          7520 => x"3a3b3c3d",
          7521 => x"3e3f5b5d",
          7522 => x"7c7f0000",
          7523 => x"46415400",
          7524 => x"46415433",
          7525 => x"32000000",
          7526 => x"ebfe904d",
          7527 => x"53444f53",
          7528 => x"352e3000",
          7529 => x"4e4f204e",
          7530 => x"414d4520",
          7531 => x"20202046",
          7532 => x"41543332",
          7533 => x"20202000",
          7534 => x"4e4f204e",
          7535 => x"414d4520",
          7536 => x"20202046",
          7537 => x"41542020",
          7538 => x"20202000",
          7539 => x"00007578",
          7540 => x"00000000",
          7541 => x"00000000",
          7542 => x"00000000",
          7543 => x"809a4541",
          7544 => x"8e418f80",
          7545 => x"45454549",
          7546 => x"49498e8f",
          7547 => x"9092924f",
          7548 => x"994f5555",
          7549 => x"59999a9b",
          7550 => x"9c9d9e9f",
          7551 => x"41494f55",
          7552 => x"a5a5a6a7",
          7553 => x"a8a9aaab",
          7554 => x"acadaeaf",
          7555 => x"b0b1b2b3",
          7556 => x"b4b5b6b7",
          7557 => x"b8b9babb",
          7558 => x"bcbdbebf",
          7559 => x"c0c1c2c3",
          7560 => x"c4c5c6c7",
          7561 => x"c8c9cacb",
          7562 => x"cccdcecf",
          7563 => x"d0d1d2d3",
          7564 => x"d4d5d6d7",
          7565 => x"d8d9dadb",
          7566 => x"dcdddedf",
          7567 => x"e0e1e2e3",
          7568 => x"e4e5e6e7",
          7569 => x"e8e9eaeb",
          7570 => x"ecedeeef",
          7571 => x"f0f1f2f3",
          7572 => x"f4f5f6f7",
          7573 => x"f8f9fafb",
          7574 => x"fcfdfeff",
          7575 => x"2b2e2c3b",
          7576 => x"3d5b5d2f",
          7577 => x"5c222a3a",
          7578 => x"3c3e3f7c",
          7579 => x"7f000000",
          7580 => x"00010004",
          7581 => x"00100040",
          7582 => x"01000200",
          7583 => x"00000000",
          7584 => x"00010002",
          7585 => x"00040008",
          7586 => x"00100020",
          7587 => x"00000000",
          7588 => x"64696e69",
          7589 => x"74000000",
          7590 => x"64696f63",
          7591 => x"746c0000",
          7592 => x"66696e69",
          7593 => x"74000000",
          7594 => x"666c6f61",
          7595 => x"64000000",
          7596 => x"66657865",
          7597 => x"63000000",
          7598 => x"6d636c65",
          7599 => x"61720000",
          7600 => x"6d636f70",
          7601 => x"79000000",
          7602 => x"6d646966",
          7603 => x"66000000",
          7604 => x"6d64756d",
          7605 => x"70000000",
          7606 => x"6d656200",
          7607 => x"6d656800",
          7608 => x"6d657700",
          7609 => x"68696400",
          7610 => x"68696500",
          7611 => x"68666400",
          7612 => x"68666500",
          7613 => x"63616c6c",
          7614 => x"00000000",
          7615 => x"6a6d7000",
          7616 => x"72657374",
          7617 => x"61727400",
          7618 => x"72657365",
          7619 => x"74000000",
          7620 => x"696e666f",
          7621 => x"00000000",
          7622 => x"74657374",
          7623 => x"00000000",
          7624 => x"74626173",
          7625 => x"69630000",
          7626 => x"6d626173",
          7627 => x"69630000",
          7628 => x"6b696c6f",
          7629 => x"00000000",
          7630 => x"4469736b",
          7631 => x"20457272",
          7632 => x"6f720a00",
          7633 => x"496e7465",
          7634 => x"726e616c",
          7635 => x"20657272",
          7636 => x"6f722e0a",
          7637 => x"00000000",
          7638 => x"4469736b",
          7639 => x"206e6f74",
          7640 => x"20726561",
          7641 => x"64792e0a",
          7642 => x"00000000",
          7643 => x"4e6f2066",
          7644 => x"696c6520",
          7645 => x"666f756e",
          7646 => x"642e0a00",
          7647 => x"4e6f2070",
          7648 => x"61746820",
          7649 => x"666f756e",
          7650 => x"642e0a00",
          7651 => x"496e7661",
          7652 => x"6c696420",
          7653 => x"66696c65",
          7654 => x"6e616d65",
          7655 => x"2e0a0000",
          7656 => x"41636365",
          7657 => x"73732064",
          7658 => x"656e6965",
          7659 => x"642e0a00",
          7660 => x"46696c65",
          7661 => x"20616c72",
          7662 => x"65616479",
          7663 => x"20657869",
          7664 => x"7374732e",
          7665 => x"0a000000",
          7666 => x"46696c65",
          7667 => x"2068616e",
          7668 => x"646c6520",
          7669 => x"696e7661",
          7670 => x"6c69642e",
          7671 => x"0a000000",
          7672 => x"53442069",
          7673 => x"73207772",
          7674 => x"69746520",
          7675 => x"70726f74",
          7676 => x"65637465",
          7677 => x"642e0a00",
          7678 => x"44726976",
          7679 => x"65206e75",
          7680 => x"6d626572",
          7681 => x"20697320",
          7682 => x"696e7661",
          7683 => x"6c69642e",
          7684 => x"0a000000",
          7685 => x"4469736b",
          7686 => x"206e6f74",
          7687 => x"20656e61",
          7688 => x"626c6564",
          7689 => x"2e0a0000",
          7690 => x"4e6f2063",
          7691 => x"6f6d7061",
          7692 => x"7469626c",
          7693 => x"65206669",
          7694 => x"6c657379",
          7695 => x"7374656d",
          7696 => x"20666f75",
          7697 => x"6e64206f",
          7698 => x"6e206469",
          7699 => x"736b2e0a",
          7700 => x"00000000",
          7701 => x"466f726d",
          7702 => x"61742061",
          7703 => x"626f7274",
          7704 => x"65642e0a",
          7705 => x"00000000",
          7706 => x"54696d65",
          7707 => x"6f75742c",
          7708 => x"206f7065",
          7709 => x"72617469",
          7710 => x"6f6e2063",
          7711 => x"616e6365",
          7712 => x"6c6c6564",
          7713 => x"2e0a0000",
          7714 => x"46696c65",
          7715 => x"20697320",
          7716 => x"6c6f636b",
          7717 => x"65642e0a",
          7718 => x"00000000",
          7719 => x"496e7375",
          7720 => x"66666963",
          7721 => x"69656e74",
          7722 => x"206d656d",
          7723 => x"6f72792e",
          7724 => x"0a000000",
          7725 => x"546f6f20",
          7726 => x"6d616e79",
          7727 => x"206f7065",
          7728 => x"6e206669",
          7729 => x"6c65732e",
          7730 => x"0a000000",
          7731 => x"50617261",
          7732 => x"6d657465",
          7733 => x"72732069",
          7734 => x"6e636f72",
          7735 => x"72656374",
          7736 => x"2e0a0000",
          7737 => x"53756363",
          7738 => x"6573732e",
          7739 => x"0a000000",
          7740 => x"556e6b6e",
          7741 => x"6f776e20",
          7742 => x"6572726f",
          7743 => x"722e0a00",
          7744 => x"0a256c75",
          7745 => x"20627974",
          7746 => x"65732025",
          7747 => x"73206174",
          7748 => x"20256c75",
          7749 => x"20627974",
          7750 => x"65732f73",
          7751 => x"65632e0a",
          7752 => x"00000000",
          7753 => x"72656164",
          7754 => x"00000000",
          7755 => x"25303858",
          7756 => x"00000000",
          7757 => x"3a202000",
          7758 => x"25303458",
          7759 => x"00000000",
          7760 => x"20202020",
          7761 => x"20202020",
          7762 => x"00000000",
          7763 => x"25303258",
          7764 => x"00000000",
          7765 => x"20200000",
          7766 => x"207c0000",
          7767 => x"7c0d0a00",
          7768 => x"5a505554",
          7769 => x"41000000",
          7770 => x"0a2a2a20",
          7771 => x"25732028",
          7772 => x"00000000",
          7773 => x"32312f30",
          7774 => x"342f3230",
          7775 => x"32300000",
          7776 => x"76312e35",
          7777 => x"31000000",
          7778 => x"205a5055",
          7779 => x"2c207265",
          7780 => x"76202530",
          7781 => x"32782920",
          7782 => x"25732025",
          7783 => x"73202a2a",
          7784 => x"0a0a0000",
          7785 => x"5a505554",
          7786 => x"4120496e",
          7787 => x"74657272",
          7788 => x"75707420",
          7789 => x"48616e64",
          7790 => x"6c65720a",
          7791 => x"00000000",
          7792 => x"54696d65",
          7793 => x"7220696e",
          7794 => x"74657272",
          7795 => x"7570740a",
          7796 => x"00000000",
          7797 => x"50533220",
          7798 => x"696e7465",
          7799 => x"72727570",
          7800 => x"740a0000",
          7801 => x"494f4354",
          7802 => x"4c205244",
          7803 => x"20696e74",
          7804 => x"65727275",
          7805 => x"70740a00",
          7806 => x"494f4354",
          7807 => x"4c205752",
          7808 => x"20696e74",
          7809 => x"65727275",
          7810 => x"70740a00",
          7811 => x"55415254",
          7812 => x"30205258",
          7813 => x"20696e74",
          7814 => x"65727275",
          7815 => x"70740a00",
          7816 => x"55415254",
          7817 => x"30205458",
          7818 => x"20696e74",
          7819 => x"65727275",
          7820 => x"70740a00",
          7821 => x"55415254",
          7822 => x"31205258",
          7823 => x"20696e74",
          7824 => x"65727275",
          7825 => x"70740a00",
          7826 => x"55415254",
          7827 => x"31205458",
          7828 => x"20696e74",
          7829 => x"65727275",
          7830 => x"70740a00",
          7831 => x"53657474",
          7832 => x"696e6720",
          7833 => x"75702074",
          7834 => x"696d6572",
          7835 => x"2e2e2e0a",
          7836 => x"00000000",
          7837 => x"456e6162",
          7838 => x"6c696e67",
          7839 => x"2074696d",
          7840 => x"65722e2e",
          7841 => x"2e0a0000",
          7842 => x"6175746f",
          7843 => x"65786563",
          7844 => x"2e626174",
          7845 => x"00000000",
          7846 => x"303a0000",
          7847 => x"4661696c",
          7848 => x"65642074",
          7849 => x"6f20696e",
          7850 => x"69746961",
          7851 => x"6c697365",
          7852 => x"20736420",
          7853 => x"63617264",
          7854 => x"20302c20",
          7855 => x"706c6561",
          7856 => x"73652069",
          7857 => x"6e697420",
          7858 => x"6d616e75",
          7859 => x"616c6c79",
          7860 => x"2e0a0000",
          7861 => x"2a200000",
          7862 => x"42616420",
          7863 => x"6469736b",
          7864 => x"20696421",
          7865 => x"0a000000",
          7866 => x"496e6974",
          7867 => x"69616c69",
          7868 => x"7365642e",
          7869 => x"0a000000",
          7870 => x"4661696c",
          7871 => x"65642074",
          7872 => x"6f20696e",
          7873 => x"69746961",
          7874 => x"6c697365",
          7875 => x"2e0a0000",
          7876 => x"72633d25",
          7877 => x"640a0000",
          7878 => x"25753a00",
          7879 => x"436c6561",
          7880 => x"72696e67",
          7881 => x"2e2e2e2e",
          7882 => x"00000000",
          7883 => x"436f7079",
          7884 => x"696e672e",
          7885 => x"2e2e0000",
          7886 => x"436f6d70",
          7887 => x"6172696e",
          7888 => x"672e2e2e",
          7889 => x"00000000",
          7890 => x"2530386c",
          7891 => x"78282530",
          7892 => x"3878292d",
          7893 => x"3e253038",
          7894 => x"6c782825",
          7895 => x"30387829",
          7896 => x"0a000000",
          7897 => x"44756d70",
          7898 => x"204d656d",
          7899 => x"6f72790a",
          7900 => x"00000000",
          7901 => x"0a436f6d",
          7902 => x"706c6574",
          7903 => x"652e0a00",
          7904 => x"25303858",
          7905 => x"20253032",
          7906 => x"582d0000",
          7907 => x"3f3f3f0a",
          7908 => x"00000000",
          7909 => x"25303858",
          7910 => x"20253034",
          7911 => x"582d0000",
          7912 => x"25303858",
          7913 => x"20253038",
          7914 => x"582d0000",
          7915 => x"44697361",
          7916 => x"626c696e",
          7917 => x"6720696e",
          7918 => x"74657272",
          7919 => x"75707473",
          7920 => x"0a000000",
          7921 => x"456e6162",
          7922 => x"6c696e67",
          7923 => x"20696e74",
          7924 => x"65727275",
          7925 => x"7074730a",
          7926 => x"00000000",
          7927 => x"44697361",
          7928 => x"626c6564",
          7929 => x"20756172",
          7930 => x"74206669",
          7931 => x"666f0a00",
          7932 => x"456e6162",
          7933 => x"6c696e67",
          7934 => x"20756172",
          7935 => x"74206669",
          7936 => x"666f0a00",
          7937 => x"45786563",
          7938 => x"7574696e",
          7939 => x"6720636f",
          7940 => x"64652040",
          7941 => x"20253038",
          7942 => x"78202e2e",
          7943 => x"2e0a0000",
          7944 => x"43616c6c",
          7945 => x"696e6720",
          7946 => x"636f6465",
          7947 => x"20402025",
          7948 => x"30387820",
          7949 => x"2e2e2e0a",
          7950 => x"00000000",
          7951 => x"43616c6c",
          7952 => x"20726574",
          7953 => x"75726e65",
          7954 => x"6420636f",
          7955 => x"64652028",
          7956 => x"2564292e",
          7957 => x"0a000000",
          7958 => x"52657374",
          7959 => x"61727469",
          7960 => x"6e672061",
          7961 => x"70706c69",
          7962 => x"63617469",
          7963 => x"6f6e2e2e",
          7964 => x"2e0a0000",
          7965 => x"436f6c64",
          7966 => x"20726562",
          7967 => x"6f6f7469",
          7968 => x"6e672e2e",
          7969 => x"2e0a0000",
          7970 => x"5a505500",
          7971 => x"62696e00",
          7972 => x"25643a5c",
          7973 => x"25735c25",
          7974 => x"732e2573",
          7975 => x"00000000",
          7976 => x"25643a5c",
          7977 => x"25735c25",
          7978 => x"73000000",
          7979 => x"25643a5c",
          7980 => x"25730000",
          7981 => x"42616420",
          7982 => x"636f6d6d",
          7983 => x"616e642e",
          7984 => x"0a000000",
          7985 => x"52756e6e",
          7986 => x"696e672e",
          7987 => x"2e2e0a00",
          7988 => x"456e6162",
          7989 => x"6c696e67",
          7990 => x"20696e74",
          7991 => x"65727275",
          7992 => x"7074732e",
          7993 => x"2e2e0a00",
          7994 => x"00000000",
          7995 => x"00000000",
          7996 => x"00007fff",
          7997 => x"00000000",
          7998 => x"00007fff",
          7999 => x"00010000",
          8000 => x"00007fff",
          8001 => x"00010000",
          8002 => x"00810000",
          8003 => x"01000000",
          8004 => x"017fffff",
          8005 => x"00000000",
          8006 => x"00000000",
          8007 => x"00007800",
          8008 => x"00000000",
          8009 => x"05f5e100",
          8010 => x"05f5e100",
          8011 => x"05f5e100",
          8012 => x"00000000",
          8013 => x"01010101",
          8014 => x"01010101",
          8015 => x"01011001",
          8016 => x"01000000",
          8017 => x"00000000",
          8018 => x"00000002",
          8019 => x"00000000",
          8020 => x"00007d48",
          8021 => x"00007d48",
          8022 => x"00007d48",
          8023 => x"00007d48",
          8024 => x"00007440",
          8025 => x"00000000",
          8026 => x"00000000",
          8027 => x"00000000",
          8028 => x"00000000",
          8029 => x"00000000",
          8030 => x"00000000",
          8031 => x"00000000",
          8032 => x"00000000",
          8033 => x"00000000",
          8034 => x"00000000",
          8035 => x"00000000",
          8036 => x"00000000",
          8037 => x"00000000",
          8038 => x"00000000",
          8039 => x"00000000",
          8040 => x"00000000",
          8041 => x"00000000",
          8042 => x"00000000",
          8043 => x"00000000",
          8044 => x"00000000",
          8045 => x"00000000",
          8046 => x"00000000",
          8047 => x"00000000",
          8048 => x"0000744c",
          8049 => x"01000000",
          8050 => x"00007454",
          8051 => x"01000000",
          8052 => x"0000745c",
          8053 => x"02000000",
          8054 => x"01000000",
          8055 => x"00000000",
          8056 => x"00007690",
          8057 => x"01020100",
          8058 => x"00000000",
          8059 => x"00000000",
          8060 => x"00007698",
          8061 => x"01040100",
          8062 => x"00000000",
          8063 => x"00000000",
          8064 => x"000076a0",
          8065 => x"01140300",
          8066 => x"00000000",
          8067 => x"00000000",
          8068 => x"000076a8",
          8069 => x"012b0300",
          8070 => x"00000000",
          8071 => x"00000000",
          8072 => x"000076b0",
          8073 => x"01300300",
          8074 => x"00000000",
          8075 => x"00000000",
          8076 => x"000076b8",
          8077 => x"013c0400",
          8078 => x"00000000",
          8079 => x"00000000",
          8080 => x"000076c0",
          8081 => x"013d0400",
          8082 => x"00000000",
          8083 => x"00000000",
          8084 => x"000076c8",
          8085 => x"013f0400",
          8086 => x"00000000",
          8087 => x"00000000",
          8088 => x"000076d0",
          8089 => x"01400400",
          8090 => x"00000000",
          8091 => x"00000000",
          8092 => x"000076d8",
          8093 => x"01410400",
          8094 => x"00000000",
          8095 => x"00000000",
          8096 => x"000076dc",
          8097 => x"01420400",
          8098 => x"00000000",
          8099 => x"00000000",
          8100 => x"000076e0",
          8101 => x"01430400",
          8102 => x"00000000",
          8103 => x"00000000",
          8104 => x"000076e4",
          8105 => x"01500500",
          8106 => x"00000000",
          8107 => x"00000000",
          8108 => x"000076e8",
          8109 => x"01510500",
          8110 => x"00000000",
          8111 => x"00000000",
          8112 => x"000076ec",
          8113 => x"01540500",
          8114 => x"00000000",
          8115 => x"00000000",
          8116 => x"000076f0",
          8117 => x"01550500",
          8118 => x"00000000",
          8119 => x"00000000",
          8120 => x"000076f4",
          8121 => x"01790700",
          8122 => x"00000000",
          8123 => x"00000000",
          8124 => x"000076fc",
          8125 => x"01780700",
          8126 => x"00000000",
          8127 => x"00000000",
          8128 => x"00007700",
          8129 => x"01820800",
          8130 => x"00000000",
          8131 => x"00000000",
          8132 => x"00007708",
          8133 => x"01830800",
          8134 => x"00000000",
          8135 => x"00000000",
          8136 => x"00007710",
          8137 => x"01850800",
          8138 => x"00000000",
          8139 => x"00000000",
          8140 => x"00007718",
          8141 => x"01870800",
          8142 => x"00000000",
          8143 => x"00000000",
          8144 => x"00007720",
          8145 => x"018c0900",
          8146 => x"00000000",
          8147 => x"00000000",
          8148 => x"00007728",
          8149 => x"018d0900",
          8150 => x"00000000",
          8151 => x"00000000",
          8152 => x"00007730",
          8153 => x"018e0900",
          8154 => x"00000000",
          8155 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

