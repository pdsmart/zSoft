-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b0b93",
          2049 => x"8c040000",
          2050 => x"00000000",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b92",
          2121 => x"f0040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b92d3",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b81dc",
          2210 => x"ac738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"92d80400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b0b94",
          2219 => x"912d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b0b95",
          2227 => x"fd2d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"94040b0b",
          2317 => x"0b8ca304",
          2318 => x"0b0b0b8c",
          2319 => x"b2040b0b",
          2320 => x"0b8cc104",
          2321 => x"0b0b0b8c",
          2322 => x"d0040b0b",
          2323 => x"0b8cdf04",
          2324 => x"0b0b0b8c",
          2325 => x"ee040b0b",
          2326 => x"0b8cfd04",
          2327 => x"0b0b0b8d",
          2328 => x"8c040b0b",
          2329 => x"0b8d9b04",
          2330 => x"0b0b0b8d",
          2331 => x"aa040b0b",
          2332 => x"0b8db904",
          2333 => x"0b0b0b8d",
          2334 => x"c8040b0b",
          2335 => x"0b8dd704",
          2336 => x"0b0b0b8d",
          2337 => x"e6040b0b",
          2338 => x"0b8df504",
          2339 => x"0b0b0b8e",
          2340 => x"84040b0b",
          2341 => x"0b8e9304",
          2342 => x"0b0b0b8e",
          2343 => x"a3040b0b",
          2344 => x"0b8eb304",
          2345 => x"0b0b0b8e",
          2346 => x"c3040b0b",
          2347 => x"0b8ed304",
          2348 => x"0b0b0b8e",
          2349 => x"e3040b0b",
          2350 => x"0b8ef304",
          2351 => x"0b0b0b8f",
          2352 => x"83040b0b",
          2353 => x"0b8f9304",
          2354 => x"0b0b0b8f",
          2355 => x"a3040b0b",
          2356 => x"0b8fb304",
          2357 => x"0b0b0b8f",
          2358 => x"c3040b0b",
          2359 => x"0b8fd304",
          2360 => x"0b0b0b8f",
          2361 => x"e3040b0b",
          2362 => x"0b8ff304",
          2363 => x"0b0b0b90",
          2364 => x"83040b0b",
          2365 => x"0b909304",
          2366 => x"0b0b0b90",
          2367 => x"a3040b0b",
          2368 => x"0b90b304",
          2369 => x"0b0b0b90",
          2370 => x"c3040b0b",
          2371 => x"0b90d304",
          2372 => x"0b0b0b90",
          2373 => x"e3040b0b",
          2374 => x"0b90f304",
          2375 => x"0b0b0b91",
          2376 => x"83040b0b",
          2377 => x"0b919304",
          2378 => x"0b0b0b91",
          2379 => x"a3040b0b",
          2380 => x"0b91b304",
          2381 => x"0b0b0b91",
          2382 => x"c3040b0b",
          2383 => x"0b91d304",
          2384 => x"0b0b0b91",
          2385 => x"e3040b0b",
          2386 => x"0b91f304",
          2387 => x"0b0b0b92",
          2388 => x"82040b0b",
          2389 => x"0b929104",
          2390 => x"0b0b0b92",
          2391 => x"a004ffff",
          2392 => x"ffffffff",
          2393 => x"ffffffff",
          2394 => x"ffffffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0481f8d4",
          2434 => x"0ca3ff2d",
          2435 => x"81f8d408",
          2436 => x"83809004",
          2437 => x"81f8d40c",
          2438 => x"b5872d81",
          2439 => x"f8d40883",
          2440 => x"80900481",
          2441 => x"f8d40cb5",
          2442 => x"c62d81f8",
          2443 => x"d4088380",
          2444 => x"900481f8",
          2445 => x"d40cb5e4",
          2446 => x"2d81f8d4",
          2447 => x"08838090",
          2448 => x"0481f8d4",
          2449 => x"0cbca22d",
          2450 => x"81f8d408",
          2451 => x"83809004",
          2452 => x"81f8d40c",
          2453 => x"bda02d81",
          2454 => x"f8d40883",
          2455 => x"80900481",
          2456 => x"f8d40cb6",
          2457 => x"872d81f8",
          2458 => x"d4088380",
          2459 => x"900481f8",
          2460 => x"d40cbdbd",
          2461 => x"2d81f8d4",
          2462 => x"08838090",
          2463 => x"0481f8d4",
          2464 => x"0cbfaf2d",
          2465 => x"81f8d408",
          2466 => x"83809004",
          2467 => x"81f8d40c",
          2468 => x"bbc82d81",
          2469 => x"f8d40883",
          2470 => x"80900481",
          2471 => x"f8d40cb6",
          2472 => x"b92d81f8",
          2473 => x"d4088380",
          2474 => x"900481f8",
          2475 => x"d40cbbde",
          2476 => x"2d81f8d4",
          2477 => x"08838090",
          2478 => x"0481f8d4",
          2479 => x"0cbc822d",
          2480 => x"81f8d408",
          2481 => x"83809004",
          2482 => x"81f8d40c",
          2483 => x"a68c2d81",
          2484 => x"f8d40883",
          2485 => x"80900481",
          2486 => x"f8d40ca6",
          2487 => x"dd2d81f8",
          2488 => x"d4088380",
          2489 => x"900481f8",
          2490 => x"d40c9ef9",
          2491 => x"2d81f8d4",
          2492 => x"08838090",
          2493 => x"0481f8d4",
          2494 => x"0ca0ae2d",
          2495 => x"81f8d408",
          2496 => x"83809004",
          2497 => x"81f8d40c",
          2498 => x"a1e12d81",
          2499 => x"f8d40883",
          2500 => x"80900481",
          2501 => x"f8d40c81",
          2502 => x"84822d81",
          2503 => x"f8d40883",
          2504 => x"80900481",
          2505 => x"f8d40c81",
          2506 => x"90f32d81",
          2507 => x"f8d40883",
          2508 => x"80900481",
          2509 => x"f8d40c81",
          2510 => x"88e72d81",
          2511 => x"f8d40883",
          2512 => x"80900481",
          2513 => x"f8d40c81",
          2514 => x"8be42d81",
          2515 => x"f8d40883",
          2516 => x"80900481",
          2517 => x"f8d40c81",
          2518 => x"96822d81",
          2519 => x"f8d40883",
          2520 => x"80900481",
          2521 => x"f8d40c81",
          2522 => x"9ee22d81",
          2523 => x"f8d40883",
          2524 => x"80900481",
          2525 => x"f8d40c81",
          2526 => x"8fd52d81",
          2527 => x"f8d40883",
          2528 => x"80900481",
          2529 => x"f8d40c81",
          2530 => x"99a12d81",
          2531 => x"f8d40883",
          2532 => x"80900481",
          2533 => x"f8d40c81",
          2534 => x"9ac02d81",
          2535 => x"f8d40883",
          2536 => x"80900481",
          2537 => x"f8d40c81",
          2538 => x"9adf2d81",
          2539 => x"f8d40883",
          2540 => x"80900481",
          2541 => x"f8d40c81",
          2542 => x"a2c92d81",
          2543 => x"f8d40883",
          2544 => x"80900481",
          2545 => x"f8d40c81",
          2546 => x"a0af2d81",
          2547 => x"f8d40883",
          2548 => x"80900481",
          2549 => x"f8d40c81",
          2550 => x"a59d2d81",
          2551 => x"f8d40883",
          2552 => x"80900481",
          2553 => x"f8d40c81",
          2554 => x"9be32d81",
          2555 => x"f8d40883",
          2556 => x"80900481",
          2557 => x"f8d40c81",
          2558 => x"a89d2d81",
          2559 => x"f8d40883",
          2560 => x"80900481",
          2561 => x"f8d40c81",
          2562 => x"a99e2d81",
          2563 => x"f8d40883",
          2564 => x"80900481",
          2565 => x"f8d40c81",
          2566 => x"91d32d81",
          2567 => x"f8d40883",
          2568 => x"80900481",
          2569 => x"f8d40c81",
          2570 => x"91ac2d81",
          2571 => x"f8d40883",
          2572 => x"80900481",
          2573 => x"f8d40c81",
          2574 => x"92d72d81",
          2575 => x"f8d40883",
          2576 => x"80900481",
          2577 => x"f8d40c81",
          2578 => x"9cba2d81",
          2579 => x"f8d40883",
          2580 => x"80900481",
          2581 => x"f8d40c81",
          2582 => x"aa8f2d81",
          2583 => x"f8d40883",
          2584 => x"80900481",
          2585 => x"f8d40c81",
          2586 => x"ac992d81",
          2587 => x"f8d40883",
          2588 => x"80900481",
          2589 => x"f8d40c81",
          2590 => x"afdb2d81",
          2591 => x"f8d40883",
          2592 => x"80900481",
          2593 => x"f8d40c81",
          2594 => x"83a12d81",
          2595 => x"f8d40883",
          2596 => x"80900481",
          2597 => x"f8d40c81",
          2598 => x"b2c72d81",
          2599 => x"f8d40883",
          2600 => x"80900481",
          2601 => x"f8d40c81",
          2602 => x"c0fc2d81",
          2603 => x"f8d40883",
          2604 => x"80900481",
          2605 => x"f8d40c81",
          2606 => x"bee82d81",
          2607 => x"f8d40883",
          2608 => x"80900481",
          2609 => x"f8d40c80",
          2610 => x"d4dc2d81",
          2611 => x"f8d40883",
          2612 => x"80900481",
          2613 => x"f8d40c80",
          2614 => x"d6c62d81",
          2615 => x"f8d40883",
          2616 => x"80900481",
          2617 => x"f8d40c80",
          2618 => x"d8aa2d81",
          2619 => x"f8d40883",
          2620 => x"80900481",
          2621 => x"f8d40c9f",
          2622 => x"a22d81f8",
          2623 => x"d4088380",
          2624 => x"900481f8",
          2625 => x"d40ca084",
          2626 => x"2d81f8d4",
          2627 => x"08838090",
          2628 => x"0481f8d4",
          2629 => x"0ca2f12d",
          2630 => x"81f8d408",
          2631 => x"83809004",
          2632 => x"81f8d40c",
          2633 => x"81c2972d",
          2634 => x"81f8d408",
          2635 => x"83809004",
          2636 => x"3c040000",
          2637 => x"10101010",
          2638 => x"10101010",
          2639 => x"10101010",
          2640 => x"10101010",
          2641 => x"10101010",
          2642 => x"10101010",
          2643 => x"10101010",
          2644 => x"10101053",
          2645 => x"51040000",
          2646 => x"7381ff06",
          2647 => x"73830609",
          2648 => x"81058305",
          2649 => x"1010102b",
          2650 => x"0772fc06",
          2651 => x"0c515104",
          2652 => x"72728072",
          2653 => x"8106ff05",
          2654 => x"09720605",
          2655 => x"71105272",
          2656 => x"0a100a53",
          2657 => x"72ed3851",
          2658 => x"51535104",
          2659 => x"81f8c870",
          2660 => x"82908827",
          2661 => x"8e388071",
          2662 => x"70840553",
          2663 => x"0c0b0b0b",
          2664 => x"938f048c",
          2665 => x"815181da",
          2666 => x"fd040081",
          2667 => x"f8d40802",
          2668 => x"81f8d40c",
          2669 => x"fd3d0d80",
          2670 => x"5381f8d4",
          2671 => x"088c0508",
          2672 => x"5281f8d4",
          2673 => x"08880508",
          2674 => x"5183d43f",
          2675 => x"81f8c808",
          2676 => x"7081f8c8",
          2677 => x"0c54853d",
          2678 => x"0d81f8d4",
          2679 => x"0c0481f8",
          2680 => x"d4080281",
          2681 => x"f8d40cfd",
          2682 => x"3d0d8153",
          2683 => x"81f8d408",
          2684 => x"8c050852",
          2685 => x"81f8d408",
          2686 => x"88050851",
          2687 => x"83a13f81",
          2688 => x"f8c80870",
          2689 => x"81f8c80c",
          2690 => x"54853d0d",
          2691 => x"81f8d40c",
          2692 => x"0481f8d4",
          2693 => x"080281f8",
          2694 => x"d40cf93d",
          2695 => x"0d800b81",
          2696 => x"f8d408fc",
          2697 => x"050c81f8",
          2698 => x"d4088805",
          2699 => x"088025b9",
          2700 => x"3881f8d4",
          2701 => x"08880508",
          2702 => x"3081f8d4",
          2703 => x"0888050c",
          2704 => x"800b81f8",
          2705 => x"d408f405",
          2706 => x"0c81f8d4",
          2707 => x"08fc0508",
          2708 => x"8a38810b",
          2709 => x"81f8d408",
          2710 => x"f4050c81",
          2711 => x"f8d408f4",
          2712 => x"050881f8",
          2713 => x"d408fc05",
          2714 => x"0c81f8d4",
          2715 => x"088c0508",
          2716 => x"8025b938",
          2717 => x"81f8d408",
          2718 => x"8c050830",
          2719 => x"81f8d408",
          2720 => x"8c050c80",
          2721 => x"0b81f8d4",
          2722 => x"08f0050c",
          2723 => x"81f8d408",
          2724 => x"fc05088a",
          2725 => x"38810b81",
          2726 => x"f8d408f0",
          2727 => x"050c81f8",
          2728 => x"d408f005",
          2729 => x"0881f8d4",
          2730 => x"08fc050c",
          2731 => x"805381f8",
          2732 => x"d4088c05",
          2733 => x"085281f8",
          2734 => x"d4088805",
          2735 => x"085181df",
          2736 => x"3f81f8c8",
          2737 => x"087081f8",
          2738 => x"d408f805",
          2739 => x"0c5481f8",
          2740 => x"d408fc05",
          2741 => x"08802e90",
          2742 => x"3881f8d4",
          2743 => x"08f80508",
          2744 => x"3081f8d4",
          2745 => x"08f8050c",
          2746 => x"81f8d408",
          2747 => x"f8050870",
          2748 => x"81f8c80c",
          2749 => x"54893d0d",
          2750 => x"81f8d40c",
          2751 => x"0481f8d4",
          2752 => x"080281f8",
          2753 => x"d40cfb3d",
          2754 => x"0d800b81",
          2755 => x"f8d408fc",
          2756 => x"050c81f8",
          2757 => x"d4088805",
          2758 => x"08802599",
          2759 => x"3881f8d4",
          2760 => x"08880508",
          2761 => x"3081f8d4",
          2762 => x"0888050c",
          2763 => x"810b81f8",
          2764 => x"d408fc05",
          2765 => x"0c81f8d4",
          2766 => x"088c0508",
          2767 => x"80259038",
          2768 => x"81f8d408",
          2769 => x"8c050830",
          2770 => x"81f8d408",
          2771 => x"8c050c81",
          2772 => x"5381f8d4",
          2773 => x"088c0508",
          2774 => x"5281f8d4",
          2775 => x"08880508",
          2776 => x"51bd3f81",
          2777 => x"f8c80870",
          2778 => x"81f8d408",
          2779 => x"f8050c54",
          2780 => x"81f8d408",
          2781 => x"fc050880",
          2782 => x"2e903881",
          2783 => x"f8d408f8",
          2784 => x"05083081",
          2785 => x"f8d408f8",
          2786 => x"050c81f8",
          2787 => x"d408f805",
          2788 => x"087081f8",
          2789 => x"c80c5487",
          2790 => x"3d0d81f8",
          2791 => x"d40c0481",
          2792 => x"f8d40802",
          2793 => x"81f8d40c",
          2794 => x"fd3d0d81",
          2795 => x"0b81f8d4",
          2796 => x"08fc050c",
          2797 => x"800b81f8",
          2798 => x"d408f805",
          2799 => x"0c81f8d4",
          2800 => x"088c0508",
          2801 => x"81f8d408",
          2802 => x"88050827",
          2803 => x"b93881f8",
          2804 => x"d408fc05",
          2805 => x"08802eae",
          2806 => x"38800b81",
          2807 => x"f8d4088c",
          2808 => x"050824a2",
          2809 => x"3881f8d4",
          2810 => x"088c0508",
          2811 => x"1081f8d4",
          2812 => x"088c050c",
          2813 => x"81f8d408",
          2814 => x"fc050810",
          2815 => x"81f8d408",
          2816 => x"fc050cff",
          2817 => x"b83981f8",
          2818 => x"d408fc05",
          2819 => x"08802e80",
          2820 => x"e13881f8",
          2821 => x"d4088c05",
          2822 => x"0881f8d4",
          2823 => x"08880508",
          2824 => x"26ad3881",
          2825 => x"f8d40888",
          2826 => x"050881f8",
          2827 => x"d4088c05",
          2828 => x"083181f8",
          2829 => x"d4088805",
          2830 => x"0c81f8d4",
          2831 => x"08f80508",
          2832 => x"81f8d408",
          2833 => x"fc050807",
          2834 => x"81f8d408",
          2835 => x"f8050c81",
          2836 => x"f8d408fc",
          2837 => x"0508812a",
          2838 => x"81f8d408",
          2839 => x"fc050c81",
          2840 => x"f8d4088c",
          2841 => x"0508812a",
          2842 => x"81f8d408",
          2843 => x"8c050cff",
          2844 => x"953981f8",
          2845 => x"d4089005",
          2846 => x"08802e93",
          2847 => x"3881f8d4",
          2848 => x"08880508",
          2849 => x"7081f8d4",
          2850 => x"08f4050c",
          2851 => x"51913981",
          2852 => x"f8d408f8",
          2853 => x"05087081",
          2854 => x"f8d408f4",
          2855 => x"050c5181",
          2856 => x"f8d408f4",
          2857 => x"050881f8",
          2858 => x"c80c853d",
          2859 => x"0d81f8d4",
          2860 => x"0c04fc3d",
          2861 => x"0d767079",
          2862 => x"7b555555",
          2863 => x"558f7227",
          2864 => x"8c387275",
          2865 => x"07830651",
          2866 => x"70802ea9",
          2867 => x"38ff1252",
          2868 => x"71ff2e98",
          2869 => x"38727081",
          2870 => x"05543374",
          2871 => x"70810556",
          2872 => x"34ff1252",
          2873 => x"71ff2e09",
          2874 => x"8106ea38",
          2875 => x"7481f8c8",
          2876 => x"0c863d0d",
          2877 => x"04745172",
          2878 => x"70840554",
          2879 => x"08717084",
          2880 => x"05530c72",
          2881 => x"70840554",
          2882 => x"08717084",
          2883 => x"05530c72",
          2884 => x"70840554",
          2885 => x"08717084",
          2886 => x"05530c72",
          2887 => x"70840554",
          2888 => x"08717084",
          2889 => x"05530cf0",
          2890 => x"1252718f",
          2891 => x"26c93883",
          2892 => x"72279538",
          2893 => x"72708405",
          2894 => x"54087170",
          2895 => x"8405530c",
          2896 => x"fc125271",
          2897 => x"8326ed38",
          2898 => x"7054ff81",
          2899 => x"39fc3d0d",
          2900 => x"76797102",
          2901 => x"8c059f05",
          2902 => x"33575553",
          2903 => x"55837227",
          2904 => x"8a387483",
          2905 => x"06517080",
          2906 => x"2ea438ff",
          2907 => x"125271ff",
          2908 => x"2e933873",
          2909 => x"73708105",
          2910 => x"5534ff12",
          2911 => x"5271ff2e",
          2912 => x"098106ef",
          2913 => x"387481f8",
          2914 => x"c80c863d",
          2915 => x"0d047474",
          2916 => x"882b7507",
          2917 => x"7071902b",
          2918 => x"07515451",
          2919 => x"8f7227a5",
          2920 => x"38727170",
          2921 => x"8405530c",
          2922 => x"72717084",
          2923 => x"05530c72",
          2924 => x"71708405",
          2925 => x"530c7271",
          2926 => x"70840553",
          2927 => x"0cf01252",
          2928 => x"718f26dd",
          2929 => x"38837227",
          2930 => x"90387271",
          2931 => x"70840553",
          2932 => x"0cfc1252",
          2933 => x"718326f2",
          2934 => x"387053ff",
          2935 => x"8e39fc3d",
          2936 => x"0d767079",
          2937 => x"70730783",
          2938 => x"06545454",
          2939 => x"557080c3",
          2940 => x"38717008",
          2941 => x"700970f7",
          2942 => x"fbfdff13",
          2943 => x"0670f884",
          2944 => x"82818006",
          2945 => x"51515353",
          2946 => x"5470a638",
          2947 => x"84147274",
          2948 => x"70840556",
          2949 => x"0c700870",
          2950 => x"0970f7fb",
          2951 => x"fdff1306",
          2952 => x"70f88482",
          2953 => x"81800651",
          2954 => x"51535354",
          2955 => x"70802edc",
          2956 => x"38735271",
          2957 => x"70810553",
          2958 => x"33517073",
          2959 => x"70810555",
          2960 => x"3470f038",
          2961 => x"7481f8c8",
          2962 => x"0c863d0d",
          2963 => x"04fd3d0d",
          2964 => x"75707183",
          2965 => x"06535552",
          2966 => x"70b83871",
          2967 => x"70087009",
          2968 => x"f7fbfdff",
          2969 => x"120670f8",
          2970 => x"84828180",
          2971 => x"06515152",
          2972 => x"53709d38",
          2973 => x"84137008",
          2974 => x"7009f7fb",
          2975 => x"fdff1206",
          2976 => x"70f88482",
          2977 => x"81800651",
          2978 => x"51525370",
          2979 => x"802ee538",
          2980 => x"72527133",
          2981 => x"5170802e",
          2982 => x"8a388112",
          2983 => x"70335252",
          2984 => x"70f83871",
          2985 => x"743181f8",
          2986 => x"c80c853d",
          2987 => x"0d04fa3d",
          2988 => x"0d787a7c",
          2989 => x"70545555",
          2990 => x"5272802e",
          2991 => x"80d93871",
          2992 => x"74078306",
          2993 => x"5170802e",
          2994 => x"80d638ff",
          2995 => x"135372ff",
          2996 => x"2eb13871",
          2997 => x"33743356",
          2998 => x"5174712e",
          2999 => x"098106a9",
          3000 => x"3872802e",
          3001 => x"81893870",
          3002 => x"81ff0651",
          3003 => x"70802e80",
          3004 => x"fe388112",
          3005 => x"8115ff15",
          3006 => x"55555272",
          3007 => x"ff2e0981",
          3008 => x"06d13871",
          3009 => x"33743356",
          3010 => x"517081ff",
          3011 => x"067581ff",
          3012 => x"06717131",
          3013 => x"51525270",
          3014 => x"81f8c80c",
          3015 => x"883d0d04",
          3016 => x"71745755",
          3017 => x"83732788",
          3018 => x"38710874",
          3019 => x"082e8838",
          3020 => x"74765552",
          3021 => x"ff9539fc",
          3022 => x"13537280",
          3023 => x"2eb13874",
          3024 => x"087009f7",
          3025 => x"fbfdff12",
          3026 => x"0670f884",
          3027 => x"82818006",
          3028 => x"51515170",
          3029 => x"9a388415",
          3030 => x"84175755",
          3031 => x"837327d0",
          3032 => x"38740876",
          3033 => x"082ed038",
          3034 => x"74765552",
          3035 => x"fedd3980",
          3036 => x"0b81f8c8",
          3037 => x"0c883d0d",
          3038 => x"04fe3d0d",
          3039 => x"80528353",
          3040 => x"71882b52",
          3041 => x"87863f81",
          3042 => x"f8c80881",
          3043 => x"ff067207",
          3044 => x"ff145452",
          3045 => x"728025e8",
          3046 => x"387181f8",
          3047 => x"c80c843d",
          3048 => x"0d04fb3d",
          3049 => x"0d777008",
          3050 => x"70535356",
          3051 => x"71802e80",
          3052 => x"ca387133",
          3053 => x"5170a02e",
          3054 => x"09810686",
          3055 => x"38811252",
          3056 => x"f1397153",
          3057 => x"84398113",
          3058 => x"53807333",
          3059 => x"7081ff06",
          3060 => x"53555570",
          3061 => x"a02e8338",
          3062 => x"81557080",
          3063 => x"2e843874",
          3064 => x"e5387381",
          3065 => x"ff065170",
          3066 => x"a02e0981",
          3067 => x"06883880",
          3068 => x"73708105",
          3069 => x"55347276",
          3070 => x"0c715170",
          3071 => x"81f8c80c",
          3072 => x"873d0d04",
          3073 => x"fc3d0d76",
          3074 => x"53720880",
          3075 => x"2e913886",
          3076 => x"3dfc0552",
          3077 => x"72519f97",
          3078 => x"3f81f8c8",
          3079 => x"08853880",
          3080 => x"53833974",
          3081 => x"537281f8",
          3082 => x"c80c863d",
          3083 => x"0d04fc3d",
          3084 => x"0d768211",
          3085 => x"33ff0552",
          3086 => x"53815270",
          3087 => x"8b268198",
          3088 => x"38831333",
          3089 => x"ff055182",
          3090 => x"52709e26",
          3091 => x"818a3884",
          3092 => x"13335183",
          3093 => x"52709726",
          3094 => x"80fe3885",
          3095 => x"13335184",
          3096 => x"5270bb26",
          3097 => x"80f23886",
          3098 => x"13335185",
          3099 => x"5270bb26",
          3100 => x"80e63888",
          3101 => x"13225586",
          3102 => x"527487e7",
          3103 => x"2680d938",
          3104 => x"8a132254",
          3105 => x"87527387",
          3106 => x"e72680cc",
          3107 => x"38810b87",
          3108 => x"c0989c0c",
          3109 => x"722287c0",
          3110 => x"98bc0c82",
          3111 => x"133387c0",
          3112 => x"98b80c83",
          3113 => x"133387c0",
          3114 => x"98b40c84",
          3115 => x"133387c0",
          3116 => x"98b00c85",
          3117 => x"133387c0",
          3118 => x"98ac0c86",
          3119 => x"133387c0",
          3120 => x"98a80c74",
          3121 => x"87c098a4",
          3122 => x"0c7387c0",
          3123 => x"98a00c80",
          3124 => x"0b87c098",
          3125 => x"9c0c8052",
          3126 => x"7181f8c8",
          3127 => x"0c863d0d",
          3128 => x"04f33d0d",
          3129 => x"7f5b87c0",
          3130 => x"989c5d81",
          3131 => x"7d0c87c0",
          3132 => x"98bc085e",
          3133 => x"7d7b2387",
          3134 => x"c098b808",
          3135 => x"5a79821c",
          3136 => x"3487c098",
          3137 => x"b4085a79",
          3138 => x"831c3487",
          3139 => x"c098b008",
          3140 => x"5a79841c",
          3141 => x"3487c098",
          3142 => x"ac085a79",
          3143 => x"851c3487",
          3144 => x"c098a808",
          3145 => x"5a79861c",
          3146 => x"3487c098",
          3147 => x"a4085c7b",
          3148 => x"881c2387",
          3149 => x"c098a008",
          3150 => x"5a798a1c",
          3151 => x"23807d0c",
          3152 => x"7983ffff",
          3153 => x"06597b83",
          3154 => x"ffff0658",
          3155 => x"861b3357",
          3156 => x"851b3356",
          3157 => x"841b3355",
          3158 => x"831b3354",
          3159 => x"821b3353",
          3160 => x"7d83ffff",
          3161 => x"065281dd",
          3162 => x"d05198dc",
          3163 => x"3f8f3d0d",
          3164 => x"04ff3d0d",
          3165 => x"028f0533",
          3166 => x"7030709f",
          3167 => x"2a515252",
          3168 => x"700b0b81",
          3169 => x"f3c03483",
          3170 => x"3d0d04fb",
          3171 => x"3d0d770b",
          3172 => x"0b81f3c0",
          3173 => x"337081ff",
          3174 => x"06575556",
          3175 => x"87c09484",
          3176 => x"5174802e",
          3177 => x"863887c0",
          3178 => x"94945170",
          3179 => x"0870962a",
          3180 => x"70810653",
          3181 => x"54527080",
          3182 => x"2e8c3871",
          3183 => x"912a7081",
          3184 => x"06515170",
          3185 => x"d7387281",
          3186 => x"32708106",
          3187 => x"51517080",
          3188 => x"2e8d3871",
          3189 => x"932a7081",
          3190 => x"06515170",
          3191 => x"ffbe3873",
          3192 => x"81ff0651",
          3193 => x"87c09480",
          3194 => x"5270802e",
          3195 => x"863887c0",
          3196 => x"94905275",
          3197 => x"720c7581",
          3198 => x"f8c80c87",
          3199 => x"3d0d04fb",
          3200 => x"3d0d029f",
          3201 => x"05330b0b",
          3202 => x"81f3c033",
          3203 => x"7081ff06",
          3204 => x"57555687",
          3205 => x"c0948451",
          3206 => x"74802e86",
          3207 => x"3887c094",
          3208 => x"94517008",
          3209 => x"70962a70",
          3210 => x"81065354",
          3211 => x"5270802e",
          3212 => x"8c387191",
          3213 => x"2a708106",
          3214 => x"515170d7",
          3215 => x"38728132",
          3216 => x"70810651",
          3217 => x"5170802e",
          3218 => x"8d387193",
          3219 => x"2a708106",
          3220 => x"515170ff",
          3221 => x"be387381",
          3222 => x"ff065187",
          3223 => x"c0948052",
          3224 => x"70802e86",
          3225 => x"3887c094",
          3226 => x"90527572",
          3227 => x"0c873d0d",
          3228 => x"04f93d0d",
          3229 => x"79548074",
          3230 => x"337081ff",
          3231 => x"06535357",
          3232 => x"70772e80",
          3233 => x"fe387181",
          3234 => x"ff068115",
          3235 => x"0b0b81f3",
          3236 => x"c0337081",
          3237 => x"ff065957",
          3238 => x"555887c0",
          3239 => x"94845175",
          3240 => x"802e8638",
          3241 => x"87c09494",
          3242 => x"51700870",
          3243 => x"962a7081",
          3244 => x"06535452",
          3245 => x"70802e8c",
          3246 => x"3871912a",
          3247 => x"70810651",
          3248 => x"5170d738",
          3249 => x"72813270",
          3250 => x"81065151",
          3251 => x"70802e8d",
          3252 => x"3871932a",
          3253 => x"70810651",
          3254 => x"5170ffbe",
          3255 => x"387481ff",
          3256 => x"065187c0",
          3257 => x"94805270",
          3258 => x"802e8638",
          3259 => x"87c09490",
          3260 => x"5277720c",
          3261 => x"81177433",
          3262 => x"7081ff06",
          3263 => x"53535770",
          3264 => x"ff843876",
          3265 => x"81f8c80c",
          3266 => x"893d0d04",
          3267 => x"fe3d0d0b",
          3268 => x"0b81f3c0",
          3269 => x"337081ff",
          3270 => x"06545287",
          3271 => x"c0948451",
          3272 => x"72802e86",
          3273 => x"3887c094",
          3274 => x"94517008",
          3275 => x"70822a70",
          3276 => x"81065151",
          3277 => x"5170802e",
          3278 => x"e2387181",
          3279 => x"ff065187",
          3280 => x"c0948052",
          3281 => x"70802e86",
          3282 => x"3887c094",
          3283 => x"90527108",
          3284 => x"7081ff06",
          3285 => x"81f8c80c",
          3286 => x"51843d0d",
          3287 => x"04fe3d0d",
          3288 => x"0b0b81f3",
          3289 => x"c0337081",
          3290 => x"ff065253",
          3291 => x"87c09484",
          3292 => x"5270802e",
          3293 => x"863887c0",
          3294 => x"94945271",
          3295 => x"0870822a",
          3296 => x"70810651",
          3297 => x"5151ff52",
          3298 => x"70802ea0",
          3299 => x"387281ff",
          3300 => x"065187c0",
          3301 => x"94805270",
          3302 => x"802e8638",
          3303 => x"87c09490",
          3304 => x"52710870",
          3305 => x"982b7098",
          3306 => x"2c515351",
          3307 => x"7181f8c8",
          3308 => x"0c843d0d",
          3309 => x"04ff3d0d",
          3310 => x"87c09e80",
          3311 => x"08709c2a",
          3312 => x"8a065151",
          3313 => x"70802e84",
          3314 => x"b43887c0",
          3315 => x"9ea40881",
          3316 => x"f3c40c87",
          3317 => x"c09ea808",
          3318 => x"81f3c80c",
          3319 => x"87c09e94",
          3320 => x"0881f3cc",
          3321 => x"0c87c09e",
          3322 => x"980881f3",
          3323 => x"d00c87c0",
          3324 => x"9e9c0881",
          3325 => x"f3d40c87",
          3326 => x"c09ea008",
          3327 => x"81f3d80c",
          3328 => x"87c09eac",
          3329 => x"0881f3dc",
          3330 => x"0c87c09e",
          3331 => x"b00881f3",
          3332 => x"e00c87c0",
          3333 => x"9eb40881",
          3334 => x"f3e40c87",
          3335 => x"c09eb808",
          3336 => x"81f3e80c",
          3337 => x"87c09ebc",
          3338 => x"0881f3ec",
          3339 => x"0c87c09e",
          3340 => x"c00881f3",
          3341 => x"f00c87c0",
          3342 => x"9ec40881",
          3343 => x"f3f40c87",
          3344 => x"c09e8008",
          3345 => x"517081f3",
          3346 => x"f82387c0",
          3347 => x"9e840881",
          3348 => x"f3fc0c87",
          3349 => x"c09e8808",
          3350 => x"81f4800c",
          3351 => x"87c09e8c",
          3352 => x"0881f484",
          3353 => x"0c810b81",
          3354 => x"f4883480",
          3355 => x"0b87c09e",
          3356 => x"90087084",
          3357 => x"800a0651",
          3358 => x"52527080",
          3359 => x"2e833881",
          3360 => x"527181f4",
          3361 => x"8934800b",
          3362 => x"87c09e90",
          3363 => x"08708880",
          3364 => x"0a065152",
          3365 => x"5270802e",
          3366 => x"83388152",
          3367 => x"7181f48a",
          3368 => x"34800b87",
          3369 => x"c09e9008",
          3370 => x"7090800a",
          3371 => x"06515252",
          3372 => x"70802e83",
          3373 => x"38815271",
          3374 => x"81f48b34",
          3375 => x"800b87c0",
          3376 => x"9e900870",
          3377 => x"88808006",
          3378 => x"51525270",
          3379 => x"802e8338",
          3380 => x"81527181",
          3381 => x"f48c3480",
          3382 => x"0b87c09e",
          3383 => x"900870a0",
          3384 => x"80800651",
          3385 => x"52527080",
          3386 => x"2e833881",
          3387 => x"527181f4",
          3388 => x"8d34800b",
          3389 => x"87c09e90",
          3390 => x"08709080",
          3391 => x"80065152",
          3392 => x"5270802e",
          3393 => x"83388152",
          3394 => x"7181f48e",
          3395 => x"34800b87",
          3396 => x"c09e9008",
          3397 => x"70848080",
          3398 => x"06515252",
          3399 => x"70802e83",
          3400 => x"38815271",
          3401 => x"81f48f34",
          3402 => x"800b87c0",
          3403 => x"9e900870",
          3404 => x"82808006",
          3405 => x"51525270",
          3406 => x"802e8338",
          3407 => x"81527181",
          3408 => x"f4903480",
          3409 => x"0b87c09e",
          3410 => x"90087081",
          3411 => x"80800651",
          3412 => x"52527080",
          3413 => x"2e833881",
          3414 => x"527181f4",
          3415 => x"9134800b",
          3416 => x"87c09e90",
          3417 => x"087080c0",
          3418 => x"80065152",
          3419 => x"5270802e",
          3420 => x"83388152",
          3421 => x"7181f492",
          3422 => x"34800b87",
          3423 => x"c09e9008",
          3424 => x"70a08006",
          3425 => x"51525270",
          3426 => x"802e8338",
          3427 => x"81527181",
          3428 => x"f4933487",
          3429 => x"c09e9008",
          3430 => x"70988006",
          3431 => x"708a2a51",
          3432 => x"51517081",
          3433 => x"f4943480",
          3434 => x"0b87c09e",
          3435 => x"90087084",
          3436 => x"80065152",
          3437 => x"5270802e",
          3438 => x"83388152",
          3439 => x"7181f495",
          3440 => x"3487c09e",
          3441 => x"90087083",
          3442 => x"f0067084",
          3443 => x"2a515151",
          3444 => x"7081f496",
          3445 => x"34800b87",
          3446 => x"c09e9008",
          3447 => x"70880651",
          3448 => x"52527080",
          3449 => x"2e833881",
          3450 => x"527181f4",
          3451 => x"973487c0",
          3452 => x"9e900870",
          3453 => x"87065151",
          3454 => x"7081f498",
          3455 => x"34833d0d",
          3456 => x"04fb3d0d",
          3457 => x"81dde851",
          3458 => x"89da3f81",
          3459 => x"f4883354",
          3460 => x"73802e88",
          3461 => x"3881ddfc",
          3462 => x"5189c93f",
          3463 => x"81de9051",
          3464 => x"89c23f81",
          3465 => x"f48a3354",
          3466 => x"73802e93",
          3467 => x"3881f3e4",
          3468 => x"0881f3e8",
          3469 => x"08115452",
          3470 => x"81dea851",
          3471 => x"8f8a3f81",
          3472 => x"f48f3354",
          3473 => x"73802e93",
          3474 => x"3881f3dc",
          3475 => x"0881f3e0",
          3476 => x"08115452",
          3477 => x"81dec451",
          3478 => x"8eee3f81",
          3479 => x"f48c3354",
          3480 => x"73802e93",
          3481 => x"3881f3c4",
          3482 => x"0881f3c8",
          3483 => x"08115452",
          3484 => x"81dee051",
          3485 => x"8ed23f81",
          3486 => x"f48d3354",
          3487 => x"73802e93",
          3488 => x"3881f3cc",
          3489 => x"0881f3d0",
          3490 => x"08115452",
          3491 => x"81defc51",
          3492 => x"8eb63f81",
          3493 => x"f48e3354",
          3494 => x"73802e93",
          3495 => x"3881f3d4",
          3496 => x"0881f3d8",
          3497 => x"08115452",
          3498 => x"81df9851",
          3499 => x"8e9a3f81",
          3500 => x"f4933354",
          3501 => x"73802e8d",
          3502 => x"3881f494",
          3503 => x"335281df",
          3504 => x"b4518e84",
          3505 => x"3f81f497",
          3506 => x"33547380",
          3507 => x"2e8d3881",
          3508 => x"f4983352",
          3509 => x"81dfd451",
          3510 => x"8dee3f81",
          3511 => x"f4953354",
          3512 => x"73802e8d",
          3513 => x"3881f496",
          3514 => x"335281df",
          3515 => x"f4518dd8",
          3516 => x"3f81f489",
          3517 => x"33547380",
          3518 => x"2e883881",
          3519 => x"e0945187",
          3520 => x"e33f81f4",
          3521 => x"8b335473",
          3522 => x"802e8838",
          3523 => x"81e0a851",
          3524 => x"87d23f81",
          3525 => x"f4903354",
          3526 => x"73802e88",
          3527 => x"3881e0b4",
          3528 => x"5187c13f",
          3529 => x"81f49133",
          3530 => x"5473802e",
          3531 => x"883881e0",
          3532 => x"c05187b0",
          3533 => x"3f81f492",
          3534 => x"33547380",
          3535 => x"2e883881",
          3536 => x"e0cc5187",
          3537 => x"9f3f81e0",
          3538 => x"d8518798",
          3539 => x"3f81f3ec",
          3540 => x"085281e0",
          3541 => x"e4518cf0",
          3542 => x"3f81f3f0",
          3543 => x"085281e1",
          3544 => x"8c518ce4",
          3545 => x"3f81f3f4",
          3546 => x"085281e1",
          3547 => x"b4518cd8",
          3548 => x"3f81e1dc",
          3549 => x"5186ed3f",
          3550 => x"81f3f822",
          3551 => x"5281e1e4",
          3552 => x"518cc53f",
          3553 => x"81f3fc08",
          3554 => x"56bd84c0",
          3555 => x"527551e4",
          3556 => x"9a3f81f8",
          3557 => x"c808bd84",
          3558 => x"c0297671",
          3559 => x"31545481",
          3560 => x"f8c80852",
          3561 => x"81e28c51",
          3562 => x"8c9e3f81",
          3563 => x"f48f3354",
          3564 => x"73802ea8",
          3565 => x"3881f480",
          3566 => x"0856bd84",
          3567 => x"c0527551",
          3568 => x"e3e93f81",
          3569 => x"f8c808bd",
          3570 => x"84c02976",
          3571 => x"71315454",
          3572 => x"81f8c808",
          3573 => x"5281e2b8",
          3574 => x"518bed3f",
          3575 => x"81f48a33",
          3576 => x"5473802e",
          3577 => x"a83881f4",
          3578 => x"840856bd",
          3579 => x"84c05275",
          3580 => x"51e3b83f",
          3581 => x"81f8c808",
          3582 => x"bd84c029",
          3583 => x"76713154",
          3584 => x"5481f8c8",
          3585 => x"085281e2",
          3586 => x"e4518bbc",
          3587 => x"3f81f190",
          3588 => x"5185d13f",
          3589 => x"873d0d04",
          3590 => x"fe3d0d02",
          3591 => x"920533ff",
          3592 => x"05527184",
          3593 => x"26aa3871",
          3594 => x"842981dc",
          3595 => x"bc055271",
          3596 => x"080481e3",
          3597 => x"90519d39",
          3598 => x"81e39851",
          3599 => x"973981e3",
          3600 => x"a0519139",
          3601 => x"81e3a851",
          3602 => x"8b3981e3",
          3603 => x"ac518539",
          3604 => x"81e3b451",
          3605 => x"858e3f84",
          3606 => x"3d0d0471",
          3607 => x"88800c04",
          3608 => x"800b87c0",
          3609 => x"96840c04",
          3610 => x"81f49c08",
          3611 => x"87c09684",
          3612 => x"0c04fe3d",
          3613 => x"0d81f8d8",
          3614 => x"08893882",
          3615 => x"90880b81",
          3616 => x"f8d80c81",
          3617 => x"f8d80875",
          3618 => x"115252ff",
          3619 => x"537083b7",
          3620 => x"f8268838",
          3621 => x"7081f8d8",
          3622 => x"0c715372",
          3623 => x"81f8c80c",
          3624 => x"843d0d04",
          3625 => x"f93d0d79",
          3626 => x"7b841208",
          3627 => x"a0129014",
          3628 => x"08941508",
          3629 => x"90165e5a",
          3630 => x"58545957",
          3631 => x"53707726",
          3632 => x"ba387513",
          3633 => x"88140853",
          3634 => x"5181710c",
          3635 => x"76763184",
          3636 => x"120c8073",
          3637 => x"0c758414",
          3638 => x"0c728c12",
          3639 => x"0c718812",
          3640 => x"0c708c13",
          3641 => x"0c708814",
          3642 => x"0c739012",
          3643 => x"0c749412",
          3644 => x"0c709415",
          3645 => x"0c709016",
          3646 => x"0c8c3980",
          3647 => x"730c7390",
          3648 => x"160c7494",
          3649 => x"150c7781",
          3650 => x"f8c80c89",
          3651 => x"3d0d04fc",
          3652 => x"3d0d768c",
          3653 => x"11088812",
          3654 => x"08565353",
          3655 => x"7108812e",
          3656 => x"098106a3",
          3657 => x"38841208",
          3658 => x"70135255",
          3659 => x"70732e09",
          3660 => x"81069438",
          3661 => x"84130815",
          3662 => x"84130c73",
          3663 => x"88130c71",
          3664 => x"8c150c71",
          3665 => x"539f3981",
          3666 => x"730c81f4",
          3667 => x"b0089014",
          3668 => x"0c81f4a0",
          3669 => x"0b94140c",
          3670 => x"7281f4b0",
          3671 => x"0c901308",
          3672 => x"7394120c",
          3673 => x"51730881",
          3674 => x"2e098106",
          3675 => x"b3388413",
          3676 => x"08701452",
          3677 => x"5270742e",
          3678 => x"098106a4",
          3679 => x"38841408",
          3680 => x"1284140c",
          3681 => x"94140890",
          3682 => x"15087090",
          3683 => x"130c5294",
          3684 => x"120c8c14",
          3685 => x"08881508",
          3686 => x"7088130c",
          3687 => x"528c120c",
          3688 => x"7281f8c8",
          3689 => x"0c863d0d",
          3690 => x"04f93d0d",
          3691 => x"79705557",
          3692 => x"76802e81",
          3693 => x"b5389f17",
          3694 => x"f00681f4",
          3695 => x"b0085757",
          3696 => x"7508822e",
          3697 => x"8f388416",
          3698 => x"08772780",
          3699 => x"c7389016",
          3700 => x"0856ed39",
          3701 => x"83ffff17",
          3702 => x"fc808006",
          3703 => x"705258fd",
          3704 => x"913f81f8",
          3705 => x"c80881f8",
          3706 => x"c8083070",
          3707 => x"81f8c808",
          3708 => x"07802581",
          3709 => x"f8c80809",
          3710 => x"70307072",
          3711 => x"07802573",
          3712 => x"07535858",
          3713 => x"51545680",
          3714 => x"5472742e",
          3715 => x"09810680",
          3716 => x"d9388839",
          3717 => x"76527551",
          3718 => x"80c83981",
          3719 => x"0b81f8c8",
          3720 => x"080c7781",
          3721 => x"f8c80884",
          3722 => x"050c81f4",
          3723 => x"ac085372",
          3724 => x"08822e8c",
          3725 => x"38757326",
          3726 => x"87388c13",
          3727 => x"0853f039",
          3728 => x"88130888",
          3729 => x"170c728c",
          3730 => x"170c7588",
          3731 => x"140c8816",
          3732 => x"08768c12",
          3733 => x"0c537551",
          3734 => x"fdb53f76",
          3735 => x"5281f8c8",
          3736 => x"0851fcc0",
          3737 => x"3f81f8c8",
          3738 => x"08547381",
          3739 => x"f8c80c89",
          3740 => x"3d0d04ff",
          3741 => x"3d0d7352",
          3742 => x"71802e87",
          3743 => x"38f01251",
          3744 => x"fd8d3f83",
          3745 => x"3d0d04fe",
          3746 => x"3d0d0293",
          3747 => x"05335372",
          3748 => x"8a2e0981",
          3749 => x"0685388d",
          3750 => x"51ed3f81",
          3751 => x"f8e40852",
          3752 => x"71802e90",
          3753 => x"38727234",
          3754 => x"81f8e408",
          3755 => x"810581f8",
          3756 => x"e40c8f39",
          3757 => x"81f8dc08",
          3758 => x"5271802e",
          3759 => x"85387251",
          3760 => x"712d843d",
          3761 => x"0d04fe3d",
          3762 => x"0d029705",
          3763 => x"3381f8dc",
          3764 => x"087681f8",
          3765 => x"dc0c5451",
          3766 => x"ffad3f72",
          3767 => x"81f8dc0c",
          3768 => x"843d0d04",
          3769 => x"fd3d0d75",
          3770 => x"54733370",
          3771 => x"81ff0653",
          3772 => x"5371802e",
          3773 => x"8e387281",
          3774 => x"ff065181",
          3775 => x"1454ff87",
          3776 => x"3fe73985",
          3777 => x"3d0d04fc",
          3778 => x"3d0d7781",
          3779 => x"f8dc0878",
          3780 => x"81f8dc0c",
          3781 => x"56547333",
          3782 => x"7081ff06",
          3783 => x"53537180",
          3784 => x"2e8e3872",
          3785 => x"81ff0651",
          3786 => x"811454fe",
          3787 => x"da3fe739",
          3788 => x"7481f8dc",
          3789 => x"0c863d0d",
          3790 => x"04ec3d0d",
          3791 => x"66685959",
          3792 => x"78708105",
          3793 => x"5a335675",
          3794 => x"802e84f8",
          3795 => x"3875a52e",
          3796 => x"09810682",
          3797 => x"de388070",
          3798 => x"7a708105",
          3799 => x"5c33585b",
          3800 => x"5b75b02e",
          3801 => x"09810685",
          3802 => x"38815a8b",
          3803 => x"3975ad2e",
          3804 => x"0981068a",
          3805 => x"38825a78",
          3806 => x"7081055a",
          3807 => x"335675aa",
          3808 => x"2e098106",
          3809 => x"92387784",
          3810 => x"1971087b",
          3811 => x"7081055d",
          3812 => x"33595d59",
          3813 => x"539d39d0",
          3814 => x"16537289",
          3815 => x"2695387a",
          3816 => x"88297b10",
          3817 => x"057605d0",
          3818 => x"05797081",
          3819 => x"055b3357",
          3820 => x"5be53975",
          3821 => x"80ec3270",
          3822 => x"30707207",
          3823 => x"80257880",
          3824 => x"cc327030",
          3825 => x"70720780",
          3826 => x"25730753",
          3827 => x"54585155",
          3828 => x"5373802e",
          3829 => x"8c387984",
          3830 => x"07797081",
          3831 => x"055b3357",
          3832 => x"5a75802e",
          3833 => x"83de3875",
          3834 => x"5480e076",
          3835 => x"278938e0",
          3836 => x"167081ff",
          3837 => x"06555373",
          3838 => x"80cf2e81",
          3839 => x"aa387380",
          3840 => x"cf24a238",
          3841 => x"7380c32e",
          3842 => x"818e3873",
          3843 => x"80c3248b",
          3844 => x"387380c2",
          3845 => x"2e818c38",
          3846 => x"81993973",
          3847 => x"80c42e81",
          3848 => x"8a38818f",
          3849 => x"397380d5",
          3850 => x"2e818038",
          3851 => x"7380d524",
          3852 => x"8a387380",
          3853 => x"d32e8e38",
          3854 => x"80f93973",
          3855 => x"80d82e80",
          3856 => x"ee3880ef",
          3857 => x"39778419",
          3858 => x"71085659",
          3859 => x"53807433",
          3860 => x"54557275",
          3861 => x"2e8d3881",
          3862 => x"15701570",
          3863 => x"33515455",
          3864 => x"72f53879",
          3865 => x"812a5690",
          3866 => x"39748116",
          3867 => x"5653727b",
          3868 => x"278f38a0",
          3869 => x"51fc903f",
          3870 => x"75810653",
          3871 => x"72802ee9",
          3872 => x"387351fc",
          3873 => x"df3f7481",
          3874 => x"16565372",
          3875 => x"7b27fdb0",
          3876 => x"38a051fb",
          3877 => x"f23fef39",
          3878 => x"77841983",
          3879 => x"12335359",
          3880 => x"53933982",
          3881 => x"5c953988",
          3882 => x"5c91398a",
          3883 => x"5c8d3990",
          3884 => x"5c893975",
          3885 => x"51fbd03f",
          3886 => x"fd863979",
          3887 => x"822a7081",
          3888 => x"06515372",
          3889 => x"802e8838",
          3890 => x"77841959",
          3891 => x"53863984",
          3892 => x"18785458",
          3893 => x"72087480",
          3894 => x"c4327030",
          3895 => x"70720780",
          3896 => x"25515555",
          3897 => x"55748025",
          3898 => x"8d387280",
          3899 => x"2e883874",
          3900 => x"307a9007",
          3901 => x"5b55800b",
          3902 => x"8f3d5e57",
          3903 => x"7b527451",
          3904 => x"d9dc3f81",
          3905 => x"f8c80881",
          3906 => x"ff067c53",
          3907 => x"755254d9",
          3908 => x"9a3f81f8",
          3909 => x"c8085589",
          3910 => x"74279238",
          3911 => x"a7145375",
          3912 => x"80f82e84",
          3913 => x"38871453",
          3914 => x"7281ff06",
          3915 => x"54b01453",
          3916 => x"727d7081",
          3917 => x"055f3481",
          3918 => x"17753070",
          3919 => x"77079f2a",
          3920 => x"51545776",
          3921 => x"9f268538",
          3922 => x"72ffb138",
          3923 => x"79842a70",
          3924 => x"81065153",
          3925 => x"72802e8e",
          3926 => x"38963d77",
          3927 => x"05e00553",
          3928 => x"ad733481",
          3929 => x"1757767a",
          3930 => x"81065455",
          3931 => x"b0547283",
          3932 => x"38a05479",
          3933 => x"812a7081",
          3934 => x"06545672",
          3935 => x"9f388117",
          3936 => x"55767b27",
          3937 => x"97387351",
          3938 => x"f9fd3f75",
          3939 => x"81065372",
          3940 => x"8b387481",
          3941 => x"1656537a",
          3942 => x"7326eb38",
          3943 => x"963d7705",
          3944 => x"e00553ff",
          3945 => x"17ff1470",
          3946 => x"33535457",
          3947 => x"f9d93f76",
          3948 => x"f2387481",
          3949 => x"16565372",
          3950 => x"7b27fb84",
          3951 => x"38a051f9",
          3952 => x"c63fef39",
          3953 => x"963d0d04",
          3954 => x"fd3d0d86",
          3955 => x"3d707084",
          3956 => x"05520855",
          3957 => x"527351fa",
          3958 => x"e03f853d",
          3959 => x"0d04fe3d",
          3960 => x"0d7481f8",
          3961 => x"e40c853d",
          3962 => x"88055275",
          3963 => x"51faca3f",
          3964 => x"81f8e408",
          3965 => x"53807334",
          3966 => x"800b81f8",
          3967 => x"e40c843d",
          3968 => x"0d04fd3d",
          3969 => x"0d81f8dc",
          3970 => x"087681f8",
          3971 => x"dc0c873d",
          3972 => x"88055377",
          3973 => x"5253faa1",
          3974 => x"3f7281f8",
          3975 => x"dc0c853d",
          3976 => x"0d04fb3d",
          3977 => x"0d777981",
          3978 => x"f8e00870",
          3979 => x"56545755",
          3980 => x"80547180",
          3981 => x"2e80e038",
          3982 => x"81f8e008",
          3983 => x"52712d81",
          3984 => x"f8c80881",
          3985 => x"ff065372",
          3986 => x"802e80cb",
          3987 => x"38728d2e",
          3988 => x"b9387288",
          3989 => x"32703070",
          3990 => x"80255151",
          3991 => x"5273802e",
          3992 => x"8b387180",
          3993 => x"2e8638ff",
          3994 => x"14549739",
          3995 => x"9f7325c8",
          3996 => x"38ff1652",
          3997 => x"737225c0",
          3998 => x"38741452",
          3999 => x"72723481",
          4000 => x"14547251",
          4001 => x"f8813fff",
          4002 => x"af397315",
          4003 => x"52807234",
          4004 => x"8a51f7f3",
          4005 => x"3f815372",
          4006 => x"81f8c80c",
          4007 => x"873d0d04",
          4008 => x"fe3d0d81",
          4009 => x"f8e00875",
          4010 => x"81f8e00c",
          4011 => x"77537652",
          4012 => x"53feef3f",
          4013 => x"7281f8e0",
          4014 => x"0c843d0d",
          4015 => x"04f83d0d",
          4016 => x"7a7c5a56",
          4017 => x"80707a0c",
          4018 => x"58750870",
          4019 => x"33555373",
          4020 => x"a02e0981",
          4021 => x"06873881",
          4022 => x"13760ced",
          4023 => x"3973ad2e",
          4024 => x"0981068e",
          4025 => x"38817608",
          4026 => x"11770c76",
          4027 => x"08703356",
          4028 => x"545873b0",
          4029 => x"2e098106",
          4030 => x"80c23875",
          4031 => x"08810576",
          4032 => x"0c750870",
          4033 => x"33555373",
          4034 => x"80e22e8b",
          4035 => x"38905773",
          4036 => x"80f82e85",
          4037 => x"388f3982",
          4038 => x"57811376",
          4039 => x"0c750870",
          4040 => x"335553ac",
          4041 => x"398155a0",
          4042 => x"742780fa",
          4043 => x"38d01453",
          4044 => x"80558857",
          4045 => x"89732798",
          4046 => x"3880eb39",
          4047 => x"d0145380",
          4048 => x"55728926",
          4049 => x"80e03886",
          4050 => x"39805580",
          4051 => x"d9398a57",
          4052 => x"8055a074",
          4053 => x"2780c238",
          4054 => x"80e07427",
          4055 => x"8938e014",
          4056 => x"7081ff06",
          4057 => x"5553d014",
          4058 => x"7081ff06",
          4059 => x"55539074",
          4060 => x"278e38f9",
          4061 => x"147081ff",
          4062 => x"06555389",
          4063 => x"7427ca38",
          4064 => x"737727c5",
          4065 => x"38747729",
          4066 => x"14760881",
          4067 => x"05770c76",
          4068 => x"08703356",
          4069 => x"5455ffba",
          4070 => x"3977802e",
          4071 => x"84387430",
          4072 => x"5574790c",
          4073 => x"81557481",
          4074 => x"f8c80c8a",
          4075 => x"3d0d04f8",
          4076 => x"3d0d7a7c",
          4077 => x"5a568070",
          4078 => x"7a0c5875",
          4079 => x"08703355",
          4080 => x"5373a02e",
          4081 => x"09810687",
          4082 => x"38811376",
          4083 => x"0ced3973",
          4084 => x"ad2e0981",
          4085 => x"068e3881",
          4086 => x"76081177",
          4087 => x"0c760870",
          4088 => x"33565458",
          4089 => x"73b02e09",
          4090 => x"810680c2",
          4091 => x"38750881",
          4092 => x"05760c75",
          4093 => x"08703355",
          4094 => x"537380e2",
          4095 => x"2e8b3890",
          4096 => x"577380f8",
          4097 => x"2e85388f",
          4098 => x"39825781",
          4099 => x"13760c75",
          4100 => x"08703355",
          4101 => x"53ac3981",
          4102 => x"55a07427",
          4103 => x"80fa38d0",
          4104 => x"14538055",
          4105 => x"88578973",
          4106 => x"27983880",
          4107 => x"eb39d014",
          4108 => x"53805572",
          4109 => x"892680e0",
          4110 => x"38863980",
          4111 => x"5580d939",
          4112 => x"8a578055",
          4113 => x"a0742780",
          4114 => x"c23880e0",
          4115 => x"74278938",
          4116 => x"e0147081",
          4117 => x"ff065553",
          4118 => x"d0147081",
          4119 => x"ff065553",
          4120 => x"9074278e",
          4121 => x"38f91470",
          4122 => x"81ff0655",
          4123 => x"53897427",
          4124 => x"ca387377",
          4125 => x"27c53874",
          4126 => x"77291476",
          4127 => x"08810577",
          4128 => x"0c760870",
          4129 => x"33565455",
          4130 => x"ffba3977",
          4131 => x"802e8438",
          4132 => x"74305574",
          4133 => x"790c8155",
          4134 => x"7481f8c8",
          4135 => x"0c8a3d0d",
          4136 => x"04fd3d0d",
          4137 => x"76982b70",
          4138 => x"982c7998",
          4139 => x"2b70982c",
          4140 => x"72101370",
          4141 => x"822b5153",
          4142 => x"51545151",
          4143 => x"800b81e4",
          4144 => x"c8123355",
          4145 => x"53717425",
          4146 => x"9c3881e4",
          4147 => x"c4110812",
          4148 => x"02840597",
          4149 => x"05337133",
          4150 => x"52525270",
          4151 => x"722e0981",
          4152 => x"06833881",
          4153 => x"537281f8",
          4154 => x"c80c853d",
          4155 => x"0d04fc3d",
          4156 => x"0d780284",
          4157 => x"059f0533",
          4158 => x"71335455",
          4159 => x"5371802e",
          4160 => x"9f388851",
          4161 => x"f3813fa0",
          4162 => x"51f2fc3f",
          4163 => x"8851f2f7",
          4164 => x"3f7233ff",
          4165 => x"05527173",
          4166 => x"347181ff",
          4167 => x"0652de39",
          4168 => x"7651f3c0",
          4169 => x"3f737334",
          4170 => x"863d0d04",
          4171 => x"f63d0d7c",
          4172 => x"028405b7",
          4173 => x"05330288",
          4174 => x"05bb0533",
          4175 => x"81f59433",
          4176 => x"70842981",
          4177 => x"f4bc0570",
          4178 => x"08515959",
          4179 => x"5a585974",
          4180 => x"802e8638",
          4181 => x"7451f29b",
          4182 => x"3f81f594",
          4183 => x"33708429",
          4184 => x"81f4bc05",
          4185 => x"81197054",
          4186 => x"58565af0",
          4187 => x"bc3f81f8",
          4188 => x"c808750c",
          4189 => x"81f59433",
          4190 => x"70842981",
          4191 => x"f4bc0570",
          4192 => x"0851565a",
          4193 => x"74802ea6",
          4194 => x"38755378",
          4195 => x"527451d6",
          4196 => x"a13f81f5",
          4197 => x"94338105",
          4198 => x"557481f5",
          4199 => x"94347481",
          4200 => x"ff065593",
          4201 => x"75278738",
          4202 => x"800b81f5",
          4203 => x"94347780",
          4204 => x"2eb63881",
          4205 => x"f5900856",
          4206 => x"75802eac",
          4207 => x"3881f58c",
          4208 => x"335574a4",
          4209 => x"388c3dfc",
          4210 => x"05547653",
          4211 => x"78527551",
          4212 => x"80c8913f",
          4213 => x"81f59008",
          4214 => x"528a5180",
          4215 => x"fd9e3f81",
          4216 => x"f5900851",
          4217 => x"80cbee3f",
          4218 => x"8c3d0d04",
          4219 => x"dc3d0d81",
          4220 => x"57805281",
          4221 => x"f5900851",
          4222 => x"80d2873f",
          4223 => x"81f8c808",
          4224 => x"80d13881",
          4225 => x"f5900853",
          4226 => x"80f85288",
          4227 => x"3d705256",
          4228 => x"80fad53f",
          4229 => x"81f8c808",
          4230 => x"802eb838",
          4231 => x"7551d8ad",
          4232 => x"3f81f8c8",
          4233 => x"0855800b",
          4234 => x"81f8c808",
          4235 => x"259c3881",
          4236 => x"f8c808ff",
          4237 => x"05701755",
          4238 => x"55807434",
          4239 => x"75537652",
          4240 => x"811781e3",
          4241 => x"dc5257f6",
          4242 => x"ff3f74ff",
          4243 => x"2e098106",
          4244 => x"ffb138a6",
          4245 => x"3d0d04d9",
          4246 => x"3d0daa3d",
          4247 => x"08ad3d08",
          4248 => x"5a5a8170",
          4249 => x"58588052",
          4250 => x"81f59008",
          4251 => x"5180d192",
          4252 => x"3f81f8c8",
          4253 => x"08819138",
          4254 => x"ff0b81f5",
          4255 => x"90085455",
          4256 => x"80f8528b",
          4257 => x"3d705256",
          4258 => x"80f9dd3f",
          4259 => x"81f8c808",
          4260 => x"802ea438",
          4261 => x"7551d7b5",
          4262 => x"3f81f8c8",
          4263 => x"08811858",
          4264 => x"55800b81",
          4265 => x"f8c80825",
          4266 => x"8e3881f8",
          4267 => x"c808ff05",
          4268 => x"70175555",
          4269 => x"80743474",
          4270 => x"09703070",
          4271 => x"72079f2a",
          4272 => x"51555578",
          4273 => x"772e8538",
          4274 => x"73ffad38",
          4275 => x"81f59008",
          4276 => x"8c110853",
          4277 => x"5180d0aa",
          4278 => x"3f81f8c8",
          4279 => x"08802e88",
          4280 => x"3881e3e8",
          4281 => x"51effd3f",
          4282 => x"78772e09",
          4283 => x"81069938",
          4284 => x"75527951",
          4285 => x"d5e83f79",
          4286 => x"51d6d23f",
          4287 => x"ab3d0854",
          4288 => x"81f8c808",
          4289 => x"74348058",
          4290 => x"7781f8c8",
          4291 => x"0ca93d0d",
          4292 => x"04f63d0d",
          4293 => x"7c7e715c",
          4294 => x"71723357",
          4295 => x"595a5873",
          4296 => x"a02e0981",
          4297 => x"06a23878",
          4298 => x"33780556",
          4299 => x"77762798",
          4300 => x"38811770",
          4301 => x"5b707133",
          4302 => x"56585573",
          4303 => x"a02e0981",
          4304 => x"06863875",
          4305 => x"7526ea38",
          4306 => x"80547388",
          4307 => x"2981f598",
          4308 => x"05700852",
          4309 => x"55d5f63f",
          4310 => x"81f8c808",
          4311 => x"53795274",
          4312 => x"0851d6ca",
          4313 => x"3f81f8c8",
          4314 => x"0880c438",
          4315 => x"84153355",
          4316 => x"74812e88",
          4317 => x"3874822e",
          4318 => x"8838b439",
          4319 => x"fcee3fab",
          4320 => x"39811a5a",
          4321 => x"8c3dfc11",
          4322 => x"53f80551",
          4323 => x"f6af3f81",
          4324 => x"f8c80880",
          4325 => x"2e99387a",
          4326 => x"53785277",
          4327 => x"51fdb83f",
          4328 => x"81f8c808",
          4329 => x"81ff0655",
          4330 => x"74853874",
          4331 => x"54913981",
          4332 => x"147081ff",
          4333 => x"06515482",
          4334 => x"7427ff8e",
          4335 => x"38805473",
          4336 => x"81f8c80c",
          4337 => x"8c3d0d04",
          4338 => x"d33d0db0",
          4339 => x"3d080284",
          4340 => x"0581c305",
          4341 => x"335f5a80",
          4342 => x"0baf3d34",
          4343 => x"81f59433",
          4344 => x"5b81f590",
          4345 => x"0881a338",
          4346 => x"81f58c33",
          4347 => x"5473819a",
          4348 => x"38a851eb",
          4349 => x"b43f81f8",
          4350 => x"c80881f5",
          4351 => x"900c81f8",
          4352 => x"c808802e",
          4353 => x"80fe3893",
          4354 => x"5381f4b8",
          4355 => x"085281f8",
          4356 => x"c80851bb",
          4357 => x"ed3f81f8",
          4358 => x"c808802e",
          4359 => x"8b3881e4",
          4360 => x"9451f3a4",
          4361 => x"3f80e339",
          4362 => x"81f59008",
          4363 => x"5380f852",
          4364 => x"903d7052",
          4365 => x"5480f6b0",
          4366 => x"3f81f8c8",
          4367 => x"085681f8",
          4368 => x"c808742e",
          4369 => x"09810680",
          4370 => x"c13881f8",
          4371 => x"c80851d3",
          4372 => x"fc3f81f8",
          4373 => x"c8085580",
          4374 => x"0b81f8c8",
          4375 => x"08259a38",
          4376 => x"81f8c808",
          4377 => x"ff057017",
          4378 => x"55558074",
          4379 => x"34805374",
          4380 => x"81ff0652",
          4381 => x"7551f9b4",
          4382 => x"3f74ff2e",
          4383 => x"098106ff",
          4384 => x"a7388739",
          4385 => x"810b81f5",
          4386 => x"8c348f3d",
          4387 => x"5dddce3f",
          4388 => x"81f8c808",
          4389 => x"982b7098",
          4390 => x"2c515978",
          4391 => x"ff2eee38",
          4392 => x"7881ff06",
          4393 => x"81f8ec33",
          4394 => x"70982b70",
          4395 => x"982c81f8",
          4396 => x"e8337098",
          4397 => x"2b70972c",
          4398 => x"71982c05",
          4399 => x"70842981",
          4400 => x"e4c40570",
          4401 => x"08157033",
          4402 => x"51515151",
          4403 => x"59595159",
          4404 => x"5d588156",
          4405 => x"73782e80",
          4406 => x"e9387774",
          4407 => x"27b43874",
          4408 => x"81800a29",
          4409 => x"81ff0a05",
          4410 => x"70982c51",
          4411 => x"55807524",
          4412 => x"80ce3876",
          4413 => x"53745277",
          4414 => x"51f7a63f",
          4415 => x"81f8c808",
          4416 => x"81ff0654",
          4417 => x"73802ed7",
          4418 => x"387481f8",
          4419 => x"e8348156",
          4420 => x"b1397481",
          4421 => x"800a2981",
          4422 => x"800a0570",
          4423 => x"982c7081",
          4424 => x"ff065651",
          4425 => x"55738a26",
          4426 => x"97387653",
          4427 => x"74527751",
          4428 => x"f6ef3f81",
          4429 => x"f8c80881",
          4430 => x"ff065473",
          4431 => x"cc38d339",
          4432 => x"80567580",
          4433 => x"2e80ca38",
          4434 => x"811c5574",
          4435 => x"81f8ec34",
          4436 => x"74982b70",
          4437 => x"982c81f8",
          4438 => x"e8337098",
          4439 => x"2b70982c",
          4440 => x"70101170",
          4441 => x"822b81e4",
          4442 => x"c811335e",
          4443 => x"51515157",
          4444 => x"58515574",
          4445 => x"772e0981",
          4446 => x"06fe9238",
          4447 => x"81e4cc14",
          4448 => x"087d0c80",
          4449 => x"0b81f8ec",
          4450 => x"34800b81",
          4451 => x"f8e83492",
          4452 => x"397581f8",
          4453 => x"ec347581",
          4454 => x"f8e83478",
          4455 => x"af3d3475",
          4456 => x"7d0c7e54",
          4457 => x"738b26fd",
          4458 => x"e1387384",
          4459 => x"2981dcd0",
          4460 => x"05547308",
          4461 => x"0481f8f4",
          4462 => x"3354737e",
          4463 => x"2efdcb38",
          4464 => x"81f8f033",
          4465 => x"55737527",
          4466 => x"ab387498",
          4467 => x"2b70982c",
          4468 => x"51557375",
          4469 => x"249e3874",
          4470 => x"1a547333",
          4471 => x"81153474",
          4472 => x"81800a29",
          4473 => x"81ff0a05",
          4474 => x"70982c81",
          4475 => x"f8f43356",
          4476 => x"5155df39",
          4477 => x"81f8f433",
          4478 => x"81115654",
          4479 => x"7481f8f4",
          4480 => x"34731a54",
          4481 => x"ae3d3374",
          4482 => x"3481f8f0",
          4483 => x"3354737e",
          4484 => x"27893881",
          4485 => x"14547381",
          4486 => x"f8f03481",
          4487 => x"f8f43370",
          4488 => x"81800a29",
          4489 => x"81ff0a05",
          4490 => x"70982c81",
          4491 => x"f8f0335a",
          4492 => x"51565674",
          4493 => x"7725a238",
          4494 => x"741a7033",
          4495 => x"5254e8c7",
          4496 => x"3f748180",
          4497 => x"0a298180",
          4498 => x"0a057098",
          4499 => x"2c81f8f0",
          4500 => x"33565155",
          4501 => x"737524e0",
          4502 => x"3881f8f4",
          4503 => x"3370982b",
          4504 => x"70982c81",
          4505 => x"f8f0335a",
          4506 => x"51565674",
          4507 => x"7725fc9a",
          4508 => x"388851e8",
          4509 => x"923f7481",
          4510 => x"800a2981",
          4511 => x"800a0570",
          4512 => x"982c81f8",
          4513 => x"f0335651",
          4514 => x"55737524",
          4515 => x"e438fbfa",
          4516 => x"3981f8f4",
          4517 => x"337081ff",
          4518 => x"06555573",
          4519 => x"802efbea",
          4520 => x"3881f8f0",
          4521 => x"33ff0554",
          4522 => x"7381f8f0",
          4523 => x"34ff1554",
          4524 => x"7381f8f4",
          4525 => x"348851e7",
          4526 => x"ce3f81f8",
          4527 => x"f4337098",
          4528 => x"2b70982c",
          4529 => x"81f8f033",
          4530 => x"57515657",
          4531 => x"747425a7",
          4532 => x"38741a54",
          4533 => x"81143374",
          4534 => x"34733351",
          4535 => x"e7a93f74",
          4536 => x"81800a29",
          4537 => x"81800a05",
          4538 => x"70982c81",
          4539 => x"f8f03358",
          4540 => x"51557575",
          4541 => x"24db38a0",
          4542 => x"51e78c3f",
          4543 => x"81f8f433",
          4544 => x"70982b70",
          4545 => x"982c81f8",
          4546 => x"f0335751",
          4547 => x"56577474",
          4548 => x"24faf738",
          4549 => x"8851e6ef",
          4550 => x"3f748180",
          4551 => x"0a298180",
          4552 => x"0a057098",
          4553 => x"2c81f8f0",
          4554 => x"33585155",
          4555 => x"757525e4",
          4556 => x"38fad739",
          4557 => x"81f8f033",
          4558 => x"7a055480",
          4559 => x"74348a51",
          4560 => x"e6c53f81",
          4561 => x"f8f05279",
          4562 => x"51f7c63f",
          4563 => x"81f8c808",
          4564 => x"81ff0654",
          4565 => x"73983881",
          4566 => x"f8f03354",
          4567 => x"73802e84",
          4568 => x"c9388153",
          4569 => x"73527951",
          4570 => x"f3c23f84",
          4571 => x"bd39807a",
          4572 => x"3484b739",
          4573 => x"81f8f433",
          4574 => x"5473802e",
          4575 => x"fa8c3888",
          4576 => x"51e6843f",
          4577 => x"81f8f433",
          4578 => x"ff055473",
          4579 => x"81f8f434",
          4580 => x"7381ff06",
          4581 => x"54e33981",
          4582 => x"f8f43381",
          4583 => x"f8f03355",
          4584 => x"5573752e",
          4585 => x"f9e438ff",
          4586 => x"14547381",
          4587 => x"f8f03474",
          4588 => x"982b7098",
          4589 => x"2c7581ff",
          4590 => x"06565155",
          4591 => x"747425a7",
          4592 => x"38741a54",
          4593 => x"81143374",
          4594 => x"34733351",
          4595 => x"e5b93f74",
          4596 => x"81800a29",
          4597 => x"81800a05",
          4598 => x"70982c81",
          4599 => x"f8f03358",
          4600 => x"51557575",
          4601 => x"24db38a0",
          4602 => x"51e59c3f",
          4603 => x"81f8f433",
          4604 => x"70982b70",
          4605 => x"982c81f8",
          4606 => x"f0335751",
          4607 => x"56577474",
          4608 => x"24f98738",
          4609 => x"8851e4ff",
          4610 => x"3f748180",
          4611 => x"0a298180",
          4612 => x"0a057098",
          4613 => x"2c81f8f0",
          4614 => x"33585155",
          4615 => x"757525e4",
          4616 => x"38f8e739",
          4617 => x"81f8f433",
          4618 => x"7081ff06",
          4619 => x"81f8f033",
          4620 => x"59565474",
          4621 => x"7727f8d2",
          4622 => x"38811454",
          4623 => x"7381f8f4",
          4624 => x"34741a70",
          4625 => x"335254e4",
          4626 => x"be3f81f8",
          4627 => x"f4337081",
          4628 => x"ff0681f8",
          4629 => x"f0335856",
          4630 => x"54757526",
          4631 => x"dc38f8aa",
          4632 => x"397aae38",
          4633 => x"81f58808",
          4634 => x"5574802e",
          4635 => x"a4387451",
          4636 => x"cbdb3f81",
          4637 => x"f8c80881",
          4638 => x"f8f03481",
          4639 => x"f8c80881",
          4640 => x"ff068105",
          4641 => x"53745279",
          4642 => x"51c8a73f",
          4643 => x"935b81c1",
          4644 => x"397a8429",
          4645 => x"81f4bc05",
          4646 => x"fc110856",
          4647 => x"5474802e",
          4648 => x"a5387451",
          4649 => x"cba73f81",
          4650 => x"f8c80881",
          4651 => x"f8f03481",
          4652 => x"f8c80881",
          4653 => x"ff068105",
          4654 => x"53745279",
          4655 => x"51c7f33f",
          4656 => x"ff1b5480",
          4657 => x"de397308",
          4658 => x"5574802e",
          4659 => x"f7bc3874",
          4660 => x"51cafa3f",
          4661 => x"80e2397a",
          4662 => x"932e0981",
          4663 => x"06933881",
          4664 => x"f4bc0855",
          4665 => x"74802e89",
          4666 => x"387451ca",
          4667 => x"e03f80c8",
          4668 => x"397a8429",
          4669 => x"81f4bc05",
          4670 => x"84110856",
          4671 => x"5474802e",
          4672 => x"a9387451",
          4673 => x"cac73f81",
          4674 => x"f8c80881",
          4675 => x"f8f03481",
          4676 => x"f8c80881",
          4677 => x"ff068105",
          4678 => x"53745279",
          4679 => x"51c7933f",
          4680 => x"811b5473",
          4681 => x"81ff065b",
          4682 => x"a8397308",
          4683 => x"5574802e",
          4684 => x"f6d83874",
          4685 => x"51ca963f",
          4686 => x"81f8c808",
          4687 => x"81f8f034",
          4688 => x"81f8c808",
          4689 => x"81ff0681",
          4690 => x"05537452",
          4691 => x"7951c6e2",
          4692 => x"3f81f8f4",
          4693 => x"5381f8f0",
          4694 => x"33527951",
          4695 => x"ef903ff6",
          4696 => x"a93981f8",
          4697 => x"f4337081",
          4698 => x"ff0681f8",
          4699 => x"f0335956",
          4700 => x"54747727",
          4701 => x"f6943881",
          4702 => x"14547381",
          4703 => x"f8f43474",
          4704 => x"1a703352",
          4705 => x"54e2803f",
          4706 => x"f6803981",
          4707 => x"f8f43354",
          4708 => x"73802ef5",
          4709 => x"f5388851",
          4710 => x"e1ed3f81",
          4711 => x"f8f433ff",
          4712 => x"05547381",
          4713 => x"f8f434f5",
          4714 => x"e139800b",
          4715 => x"81f8f434",
          4716 => x"800b81f8",
          4717 => x"f0347981",
          4718 => x"f8c80caf",
          4719 => x"3d0d04ff",
          4720 => x"3d0d028f",
          4721 => x"05335181",
          4722 => x"52707226",
          4723 => x"873881f5",
          4724 => x"b0113352",
          4725 => x"7181f8c8",
          4726 => x"0c833d0d",
          4727 => x"04fc3d0d",
          4728 => x"029b0533",
          4729 => x"0284059f",
          4730 => x"05335653",
          4731 => x"83517281",
          4732 => x"2680e038",
          4733 => x"72842b87",
          4734 => x"c0928c11",
          4735 => x"53518854",
          4736 => x"74802e84",
          4737 => x"38818854",
          4738 => x"73720c87",
          4739 => x"c0928c11",
          4740 => x"5181710c",
          4741 => x"850b87c0",
          4742 => x"988c0c70",
          4743 => x"52710870",
          4744 => x"82065151",
          4745 => x"70802e8a",
          4746 => x"3887c098",
          4747 => x"8c085170",
          4748 => x"ec387108",
          4749 => x"fc808006",
          4750 => x"52719238",
          4751 => x"87c0988c",
          4752 => x"08517080",
          4753 => x"2e873871",
          4754 => x"81f5b014",
          4755 => x"3481f5b0",
          4756 => x"13335170",
          4757 => x"81f8c80c",
          4758 => x"863d0d04",
          4759 => x"f33d0d60",
          4760 => x"6264028c",
          4761 => x"05bf0533",
          4762 => x"5740585b",
          4763 => x"8374525a",
          4764 => x"fecd3f81",
          4765 => x"f8c80881",
          4766 => x"067a5452",
          4767 => x"7181be38",
          4768 => x"71727584",
          4769 => x"2b87c092",
          4770 => x"801187c0",
          4771 => x"928c1287",
          4772 => x"c0928413",
          4773 => x"415a4057",
          4774 => x"5a58850b",
          4775 => x"87c0988c",
          4776 => x"0c767d0c",
          4777 => x"84760c75",
          4778 => x"0870852a",
          4779 => x"70810651",
          4780 => x"53547180",
          4781 => x"2e8e387b",
          4782 => x"0852717b",
          4783 => x"7081055d",
          4784 => x"34811959",
          4785 => x"8074a206",
          4786 => x"53537173",
          4787 => x"2e833881",
          4788 => x"537883ff",
          4789 => x"268f3872",
          4790 => x"802e8a38",
          4791 => x"87c0988c",
          4792 => x"085271c3",
          4793 => x"3887c098",
          4794 => x"8c085271",
          4795 => x"802e8738",
          4796 => x"7884802e",
          4797 => x"99388176",
          4798 => x"0c87c092",
          4799 => x"8c155372",
          4800 => x"08708206",
          4801 => x"515271f7",
          4802 => x"38ff1a5a",
          4803 => x"8d398480",
          4804 => x"17811970",
          4805 => x"81ff065a",
          4806 => x"53577980",
          4807 => x"2e903873",
          4808 => x"fc808006",
          4809 => x"52718738",
          4810 => x"7d7826fe",
          4811 => x"ed3873fc",
          4812 => x"80800652",
          4813 => x"71802e83",
          4814 => x"38815271",
          4815 => x"537281f8",
          4816 => x"c80c8f3d",
          4817 => x"0d04f33d",
          4818 => x"0d606264",
          4819 => x"028c05bf",
          4820 => x"05335740",
          4821 => x"585b8359",
          4822 => x"80745258",
          4823 => x"fce13f81",
          4824 => x"f8c80881",
          4825 => x"06795452",
          4826 => x"71782e09",
          4827 => x"810681b1",
          4828 => x"38777484",
          4829 => x"2b87c092",
          4830 => x"801187c0",
          4831 => x"928c1287",
          4832 => x"c0928413",
          4833 => x"40595f56",
          4834 => x"5a850b87",
          4835 => x"c0988c0c",
          4836 => x"767d0c82",
          4837 => x"760c8058",
          4838 => x"75087084",
          4839 => x"2a708106",
          4840 => x"51535471",
          4841 => x"802e8c38",
          4842 => x"7a708105",
          4843 => x"5c337c0c",
          4844 => x"81185873",
          4845 => x"812a7081",
          4846 => x"06515271",
          4847 => x"802e8a38",
          4848 => x"87c0988c",
          4849 => x"085271d0",
          4850 => x"3887c098",
          4851 => x"8c085271",
          4852 => x"802e8738",
          4853 => x"7784802e",
          4854 => x"99388176",
          4855 => x"0c87c092",
          4856 => x"8c155372",
          4857 => x"08708206",
          4858 => x"515271f7",
          4859 => x"38ff1959",
          4860 => x"8d39811a",
          4861 => x"7081ff06",
          4862 => x"84801959",
          4863 => x"5b527880",
          4864 => x"2e903873",
          4865 => x"fc808006",
          4866 => x"52718738",
          4867 => x"7d7a26fe",
          4868 => x"f83873fc",
          4869 => x"80800652",
          4870 => x"71802e83",
          4871 => x"38815271",
          4872 => x"537281f8",
          4873 => x"c80c8f3d",
          4874 => x"0d04fa3d",
          4875 => x"0d7a0284",
          4876 => x"05a30533",
          4877 => x"028805a7",
          4878 => x"05337154",
          4879 => x"545657fa",
          4880 => x"fe3f81f8",
          4881 => x"c8088106",
          4882 => x"53835472",
          4883 => x"80fe3885",
          4884 => x"0b87c098",
          4885 => x"8c0c8156",
          4886 => x"71762e80",
          4887 => x"dc387176",
          4888 => x"24933874",
          4889 => x"842b87c0",
          4890 => x"928c1154",
          4891 => x"5471802e",
          4892 => x"8d3880d4",
          4893 => x"3971832e",
          4894 => x"80c63880",
          4895 => x"cb397208",
          4896 => x"70812a70",
          4897 => x"81065151",
          4898 => x"5271802e",
          4899 => x"8a3887c0",
          4900 => x"988c0852",
          4901 => x"71e83887",
          4902 => x"c0988c08",
          4903 => x"52719638",
          4904 => x"81730c87",
          4905 => x"c0928c14",
          4906 => x"53720870",
          4907 => x"82065152",
          4908 => x"71f73896",
          4909 => x"39805692",
          4910 => x"3988800a",
          4911 => x"770c8539",
          4912 => x"8180770c",
          4913 => x"72568339",
          4914 => x"84567554",
          4915 => x"7381f8c8",
          4916 => x"0c883d0d",
          4917 => x"04fe3d0d",
          4918 => x"74811133",
          4919 => x"71337188",
          4920 => x"2b0781f8",
          4921 => x"c80c5351",
          4922 => x"843d0d04",
          4923 => x"fd3d0d75",
          4924 => x"83113382",
          4925 => x"12337190",
          4926 => x"2b71882b",
          4927 => x"07811433",
          4928 => x"70720788",
          4929 => x"2b753371",
          4930 => x"0781f8c8",
          4931 => x"0c525354",
          4932 => x"56545285",
          4933 => x"3d0d04ff",
          4934 => x"3d0d7302",
          4935 => x"84059205",
          4936 => x"22525270",
          4937 => x"72708105",
          4938 => x"54347088",
          4939 => x"2a517072",
          4940 => x"34833d0d",
          4941 => x"04ff3d0d",
          4942 => x"73755252",
          4943 => x"70727081",
          4944 => x"05543470",
          4945 => x"882a5170",
          4946 => x"72708105",
          4947 => x"54347088",
          4948 => x"2a517072",
          4949 => x"70810554",
          4950 => x"3470882a",
          4951 => x"51707234",
          4952 => x"833d0d04",
          4953 => x"fe3d0d76",
          4954 => x"75775454",
          4955 => x"5170802e",
          4956 => x"92387170",
          4957 => x"81055333",
          4958 => x"73708105",
          4959 => x"5534ff11",
          4960 => x"51eb3984",
          4961 => x"3d0d04fe",
          4962 => x"3d0d7577",
          4963 => x"76545253",
          4964 => x"72727081",
          4965 => x"055434ff",
          4966 => x"115170f4",
          4967 => x"38843d0d",
          4968 => x"04fc3d0d",
          4969 => x"78777956",
          4970 => x"56537470",
          4971 => x"81055633",
          4972 => x"74708105",
          4973 => x"56337171",
          4974 => x"31ff1656",
          4975 => x"52525272",
          4976 => x"802e8638",
          4977 => x"71802ee2",
          4978 => x"387181f8",
          4979 => x"c80c863d",
          4980 => x"0d04fe3d",
          4981 => x"0d747654",
          4982 => x"51893971",
          4983 => x"732e8a38",
          4984 => x"81115170",
          4985 => x"335271f3",
          4986 => x"38703381",
          4987 => x"f8c80c84",
          4988 => x"3d0d0480",
          4989 => x"0b81f8c8",
          4990 => x"0c04800b",
          4991 => x"81f8c80c",
          4992 => x"04f73d0d",
          4993 => x"7b56800b",
          4994 => x"83173356",
          4995 => x"5a747a2e",
          4996 => x"80d63881",
          4997 => x"54b01608",
          4998 => x"53b41670",
          4999 => x"53811733",
          5000 => x"5259faa2",
          5001 => x"3f81f8c8",
          5002 => x"087a2e09",
          5003 => x"8106b738",
          5004 => x"81f8c808",
          5005 => x"831734b0",
          5006 => x"160870a4",
          5007 => x"1808319c",
          5008 => x"18085956",
          5009 => x"58747727",
          5010 => x"9f388216",
          5011 => x"33557482",
          5012 => x"2e098106",
          5013 => x"93388154",
          5014 => x"76185378",
          5015 => x"52811633",
          5016 => x"51f9e33f",
          5017 => x"8339815a",
          5018 => x"7981f8c8",
          5019 => x"0c8b3d0d",
          5020 => x"04fa3d0d",
          5021 => x"787a5656",
          5022 => x"805774b0",
          5023 => x"17082eaf",
          5024 => x"387551fe",
          5025 => x"fc3f81f8",
          5026 => x"c8085781",
          5027 => x"f8c8089f",
          5028 => x"38815474",
          5029 => x"53b41652",
          5030 => x"81163351",
          5031 => x"f7be3f81",
          5032 => x"f8c80880",
          5033 => x"2e8538ff",
          5034 => x"55815774",
          5035 => x"b0170c76",
          5036 => x"81f8c80c",
          5037 => x"883d0d04",
          5038 => x"f83d0d7a",
          5039 => x"705257fe",
          5040 => x"c03f81f8",
          5041 => x"c8085881",
          5042 => x"f8c80881",
          5043 => x"91387633",
          5044 => x"5574832e",
          5045 => x"09810680",
          5046 => x"f0388417",
          5047 => x"33597881",
          5048 => x"2e098106",
          5049 => x"80e33884",
          5050 => x"805381f8",
          5051 => x"c80852b4",
          5052 => x"17705256",
          5053 => x"fd913f82",
          5054 => x"d4d55284",
          5055 => x"b21751fc",
          5056 => x"963f848b",
          5057 => x"85a4d252",
          5058 => x"7551fca9",
          5059 => x"3f868a85",
          5060 => x"e4f25284",
          5061 => x"981751fc",
          5062 => x"9c3f9017",
          5063 => x"0852849c",
          5064 => x"1751fc91",
          5065 => x"3f8c1708",
          5066 => x"5284a017",
          5067 => x"51fc863f",
          5068 => x"a0170881",
          5069 => x"0570b019",
          5070 => x"0c795553",
          5071 => x"75528117",
          5072 => x"3351f882",
          5073 => x"3f778418",
          5074 => x"34805380",
          5075 => x"52811733",
          5076 => x"51f9d73f",
          5077 => x"81f8c808",
          5078 => x"802e8338",
          5079 => x"81587781",
          5080 => x"f8c80c8a",
          5081 => x"3d0d04fb",
          5082 => x"3d0d77fe",
          5083 => x"1a981208",
          5084 => x"fe055556",
          5085 => x"54805674",
          5086 => x"73278d38",
          5087 => x"8a142275",
          5088 => x"7129ac16",
          5089 => x"08055753",
          5090 => x"7581f8c8",
          5091 => x"0c873d0d",
          5092 => x"04f93d0d",
          5093 => x"7a7a7008",
          5094 => x"56545781",
          5095 => x"772781df",
          5096 => x"38769815",
          5097 => x"082781d7",
          5098 => x"38ff7433",
          5099 => x"54587282",
          5100 => x"2e80f538",
          5101 => x"72822489",
          5102 => x"3872812e",
          5103 => x"8d3881bf",
          5104 => x"3972832e",
          5105 => x"818e3881",
          5106 => x"b6397681",
          5107 => x"2a177089",
          5108 => x"2aa41608",
          5109 => x"05537452",
          5110 => x"55fd963f",
          5111 => x"81f8c808",
          5112 => x"819f3874",
          5113 => x"83ff0614",
          5114 => x"b4113381",
          5115 => x"1770892a",
          5116 => x"a4180805",
          5117 => x"55765457",
          5118 => x"5753fcf5",
          5119 => x"3f81f8c8",
          5120 => x"0880fe38",
          5121 => x"7483ff06",
          5122 => x"14b41133",
          5123 => x"70882b78",
          5124 => x"07798106",
          5125 => x"71842a5c",
          5126 => x"52585153",
          5127 => x"7280e238",
          5128 => x"759fff06",
          5129 => x"5880da39",
          5130 => x"76882aa4",
          5131 => x"15080552",
          5132 => x"7351fcbd",
          5133 => x"3f81f8c8",
          5134 => x"0880c638",
          5135 => x"761083fe",
          5136 => x"067405b4",
          5137 => x"0551f98d",
          5138 => x"3f81f8c8",
          5139 => x"0883ffff",
          5140 => x"0658ae39",
          5141 => x"76872aa4",
          5142 => x"15080552",
          5143 => x"7351fc91",
          5144 => x"3f81f8c8",
          5145 => x"089b3876",
          5146 => x"822b83fc",
          5147 => x"067405b4",
          5148 => x"0551f8f8",
          5149 => x"3f81f8c8",
          5150 => x"08f00a06",
          5151 => x"58833981",
          5152 => x"587781f8",
          5153 => x"c80c893d",
          5154 => x"0d04f83d",
          5155 => x"0d7a7c7e",
          5156 => x"5a585682",
          5157 => x"59817727",
          5158 => x"829e3876",
          5159 => x"98170827",
          5160 => x"82963875",
          5161 => x"33537279",
          5162 => x"2e819d38",
          5163 => x"72792489",
          5164 => x"3872812e",
          5165 => x"8d388280",
          5166 => x"3972832e",
          5167 => x"81b83881",
          5168 => x"f7397681",
          5169 => x"2a177089",
          5170 => x"2aa41808",
          5171 => x"05537652",
          5172 => x"55fb9e3f",
          5173 => x"81f8c808",
          5174 => x"5981f8c8",
          5175 => x"0881d938",
          5176 => x"7483ff06",
          5177 => x"16b40581",
          5178 => x"16788106",
          5179 => x"59565477",
          5180 => x"5376802e",
          5181 => x"8f387784",
          5182 => x"2b9ff006",
          5183 => x"74338f06",
          5184 => x"71075153",
          5185 => x"72743481",
          5186 => x"0b831734",
          5187 => x"74892aa4",
          5188 => x"17080552",
          5189 => x"7551fad9",
          5190 => x"3f81f8c8",
          5191 => x"085981f8",
          5192 => x"c8088194",
          5193 => x"387483ff",
          5194 => x"0616b405",
          5195 => x"78842a54",
          5196 => x"54768f38",
          5197 => x"77882a74",
          5198 => x"3381f006",
          5199 => x"718f0607",
          5200 => x"51537274",
          5201 => x"3480ec39",
          5202 => x"76882aa4",
          5203 => x"17080552",
          5204 => x"7551fa9d",
          5205 => x"3f81f8c8",
          5206 => x"085981f8",
          5207 => x"c80880d8",
          5208 => x"387783ff",
          5209 => x"ff065276",
          5210 => x"1083fe06",
          5211 => x"7605b405",
          5212 => x"51f7a43f",
          5213 => x"be397687",
          5214 => x"2aa41708",
          5215 => x"05527551",
          5216 => x"f9ef3f81",
          5217 => x"f8c80859",
          5218 => x"81f8c808",
          5219 => x"ab3877f0",
          5220 => x"0a067782",
          5221 => x"2b83fc06",
          5222 => x"7018b405",
          5223 => x"70545154",
          5224 => x"54f6c93f",
          5225 => x"81f8c808",
          5226 => x"8f0a0674",
          5227 => x"07527251",
          5228 => x"f7833f81",
          5229 => x"0b831734",
          5230 => x"7881f8c8",
          5231 => x"0c8a3d0d",
          5232 => x"04f83d0d",
          5233 => x"7a7c7e72",
          5234 => x"08595656",
          5235 => x"59817527",
          5236 => x"a4387498",
          5237 => x"1708279d",
          5238 => x"3873802e",
          5239 => x"aa38ff53",
          5240 => x"73527551",
          5241 => x"fda43f81",
          5242 => x"f8c80854",
          5243 => x"81f8c808",
          5244 => x"80f23893",
          5245 => x"39825480",
          5246 => x"eb398154",
          5247 => x"80e63981",
          5248 => x"f8c80854",
          5249 => x"80de3974",
          5250 => x"527851fb",
          5251 => x"843f81f8",
          5252 => x"c8085881",
          5253 => x"f8c80880",
          5254 => x"2e80c738",
          5255 => x"81f8c808",
          5256 => x"812ed238",
          5257 => x"81f8c808",
          5258 => x"ff2ecf38",
          5259 => x"80537452",
          5260 => x"7551fcd6",
          5261 => x"3f81f8c8",
          5262 => x"08c53898",
          5263 => x"1608fe11",
          5264 => x"90180857",
          5265 => x"55577474",
          5266 => x"27903881",
          5267 => x"1590170c",
          5268 => x"84163381",
          5269 => x"07547384",
          5270 => x"17347755",
          5271 => x"767826ff",
          5272 => x"a6388054",
          5273 => x"7381f8c8",
          5274 => x"0c8a3d0d",
          5275 => x"04f63d0d",
          5276 => x"7c7e7108",
          5277 => x"595b5b79",
          5278 => x"95388c17",
          5279 => x"08587780",
          5280 => x"2e883898",
          5281 => x"17087826",
          5282 => x"b2388158",
          5283 => x"ae397952",
          5284 => x"7a51f9fd",
          5285 => x"3f815574",
          5286 => x"81f8c808",
          5287 => x"2782e038",
          5288 => x"81f8c808",
          5289 => x"5581f8c8",
          5290 => x"08ff2e82",
          5291 => x"d2389817",
          5292 => x"0881f8c8",
          5293 => x"082682c7",
          5294 => x"38795890",
          5295 => x"17087056",
          5296 => x"5473802e",
          5297 => x"82b93877",
          5298 => x"7a2e0981",
          5299 => x"0680e238",
          5300 => x"811a5698",
          5301 => x"17087626",
          5302 => x"83388256",
          5303 => x"75527a51",
          5304 => x"f9af3f80",
          5305 => x"5981f8c8",
          5306 => x"08812e09",
          5307 => x"81068638",
          5308 => x"81f8c808",
          5309 => x"5981f8c8",
          5310 => x"08097030",
          5311 => x"70720780",
          5312 => x"25707c07",
          5313 => x"81f8c808",
          5314 => x"54515155",
          5315 => x"557381ef",
          5316 => x"3881f8c8",
          5317 => x"08802e95",
          5318 => x"388c1708",
          5319 => x"54817427",
          5320 => x"90387398",
          5321 => x"18082789",
          5322 => x"38735885",
          5323 => x"397580db",
          5324 => x"38775681",
          5325 => x"16569817",
          5326 => x"08762689",
          5327 => x"38825675",
          5328 => x"782681ac",
          5329 => x"3875527a",
          5330 => x"51f8c63f",
          5331 => x"81f8c808",
          5332 => x"802eb838",
          5333 => x"805981f8",
          5334 => x"c808812e",
          5335 => x"09810686",
          5336 => x"3881f8c8",
          5337 => x"085981f8",
          5338 => x"c8080970",
          5339 => x"30707207",
          5340 => x"8025707c",
          5341 => x"07515155",
          5342 => x"557380f8",
          5343 => x"3875782e",
          5344 => x"098106ff",
          5345 => x"ae387355",
          5346 => x"80f539ff",
          5347 => x"53755276",
          5348 => x"51f9f73f",
          5349 => x"81f8c808",
          5350 => x"81f8c808",
          5351 => x"307081f8",
          5352 => x"c8080780",
          5353 => x"25515555",
          5354 => x"79802e94",
          5355 => x"3873802e",
          5356 => x"8f387553",
          5357 => x"79527651",
          5358 => x"f9d03f81",
          5359 => x"f8c80855",
          5360 => x"74a53875",
          5361 => x"8c180c98",
          5362 => x"1708fe05",
          5363 => x"90180856",
          5364 => x"54747426",
          5365 => x"8638ff15",
          5366 => x"90180c84",
          5367 => x"17338107",
          5368 => x"54738418",
          5369 => x"349739ff",
          5370 => x"5674812e",
          5371 => x"90388c39",
          5372 => x"80558c39",
          5373 => x"81f8c808",
          5374 => x"55853981",
          5375 => x"56755574",
          5376 => x"81f8c80c",
          5377 => x"8c3d0d04",
          5378 => x"f83d0d7a",
          5379 => x"705255f3",
          5380 => x"f03f81f8",
          5381 => x"c8085881",
          5382 => x"5681f8c8",
          5383 => x"0880d838",
          5384 => x"7b527451",
          5385 => x"f6c13f81",
          5386 => x"f8c80881",
          5387 => x"f8c808b0",
          5388 => x"170c5984",
          5389 => x"80537752",
          5390 => x"b4157052",
          5391 => x"57f2c83f",
          5392 => x"77568439",
          5393 => x"8116568a",
          5394 => x"15225875",
          5395 => x"78279738",
          5396 => x"81547519",
          5397 => x"53765281",
          5398 => x"153351ed",
          5399 => x"e93f81f8",
          5400 => x"c808802e",
          5401 => x"df388a15",
          5402 => x"22763270",
          5403 => x"30707207",
          5404 => x"709f2a53",
          5405 => x"51565675",
          5406 => x"81f8c80c",
          5407 => x"8a3d0d04",
          5408 => x"f83d0d7a",
          5409 => x"7c710858",
          5410 => x"565774f0",
          5411 => x"800a2680",
          5412 => x"f138749f",
          5413 => x"06537280",
          5414 => x"e9387490",
          5415 => x"180c8817",
          5416 => x"085473aa",
          5417 => x"38753353",
          5418 => x"82732788",
          5419 => x"38a81608",
          5420 => x"54739b38",
          5421 => x"74852a53",
          5422 => x"820b8817",
          5423 => x"225a5872",
          5424 => x"792780fe",
          5425 => x"38a81608",
          5426 => x"98180c80",
          5427 => x"cd398a16",
          5428 => x"2270892b",
          5429 => x"54587275",
          5430 => x"26b23873",
          5431 => x"527651f5",
          5432 => x"b03f81f8",
          5433 => x"c8085481",
          5434 => x"f8c808ff",
          5435 => x"2ebd3881",
          5436 => x"0b81f8c8",
          5437 => x"08278b38",
          5438 => x"98160881",
          5439 => x"f8c80826",
          5440 => x"85388258",
          5441 => x"bd397473",
          5442 => x"3155cb39",
          5443 => x"73527551",
          5444 => x"f4d53f81",
          5445 => x"f8c80898",
          5446 => x"180c7394",
          5447 => x"180c9817",
          5448 => x"08538258",
          5449 => x"72802e9a",
          5450 => x"38853981",
          5451 => x"58943974",
          5452 => x"892a1398",
          5453 => x"180c7483",
          5454 => x"ff0616b4",
          5455 => x"059c180c",
          5456 => x"80587781",
          5457 => x"f8c80c8a",
          5458 => x"3d0d04f8",
          5459 => x"3d0d7a70",
          5460 => x"08901208",
          5461 => x"a0055957",
          5462 => x"54f0800a",
          5463 => x"77278638",
          5464 => x"800b9815",
          5465 => x"0c981408",
          5466 => x"53845572",
          5467 => x"802e81cb",
          5468 => x"387683ff",
          5469 => x"06587781",
          5470 => x"b5388113",
          5471 => x"98150c94",
          5472 => x"14085574",
          5473 => x"92387685",
          5474 => x"2a881722",
          5475 => x"56537473",
          5476 => x"26819b38",
          5477 => x"80c0398a",
          5478 => x"1622ff05",
          5479 => x"77892a06",
          5480 => x"5372818a",
          5481 => x"38745273",
          5482 => x"51f3e63f",
          5483 => x"81f8c808",
          5484 => x"53825581",
          5485 => x"0b81f8c8",
          5486 => x"082780ff",
          5487 => x"38815581",
          5488 => x"f8c808ff",
          5489 => x"2e80f438",
          5490 => x"98160881",
          5491 => x"f8c80826",
          5492 => x"80ca387b",
          5493 => x"8a387798",
          5494 => x"150c8455",
          5495 => x"80dd3994",
          5496 => x"14085273",
          5497 => x"51f9863f",
          5498 => x"81f8c808",
          5499 => x"53875581",
          5500 => x"f8c80880",
          5501 => x"2e80c438",
          5502 => x"825581f8",
          5503 => x"c808812e",
          5504 => x"ba388155",
          5505 => x"81f8c808",
          5506 => x"ff2eb038",
          5507 => x"81f8c808",
          5508 => x"527551fb",
          5509 => x"f33f81f8",
          5510 => x"c808a038",
          5511 => x"7294150c",
          5512 => x"72527551",
          5513 => x"f2c13f81",
          5514 => x"f8c80898",
          5515 => x"150c7690",
          5516 => x"150c7716",
          5517 => x"b4059c15",
          5518 => x"0c805574",
          5519 => x"81f8c80c",
          5520 => x"8a3d0d04",
          5521 => x"f73d0d7b",
          5522 => x"7d71085b",
          5523 => x"5b578052",
          5524 => x"7651fcac",
          5525 => x"3f81f8c8",
          5526 => x"085481f8",
          5527 => x"c80880ec",
          5528 => x"3881f8c8",
          5529 => x"08569817",
          5530 => x"08527851",
          5531 => x"f0833f81",
          5532 => x"f8c80854",
          5533 => x"81f8c808",
          5534 => x"80d23881",
          5535 => x"f8c8089c",
          5536 => x"18087033",
          5537 => x"51545872",
          5538 => x"81e52e09",
          5539 => x"81068338",
          5540 => x"815881f8",
          5541 => x"c8085572",
          5542 => x"83388155",
          5543 => x"77750753",
          5544 => x"72802e8e",
          5545 => x"38811656",
          5546 => x"757a2e09",
          5547 => x"81068838",
          5548 => x"a53981f8",
          5549 => x"c8085681",
          5550 => x"527651fd",
          5551 => x"8e3f81f8",
          5552 => x"c8085481",
          5553 => x"f8c80880",
          5554 => x"2eff9b38",
          5555 => x"73842e09",
          5556 => x"81068338",
          5557 => x"87547381",
          5558 => x"f8c80c8b",
          5559 => x"3d0d04fd",
          5560 => x"3d0d769a",
          5561 => x"115254eb",
          5562 => x"ec3f81f8",
          5563 => x"c80883ff",
          5564 => x"ff067670",
          5565 => x"33515353",
          5566 => x"71832e09",
          5567 => x"81069038",
          5568 => x"941451eb",
          5569 => x"d03f81f8",
          5570 => x"c808902b",
          5571 => x"73075372",
          5572 => x"81f8c80c",
          5573 => x"853d0d04",
          5574 => x"fc3d0d77",
          5575 => x"797083ff",
          5576 => x"ff06549a",
          5577 => x"12535555",
          5578 => x"ebed3f76",
          5579 => x"70335153",
          5580 => x"72832e09",
          5581 => x"81068b38",
          5582 => x"73902a52",
          5583 => x"941551eb",
          5584 => x"d63f863d",
          5585 => x"0d04f73d",
          5586 => x"0d7b7d5b",
          5587 => x"55847508",
          5588 => x"5a589815",
          5589 => x"08802e81",
          5590 => x"8a389815",
          5591 => x"08527851",
          5592 => x"ee8f3f81",
          5593 => x"f8c80858",
          5594 => x"81f8c808",
          5595 => x"80f5389c",
          5596 => x"15087033",
          5597 => x"55537386",
          5598 => x"38845880",
          5599 => x"e6398b13",
          5600 => x"3370bf06",
          5601 => x"7081ff06",
          5602 => x"58515372",
          5603 => x"86163481",
          5604 => x"f8c80853",
          5605 => x"7381e52e",
          5606 => x"83388153",
          5607 => x"73ae2ea9",
          5608 => x"38817074",
          5609 => x"06545772",
          5610 => x"802e9e38",
          5611 => x"758f2e99",
          5612 => x"3881f8c8",
          5613 => x"0876df06",
          5614 => x"54547288",
          5615 => x"2e098106",
          5616 => x"83387654",
          5617 => x"737a2ea0",
          5618 => x"38805274",
          5619 => x"51fafc3f",
          5620 => x"81f8c808",
          5621 => x"5881f8c8",
          5622 => x"08893898",
          5623 => x"1508fefa",
          5624 => x"38863980",
          5625 => x"0b98160c",
          5626 => x"7781f8c8",
          5627 => x"0c8b3d0d",
          5628 => x"04fb3d0d",
          5629 => x"77700857",
          5630 => x"54815273",
          5631 => x"51fcc53f",
          5632 => x"81f8c808",
          5633 => x"5581f8c8",
          5634 => x"08b43898",
          5635 => x"14085275",
          5636 => x"51ecde3f",
          5637 => x"81f8c808",
          5638 => x"5581f8c8",
          5639 => x"08a038a0",
          5640 => x"5381f8c8",
          5641 => x"08529c14",
          5642 => x"0851eadb",
          5643 => x"3f8b53a0",
          5644 => x"14529c14",
          5645 => x"0851eaac",
          5646 => x"3f810b83",
          5647 => x"17347481",
          5648 => x"f8c80c87",
          5649 => x"3d0d04fd",
          5650 => x"3d0d7570",
          5651 => x"08981208",
          5652 => x"54705355",
          5653 => x"53ec9a3f",
          5654 => x"81f8c808",
          5655 => x"8d389c13",
          5656 => x"0853e573",
          5657 => x"34810b83",
          5658 => x"1534853d",
          5659 => x"0d04fa3d",
          5660 => x"0d787a57",
          5661 => x"57800b89",
          5662 => x"17349817",
          5663 => x"08802e81",
          5664 => x"82388070",
          5665 => x"89185555",
          5666 => x"559c1708",
          5667 => x"14703381",
          5668 => x"16565152",
          5669 => x"71a02ea8",
          5670 => x"3871852e",
          5671 => x"09810684",
          5672 => x"3881e552",
          5673 => x"73892e09",
          5674 => x"81068b38",
          5675 => x"ae737081",
          5676 => x"05553481",
          5677 => x"15557173",
          5678 => x"70810555",
          5679 => x"34811555",
          5680 => x"8a7427c5",
          5681 => x"38751588",
          5682 => x"0552800b",
          5683 => x"8113349c",
          5684 => x"1708528b",
          5685 => x"12338817",
          5686 => x"349c1708",
          5687 => x"9c115252",
          5688 => x"e88a3f81",
          5689 => x"f8c80876",
          5690 => x"0c961251",
          5691 => x"e7e73f81",
          5692 => x"f8c80886",
          5693 => x"17239812",
          5694 => x"51e7da3f",
          5695 => x"81f8c808",
          5696 => x"84172388",
          5697 => x"3d0d04f3",
          5698 => x"3d0d7f70",
          5699 => x"085e5b80",
          5700 => x"61703351",
          5701 => x"555573af",
          5702 => x"2e833881",
          5703 => x"557380dc",
          5704 => x"2e913874",
          5705 => x"802e8c38",
          5706 => x"941d0888",
          5707 => x"1c0caa39",
          5708 => x"81154180",
          5709 => x"61703356",
          5710 => x"565673af",
          5711 => x"2e098106",
          5712 => x"83388156",
          5713 => x"7380dc32",
          5714 => x"70307080",
          5715 => x"25780751",
          5716 => x"515473dc",
          5717 => x"3873881c",
          5718 => x"0c607033",
          5719 => x"5154739f",
          5720 => x"269638ff",
          5721 => x"800bab1c",
          5722 => x"3480527a",
          5723 => x"51f6913f",
          5724 => x"81f8c808",
          5725 => x"55859839",
          5726 => x"913d61a0",
          5727 => x"1d5c5a5e",
          5728 => x"8b53a052",
          5729 => x"7951e7ff",
          5730 => x"3f807059",
          5731 => x"57887933",
          5732 => x"555c73ae",
          5733 => x"2e098106",
          5734 => x"80d43878",
          5735 => x"18703381",
          5736 => x"1a71ae32",
          5737 => x"7030709f",
          5738 => x"2a738226",
          5739 => x"07515153",
          5740 => x"5a575473",
          5741 => x"8c387917",
          5742 => x"54757434",
          5743 => x"811757db",
          5744 => x"3975af32",
          5745 => x"7030709f",
          5746 => x"2a515154",
          5747 => x"7580dc2e",
          5748 => x"8c387380",
          5749 => x"2e873875",
          5750 => x"a02682bd",
          5751 => x"3877197e",
          5752 => x"0ca454a0",
          5753 => x"762782bd",
          5754 => x"38a05482",
          5755 => x"b8397818",
          5756 => x"7033811a",
          5757 => x"5a5754a0",
          5758 => x"762781fc",
          5759 => x"3875af32",
          5760 => x"70307780",
          5761 => x"dc327030",
          5762 => x"72802571",
          5763 => x"80250751",
          5764 => x"51565155",
          5765 => x"73802eac",
          5766 => x"38843981",
          5767 => x"18588078",
          5768 => x"1a703351",
          5769 => x"555573af",
          5770 => x"2e098106",
          5771 => x"83388155",
          5772 => x"7380dc32",
          5773 => x"70307080",
          5774 => x"25770751",
          5775 => x"515473db",
          5776 => x"3881b539",
          5777 => x"75ae2e09",
          5778 => x"81068338",
          5779 => x"8154767c",
          5780 => x"27740754",
          5781 => x"73802ea2",
          5782 => x"387b8b32",
          5783 => x"703077ae",
          5784 => x"32703072",
          5785 => x"8025719f",
          5786 => x"2a075351",
          5787 => x"56515574",
          5788 => x"81a73888",
          5789 => x"578b5cfe",
          5790 => x"f5397598",
          5791 => x"2b547380",
          5792 => x"258c3875",
          5793 => x"80ff0681",
          5794 => x"e6d81133",
          5795 => x"57547551",
          5796 => x"e6e13f81",
          5797 => x"f8c80880",
          5798 => x"2eb23878",
          5799 => x"18703381",
          5800 => x"1a71545a",
          5801 => x"5654e6d2",
          5802 => x"3f81f8c8",
          5803 => x"08802e80",
          5804 => x"e838ff1c",
          5805 => x"54767427",
          5806 => x"80df3879",
          5807 => x"17547574",
          5808 => x"3481177a",
          5809 => x"11555774",
          5810 => x"7434a739",
          5811 => x"755281e5",
          5812 => x"f851e5fe",
          5813 => x"3f81f8c8",
          5814 => x"08bf38ff",
          5815 => x"9f165473",
          5816 => x"99268938",
          5817 => x"e0167081",
          5818 => x"ff065754",
          5819 => x"79175475",
          5820 => x"74348117",
          5821 => x"57fdf739",
          5822 => x"77197e0c",
          5823 => x"76802e99",
          5824 => x"38793354",
          5825 => x"7381e52e",
          5826 => x"09810684",
          5827 => x"38857a34",
          5828 => x"8454a076",
          5829 => x"278f388b",
          5830 => x"39865581",
          5831 => x"f2398456",
          5832 => x"80f33980",
          5833 => x"54738b1b",
          5834 => x"34807b08",
          5835 => x"58527a51",
          5836 => x"f2ce3f81",
          5837 => x"f8c80856",
          5838 => x"81f8c808",
          5839 => x"80d73898",
          5840 => x"1b085276",
          5841 => x"51e6aa3f",
          5842 => x"81f8c808",
          5843 => x"5681f8c8",
          5844 => x"0880c238",
          5845 => x"9c1b0870",
          5846 => x"33555573",
          5847 => x"802effbe",
          5848 => x"388b1533",
          5849 => x"bf065473",
          5850 => x"861c348b",
          5851 => x"15337083",
          5852 => x"2a708106",
          5853 => x"51555873",
          5854 => x"92388b53",
          5855 => x"79527451",
          5856 => x"e49f3f81",
          5857 => x"f8c80880",
          5858 => x"2e8b3875",
          5859 => x"527a51f3",
          5860 => x"ba3fff9f",
          5861 => x"3975ab1c",
          5862 => x"33575574",
          5863 => x"802ebb38",
          5864 => x"74842e09",
          5865 => x"810680e7",
          5866 => x"3875852a",
          5867 => x"70810677",
          5868 => x"822a5851",
          5869 => x"5473802e",
          5870 => x"96387581",
          5871 => x"06547380",
          5872 => x"2efbb538",
          5873 => x"ff800bab",
          5874 => x"1c348055",
          5875 => x"80c13975",
          5876 => x"81065473",
          5877 => x"ba388555",
          5878 => x"b6397582",
          5879 => x"2a708106",
          5880 => x"515473ab",
          5881 => x"38861b33",
          5882 => x"70842a70",
          5883 => x"81065155",
          5884 => x"5573802e",
          5885 => x"e138901b",
          5886 => x"0883ff06",
          5887 => x"1db40552",
          5888 => x"7c51f5db",
          5889 => x"3f81f8c8",
          5890 => x"08881c0c",
          5891 => x"faea3974",
          5892 => x"81f8c80c",
          5893 => x"8f3d0d04",
          5894 => x"f63d0d7c",
          5895 => x"5bff7b08",
          5896 => x"70717355",
          5897 => x"595c5559",
          5898 => x"73802e81",
          5899 => x"c6387570",
          5900 => x"81055733",
          5901 => x"70a02652",
          5902 => x"5271ba2e",
          5903 => x"8d3870ee",
          5904 => x"3871ba2e",
          5905 => x"09810681",
          5906 => x"a5387333",
          5907 => x"d0117081",
          5908 => x"ff065152",
          5909 => x"53708926",
          5910 => x"91388214",
          5911 => x"7381ff06",
          5912 => x"d0055652",
          5913 => x"71762e80",
          5914 => x"f738800b",
          5915 => x"81e6c859",
          5916 => x"5577087a",
          5917 => x"55577670",
          5918 => x"81055833",
          5919 => x"74708105",
          5920 => x"5633ff9f",
          5921 => x"12535353",
          5922 => x"70992689",
          5923 => x"38e01370",
          5924 => x"81ff0654",
          5925 => x"51ff9f12",
          5926 => x"51709926",
          5927 => x"8938e012",
          5928 => x"7081ff06",
          5929 => x"53517230",
          5930 => x"709f2a51",
          5931 => x"5172722e",
          5932 => x"09810685",
          5933 => x"3870ffbe",
          5934 => x"38723074",
          5935 => x"77327030",
          5936 => x"7072079f",
          5937 => x"2a739f2a",
          5938 => x"07535454",
          5939 => x"5170802e",
          5940 => x"8f388115",
          5941 => x"84195955",
          5942 => x"837525ff",
          5943 => x"94388b39",
          5944 => x"74832486",
          5945 => x"3874767c",
          5946 => x"0c597851",
          5947 => x"863981f9",
          5948 => x"8c335170",
          5949 => x"81f8c80c",
          5950 => x"8c3d0d04",
          5951 => x"fa3d0d78",
          5952 => x"56800b83",
          5953 => x"1734ff0b",
          5954 => x"b0170c79",
          5955 => x"527551e2",
          5956 => x"e03f8455",
          5957 => x"81f8c808",
          5958 => x"81803884",
          5959 => x"b21651df",
          5960 => x"b43f81f8",
          5961 => x"c80883ff",
          5962 => x"ff065483",
          5963 => x"557382d4",
          5964 => x"d52e0981",
          5965 => x"0680e338",
          5966 => x"800bb417",
          5967 => x"33565774",
          5968 => x"81e92e09",
          5969 => x"81068338",
          5970 => x"81577481",
          5971 => x"eb327030",
          5972 => x"70802579",
          5973 => x"07515154",
          5974 => x"738a3874",
          5975 => x"81e82e09",
          5976 => x"8106b538",
          5977 => x"835381e6",
          5978 => x"885280ea",
          5979 => x"1651e0b1",
          5980 => x"3f81f8c8",
          5981 => x"085581f8",
          5982 => x"c808802e",
          5983 => x"9d388553",
          5984 => x"81e68c52",
          5985 => x"81861651",
          5986 => x"e0973f81",
          5987 => x"f8c80855",
          5988 => x"81f8c808",
          5989 => x"802e8338",
          5990 => x"82557481",
          5991 => x"f8c80c88",
          5992 => x"3d0d04f2",
          5993 => x"3d0d6102",
          5994 => x"840580cb",
          5995 => x"05335855",
          5996 => x"80750c60",
          5997 => x"51fce13f",
          5998 => x"81f8c808",
          5999 => x"588b5680",
          6000 => x"0b81f8c8",
          6001 => x"082486fc",
          6002 => x"3881f8c8",
          6003 => x"08842981",
          6004 => x"f8f80570",
          6005 => x"0855538c",
          6006 => x"5673802e",
          6007 => x"86e63873",
          6008 => x"750c7681",
          6009 => x"fe067433",
          6010 => x"54577280",
          6011 => x"2eae3881",
          6012 => x"143351d7",
          6013 => x"ca3f81f8",
          6014 => x"c80881ff",
          6015 => x"06708106",
          6016 => x"54557298",
          6017 => x"3876802e",
          6018 => x"86b83874",
          6019 => x"822a7081",
          6020 => x"0651538a",
          6021 => x"567286ac",
          6022 => x"3886a739",
          6023 => x"80743477",
          6024 => x"81153481",
          6025 => x"52811433",
          6026 => x"51d7b23f",
          6027 => x"81f8c808",
          6028 => x"81ff0670",
          6029 => x"81065455",
          6030 => x"83567286",
          6031 => x"87387680",
          6032 => x"2e8f3874",
          6033 => x"822a7081",
          6034 => x"0651538a",
          6035 => x"567285f4",
          6036 => x"38807053",
          6037 => x"74525bfd",
          6038 => x"a33f81f8",
          6039 => x"c80881ff",
          6040 => x"06577682",
          6041 => x"2e098106",
          6042 => x"80e2388c",
          6043 => x"3d745658",
          6044 => x"835683f6",
          6045 => x"15337058",
          6046 => x"5372802e",
          6047 => x"8d3883fa",
          6048 => x"1551dce8",
          6049 => x"3f81f8c8",
          6050 => x"08577678",
          6051 => x"7084055a",
          6052 => x"0cff1690",
          6053 => x"16565675",
          6054 => x"8025d738",
          6055 => x"800b8d3d",
          6056 => x"54567270",
          6057 => x"84055408",
          6058 => x"5b83577a",
          6059 => x"802e9538",
          6060 => x"7a527351",
          6061 => x"fcc63f81",
          6062 => x"f8c80881",
          6063 => x"ff065781",
          6064 => x"77278938",
          6065 => x"81165683",
          6066 => x"7627d738",
          6067 => x"81567684",
          6068 => x"2e84f138",
          6069 => x"8d567681",
          6070 => x"2684e938",
          6071 => x"bf1451db",
          6072 => x"f43f81f8",
          6073 => x"c80883ff",
          6074 => x"ff065372",
          6075 => x"84802e09",
          6076 => x"810684d0",
          6077 => x"3880ca14",
          6078 => x"51dbda3f",
          6079 => x"81f8c808",
          6080 => x"83ffff06",
          6081 => x"58778d38",
          6082 => x"80d81451",
          6083 => x"dbde3f81",
          6084 => x"f8c80858",
          6085 => x"779c150c",
          6086 => x"80c41433",
          6087 => x"82153480",
          6088 => x"c41433ff",
          6089 => x"117081ff",
          6090 => x"06515455",
          6091 => x"8d567281",
          6092 => x"26849138",
          6093 => x"7481ff06",
          6094 => x"78712980",
          6095 => x"c1163352",
          6096 => x"5953728a",
          6097 => x"15237280",
          6098 => x"2e8b38ff",
          6099 => x"13730653",
          6100 => x"72802e86",
          6101 => x"388d5683",
          6102 => x"eb3980c5",
          6103 => x"1451daf5",
          6104 => x"3f81f8c8",
          6105 => x"085381f8",
          6106 => x"c8088815",
          6107 => x"23728f06",
          6108 => x"578d5676",
          6109 => x"83ce3880",
          6110 => x"c71451da",
          6111 => x"d83f81f8",
          6112 => x"c80883ff",
          6113 => x"ff065574",
          6114 => x"8d3880d4",
          6115 => x"1451dadc",
          6116 => x"3f81f8c8",
          6117 => x"085580c2",
          6118 => x"1451dab9",
          6119 => x"3f81f8c8",
          6120 => x"0883ffff",
          6121 => x"06538d56",
          6122 => x"72802e83",
          6123 => x"97388814",
          6124 => x"22781471",
          6125 => x"842a055a",
          6126 => x"5a787526",
          6127 => x"8386388a",
          6128 => x"14225274",
          6129 => x"793151ff",
          6130 => x"93e13f81",
          6131 => x"f8c80855",
          6132 => x"81f8c808",
          6133 => x"802e82ec",
          6134 => x"3881f8c8",
          6135 => x"0880ffff",
          6136 => x"fff52683",
          6137 => x"38835774",
          6138 => x"83fff526",
          6139 => x"83388257",
          6140 => x"749ff526",
          6141 => x"85388157",
          6142 => x"89398d56",
          6143 => x"76802e82",
          6144 => x"c3388215",
          6145 => x"7098160c",
          6146 => x"7ba0160c",
          6147 => x"731c70a4",
          6148 => x"170c7a1d",
          6149 => x"ac170c54",
          6150 => x"5576832e",
          6151 => x"098106af",
          6152 => x"3880de14",
          6153 => x"51d9ae3f",
          6154 => x"81f8c808",
          6155 => x"83ffff06",
          6156 => x"538d5672",
          6157 => x"828e3879",
          6158 => x"828a3880",
          6159 => x"e01451d9",
          6160 => x"ab3f81f8",
          6161 => x"c808a815",
          6162 => x"0c74822b",
          6163 => x"53a2398d",
          6164 => x"5679802e",
          6165 => x"81ee3877",
          6166 => x"13a8150c",
          6167 => x"74155376",
          6168 => x"822e8d38",
          6169 => x"74101570",
          6170 => x"812a7681",
          6171 => x"06055153",
          6172 => x"83ff1389",
          6173 => x"2a538d56",
          6174 => x"729c1508",
          6175 => x"2681c538",
          6176 => x"ff0b9015",
          6177 => x"0cff0b8c",
          6178 => x"150cff80",
          6179 => x"0b841534",
          6180 => x"76832e09",
          6181 => x"81068192",
          6182 => x"3880e414",
          6183 => x"51d8b63f",
          6184 => x"81f8c808",
          6185 => x"83ffff06",
          6186 => x"5372812e",
          6187 => x"09810680",
          6188 => x"f938811b",
          6189 => x"527351db",
          6190 => x"b83f81f8",
          6191 => x"c80880ea",
          6192 => x"3881f8c8",
          6193 => x"08841534",
          6194 => x"84b21451",
          6195 => x"d8873f81",
          6196 => x"f8c80883",
          6197 => x"ffff0653",
          6198 => x"7282d4d5",
          6199 => x"2e098106",
          6200 => x"80c838b4",
          6201 => x"1451d884",
          6202 => x"3f81f8c8",
          6203 => x"08848b85",
          6204 => x"a4d22e09",
          6205 => x"8106b338",
          6206 => x"84981451",
          6207 => x"d7ee3f81",
          6208 => x"f8c80886",
          6209 => x"8a85e4f2",
          6210 => x"2e098106",
          6211 => x"9d38849c",
          6212 => x"1451d7d8",
          6213 => x"3f81f8c8",
          6214 => x"0890150c",
          6215 => x"84a01451",
          6216 => x"d7ca3f81",
          6217 => x"f8c8088c",
          6218 => x"150c7674",
          6219 => x"3481f988",
          6220 => x"22810553",
          6221 => x"7281f988",
          6222 => x"23728615",
          6223 => x"23800b94",
          6224 => x"150c8056",
          6225 => x"7581f8c8",
          6226 => x"0c903d0d",
          6227 => x"04fb3d0d",
          6228 => x"77548955",
          6229 => x"73802eb9",
          6230 => x"38730853",
          6231 => x"72802eb1",
          6232 => x"38723352",
          6233 => x"71802ea9",
          6234 => x"38861322",
          6235 => x"84152257",
          6236 => x"5271762e",
          6237 => x"09810699",
          6238 => x"38811333",
          6239 => x"51d0c03f",
          6240 => x"81f8c808",
          6241 => x"81065271",
          6242 => x"88387174",
          6243 => x"08545583",
          6244 => x"39805378",
          6245 => x"73710c52",
          6246 => x"7481f8c8",
          6247 => x"0c873d0d",
          6248 => x"04fa3d0d",
          6249 => x"02ab0533",
          6250 => x"7a58893d",
          6251 => x"fc055256",
          6252 => x"f4e63f8b",
          6253 => x"54800b81",
          6254 => x"f8c80824",
          6255 => x"bc3881f8",
          6256 => x"c8088429",
          6257 => x"81f8f805",
          6258 => x"70085555",
          6259 => x"73802e84",
          6260 => x"38807434",
          6261 => x"78547380",
          6262 => x"2e843880",
          6263 => x"74347875",
          6264 => x"0c755475",
          6265 => x"802e9238",
          6266 => x"8053893d",
          6267 => x"70538405",
          6268 => x"51f7b03f",
          6269 => x"81f8c808",
          6270 => x"547381f8",
          6271 => x"c80c883d",
          6272 => x"0d04eb3d",
          6273 => x"0d670284",
          6274 => x"0580e705",
          6275 => x"33595989",
          6276 => x"5478802e",
          6277 => x"84c83877",
          6278 => x"bf067054",
          6279 => x"983dd005",
          6280 => x"53993d84",
          6281 => x"055258f6",
          6282 => x"fa3f81f8",
          6283 => x"c8085581",
          6284 => x"f8c80884",
          6285 => x"a4387a5c",
          6286 => x"68528c3d",
          6287 => x"705256ed",
          6288 => x"c63f81f8",
          6289 => x"c8085581",
          6290 => x"f8c80892",
          6291 => x"380280d7",
          6292 => x"05337098",
          6293 => x"2b555773",
          6294 => x"80258338",
          6295 => x"8655779c",
          6296 => x"06547380",
          6297 => x"2e81ab38",
          6298 => x"74802e95",
          6299 => x"3874842e",
          6300 => x"098106aa",
          6301 => x"387551ea",
          6302 => x"f83f81f8",
          6303 => x"c808559e",
          6304 => x"3902b205",
          6305 => x"33910654",
          6306 => x"7381b838",
          6307 => x"77822a70",
          6308 => x"81065154",
          6309 => x"73802e8e",
          6310 => x"38885583",
          6311 => x"bc397788",
          6312 => x"07587483",
          6313 => x"b4387783",
          6314 => x"2a708106",
          6315 => x"51547380",
          6316 => x"2e81af38",
          6317 => x"62527a51",
          6318 => x"e8a53f81",
          6319 => x"f8c80856",
          6320 => x"8288b20a",
          6321 => x"52628e05",
          6322 => x"51d4ea3f",
          6323 => x"6254a00b",
          6324 => x"8b153480",
          6325 => x"5362527a",
          6326 => x"51e8bd3f",
          6327 => x"8052629c",
          6328 => x"0551d4d1",
          6329 => x"3f7a5481",
          6330 => x"0b831534",
          6331 => x"75802e80",
          6332 => x"f1387ab0",
          6333 => x"11085154",
          6334 => x"80537552",
          6335 => x"973dd405",
          6336 => x"51ddbe3f",
          6337 => x"81f8c808",
          6338 => x"5581f8c8",
          6339 => x"0882ca38",
          6340 => x"b7397482",
          6341 => x"c43802b2",
          6342 => x"05337084",
          6343 => x"2a708106",
          6344 => x"51555673",
          6345 => x"802e8638",
          6346 => x"845582ad",
          6347 => x"3977812a",
          6348 => x"70810651",
          6349 => x"5473802e",
          6350 => x"a9387581",
          6351 => x"06547380",
          6352 => x"2ea03887",
          6353 => x"55829239",
          6354 => x"73527a51",
          6355 => x"d6a33f81",
          6356 => x"f8c8087b",
          6357 => x"ff188c12",
          6358 => x"0c555581",
          6359 => x"f8c80881",
          6360 => x"f8387783",
          6361 => x"2a708106",
          6362 => x"51547380",
          6363 => x"2e863877",
          6364 => x"80c00758",
          6365 => x"7ab01108",
          6366 => x"a01b0c63",
          6367 => x"a41b0c63",
          6368 => x"53705257",
          6369 => x"e6d93f81",
          6370 => x"f8c80881",
          6371 => x"f8c80888",
          6372 => x"1b0c639c",
          6373 => x"05525ad2",
          6374 => x"d33f81f8",
          6375 => x"c80881f8",
          6376 => x"c8088c1b",
          6377 => x"0c777a0c",
          6378 => x"56861722",
          6379 => x"841a2377",
          6380 => x"901a3480",
          6381 => x"0b911a34",
          6382 => x"800b9c1a",
          6383 => x"0c800b94",
          6384 => x"1a0c7785",
          6385 => x"2a708106",
          6386 => x"51547380",
          6387 => x"2e818d38",
          6388 => x"81f8c808",
          6389 => x"802e8184",
          6390 => x"3881f8c8",
          6391 => x"08941a0c",
          6392 => x"8a172270",
          6393 => x"892b7b52",
          6394 => x"5957a839",
          6395 => x"76527851",
          6396 => x"d79f3f81",
          6397 => x"f8c80857",
          6398 => x"81f8c808",
          6399 => x"81268338",
          6400 => x"825581f8",
          6401 => x"c808ff2e",
          6402 => x"09810683",
          6403 => x"38795575",
          6404 => x"78315674",
          6405 => x"30707607",
          6406 => x"80255154",
          6407 => x"7776278a",
          6408 => x"38817075",
          6409 => x"06555a73",
          6410 => x"c3387698",
          6411 => x"1a0c74a9",
          6412 => x"387583ff",
          6413 => x"06547380",
          6414 => x"2ea23876",
          6415 => x"527a51d6",
          6416 => x"a63f81f8",
          6417 => x"c8088538",
          6418 => x"82558e39",
          6419 => x"75892a81",
          6420 => x"f8c80805",
          6421 => x"9c1a0c84",
          6422 => x"3980790c",
          6423 => x"74547381",
          6424 => x"f8c80c97",
          6425 => x"3d0d04f2",
          6426 => x"3d0d6063",
          6427 => x"65644040",
          6428 => x"5d59807e",
          6429 => x"0c903dfc",
          6430 => x"05527851",
          6431 => x"f9cf3f81",
          6432 => x"f8c80855",
          6433 => x"81f8c808",
          6434 => x"8a389119",
          6435 => x"33557480",
          6436 => x"2e863874",
          6437 => x"5682c439",
          6438 => x"90193381",
          6439 => x"06558756",
          6440 => x"74802e82",
          6441 => x"b6389539",
          6442 => x"820b911a",
          6443 => x"34825682",
          6444 => x"aa39810b",
          6445 => x"911a3481",
          6446 => x"5682a039",
          6447 => x"8c190894",
          6448 => x"1a083155",
          6449 => x"747c2783",
          6450 => x"38745c7b",
          6451 => x"802e8289",
          6452 => x"38941908",
          6453 => x"7083ff06",
          6454 => x"56567481",
          6455 => x"b2387e8a",
          6456 => x"1122ff05",
          6457 => x"77892a06",
          6458 => x"5b5579a8",
          6459 => x"38758738",
          6460 => x"88190855",
          6461 => x"8f399819",
          6462 => x"08527851",
          6463 => x"d5933f81",
          6464 => x"f8c80855",
          6465 => x"817527ff",
          6466 => x"9f3874ff",
          6467 => x"2effa338",
          6468 => x"74981a0c",
          6469 => x"98190852",
          6470 => x"7e51d4cb",
          6471 => x"3f81f8c8",
          6472 => x"08802eff",
          6473 => x"833881f8",
          6474 => x"c8081a7c",
          6475 => x"892a5957",
          6476 => x"77802e80",
          6477 => x"d638771a",
          6478 => x"7f8a1122",
          6479 => x"585c5575",
          6480 => x"75278538",
          6481 => x"757a3158",
          6482 => x"77547653",
          6483 => x"7c52811b",
          6484 => x"3351ca88",
          6485 => x"3f81f8c8",
          6486 => x"08fed738",
          6487 => x"7e831133",
          6488 => x"56567480",
          6489 => x"2e9f38b0",
          6490 => x"16087731",
          6491 => x"55747827",
          6492 => x"94388480",
          6493 => x"53b41652",
          6494 => x"b0160877",
          6495 => x"31892b7d",
          6496 => x"0551cfe0",
          6497 => x"3f77892b",
          6498 => x"56b93976",
          6499 => x"9c1a0c94",
          6500 => x"190883ff",
          6501 => x"06848071",
          6502 => x"3157557b",
          6503 => x"76278338",
          6504 => x"7b569c19",
          6505 => x"08527e51",
          6506 => x"d1c73f81",
          6507 => x"f8c808fe",
          6508 => x"81387553",
          6509 => x"94190883",
          6510 => x"ff061fb4",
          6511 => x"05527c51",
          6512 => x"cfa23f7b",
          6513 => x"76317e08",
          6514 => x"177f0c76",
          6515 => x"1e941b08",
          6516 => x"18941c0c",
          6517 => x"5e5cfdf3",
          6518 => x"39805675",
          6519 => x"81f8c80c",
          6520 => x"903d0d04",
          6521 => x"f23d0d60",
          6522 => x"63656440",
          6523 => x"405d5880",
          6524 => x"7e0c903d",
          6525 => x"fc055277",
          6526 => x"51f6d23f",
          6527 => x"81f8c808",
          6528 => x"5581f8c8",
          6529 => x"088a3891",
          6530 => x"18335574",
          6531 => x"802e8638",
          6532 => x"745683b8",
          6533 => x"39901833",
          6534 => x"70812a70",
          6535 => x"81065156",
          6536 => x"56875674",
          6537 => x"802e83a4",
          6538 => x"38953982",
          6539 => x"0b911934",
          6540 => x"82568398",
          6541 => x"39810b91",
          6542 => x"19348156",
          6543 => x"838e3994",
          6544 => x"18087c11",
          6545 => x"56567476",
          6546 => x"27843875",
          6547 => x"095c7b80",
          6548 => x"2e82ec38",
          6549 => x"94180870",
          6550 => x"83ff0656",
          6551 => x"567481fd",
          6552 => x"387e8a11",
          6553 => x"22ff0577",
          6554 => x"892a065c",
          6555 => x"557abf38",
          6556 => x"758c3888",
          6557 => x"18085574",
          6558 => x"9c387a52",
          6559 => x"85399818",
          6560 => x"08527751",
          6561 => x"d7e73f81",
          6562 => x"f8c80855",
          6563 => x"81f8c808",
          6564 => x"802e82ab",
          6565 => x"3874812e",
          6566 => x"ff913874",
          6567 => x"ff2eff95",
          6568 => x"38749819",
          6569 => x"0c881808",
          6570 => x"85387488",
          6571 => x"190c7e55",
          6572 => x"b015089c",
          6573 => x"19082e09",
          6574 => x"81068d38",
          6575 => x"7451cec1",
          6576 => x"3f81f8c8",
          6577 => x"08feee38",
          6578 => x"98180852",
          6579 => x"7e51d197",
          6580 => x"3f81f8c8",
          6581 => x"08802efe",
          6582 => x"d23881f8",
          6583 => x"c8081b7c",
          6584 => x"892a5a57",
          6585 => x"78802e80",
          6586 => x"d538781b",
          6587 => x"7f8a1122",
          6588 => x"585b5575",
          6589 => x"75278538",
          6590 => x"757b3159",
          6591 => x"78547653",
          6592 => x"7c52811a",
          6593 => x"3351c8be",
          6594 => x"3f81f8c8",
          6595 => x"08fea638",
          6596 => x"7eb01108",
          6597 => x"78315656",
          6598 => x"7479279b",
          6599 => x"38848053",
          6600 => x"b0160877",
          6601 => x"31892b7d",
          6602 => x"0552b416",
          6603 => x"51ccb53f",
          6604 => x"7e55800b",
          6605 => x"83163478",
          6606 => x"892b5680",
          6607 => x"db398c18",
          6608 => x"08941908",
          6609 => x"2693387e",
          6610 => x"51cdb63f",
          6611 => x"81f8c808",
          6612 => x"fde3387e",
          6613 => x"77b0120c",
          6614 => x"55769c19",
          6615 => x"0c941808",
          6616 => x"83ff0684",
          6617 => x"80713157",
          6618 => x"557b7627",
          6619 => x"83387b56",
          6620 => x"9c180852",
          6621 => x"7e51cdf9",
          6622 => x"3f81f8c8",
          6623 => x"08fdb638",
          6624 => x"75537c52",
          6625 => x"94180883",
          6626 => x"ff061fb4",
          6627 => x"0551cbd4",
          6628 => x"3f7e5581",
          6629 => x"0b831634",
          6630 => x"7b76317e",
          6631 => x"08177f0c",
          6632 => x"761e941a",
          6633 => x"08187094",
          6634 => x"1c0c8c1b",
          6635 => x"0858585e",
          6636 => x"5c747627",
          6637 => x"83387555",
          6638 => x"748c190c",
          6639 => x"fd903990",
          6640 => x"183380c0",
          6641 => x"07557490",
          6642 => x"19348056",
          6643 => x"7581f8c8",
          6644 => x"0c903d0d",
          6645 => x"04f83d0d",
          6646 => x"7a8b3dfc",
          6647 => x"05537052",
          6648 => x"56f2ea3f",
          6649 => x"81f8c808",
          6650 => x"5781f8c8",
          6651 => x"0880fb38",
          6652 => x"90163370",
          6653 => x"862a7081",
          6654 => x"06515555",
          6655 => x"73802e80",
          6656 => x"e938a016",
          6657 => x"08527851",
          6658 => x"cce73f81",
          6659 => x"f8c80857",
          6660 => x"81f8c808",
          6661 => x"80d438a4",
          6662 => x"16088b11",
          6663 => x"33a00755",
          6664 => x"55738b16",
          6665 => x"34881608",
          6666 => x"53745275",
          6667 => x"0851dde8",
          6668 => x"3f8c1608",
          6669 => x"529c1551",
          6670 => x"c9fb3f82",
          6671 => x"88b20a52",
          6672 => x"961551c9",
          6673 => x"f03f7652",
          6674 => x"921551c9",
          6675 => x"ca3f7854",
          6676 => x"810b8315",
          6677 => x"347851cc",
          6678 => x"df3f81f8",
          6679 => x"c8089017",
          6680 => x"3381bf06",
          6681 => x"55577390",
          6682 => x"17347681",
          6683 => x"f8c80c8a",
          6684 => x"3d0d04fc",
          6685 => x"3d0d7670",
          6686 => x"5254fed9",
          6687 => x"3f81f8c8",
          6688 => x"085381f8",
          6689 => x"c8089c38",
          6690 => x"863dfc05",
          6691 => x"527351f1",
          6692 => x"bc3f81f8",
          6693 => x"c8085381",
          6694 => x"f8c80887",
          6695 => x"3881f8c8",
          6696 => x"08740c72",
          6697 => x"81f8c80c",
          6698 => x"863d0d04",
          6699 => x"ff3d0d84",
          6700 => x"3d51e6e4",
          6701 => x"3f8b5280",
          6702 => x"0b81f8c8",
          6703 => x"08248b38",
          6704 => x"81f8c808",
          6705 => x"81f98c34",
          6706 => x"80527181",
          6707 => x"f8c80c83",
          6708 => x"3d0d04ef",
          6709 => x"3d0d8053",
          6710 => x"933dd005",
          6711 => x"52943d51",
          6712 => x"e9c13f81",
          6713 => x"f8c80855",
          6714 => x"81f8c808",
          6715 => x"80e03876",
          6716 => x"58635293",
          6717 => x"3dd40551",
          6718 => x"e08d3f81",
          6719 => x"f8c80855",
          6720 => x"81f8c808",
          6721 => x"bc380280",
          6722 => x"c7053370",
          6723 => x"982b5556",
          6724 => x"73802589",
          6725 => x"38767a94",
          6726 => x"120c54b2",
          6727 => x"3902a205",
          6728 => x"3370842a",
          6729 => x"70810651",
          6730 => x"55567380",
          6731 => x"2e9e3876",
          6732 => x"7f537052",
          6733 => x"54dba83f",
          6734 => x"81f8c808",
          6735 => x"94150c8e",
          6736 => x"3981f8c8",
          6737 => x"08842e09",
          6738 => x"81068338",
          6739 => x"85557481",
          6740 => x"f8c80c93",
          6741 => x"3d0d04e4",
          6742 => x"3d0d6f6f",
          6743 => x"5b5b807a",
          6744 => x"3480539e",
          6745 => x"3dffb805",
          6746 => x"529f3d51",
          6747 => x"e8b53f81",
          6748 => x"f8c80857",
          6749 => x"81f8c808",
          6750 => x"82fc387b",
          6751 => x"437a7c94",
          6752 => x"11084755",
          6753 => x"58645473",
          6754 => x"802e81ed",
          6755 => x"38a05293",
          6756 => x"3d705255",
          6757 => x"d5ea3f81",
          6758 => x"f8c80857",
          6759 => x"81f8c808",
          6760 => x"82d43868",
          6761 => x"527b51c9",
          6762 => x"c83f81f8",
          6763 => x"c8085781",
          6764 => x"f8c80882",
          6765 => x"c1386952",
          6766 => x"7b51daa3",
          6767 => x"3f81f8c8",
          6768 => x"08457652",
          6769 => x"7451d5b8",
          6770 => x"3f81f8c8",
          6771 => x"085781f8",
          6772 => x"c80882a2",
          6773 => x"38805274",
          6774 => x"51daeb3f",
          6775 => x"81f8c808",
          6776 => x"5781f8c8",
          6777 => x"08a43869",
          6778 => x"527b51d9",
          6779 => x"f23f7381",
          6780 => x"f8c8082e",
          6781 => x"a6387652",
          6782 => x"7451d6cf",
          6783 => x"3f81f8c8",
          6784 => x"085781f8",
          6785 => x"c808802e",
          6786 => x"cc387684",
          6787 => x"2e098106",
          6788 => x"86388257",
          6789 => x"81e03976",
          6790 => x"81dc389e",
          6791 => x"3dffbc05",
          6792 => x"527451dc",
          6793 => x"c93f7690",
          6794 => x"3d781181",
          6795 => x"11335156",
          6796 => x"5a567380",
          6797 => x"2e913802",
          6798 => x"b9055581",
          6799 => x"16811670",
          6800 => x"33565656",
          6801 => x"73f53881",
          6802 => x"16547378",
          6803 => x"26819038",
          6804 => x"75802e99",
          6805 => x"38781681",
          6806 => x"0555ff18",
          6807 => x"6f11ff18",
          6808 => x"ff185858",
          6809 => x"55587433",
          6810 => x"743475ee",
          6811 => x"38ff186f",
          6812 => x"115558af",
          6813 => x"7434fe8d",
          6814 => x"39777b2e",
          6815 => x"0981068a",
          6816 => x"38ff186f",
          6817 => x"115558af",
          6818 => x"7434800b",
          6819 => x"81f98c33",
          6820 => x"70842981",
          6821 => x"e6c80570",
          6822 => x"08703352",
          6823 => x"5c565656",
          6824 => x"73762e8d",
          6825 => x"38811670",
          6826 => x"1a703351",
          6827 => x"555673f5",
          6828 => x"38821654",
          6829 => x"737826a7",
          6830 => x"38805574",
          6831 => x"76279138",
          6832 => x"74195473",
          6833 => x"337a7081",
          6834 => x"055c3481",
          6835 => x"1555ec39",
          6836 => x"ba7a7081",
          6837 => x"055c3474",
          6838 => x"ff2e0981",
          6839 => x"06853891",
          6840 => x"5794396e",
          6841 => x"18811959",
          6842 => x"5473337a",
          6843 => x"7081055c",
          6844 => x"347a7826",
          6845 => x"ee38807a",
          6846 => x"347681f8",
          6847 => x"c80c9e3d",
          6848 => x"0d04f73d",
          6849 => x"0d7b7d8d",
          6850 => x"3dfc0554",
          6851 => x"71535755",
          6852 => x"ecbb3f81",
          6853 => x"f8c80853",
          6854 => x"81f8c808",
          6855 => x"82fa3891",
          6856 => x"15335372",
          6857 => x"82f2388c",
          6858 => x"15085473",
          6859 => x"76279238",
          6860 => x"90153370",
          6861 => x"812a7081",
          6862 => x"06515457",
          6863 => x"72833873",
          6864 => x"56941508",
          6865 => x"54807094",
          6866 => x"170c5875",
          6867 => x"782e8297",
          6868 => x"38798a11",
          6869 => x"2270892b",
          6870 => x"59515373",
          6871 => x"782eb738",
          6872 => x"7652ff16",
          6873 => x"51fefcc3",
          6874 => x"3f81f8c8",
          6875 => x"08ff1578",
          6876 => x"54705355",
          6877 => x"53fefcb3",
          6878 => x"3f81f8c8",
          6879 => x"08732696",
          6880 => x"38763070",
          6881 => x"75067094",
          6882 => x"180c7771",
          6883 => x"31981808",
          6884 => x"57585153",
          6885 => x"b1398815",
          6886 => x"085473a6",
          6887 => x"38735274",
          6888 => x"51cdca3f",
          6889 => x"81f8c808",
          6890 => x"5481f8c8",
          6891 => x"08812e81",
          6892 => x"9a3881f8",
          6893 => x"c808ff2e",
          6894 => x"819b3881",
          6895 => x"f8c80888",
          6896 => x"160c7398",
          6897 => x"160c7380",
          6898 => x"2e819c38",
          6899 => x"76762780",
          6900 => x"dc387577",
          6901 => x"31941608",
          6902 => x"1894170c",
          6903 => x"90163370",
          6904 => x"812a7081",
          6905 => x"0651555a",
          6906 => x"5672802e",
          6907 => x"9a387352",
          6908 => x"7451ccf9",
          6909 => x"3f81f8c8",
          6910 => x"085481f8",
          6911 => x"c8089438",
          6912 => x"81f8c808",
          6913 => x"56a73973",
          6914 => x"527451c7",
          6915 => x"843f81f8",
          6916 => x"c8085473",
          6917 => x"ff2ebe38",
          6918 => x"817427af",
          6919 => x"38795373",
          6920 => x"98140827",
          6921 => x"a6387398",
          6922 => x"160cffa0",
          6923 => x"39941508",
          6924 => x"1694160c",
          6925 => x"7583ff06",
          6926 => x"5372802e",
          6927 => x"aa387352",
          6928 => x"7951c6a3",
          6929 => x"3f81f8c8",
          6930 => x"08943882",
          6931 => x"0b911634",
          6932 => x"825380c4",
          6933 => x"39810b91",
          6934 => x"16348153",
          6935 => x"bb397589",
          6936 => x"2a81f8c8",
          6937 => x"08055894",
          6938 => x"1508548c",
          6939 => x"15087427",
          6940 => x"9038738c",
          6941 => x"160c9015",
          6942 => x"3380c007",
          6943 => x"53729016",
          6944 => x"347383ff",
          6945 => x"06537280",
          6946 => x"2e8c3877",
          6947 => x"9c16082e",
          6948 => x"8538779c",
          6949 => x"160c8053",
          6950 => x"7281f8c8",
          6951 => x"0c8b3d0d",
          6952 => x"04f93d0d",
          6953 => x"79568954",
          6954 => x"75802e81",
          6955 => x"8a388053",
          6956 => x"893dfc05",
          6957 => x"528a3d84",
          6958 => x"0551e1e7",
          6959 => x"3f81f8c8",
          6960 => x"085581f8",
          6961 => x"c80880ea",
          6962 => x"3877760c",
          6963 => x"7a527551",
          6964 => x"d8b53f81",
          6965 => x"f8c80855",
          6966 => x"81f8c808",
          6967 => x"80c338ab",
          6968 => x"16337098",
          6969 => x"2b555780",
          6970 => x"7424a238",
          6971 => x"86163370",
          6972 => x"842a7081",
          6973 => x"06515557",
          6974 => x"73802ead",
          6975 => x"389c1608",
          6976 => x"527751d3",
          6977 => x"da3f81f8",
          6978 => x"c8088817",
          6979 => x"0c775486",
          6980 => x"14228417",
          6981 => x"23745275",
          6982 => x"51cee53f",
          6983 => x"81f8c808",
          6984 => x"5574842e",
          6985 => x"09810685",
          6986 => x"38855586",
          6987 => x"3974802e",
          6988 => x"84388076",
          6989 => x"0c745473",
          6990 => x"81f8c80c",
          6991 => x"893d0d04",
          6992 => x"fc3d0d76",
          6993 => x"873dfc05",
          6994 => x"53705253",
          6995 => x"e7ff3f81",
          6996 => x"f8c80887",
          6997 => x"3881f8c8",
          6998 => x"08730c86",
          6999 => x"3d0d04fb",
          7000 => x"3d0d7779",
          7001 => x"893dfc05",
          7002 => x"54715356",
          7003 => x"54e7de3f",
          7004 => x"81f8c808",
          7005 => x"5381f8c8",
          7006 => x"0880df38",
          7007 => x"74933881",
          7008 => x"f8c80852",
          7009 => x"7351cdf8",
          7010 => x"3f81f8c8",
          7011 => x"085380ca",
          7012 => x"3981f8c8",
          7013 => x"08527351",
          7014 => x"d3ac3f81",
          7015 => x"f8c80853",
          7016 => x"81f8c808",
          7017 => x"842e0981",
          7018 => x"06853880",
          7019 => x"53873981",
          7020 => x"f8c808a6",
          7021 => x"38745273",
          7022 => x"51d5b33f",
          7023 => x"72527351",
          7024 => x"cf893f81",
          7025 => x"f8c80884",
          7026 => x"32703070",
          7027 => x"72079f2c",
          7028 => x"7081f8c8",
          7029 => x"08065151",
          7030 => x"54547281",
          7031 => x"f8c80c87",
          7032 => x"3d0d04ee",
          7033 => x"3d0d6557",
          7034 => x"8053893d",
          7035 => x"7053963d",
          7036 => x"5256dfaf",
          7037 => x"3f81f8c8",
          7038 => x"085581f8",
          7039 => x"c808b238",
          7040 => x"64527551",
          7041 => x"d6813f81",
          7042 => x"f8c80855",
          7043 => x"81f8c808",
          7044 => x"a0380280",
          7045 => x"cb053370",
          7046 => x"982b5558",
          7047 => x"73802585",
          7048 => x"3886558d",
          7049 => x"3976802e",
          7050 => x"88387652",
          7051 => x"7551d4be",
          7052 => x"3f7481f8",
          7053 => x"c80c943d",
          7054 => x"0d04f03d",
          7055 => x"0d636555",
          7056 => x"5c805392",
          7057 => x"3dec0552",
          7058 => x"933d51de",
          7059 => x"d63f81f8",
          7060 => x"c8085b81",
          7061 => x"f8c80882",
          7062 => x"80387c74",
          7063 => x"0c730898",
          7064 => x"1108fe11",
          7065 => x"90130859",
          7066 => x"56585575",
          7067 => x"74269138",
          7068 => x"757c0c81",
          7069 => x"e439815b",
          7070 => x"81cc3982",
          7071 => x"5b81c739",
          7072 => x"81f8c808",
          7073 => x"75335559",
          7074 => x"73812e09",
          7075 => x"8106bf38",
          7076 => x"82755f57",
          7077 => x"7652923d",
          7078 => x"f00551c1",
          7079 => x"f43f81f8",
          7080 => x"c808ff2e",
          7081 => x"d13881f8",
          7082 => x"c808812e",
          7083 => x"ce3881f8",
          7084 => x"c8083070",
          7085 => x"81f8c808",
          7086 => x"0780257a",
          7087 => x"0581197f",
          7088 => x"53595a54",
          7089 => x"98140877",
          7090 => x"26ca3880",
          7091 => x"f939a415",
          7092 => x"0881f8c8",
          7093 => x"08575875",
          7094 => x"98387752",
          7095 => x"81187d52",
          7096 => x"58ffbf8d",
          7097 => x"3f81f8c8",
          7098 => x"085b81f8",
          7099 => x"c80880d6",
          7100 => x"387c7033",
          7101 => x"7712ff1a",
          7102 => x"5d525654",
          7103 => x"74822e09",
          7104 => x"81069e38",
          7105 => x"b41451ff",
          7106 => x"bbcb3f81",
          7107 => x"f8c80883",
          7108 => x"ffff0670",
          7109 => x"30708025",
          7110 => x"1b821959",
          7111 => x"5b51549b",
          7112 => x"39b41451",
          7113 => x"ffbbc53f",
          7114 => x"81f8c808",
          7115 => x"f00a0670",
          7116 => x"30708025",
          7117 => x"1b841959",
          7118 => x"5b515475",
          7119 => x"83ff067a",
          7120 => x"585679ff",
          7121 => x"9238787c",
          7122 => x"0c7c7990",
          7123 => x"120c8411",
          7124 => x"33810756",
          7125 => x"54748415",
          7126 => x"347a81f8",
          7127 => x"c80c923d",
          7128 => x"0d04f93d",
          7129 => x"0d798a3d",
          7130 => x"fc055370",
          7131 => x"5257e3dd",
          7132 => x"3f81f8c8",
          7133 => x"085681f8",
          7134 => x"c80881a8",
          7135 => x"38911733",
          7136 => x"567581a0",
          7137 => x"38901733",
          7138 => x"70812a70",
          7139 => x"81065155",
          7140 => x"55875573",
          7141 => x"802e818e",
          7142 => x"38941708",
          7143 => x"54738c18",
          7144 => x"08278180",
          7145 => x"38739b38",
          7146 => x"81f8c808",
          7147 => x"53881708",
          7148 => x"527651c4",
          7149 => x"8c3f81f8",
          7150 => x"c8087488",
          7151 => x"190c5680",
          7152 => x"c9399817",
          7153 => x"08527651",
          7154 => x"ffbfc63f",
          7155 => x"81f8c808",
          7156 => x"ff2e0981",
          7157 => x"06833881",
          7158 => x"5681f8c8",
          7159 => x"08812e09",
          7160 => x"81068538",
          7161 => x"8256a339",
          7162 => x"75a03877",
          7163 => x"5481f8c8",
          7164 => x"08981508",
          7165 => x"27943898",
          7166 => x"17085381",
          7167 => x"f8c80852",
          7168 => x"7651c3bd",
          7169 => x"3f81f8c8",
          7170 => x"08569417",
          7171 => x"088c180c",
          7172 => x"90173380",
          7173 => x"c0075473",
          7174 => x"90183475",
          7175 => x"802e8538",
          7176 => x"75911834",
          7177 => x"75557481",
          7178 => x"f8c80c89",
          7179 => x"3d0d04e2",
          7180 => x"3d0d8253",
          7181 => x"a03dffa4",
          7182 => x"0552a13d",
          7183 => x"51dae43f",
          7184 => x"81f8c808",
          7185 => x"5581f8c8",
          7186 => x"0881f538",
          7187 => x"7845a13d",
          7188 => x"0852953d",
          7189 => x"705258d1",
          7190 => x"ae3f81f8",
          7191 => x"c8085581",
          7192 => x"f8c80881",
          7193 => x"db380280",
          7194 => x"fb053370",
          7195 => x"852a7081",
          7196 => x"06515556",
          7197 => x"86557381",
          7198 => x"c7387598",
          7199 => x"2b548074",
          7200 => x"2481bd38",
          7201 => x"0280d605",
          7202 => x"33708106",
          7203 => x"58548755",
          7204 => x"7681ad38",
          7205 => x"6b527851",
          7206 => x"ccc53f81",
          7207 => x"f8c80874",
          7208 => x"842a7081",
          7209 => x"06515556",
          7210 => x"73802e80",
          7211 => x"d4387854",
          7212 => x"81f8c808",
          7213 => x"9415082e",
          7214 => x"81863873",
          7215 => x"5a81f8c8",
          7216 => x"085c7652",
          7217 => x"8a3d7052",
          7218 => x"54c7b53f",
          7219 => x"81f8c808",
          7220 => x"5581f8c8",
          7221 => x"0880e938",
          7222 => x"81f8c808",
          7223 => x"527351cc",
          7224 => x"e53f81f8",
          7225 => x"c8085581",
          7226 => x"f8c80886",
          7227 => x"38875580",
          7228 => x"cf3981f8",
          7229 => x"c808842e",
          7230 => x"883881f8",
          7231 => x"c80880c0",
          7232 => x"387751ce",
          7233 => x"c23f81f8",
          7234 => x"c80881f8",
          7235 => x"c8083070",
          7236 => x"81f8c808",
          7237 => x"07802551",
          7238 => x"55557580",
          7239 => x"2e943873",
          7240 => x"802e8f38",
          7241 => x"80537552",
          7242 => x"7751c195",
          7243 => x"3f81f8c8",
          7244 => x"0855748c",
          7245 => x"387851ff",
          7246 => x"bafe3f81",
          7247 => x"f8c80855",
          7248 => x"7481f8c8",
          7249 => x"0ca03d0d",
          7250 => x"04e93d0d",
          7251 => x"8253993d",
          7252 => x"c005529a",
          7253 => x"3d51d8cb",
          7254 => x"3f81f8c8",
          7255 => x"085481f8",
          7256 => x"c80882b0",
          7257 => x"38785e69",
          7258 => x"528e3d70",
          7259 => x"5258cf97",
          7260 => x"3f81f8c8",
          7261 => x"085481f8",
          7262 => x"c8088638",
          7263 => x"88548294",
          7264 => x"3981f8c8",
          7265 => x"08842e09",
          7266 => x"81068288",
          7267 => x"380280df",
          7268 => x"05337085",
          7269 => x"2a810651",
          7270 => x"55865474",
          7271 => x"81f63878",
          7272 => x"5a74528a",
          7273 => x"3d705257",
          7274 => x"c1c33f81",
          7275 => x"f8c80875",
          7276 => x"555681f8",
          7277 => x"c8088338",
          7278 => x"875481f8",
          7279 => x"c808812e",
          7280 => x"09810683",
          7281 => x"38825481",
          7282 => x"f8c808ff",
          7283 => x"2e098106",
          7284 => x"86388154",
          7285 => x"81b43973",
          7286 => x"81b03881",
          7287 => x"f8c80852",
          7288 => x"7851c4a4",
          7289 => x"3f81f8c8",
          7290 => x"085481f8",
          7291 => x"c808819a",
          7292 => x"388b53a0",
          7293 => x"52b41951",
          7294 => x"ffb78c3f",
          7295 => x"7854ae0b",
          7296 => x"b4153478",
          7297 => x"54900bbf",
          7298 => x"15348288",
          7299 => x"b20a5280",
          7300 => x"ca1951ff",
          7301 => x"b69f3f75",
          7302 => x"5378b411",
          7303 => x"5351c9f8",
          7304 => x"3fa05378",
          7305 => x"b4115380",
          7306 => x"d40551ff",
          7307 => x"b6b63f78",
          7308 => x"54ae0b80",
          7309 => x"d515347f",
          7310 => x"537880d4",
          7311 => x"115351c9",
          7312 => x"d73f7854",
          7313 => x"810b8315",
          7314 => x"347751cb",
          7315 => x"a43f81f8",
          7316 => x"c8085481",
          7317 => x"f8c808b2",
          7318 => x"388288b2",
          7319 => x"0a526496",
          7320 => x"0551ffb5",
          7321 => x"d03f7553",
          7322 => x"64527851",
          7323 => x"c9aa3f64",
          7324 => x"54900b8b",
          7325 => x"15347854",
          7326 => x"810b8315",
          7327 => x"347851ff",
          7328 => x"b8b63f81",
          7329 => x"f8c80854",
          7330 => x"8b398053",
          7331 => x"75527651",
          7332 => x"ffbeae3f",
          7333 => x"7381f8c8",
          7334 => x"0c993d0d",
          7335 => x"04da3d0d",
          7336 => x"a93d8405",
          7337 => x"51d2f13f",
          7338 => x"8253a83d",
          7339 => x"ff840552",
          7340 => x"a93d51d5",
          7341 => x"ee3f81f8",
          7342 => x"c8085581",
          7343 => x"f8c80882",
          7344 => x"d338784d",
          7345 => x"a93d0852",
          7346 => x"9d3d7052",
          7347 => x"58ccb83f",
          7348 => x"81f8c808",
          7349 => x"5581f8c8",
          7350 => x"0882b938",
          7351 => x"02819b05",
          7352 => x"3381a006",
          7353 => x"54865573",
          7354 => x"82aa38a0",
          7355 => x"53a43d08",
          7356 => x"52a83dff",
          7357 => x"880551ff",
          7358 => x"b4ea3fac",
          7359 => x"53775292",
          7360 => x"3d705254",
          7361 => x"ffb4dd3f",
          7362 => x"aa3d0852",
          7363 => x"7351cbf7",
          7364 => x"3f81f8c8",
          7365 => x"085581f8",
          7366 => x"c8089538",
          7367 => x"636f2e09",
          7368 => x"81068838",
          7369 => x"65a23d08",
          7370 => x"2e923888",
          7371 => x"5581e539",
          7372 => x"81f8c808",
          7373 => x"842e0981",
          7374 => x"0681b838",
          7375 => x"7351c9b1",
          7376 => x"3f81f8c8",
          7377 => x"085581f8",
          7378 => x"c80881c8",
          7379 => x"38685693",
          7380 => x"53a83dff",
          7381 => x"9505528d",
          7382 => x"1651ffb4",
          7383 => x"873f02af",
          7384 => x"05338b17",
          7385 => x"348b1633",
          7386 => x"70842a70",
          7387 => x"81065155",
          7388 => x"55738938",
          7389 => x"74a00754",
          7390 => x"738b1734",
          7391 => x"7854810b",
          7392 => x"8315348b",
          7393 => x"16337084",
          7394 => x"2a708106",
          7395 => x"51555573",
          7396 => x"802e80e5",
          7397 => x"386e642e",
          7398 => x"80df3875",
          7399 => x"527851c6",
          7400 => x"be3f81f8",
          7401 => x"c8085278",
          7402 => x"51ffb7bb",
          7403 => x"3f825581",
          7404 => x"f8c80880",
          7405 => x"2e80dd38",
          7406 => x"81f8c808",
          7407 => x"527851ff",
          7408 => x"b5af3f81",
          7409 => x"f8c80879",
          7410 => x"80d41158",
          7411 => x"585581f8",
          7412 => x"c80880c0",
          7413 => x"38811633",
          7414 => x"5473ae2e",
          7415 => x"09810699",
          7416 => x"38635375",
          7417 => x"527651c6",
          7418 => x"af3f7854",
          7419 => x"810b8315",
          7420 => x"34873981",
          7421 => x"f8c8089c",
          7422 => x"387751c8",
          7423 => x"ca3f81f8",
          7424 => x"c8085581",
          7425 => x"f8c8088c",
          7426 => x"387851ff",
          7427 => x"b5aa3f81",
          7428 => x"f8c80855",
          7429 => x"7481f8c8",
          7430 => x"0ca83d0d",
          7431 => x"04ed3d0d",
          7432 => x"0280db05",
          7433 => x"33028405",
          7434 => x"80df0533",
          7435 => x"57578253",
          7436 => x"953dd005",
          7437 => x"52963d51",
          7438 => x"d2e93f81",
          7439 => x"f8c80855",
          7440 => x"81f8c808",
          7441 => x"80cf3878",
          7442 => x"5a655295",
          7443 => x"3dd40551",
          7444 => x"c9b53f81",
          7445 => x"f8c80855",
          7446 => x"81f8c808",
          7447 => x"b8380280",
          7448 => x"cf053381",
          7449 => x"a0065486",
          7450 => x"5573aa38",
          7451 => x"75a70661",
          7452 => x"71098b12",
          7453 => x"3371067a",
          7454 => x"74060751",
          7455 => x"57555674",
          7456 => x"8b153478",
          7457 => x"54810b83",
          7458 => x"15347851",
          7459 => x"ffb4a93f",
          7460 => x"81f8c808",
          7461 => x"557481f8",
          7462 => x"c80c953d",
          7463 => x"0d04ef3d",
          7464 => x"0d645682",
          7465 => x"53933dd0",
          7466 => x"0552943d",
          7467 => x"51d1f43f",
          7468 => x"81f8c808",
          7469 => x"5581f8c8",
          7470 => x"0880cb38",
          7471 => x"76586352",
          7472 => x"933dd405",
          7473 => x"51c8c03f",
          7474 => x"81f8c808",
          7475 => x"5581f8c8",
          7476 => x"08b43802",
          7477 => x"80c70533",
          7478 => x"81a00654",
          7479 => x"865573a6",
          7480 => x"38841622",
          7481 => x"86172271",
          7482 => x"902b0753",
          7483 => x"54961f51",
          7484 => x"ffb0c23f",
          7485 => x"7654810b",
          7486 => x"83153476",
          7487 => x"51ffb3b8",
          7488 => x"3f81f8c8",
          7489 => x"08557481",
          7490 => x"f8c80c93",
          7491 => x"3d0d04ea",
          7492 => x"3d0d696b",
          7493 => x"5c5a8053",
          7494 => x"983dd005",
          7495 => x"52993d51",
          7496 => x"d1813f81",
          7497 => x"f8c80881",
          7498 => x"f8c80830",
          7499 => x"7081f8c8",
          7500 => x"08078025",
          7501 => x"51555779",
          7502 => x"802e8185",
          7503 => x"38817075",
          7504 => x"06555573",
          7505 => x"802e80f9",
          7506 => x"387b5d80",
          7507 => x"5f80528d",
          7508 => x"3d705254",
          7509 => x"ffbea93f",
          7510 => x"81f8c808",
          7511 => x"5781f8c8",
          7512 => x"0880d138",
          7513 => x"74527351",
          7514 => x"c3dc3f81",
          7515 => x"f8c80857",
          7516 => x"81f8c808",
          7517 => x"bf3881f8",
          7518 => x"c80881f8",
          7519 => x"c808655b",
          7520 => x"59567818",
          7521 => x"81197b18",
          7522 => x"56595574",
          7523 => x"33743481",
          7524 => x"16568a78",
          7525 => x"27ec388b",
          7526 => x"56751a54",
          7527 => x"80743475",
          7528 => x"802e9e38",
          7529 => x"ff16701b",
          7530 => x"70335155",
          7531 => x"5673a02e",
          7532 => x"e8388e39",
          7533 => x"76842e09",
          7534 => x"81068638",
          7535 => x"807a3480",
          7536 => x"57763070",
          7537 => x"78078025",
          7538 => x"51547a80",
          7539 => x"2e80c138",
          7540 => x"73802ebc",
          7541 => x"387ba011",
          7542 => x"085351ff",
          7543 => x"b1933f81",
          7544 => x"f8c80857",
          7545 => x"81f8c808",
          7546 => x"a7387b70",
          7547 => x"33555580",
          7548 => x"c3567383",
          7549 => x"2e8b3880",
          7550 => x"e4567384",
          7551 => x"2e8338a7",
          7552 => x"567515b4",
          7553 => x"0551ffad",
          7554 => x"e33f81f8",
          7555 => x"c8087b0c",
          7556 => x"7681f8c8",
          7557 => x"0c983d0d",
          7558 => x"04e63d0d",
          7559 => x"82539c3d",
          7560 => x"ffb80552",
          7561 => x"9d3d51ce",
          7562 => x"fa3f81f8",
          7563 => x"c80881f8",
          7564 => x"c8085654",
          7565 => x"81f8c808",
          7566 => x"8398388b",
          7567 => x"53a0528b",
          7568 => x"3d705259",
          7569 => x"ffaec03f",
          7570 => x"736d7033",
          7571 => x"7081ff06",
          7572 => x"52575557",
          7573 => x"9f742781",
          7574 => x"bc387858",
          7575 => x"7481ff06",
          7576 => x"6d81054e",
          7577 => x"705255ff",
          7578 => x"af893f81",
          7579 => x"f8c80880",
          7580 => x"2ea5386c",
          7581 => x"70337053",
          7582 => x"5754ffae",
          7583 => x"fd3f81f8",
          7584 => x"c808802e",
          7585 => x"8d387488",
          7586 => x"2b76076d",
          7587 => x"81054e55",
          7588 => x"863981f8",
          7589 => x"c80855ff",
          7590 => x"9f157083",
          7591 => x"ffff0651",
          7592 => x"54739926",
          7593 => x"8a38e015",
          7594 => x"7083ffff",
          7595 => x"06565480",
          7596 => x"ff752787",
          7597 => x"3881e5d8",
          7598 => x"15335574",
          7599 => x"802ea338",
          7600 => x"745281e7",
          7601 => x"d851ffae",
          7602 => x"893f81f8",
          7603 => x"c8089338",
          7604 => x"81ff7527",
          7605 => x"88387689",
          7606 => x"2688388b",
          7607 => x"398a7727",
          7608 => x"86388655",
          7609 => x"81ec3981",
          7610 => x"ff75278f",
          7611 => x"3874882a",
          7612 => x"54737870",
          7613 => x"81055a34",
          7614 => x"81175774",
          7615 => x"78708105",
          7616 => x"5a348117",
          7617 => x"6d703370",
          7618 => x"81ff0652",
          7619 => x"57555773",
          7620 => x"9f26fec8",
          7621 => x"388b3d33",
          7622 => x"54865573",
          7623 => x"81e52e81",
          7624 => x"b1387680",
          7625 => x"2e993802",
          7626 => x"a7055576",
          7627 => x"15703351",
          7628 => x"5473a02e",
          7629 => x"09810687",
          7630 => x"38ff1757",
          7631 => x"76ed3879",
          7632 => x"41804380",
          7633 => x"52913d70",
          7634 => x"5255ffba",
          7635 => x"b33f81f8",
          7636 => x"c8085481",
          7637 => x"f8c80880",
          7638 => x"f7388152",
          7639 => x"7451ffbf",
          7640 => x"e53f81f8",
          7641 => x"c8085481",
          7642 => x"f8c8088d",
          7643 => x"387680c4",
          7644 => x"386754e5",
          7645 => x"743480c6",
          7646 => x"3981f8c8",
          7647 => x"08842e09",
          7648 => x"810680cc",
          7649 => x"38805476",
          7650 => x"742e80c4",
          7651 => x"38815274",
          7652 => x"51ffbdb0",
          7653 => x"3f81f8c8",
          7654 => x"085481f8",
          7655 => x"c808b138",
          7656 => x"a05381f8",
          7657 => x"c8085267",
          7658 => x"51ffabdb",
          7659 => x"3f675488",
          7660 => x"0b8b1534",
          7661 => x"8b537852",
          7662 => x"6751ffab",
          7663 => x"a73f7954",
          7664 => x"810b8315",
          7665 => x"347951ff",
          7666 => x"adee3f81",
          7667 => x"f8c80854",
          7668 => x"73557481",
          7669 => x"f8c80c9c",
          7670 => x"3d0d04f2",
          7671 => x"3d0d6062",
          7672 => x"02880580",
          7673 => x"cb053393",
          7674 => x"3dfc0555",
          7675 => x"7254405e",
          7676 => x"5ad2da3f",
          7677 => x"81f8c808",
          7678 => x"5881f8c8",
          7679 => x"0882bd38",
          7680 => x"911a3358",
          7681 => x"7782b538",
          7682 => x"7c802e97",
          7683 => x"388c1a08",
          7684 => x"59789038",
          7685 => x"901a3370",
          7686 => x"812a7081",
          7687 => x"06515555",
          7688 => x"73903887",
          7689 => x"54829739",
          7690 => x"82588290",
          7691 => x"39815882",
          7692 => x"8b397e8a",
          7693 => x"11227089",
          7694 => x"2b70557f",
          7695 => x"54565656",
          7696 => x"fee2e83f",
          7697 => x"ff147d06",
          7698 => x"70307072",
          7699 => x"079f2a81",
          7700 => x"f8c80805",
          7701 => x"8c19087c",
          7702 => x"405a5d55",
          7703 => x"55817727",
          7704 => x"88389816",
          7705 => x"08772683",
          7706 => x"38825776",
          7707 => x"77565980",
          7708 => x"56745279",
          7709 => x"51ffae99",
          7710 => x"3f81157f",
          7711 => x"55559814",
          7712 => x"08752683",
          7713 => x"38825581",
          7714 => x"f8c80881",
          7715 => x"2eff9938",
          7716 => x"81f8c808",
          7717 => x"ff2eff95",
          7718 => x"3881f8c8",
          7719 => x"088e3881",
          7720 => x"1656757b",
          7721 => x"2e098106",
          7722 => x"87389339",
          7723 => x"74598056",
          7724 => x"74772e09",
          7725 => x"8106ffb9",
          7726 => x"38875880",
          7727 => x"ff397d80",
          7728 => x"2eba3878",
          7729 => x"7b55557a",
          7730 => x"802eb438",
          7731 => x"81155673",
          7732 => x"812e0981",
          7733 => x"068338ff",
          7734 => x"56755374",
          7735 => x"527e51ff",
          7736 => x"afa83f81",
          7737 => x"f8c80858",
          7738 => x"81f8c808",
          7739 => x"80ce3874",
          7740 => x"8116ff16",
          7741 => x"56565c73",
          7742 => x"d3388439",
          7743 => x"ff195c7e",
          7744 => x"7c8c120c",
          7745 => x"557d802e",
          7746 => x"b3387888",
          7747 => x"1b0c7c8c",
          7748 => x"1b0c901a",
          7749 => x"3380c007",
          7750 => x"5473901b",
          7751 => x"34981508",
          7752 => x"fe059016",
          7753 => x"08575475",
          7754 => x"74269138",
          7755 => x"757b3190",
          7756 => x"160c8415",
          7757 => x"33810754",
          7758 => x"73841634",
          7759 => x"77547381",
          7760 => x"f8c80c90",
          7761 => x"3d0d04e9",
          7762 => x"3d0d6b6d",
          7763 => x"02880580",
          7764 => x"eb05339d",
          7765 => x"3d545a5c",
          7766 => x"59c5bd3f",
          7767 => x"8b56800b",
          7768 => x"81f8c808",
          7769 => x"248bf838",
          7770 => x"81f8c808",
          7771 => x"842981f8",
          7772 => x"f8057008",
          7773 => x"51557480",
          7774 => x"2e843880",
          7775 => x"753481f8",
          7776 => x"c80881ff",
          7777 => x"065f8152",
          7778 => x"7e51ffa0",
          7779 => x"d03f81f8",
          7780 => x"c80881ff",
          7781 => x"06708106",
          7782 => x"56578356",
          7783 => x"748bc038",
          7784 => x"76822a70",
          7785 => x"81065155",
          7786 => x"8a56748b",
          7787 => x"b238993d",
          7788 => x"fc055383",
          7789 => x"527e51ff",
          7790 => x"a4f03f81",
          7791 => x"f8c80899",
          7792 => x"38675574",
          7793 => x"802e9238",
          7794 => x"74828080",
          7795 => x"268b38ff",
          7796 => x"15750655",
          7797 => x"74802e83",
          7798 => x"38814878",
          7799 => x"802e8738",
          7800 => x"84807926",
          7801 => x"92387881",
          7802 => x"800a268b",
          7803 => x"38ff1979",
          7804 => x"06557480",
          7805 => x"2e863893",
          7806 => x"568ae439",
          7807 => x"78892a6e",
          7808 => x"892a7089",
          7809 => x"2b775948",
          7810 => x"43597a83",
          7811 => x"38815661",
          7812 => x"30708025",
          7813 => x"77075155",
          7814 => x"9156748a",
          7815 => x"c238993d",
          7816 => x"f8055381",
          7817 => x"527e51ff",
          7818 => x"a4803f81",
          7819 => x"5681f8c8",
          7820 => x"088aac38",
          7821 => x"77832a70",
          7822 => x"770681f8",
          7823 => x"c8084356",
          7824 => x"45748338",
          7825 => x"bf416655",
          7826 => x"8e566075",
          7827 => x"268a9038",
          7828 => x"74613170",
          7829 => x"485580ff",
          7830 => x"75278a83",
          7831 => x"38935678",
          7832 => x"81802689",
          7833 => x"fa387781",
          7834 => x"2a708106",
          7835 => x"56437480",
          7836 => x"2e953877",
          7837 => x"87065574",
          7838 => x"822e838d",
          7839 => x"38778106",
          7840 => x"5574802e",
          7841 => x"83833877",
          7842 => x"81065593",
          7843 => x"56825e74",
          7844 => x"802e89cb",
          7845 => x"38785a7d",
          7846 => x"832e0981",
          7847 => x"0680e138",
          7848 => x"78ae3866",
          7849 => x"912a5781",
          7850 => x"0b81e7fc",
          7851 => x"22565a74",
          7852 => x"802e9d38",
          7853 => x"74772698",
          7854 => x"3881e7fc",
          7855 => x"56791082",
          7856 => x"17702257",
          7857 => x"575a7480",
          7858 => x"2e863876",
          7859 => x"7527ee38",
          7860 => x"79526651",
          7861 => x"feddd43f",
          7862 => x"81f8c808",
          7863 => x"84298487",
          7864 => x"0570892a",
          7865 => x"5e55a05c",
          7866 => x"800b81f8",
          7867 => x"c808fc80",
          7868 => x"8a055644",
          7869 => x"fdfff00a",
          7870 => x"752780ec",
          7871 => x"3888d339",
          7872 => x"78ae3866",
          7873 => x"8c2a5781",
          7874 => x"0b81e7ec",
          7875 => x"22565a74",
          7876 => x"802e9d38",
          7877 => x"74772698",
          7878 => x"3881e7ec",
          7879 => x"56791082",
          7880 => x"17702257",
          7881 => x"575a7480",
          7882 => x"2e863876",
          7883 => x"7527ee38",
          7884 => x"79526651",
          7885 => x"fedcf43f",
          7886 => x"81f8c808",
          7887 => x"10840557",
          7888 => x"81f8c808",
          7889 => x"9ff52696",
          7890 => x"38810b81",
          7891 => x"f8c80810",
          7892 => x"81f8c808",
          7893 => x"05711172",
          7894 => x"2a830559",
          7895 => x"565e83ff",
          7896 => x"17892a5d",
          7897 => x"815ca044",
          7898 => x"601c7d11",
          7899 => x"65056970",
          7900 => x"12ff0571",
          7901 => x"30707206",
          7902 => x"74315c52",
          7903 => x"59575940",
          7904 => x"7d832e09",
          7905 => x"81068938",
          7906 => x"761c6018",
          7907 => x"415c8439",
          7908 => x"761d5d79",
          7909 => x"90291870",
          7910 => x"62316858",
          7911 => x"51557476",
          7912 => x"2687af38",
          7913 => x"757c317d",
          7914 => x"317a5370",
          7915 => x"65315255",
          7916 => x"fedbf83f",
          7917 => x"81f8c808",
          7918 => x"587d832e",
          7919 => x"0981069b",
          7920 => x"3881f8c8",
          7921 => x"0883fff5",
          7922 => x"2680dd38",
          7923 => x"78878338",
          7924 => x"79812a59",
          7925 => x"78fdbe38",
          7926 => x"86f8397d",
          7927 => x"822e0981",
          7928 => x"0680c538",
          7929 => x"83fff50b",
          7930 => x"81f8c808",
          7931 => x"27a03878",
          7932 => x"8f38791a",
          7933 => x"557480c0",
          7934 => x"26863874",
          7935 => x"59fd9639",
          7936 => x"62810655",
          7937 => x"74802e8f",
          7938 => x"38835efd",
          7939 => x"883981f8",
          7940 => x"c8089ff5",
          7941 => x"26923878",
          7942 => x"86b83879",
          7943 => x"1a598180",
          7944 => x"7927fcf1",
          7945 => x"3886ab39",
          7946 => x"80557d81",
          7947 => x"2e098106",
          7948 => x"83387d55",
          7949 => x"9ff57827",
          7950 => x"8b387481",
          7951 => x"06558e56",
          7952 => x"74869c38",
          7953 => x"84805380",
          7954 => x"527a51ff",
          7955 => x"a2b93f8b",
          7956 => x"5381e694",
          7957 => x"527a51ff",
          7958 => x"a28a3f84",
          7959 => x"80528b1b",
          7960 => x"51ffa1b3",
          7961 => x"3f798d1c",
          7962 => x"347b83ff",
          7963 => x"ff06528e",
          7964 => x"1b51ffa1",
          7965 => x"a23f810b",
          7966 => x"901c347d",
          7967 => x"83327030",
          7968 => x"70962a84",
          7969 => x"80065451",
          7970 => x"55911b51",
          7971 => x"ffa1883f",
          7972 => x"66557483",
          7973 => x"ffff2690",
          7974 => x"387483ff",
          7975 => x"ff065293",
          7976 => x"1b51ffa0",
          7977 => x"f23f8a39",
          7978 => x"7452a01b",
          7979 => x"51ffa185",
          7980 => x"3ff80b95",
          7981 => x"1c34bf52",
          7982 => x"981b51ff",
          7983 => x"a0d93f81",
          7984 => x"ff529a1b",
          7985 => x"51ffa0cf",
          7986 => x"3f60529c",
          7987 => x"1b51ffa0",
          7988 => x"e43f7d83",
          7989 => x"2e098106",
          7990 => x"80cb3882",
          7991 => x"88b20a52",
          7992 => x"80c31b51",
          7993 => x"ffa0ce3f",
          7994 => x"7c52a41b",
          7995 => x"51ffa0c5",
          7996 => x"3f8252ac",
          7997 => x"1b51ffa0",
          7998 => x"bc3f8152",
          7999 => x"b01b51ff",
          8000 => x"a0953f86",
          8001 => x"52b21b51",
          8002 => x"ffa08c3f",
          8003 => x"ff800b80",
          8004 => x"c01c34a9",
          8005 => x"0b80c21c",
          8006 => x"34935381",
          8007 => x"e6a05280",
          8008 => x"c71b51ae",
          8009 => x"398288b2",
          8010 => x"0a52a71b",
          8011 => x"51ffa085",
          8012 => x"3f7c83ff",
          8013 => x"ff065296",
          8014 => x"1b51ff9f",
          8015 => x"da3fff80",
          8016 => x"0ba41c34",
          8017 => x"a90ba61c",
          8018 => x"34935381",
          8019 => x"e6b452ab",
          8020 => x"1b51ffa0",
          8021 => x"8f3f82d4",
          8022 => x"d55283fe",
          8023 => x"1b705259",
          8024 => x"ff9fb43f",
          8025 => x"81546053",
          8026 => x"7a527e51",
          8027 => x"ff9bd73f",
          8028 => x"815681f8",
          8029 => x"c80883e7",
          8030 => x"387d832e",
          8031 => x"09810680",
          8032 => x"ee387554",
          8033 => x"60860553",
          8034 => x"7a527e51",
          8035 => x"ff9bb73f",
          8036 => x"84805380",
          8037 => x"527a51ff",
          8038 => x"9fed3f84",
          8039 => x"8b85a4d2",
          8040 => x"527a51ff",
          8041 => x"9f8f3f86",
          8042 => x"8a85e4f2",
          8043 => x"5283e41b",
          8044 => x"51ff9f81",
          8045 => x"3fff1852",
          8046 => x"83e81b51",
          8047 => x"ff9ef63f",
          8048 => x"825283ec",
          8049 => x"1b51ff9e",
          8050 => x"ec3f82d4",
          8051 => x"d5527851",
          8052 => x"ff9ec43f",
          8053 => x"75546087",
          8054 => x"05537a52",
          8055 => x"7e51ff9a",
          8056 => x"e53f7554",
          8057 => x"6016537a",
          8058 => x"527e51ff",
          8059 => x"9ad83f65",
          8060 => x"5380527a",
          8061 => x"51ff9f8f",
          8062 => x"3f7f5680",
          8063 => x"587d832e",
          8064 => x"0981069a",
          8065 => x"38f8527a",
          8066 => x"51ff9ea9",
          8067 => x"3fff5284",
          8068 => x"1b51ff9e",
          8069 => x"a03ff00a",
          8070 => x"52881b51",
          8071 => x"913987ff",
          8072 => x"fff8557d",
          8073 => x"812e8338",
          8074 => x"f8557452",
          8075 => x"7a51ff9e",
          8076 => x"843f7c55",
          8077 => x"61577462",
          8078 => x"26833874",
          8079 => x"57765475",
          8080 => x"537a527e",
          8081 => x"51ff99fe",
          8082 => x"3f81f8c8",
          8083 => x"08828738",
          8084 => x"84805381",
          8085 => x"f8c80852",
          8086 => x"7a51ff9e",
          8087 => x"aa3f7616",
          8088 => x"75783156",
          8089 => x"5674cd38",
          8090 => x"81185877",
          8091 => x"802eff8d",
          8092 => x"3879557d",
          8093 => x"832e8338",
          8094 => x"63556157",
          8095 => x"74622683",
          8096 => x"38745776",
          8097 => x"5475537a",
          8098 => x"527e51ff",
          8099 => x"99b83f81",
          8100 => x"f8c80881",
          8101 => x"c1387616",
          8102 => x"75783156",
          8103 => x"5674db38",
          8104 => x"8c567d83",
          8105 => x"2e933886",
          8106 => x"566683ff",
          8107 => x"ff268a38",
          8108 => x"84567d82",
          8109 => x"2e833881",
          8110 => x"56648106",
          8111 => x"587780fe",
          8112 => x"38848053",
          8113 => x"77527a51",
          8114 => x"ff9dbc3f",
          8115 => x"82d4d552",
          8116 => x"7851ff9c",
          8117 => x"c23f83be",
          8118 => x"1b557775",
          8119 => x"34810b81",
          8120 => x"1634810b",
          8121 => x"82163477",
          8122 => x"83163475",
          8123 => x"84163460",
          8124 => x"67055680",
          8125 => x"fdc15275",
          8126 => x"51fed5af",
          8127 => x"3ffe0b85",
          8128 => x"163481f8",
          8129 => x"c808822a",
          8130 => x"bf075675",
          8131 => x"86163481",
          8132 => x"f8c80887",
          8133 => x"16346052",
          8134 => x"83c61b51",
          8135 => x"ff9c963f",
          8136 => x"665283ca",
          8137 => x"1b51ff9c",
          8138 => x"8c3f8154",
          8139 => x"77537a52",
          8140 => x"7e51ff98",
          8141 => x"913f8156",
          8142 => x"81f8c808",
          8143 => x"a2388053",
          8144 => x"80527e51",
          8145 => x"ff99e33f",
          8146 => x"815681f8",
          8147 => x"c8089038",
          8148 => x"89398e56",
          8149 => x"8a398156",
          8150 => x"863981f8",
          8151 => x"c8085675",
          8152 => x"81f8c80c",
          8153 => x"993d0d04",
          8154 => x"f53d0d7d",
          8155 => x"605b5980",
          8156 => x"7960ff05",
          8157 => x"5a575776",
          8158 => x"7825b438",
          8159 => x"8d3df811",
          8160 => x"55558153",
          8161 => x"fc155279",
          8162 => x"51c9dc3f",
          8163 => x"7a812e09",
          8164 => x"81069c38",
          8165 => x"8c3d3355",
          8166 => x"748d2edb",
          8167 => x"38747670",
          8168 => x"81055834",
          8169 => x"81175774",
          8170 => x"8a2e0981",
          8171 => x"06c93880",
          8172 => x"76347855",
          8173 => x"76833876",
          8174 => x"557481f8",
          8175 => x"c80c8d3d",
          8176 => x"0d04f73d",
          8177 => x"0d7b0284",
          8178 => x"05b30533",
          8179 => x"5957778a",
          8180 => x"2e098106",
          8181 => x"87388d52",
          8182 => x"7651e73f",
          8183 => x"84170856",
          8184 => x"807624be",
          8185 => x"38881708",
          8186 => x"77178c05",
          8187 => x"56597775",
          8188 => x"34811656",
          8189 => x"bb7625a1",
          8190 => x"388b3dfc",
          8191 => x"05547553",
          8192 => x"8c175276",
          8193 => x"0851cbdc",
          8194 => x"3f797632",
          8195 => x"70307072",
          8196 => x"079f2a70",
          8197 => x"30535156",
          8198 => x"56758418",
          8199 => x"0c811988",
          8200 => x"180c8b3d",
          8201 => x"0d04f93d",
          8202 => x"0d798411",
          8203 => x"08565680",
          8204 => x"7524a738",
          8205 => x"893dfc05",
          8206 => x"5474538c",
          8207 => x"16527508",
          8208 => x"51cba13f",
          8209 => x"81f8c808",
          8210 => x"91388416",
          8211 => x"08782e09",
          8212 => x"81068738",
          8213 => x"88160855",
          8214 => x"8339ff55",
          8215 => x"7481f8c8",
          8216 => x"0c893d0d",
          8217 => x"04fd3d0d",
          8218 => x"755480cc",
          8219 => x"53805273",
          8220 => x"51ff9a93",
          8221 => x"3f76740c",
          8222 => x"853d0d04",
          8223 => x"ea3d0d02",
          8224 => x"80e30533",
          8225 => x"6a53863d",
          8226 => x"70535454",
          8227 => x"d83f7352",
          8228 => x"7251feae",
          8229 => x"3f7251ff",
          8230 => x"8d3f983d",
          8231 => x"0d04f83d",
          8232 => x"0d7a7008",
          8233 => x"70565659",
          8234 => x"74802e80",
          8235 => x"e1388c39",
          8236 => x"7715790c",
          8237 => x"85163354",
          8238 => x"80d43974",
          8239 => x"335473a0",
          8240 => x"2e098106",
          8241 => x"86388115",
          8242 => x"55f13980",
          8243 => x"57769029",
          8244 => x"81f5b805",
          8245 => x"70085256",
          8246 => x"fedaf23f",
          8247 => x"81f8c808",
          8248 => x"81f8c808",
          8249 => x"54755376",
          8250 => x"085258fe",
          8251 => x"dbc03f81",
          8252 => x"f8c8088b",
          8253 => x"38841633",
          8254 => x"5473812e",
          8255 => x"ffb23881",
          8256 => x"177081ff",
          8257 => x"06585498",
          8258 => x"7727c238",
          8259 => x"ff547381",
          8260 => x"f8c80c8a",
          8261 => x"3d0d04ff",
          8262 => x"3d0d7352",
          8263 => x"71932681",
          8264 => x"8e387184",
          8265 => x"2981dd80",
          8266 => x"05527108",
          8267 => x"0481e9b4",
          8268 => x"51818039",
          8269 => x"81e9c051",
          8270 => x"80f93981",
          8271 => x"e9d45180",
          8272 => x"f23981e9",
          8273 => x"e85180eb",
          8274 => x"3981e9f8",
          8275 => x"5180e439",
          8276 => x"81ea8851",
          8277 => x"80dd3981",
          8278 => x"ea9c5180",
          8279 => x"d63981ea",
          8280 => x"ac5180cf",
          8281 => x"3981eac4",
          8282 => x"5180c839",
          8283 => x"81eadc51",
          8284 => x"80c13981",
          8285 => x"eaf451bb",
          8286 => x"3981eb90",
          8287 => x"51b53981",
          8288 => x"eba451af",
          8289 => x"3981ebd0",
          8290 => x"51a93981",
          8291 => x"ebe451a3",
          8292 => x"3981ec84",
          8293 => x"519d3981",
          8294 => x"ec985197",
          8295 => x"3981ecb0",
          8296 => x"51913981",
          8297 => x"ecc8518b",
          8298 => x"3981ece0",
          8299 => x"51853981",
          8300 => x"ecec51fe",
          8301 => x"f2ae3f83",
          8302 => x"3d0d04fb",
          8303 => x"3d0d7779",
          8304 => x"56567487",
          8305 => x"e7268a38",
          8306 => x"74527587",
          8307 => x"e8295191",
          8308 => x"3987e852",
          8309 => x"7451fecf",
          8310 => x"d23f81f8",
          8311 => x"c8085275",
          8312 => x"51fecfc7",
          8313 => x"3f81f8c8",
          8314 => x"08547953",
          8315 => x"755281ec",
          8316 => x"fc51fef7",
          8317 => x"d33f873d",
          8318 => x"0d04ec3d",
          8319 => x"0d660284",
          8320 => x"0580e305",
          8321 => x"335b5780",
          8322 => x"68783070",
          8323 => x"7a077325",
          8324 => x"51575959",
          8325 => x"78567787",
          8326 => x"ff268338",
          8327 => x"81567476",
          8328 => x"077081ff",
          8329 => x"06515593",
          8330 => x"56748180",
          8331 => x"38815376",
          8332 => x"528c3d70",
          8333 => x"5256ffbf",
          8334 => x"c93f81f8",
          8335 => x"c8085781",
          8336 => x"f8c808b8",
          8337 => x"3881f8c8",
          8338 => x"0887c098",
          8339 => x"880c81f8",
          8340 => x"c8085996",
          8341 => x"3dd40554",
          8342 => x"84805377",
          8343 => x"527551c4",
          8344 => x"863f81f8",
          8345 => x"c8085781",
          8346 => x"f8c80890",
          8347 => x"387a5574",
          8348 => x"802e8938",
          8349 => x"74197519",
          8350 => x"5959d839",
          8351 => x"963dd805",
          8352 => x"51cbf03f",
          8353 => x"76307078",
          8354 => x"0780257b",
          8355 => x"30709f2a",
          8356 => x"72065157",
          8357 => x"51567480",
          8358 => x"2e903881",
          8359 => x"eda05387",
          8360 => x"c0988808",
          8361 => x"527851fe",
          8362 => x"923f7656",
          8363 => x"7581f8c8",
          8364 => x"0c963d0d",
          8365 => x"04f93d0d",
          8366 => x"7b028405",
          8367 => x"b3053357",
          8368 => x"58ff5780",
          8369 => x"537a5279",
          8370 => x"51feaf3f",
          8371 => x"81f8c808",
          8372 => x"a4387580",
          8373 => x"2e883875",
          8374 => x"812e9838",
          8375 => x"98396055",
          8376 => x"7f5481f8",
          8377 => x"c8537e52",
          8378 => x"7d51772d",
          8379 => x"81f8c808",
          8380 => x"57833977",
          8381 => x"047681f8",
          8382 => x"c80c893d",
          8383 => x"0d04f33d",
          8384 => x"0d7f6163",
          8385 => x"028c0580",
          8386 => x"cf053373",
          8387 => x"73156841",
          8388 => x"5f5c5c5e",
          8389 => x"5e5e7a52",
          8390 => x"81eda851",
          8391 => x"fef5a93f",
          8392 => x"81edb051",
          8393 => x"feefbd3f",
          8394 => x"80557479",
          8395 => x"2780fc38",
          8396 => x"7b902e89",
          8397 => x"387ba02e",
          8398 => x"a73880c6",
          8399 => x"39741853",
          8400 => x"727a278e",
          8401 => x"38722252",
          8402 => x"81edb451",
          8403 => x"fef4f93f",
          8404 => x"893981ed",
          8405 => x"c051feef",
          8406 => x"8b3f8215",
          8407 => x"5580c339",
          8408 => x"74185372",
          8409 => x"7a278e38",
          8410 => x"72085281",
          8411 => x"eda851fe",
          8412 => x"f4d63f89",
          8413 => x"3981edbc",
          8414 => x"51feeee8",
          8415 => x"3f841555",
          8416 => x"a1397418",
          8417 => x"53727a27",
          8418 => x"8e387233",
          8419 => x"5281edc8",
          8420 => x"51fef4b4",
          8421 => x"3f893981",
          8422 => x"edd051fe",
          8423 => x"eec63f81",
          8424 => x"1555a051",
          8425 => x"feede03f",
          8426 => x"ff803981",
          8427 => x"edd451fe",
          8428 => x"eeb23f80",
          8429 => x"55747927",
          8430 => x"bc387418",
          8431 => x"70335553",
          8432 => x"8056727a",
          8433 => x"27833881",
          8434 => x"5680539f",
          8435 => x"74278338",
          8436 => x"81537573",
          8437 => x"067081ff",
          8438 => x"06515372",
          8439 => x"802e8b38",
          8440 => x"7380fe26",
          8441 => x"85387351",
          8442 => x"8339a051",
          8443 => x"feed983f",
          8444 => x"811555c1",
          8445 => x"3981edd8",
          8446 => x"51feede8",
          8447 => x"3f781879",
          8448 => x"1c5c58fe",
          8449 => x"ded73f81",
          8450 => x"f8c80898",
          8451 => x"2b70982c",
          8452 => x"515776a0",
          8453 => x"2e098106",
          8454 => x"ab38fede",
          8455 => x"c03f81f8",
          8456 => x"c808982b",
          8457 => x"70982c70",
          8458 => x"a0327030",
          8459 => x"729b3270",
          8460 => x"30707207",
          8461 => x"73750706",
          8462 => x"51585859",
          8463 => x"57515780",
          8464 => x"7324d738",
          8465 => x"769b2e09",
          8466 => x"81068538",
          8467 => x"80538c39",
          8468 => x"7c1e5372",
          8469 => x"7826fdbe",
          8470 => x"38ff5372",
          8471 => x"81f8c80c",
          8472 => x"8f3d0d04",
          8473 => x"fc3d0d02",
          8474 => x"9b053381",
          8475 => x"eddc5381",
          8476 => x"ede05255",
          8477 => x"fef2d13f",
          8478 => x"81f3f822",
          8479 => x"51fee798",
          8480 => x"3f81edec",
          8481 => x"5481edf8",
          8482 => x"5381f3f9",
          8483 => x"335281ee",
          8484 => x"8051fef2",
          8485 => x"b33f7480",
          8486 => x"2e8538fe",
          8487 => x"e2e33f86",
          8488 => x"3d0d04fe",
          8489 => x"3d0d87c0",
          8490 => x"96800853",
          8491 => x"fee7b13f",
          8492 => x"8151fed9",
          8493 => x"bc3f81ee",
          8494 => x"9c51fedb",
          8495 => x"b43f8051",
          8496 => x"fed9ae3f",
          8497 => x"72812a70",
          8498 => x"81065152",
          8499 => x"71802e95",
          8500 => x"388151fe",
          8501 => x"d99b3f81",
          8502 => x"eeb451fe",
          8503 => x"db933f80",
          8504 => x"51fed98d",
          8505 => x"3f72822a",
          8506 => x"70810651",
          8507 => x"5271802e",
          8508 => x"95388151",
          8509 => x"fed8fa3f",
          8510 => x"81eec851",
          8511 => x"fedaf23f",
          8512 => x"8051fed8",
          8513 => x"ec3f7283",
          8514 => x"2a708106",
          8515 => x"51527180",
          8516 => x"2e953881",
          8517 => x"51fed8d9",
          8518 => x"3f81eed8",
          8519 => x"51fedad1",
          8520 => x"3f8051fe",
          8521 => x"d8cb3f72",
          8522 => x"842a7081",
          8523 => x"06515271",
          8524 => x"802e9538",
          8525 => x"8151fed8",
          8526 => x"b83f81ee",
          8527 => x"ec51feda",
          8528 => x"b03f8051",
          8529 => x"fed8aa3f",
          8530 => x"72852a70",
          8531 => x"81065152",
          8532 => x"71802e95",
          8533 => x"388151fe",
          8534 => x"d8973f81",
          8535 => x"ef8051fe",
          8536 => x"da8f3f80",
          8537 => x"51fed889",
          8538 => x"3f72862a",
          8539 => x"70810651",
          8540 => x"5271802e",
          8541 => x"95388151",
          8542 => x"fed7f63f",
          8543 => x"81ef9451",
          8544 => x"fed9ee3f",
          8545 => x"8051fed7",
          8546 => x"e83f7287",
          8547 => x"2a708106",
          8548 => x"51527180",
          8549 => x"2e953881",
          8550 => x"51fed7d5",
          8551 => x"3f81efa8",
          8552 => x"51fed9cd",
          8553 => x"3f8051fe",
          8554 => x"d7c73f72",
          8555 => x"882a7081",
          8556 => x"06515271",
          8557 => x"802e9538",
          8558 => x"8151fed7",
          8559 => x"b43f81ef",
          8560 => x"bc51fed9",
          8561 => x"ac3f8051",
          8562 => x"fed7a63f",
          8563 => x"fee5993f",
          8564 => x"843d0d04",
          8565 => x"fb3d0d77",
          8566 => x"028405a3",
          8567 => x"05337055",
          8568 => x"56568052",
          8569 => x"7551fece",
          8570 => x"e43f81f5",
          8571 => x"b4335473",
          8572 => x"a7388153",
          8573 => x"81effc52",
          8574 => x"828fe051",
          8575 => x"ffb8833f",
          8576 => x"81f8c808",
          8577 => x"307081f8",
          8578 => x"c8080780",
          8579 => x"25827131",
          8580 => x"51515473",
          8581 => x"81f5b434",
          8582 => x"81f5b433",
          8583 => x"5473812e",
          8584 => x"098106ac",
          8585 => x"38828fe0",
          8586 => x"53745275",
          8587 => x"51f2b93f",
          8588 => x"81f8c808",
          8589 => x"802e8c38",
          8590 => x"81f8c808",
          8591 => x"51fee9a4",
          8592 => x"3f8e3982",
          8593 => x"8fe051c4",
          8594 => x"aa3f820b",
          8595 => x"81f5b434",
          8596 => x"81f5b433",
          8597 => x"5473822e",
          8598 => x"09810689",
          8599 => x"38745275",
          8600 => x"51fefae4",
          8601 => x"3f800b81",
          8602 => x"f8c80c87",
          8603 => x"3d0d04ce",
          8604 => x"3d0d8070",
          8605 => x"71828fdc",
          8606 => x"0c5f5d81",
          8607 => x"527c51ff",
          8608 => x"86db3f81",
          8609 => x"f8c80881",
          8610 => x"ff065978",
          8611 => x"7d2e0981",
          8612 => x"06a23881",
          8613 => x"f08c5296",
          8614 => x"3d705259",
          8615 => x"feeebf3f",
          8616 => x"7c537852",
          8617 => x"81fa8c51",
          8618 => x"ffb5f63f",
          8619 => x"81f8c808",
          8620 => x"7d2e8838",
          8621 => x"81f09051",
          8622 => x"8dbc3981",
          8623 => x"705f5d81",
          8624 => x"f0c851fe",
          8625 => x"e89e3f96",
          8626 => x"3d70465a",
          8627 => x"80f85279",
          8628 => x"51fe813f",
          8629 => x"b43dff84",
          8630 => x"0551f3c2",
          8631 => x"3f81f8c8",
          8632 => x"08902b70",
          8633 => x"902c5159",
          8634 => x"7880c22e",
          8635 => x"87b33878",
          8636 => x"80c224b2",
          8637 => x"3878bd2e",
          8638 => x"81d53878",
          8639 => x"bd249038",
          8640 => x"78802eff",
          8641 => x"ba3878bc",
          8642 => x"2e80da38",
          8643 => x"8ae93978",
          8644 => x"80c02e83",
          8645 => x"a1387880",
          8646 => x"c02485dd",
          8647 => x"3878bf2e",
          8648 => x"8292388a",
          8649 => x"d2397880",
          8650 => x"f92e89ea",
          8651 => x"387880f9",
          8652 => x"24923878",
          8653 => x"80c32e88",
          8654 => x"98387880",
          8655 => x"f82e89b1",
          8656 => x"388ab439",
          8657 => x"7881832e",
          8658 => x"8a993878",
          8659 => x"8183248b",
          8660 => x"38788182",
          8661 => x"2e89fd38",
          8662 => x"8a9d3978",
          8663 => x"81852e8a",
          8664 => x"8f388a93",
          8665 => x"39b43dff",
          8666 => x"801153ff",
          8667 => x"840551fe",
          8668 => x"eecb3f81",
          8669 => x"f8c80880",
          8670 => x"2efec438",
          8671 => x"b43dfefc",
          8672 => x"1153ff84",
          8673 => x"0551feee",
          8674 => x"b43f81f8",
          8675 => x"c808802e",
          8676 => x"fead38b4",
          8677 => x"3dfef811",
          8678 => x"53ff8405",
          8679 => x"51feee9d",
          8680 => x"3f81f8c8",
          8681 => x"08863881",
          8682 => x"f8c80842",
          8683 => x"81f0cc51",
          8684 => x"fee6b13f",
          8685 => x"63635c5a",
          8686 => x"797b2781",
          8687 => x"f2386159",
          8688 => x"787a7084",
          8689 => x"055c0c7a",
          8690 => x"7a26f538",
          8691 => x"81e139b4",
          8692 => x"3dff8011",
          8693 => x"53ff8405",
          8694 => x"51feede1",
          8695 => x"3f81f8c8",
          8696 => x"08802efd",
          8697 => x"da38b43d",
          8698 => x"fefc1153",
          8699 => x"ff840551",
          8700 => x"feedca3f",
          8701 => x"81f8c808",
          8702 => x"802efdc3",
          8703 => x"38b43dfe",
          8704 => x"f81153ff",
          8705 => x"840551fe",
          8706 => x"edb33f81",
          8707 => x"f8c80880",
          8708 => x"2efdac38",
          8709 => x"81f0dc51",
          8710 => x"fee5c93f",
          8711 => x"635a7963",
          8712 => x"27818c38",
          8713 => x"61597970",
          8714 => x"81055b33",
          8715 => x"79346181",
          8716 => x"0542eb39",
          8717 => x"b43dff80",
          8718 => x"1153ff84",
          8719 => x"0551feec",
          8720 => x"fc3f81f8",
          8721 => x"c808802e",
          8722 => x"fcf538b4",
          8723 => x"3dfefc11",
          8724 => x"53ff8405",
          8725 => x"51feece5",
          8726 => x"3f81f8c8",
          8727 => x"08802efc",
          8728 => x"de38b43d",
          8729 => x"fef81153",
          8730 => x"ff840551",
          8731 => x"feecce3f",
          8732 => x"81f8c808",
          8733 => x"802efcc7",
          8734 => x"3881f0e8",
          8735 => x"51fee4e4",
          8736 => x"3f635a79",
          8737 => x"6327a838",
          8738 => x"6170337b",
          8739 => x"335e5a5b",
          8740 => x"787c2e92",
          8741 => x"3878557a",
          8742 => x"54793353",
          8743 => x"795281f0",
          8744 => x"f851feea",
          8745 => x"a33f811a",
          8746 => x"62810543",
          8747 => x"5ad53981",
          8748 => x"f1905182",
          8749 => x"bd39b43d",
          8750 => x"ff801153",
          8751 => x"ff840551",
          8752 => x"feebfa3f",
          8753 => x"81f8c808",
          8754 => x"80df3881",
          8755 => x"f48c3359",
          8756 => x"78802e89",
          8757 => x"3881f3c4",
          8758 => x"084480cd",
          8759 => x"3981f48d",
          8760 => x"33597880",
          8761 => x"2e883881",
          8762 => x"f3cc0844",
          8763 => x"bc3981f4",
          8764 => x"8e335978",
          8765 => x"802e8838",
          8766 => x"81f3d408",
          8767 => x"44ab3981",
          8768 => x"f48f3359",
          8769 => x"78802e88",
          8770 => x"3881f3dc",
          8771 => x"08449a39",
          8772 => x"81f48a33",
          8773 => x"5978802e",
          8774 => x"883881f3",
          8775 => x"e4084489",
          8776 => x"3981f3f4",
          8777 => x"08fc8005",
          8778 => x"44b43dfe",
          8779 => x"fc1153ff",
          8780 => x"840551fe",
          8781 => x"eb873f81",
          8782 => x"f8c80880",
          8783 => x"de3881f4",
          8784 => x"8c335978",
          8785 => x"802e8938",
          8786 => x"81f3c808",
          8787 => x"4380cc39",
          8788 => x"81f48d33",
          8789 => x"5978802e",
          8790 => x"883881f3",
          8791 => x"d00843bb",
          8792 => x"3981f48e",
          8793 => x"33597880",
          8794 => x"2e883881",
          8795 => x"f3d80843",
          8796 => x"aa3981f4",
          8797 => x"8f335978",
          8798 => x"802e8838",
          8799 => x"81f3e008",
          8800 => x"43993981",
          8801 => x"f48a3359",
          8802 => x"78802e88",
          8803 => x"3881f3e8",
          8804 => x"08438839",
          8805 => x"81f3f408",
          8806 => x"880543b4",
          8807 => x"3dfef811",
          8808 => x"53ff8405",
          8809 => x"51feea95",
          8810 => x"3f81f8c8",
          8811 => x"08802ea7",
          8812 => x"3880625c",
          8813 => x"5c7a882e",
          8814 => x"8338815c",
          8815 => x"7a903270",
          8816 => x"30707207",
          8817 => x"9f2a707f",
          8818 => x"0651515a",
          8819 => x"5a78802e",
          8820 => x"88387aa0",
          8821 => x"2e833888",
          8822 => x"4281f194",
          8823 => x"51fee284",
          8824 => x"3fa05563",
          8825 => x"54615362",
          8826 => x"526351f2",
          8827 => x"913f81f1",
          8828 => x"a451fee1",
          8829 => x"ef3ff9c7",
          8830 => x"39b43dff",
          8831 => x"801153ff",
          8832 => x"840551fe",
          8833 => x"e9b73f81",
          8834 => x"f8c80880",
          8835 => x"2ef9b038",
          8836 => x"b43dfefc",
          8837 => x"1153ff84",
          8838 => x"0551fee9",
          8839 => x"a03f81f8",
          8840 => x"c808802e",
          8841 => x"a5386359",
          8842 => x"0280cb05",
          8843 => x"33793463",
          8844 => x"810544b4",
          8845 => x"3dfefc11",
          8846 => x"53ff8405",
          8847 => x"51fee8fd",
          8848 => x"3f81f8c8",
          8849 => x"08e038f8",
          8850 => x"f6396370",
          8851 => x"33545281",
          8852 => x"f1b051fe",
          8853 => x"e6f23f80",
          8854 => x"f8527951",
          8855 => x"fee7c33f",
          8856 => x"79457933",
          8857 => x"5978ae2e",
          8858 => x"f8d5389f",
          8859 => x"7927a038",
          8860 => x"b43dfefc",
          8861 => x"1153ff84",
          8862 => x"0551fee8",
          8863 => x"c03f81f8",
          8864 => x"c808802e",
          8865 => x"91386359",
          8866 => x"0280cb05",
          8867 => x"33793463",
          8868 => x"810544ff",
          8869 => x"b53981f1",
          8870 => x"bc51fee0",
          8871 => x"c73fffaa",
          8872 => x"39b43dfe",
          8873 => x"f41153ff",
          8874 => x"840551fe",
          8875 => x"ea813f81",
          8876 => x"f8c80880",
          8877 => x"2ef88838",
          8878 => x"b43dfef0",
          8879 => x"1153ff84",
          8880 => x"0551fee9",
          8881 => x"ea3f81f8",
          8882 => x"c808802e",
          8883 => x"a6386059",
          8884 => x"02be0522",
          8885 => x"79708205",
          8886 => x"5b237841",
          8887 => x"b43dfef0",
          8888 => x"1153ff84",
          8889 => x"0551fee9",
          8890 => x"c63f81f8",
          8891 => x"c808df38",
          8892 => x"f7cd3960",
          8893 => x"70225452",
          8894 => x"81f1c451",
          8895 => x"fee5c93f",
          8896 => x"80f85279",
          8897 => x"51fee69a",
          8898 => x"3f794579",
          8899 => x"335978ae",
          8900 => x"2ef7ac38",
          8901 => x"789f2687",
          8902 => x"38608205",
          8903 => x"41d539b4",
          8904 => x"3dfef011",
          8905 => x"53ff8405",
          8906 => x"51fee983",
          8907 => x"3f81f8c8",
          8908 => x"08802e92",
          8909 => x"38605902",
          8910 => x"be052279",
          8911 => x"7082055b",
          8912 => x"237841ff",
          8913 => x"ae3981f1",
          8914 => x"bc51fedf",
          8915 => x"973fffa3",
          8916 => x"39b43dfe",
          8917 => x"f41153ff",
          8918 => x"840551fe",
          8919 => x"e8d13f81",
          8920 => x"f8c80880",
          8921 => x"2ef6d838",
          8922 => x"b43dfef0",
          8923 => x"1153ff84",
          8924 => x"0551fee8",
          8925 => x"ba3f81f8",
          8926 => x"c808802e",
          8927 => x"a1386060",
          8928 => x"710c5960",
          8929 => x"840541b4",
          8930 => x"3dfef011",
          8931 => x"53ff8405",
          8932 => x"51fee89b",
          8933 => x"3f81f8c8",
          8934 => x"08e438f6",
          8935 => x"a2396070",
          8936 => x"08545281",
          8937 => x"f1d051fe",
          8938 => x"e49e3f80",
          8939 => x"f8527951",
          8940 => x"fee4ef3f",
          8941 => x"79457933",
          8942 => x"5978ae2e",
          8943 => x"f681389f",
          8944 => x"79279c38",
          8945 => x"b43dfef0",
          8946 => x"1153ff84",
          8947 => x"0551fee7",
          8948 => x"de3f81f8",
          8949 => x"c808802e",
          8950 => x"8d386060",
          8951 => x"710c5960",
          8952 => x"840541ff",
          8953 => x"b93981f1",
          8954 => x"bc51fedd",
          8955 => x"f73fffae",
          8956 => x"39b43dff",
          8957 => x"801153ff",
          8958 => x"840551fe",
          8959 => x"e5bf3f81",
          8960 => x"f8c80880",
          8961 => x"2ef5b838",
          8962 => x"635281f1",
          8963 => x"dc51fee3",
          8964 => x"b73f6359",
          8965 => x"7804b43d",
          8966 => x"ff801153",
          8967 => x"ff840551",
          8968 => x"fee59a3f",
          8969 => x"81f8c808",
          8970 => x"802ef593",
          8971 => x"38635281",
          8972 => x"f1f851fe",
          8973 => x"e3923f63",
          8974 => x"59782d81",
          8975 => x"f8c80880",
          8976 => x"2ef4fc38",
          8977 => x"81f8c808",
          8978 => x"5281f294",
          8979 => x"51fee2f8",
          8980 => x"3ff4ec39",
          8981 => x"81f2b051",
          8982 => x"fedd893f",
          8983 => x"febaad3f",
          8984 => x"f4dd3981",
          8985 => x"f2cc51fe",
          8986 => x"dcfa3f80",
          8987 => x"59ffa539",
          8988 => x"fed38e3f",
          8989 => x"f4c93979",
          8990 => x"45793359",
          8991 => x"78802ef4",
          8992 => x"be387d7d",
          8993 => x"06597880",
          8994 => x"2e81d338",
          8995 => x"b43dff84",
          8996 => x"0551fec6",
          8997 => x"8d3f81f8",
          8998 => x"c8085c81",
          8999 => x"5b7a822e",
          9000 => x"b2387a82",
          9001 => x"2489387a",
          9002 => x"812e8c38",
          9003 => x"80cd397a",
          9004 => x"832eb038",
          9005 => x"80c53981",
          9006 => x"f2e0567b",
          9007 => x"5581f2e4",
          9008 => x"54805381",
          9009 => x"f2e852b4",
          9010 => x"3dffb005",
          9011 => x"51fee28e",
          9012 => x"3fbb3981",
          9013 => x"f38852b4",
          9014 => x"3dffb005",
          9015 => x"51fee1fe",
          9016 => x"3fab397b",
          9017 => x"5581f2e4",
          9018 => x"54805381",
          9019 => x"f2f852b4",
          9020 => x"3dffb005",
          9021 => x"51fee1e6",
          9022 => x"3f93397b",
          9023 => x"54805381",
          9024 => x"f38452b4",
          9025 => x"3dffb005",
          9026 => x"51fee1d2",
          9027 => x"3f81f3c4",
          9028 => x"5881f990",
          9029 => x"57805664",
          9030 => x"55805483",
          9031 => x"80805383",
          9032 => x"808052b4",
          9033 => x"3dffb005",
          9034 => x"51eb8a3f",
          9035 => x"81f8c808",
          9036 => x"81f8c808",
          9037 => x"09703070",
          9038 => x"72078025",
          9039 => x"515b5b5f",
          9040 => x"805a7a83",
          9041 => x"26833881",
          9042 => x"5a787a06",
          9043 => x"5978802e",
          9044 => x"8d38811b",
          9045 => x"7081ff06",
          9046 => x"5c597afe",
          9047 => x"c0387d81",
          9048 => x"327d8132",
          9049 => x"0759788a",
          9050 => x"387eff2e",
          9051 => x"098106f2",
          9052 => x"ce3881f3",
          9053 => x"8c51fee0",
          9054 => x"cf3ff2c3",
          9055 => x"39fc3d0d",
          9056 => x"800b81f9",
          9057 => x"903487c0",
          9058 => x"948c7008",
          9059 => x"54558784",
          9060 => x"80527251",
          9061 => x"feb8943f",
          9062 => x"81f8c808",
          9063 => x"902b7508",
          9064 => x"55538784",
          9065 => x"80527351",
          9066 => x"feb8803f",
          9067 => x"7281f8c8",
          9068 => x"0807750c",
          9069 => x"87c0949c",
          9070 => x"70085455",
          9071 => x"87848052",
          9072 => x"7251feb7",
          9073 => x"e63f81f8",
          9074 => x"c808902b",
          9075 => x"75085553",
          9076 => x"87848052",
          9077 => x"7351feb7",
          9078 => x"d23f7281",
          9079 => x"f8c80807",
          9080 => x"750c8c80",
          9081 => x"830b87c0",
          9082 => x"94840c8c",
          9083 => x"80830b87",
          9084 => x"c094940c",
          9085 => x"a38b0b81",
          9086 => x"f8dc0ca6",
          9087 => x"8c0b81f8",
          9088 => x"e00cfecb",
          9089 => x"b03ffed4",
          9090 => x"d73f81f3",
          9091 => x"9c51fed9",
          9092 => x"d33f81f3",
          9093 => x"a851fed9",
          9094 => x"cb3f81c9",
          9095 => x"a351fed4",
          9096 => x"ba3f8151",
          9097 => x"ecbe3ff0",
          9098 => x"c63f8004",
          9099 => x"00ffffff",
          9100 => x"ff00ffff",
          9101 => x"ffff00ff",
          9102 => x"ffffff00",
          9103 => x"00001832",
          9104 => x"00001838",
          9105 => x"0000183e",
          9106 => x"00001844",
          9107 => x"0000184a",
          9108 => x"000025b5",
          9109 => x"00002691",
          9110 => x"00002734",
          9111 => x"00002774",
          9112 => x"00002797",
          9113 => x"00002824",
          9114 => x"0000248a",
          9115 => x"0000248a",
          9116 => x"00002861",
          9117 => x"000028d7",
          9118 => x"00002962",
          9119 => x"0000298b",
          9120 => x"000061a9",
          9121 => x"0000612d",
          9122 => x"00006134",
          9123 => x"0000613b",
          9124 => x"00006142",
          9125 => x"00006149",
          9126 => x"00006150",
          9127 => x"00006157",
          9128 => x"0000615e",
          9129 => x"00006165",
          9130 => x"0000616c",
          9131 => x"00006173",
          9132 => x"00006179",
          9133 => x"0000617f",
          9134 => x"00006185",
          9135 => x"0000618b",
          9136 => x"00006191",
          9137 => x"00006197",
          9138 => x"0000619d",
          9139 => x"000061a3",
          9140 => x"25642f25",
          9141 => x"642f2564",
          9142 => x"2025643a",
          9143 => x"25643a25",
          9144 => x"642e2564",
          9145 => x"25640a00",
          9146 => x"536f4320",
          9147 => x"436f6e66",
          9148 => x"69677572",
          9149 => x"6174696f",
          9150 => x"6e000000",
          9151 => x"20286672",
          9152 => x"6f6d2053",
          9153 => x"6f432063",
          9154 => x"6f6e6669",
          9155 => x"67290000",
          9156 => x"3a0a4465",
          9157 => x"76696365",
          9158 => x"7320696d",
          9159 => x"706c656d",
          9160 => x"656e7465",
          9161 => x"643a0a00",
          9162 => x"20202020",
          9163 => x"57422053",
          9164 => x"4452414d",
          9165 => x"20202825",
          9166 => x"3038583a",
          9167 => x"25303858",
          9168 => x"292e0a00",
          9169 => x"20202020",
          9170 => x"53445241",
          9171 => x"4d202020",
          9172 => x"20202825",
          9173 => x"3038583a",
          9174 => x"25303858",
          9175 => x"292e0a00",
          9176 => x"20202020",
          9177 => x"494e534e",
          9178 => x"20425241",
          9179 => x"4d202825",
          9180 => x"3038583a",
          9181 => x"25303858",
          9182 => x"292e0a00",
          9183 => x"20202020",
          9184 => x"4252414d",
          9185 => x"20202020",
          9186 => x"20202825",
          9187 => x"3038583a",
          9188 => x"25303858",
          9189 => x"292e0a00",
          9190 => x"20202020",
          9191 => x"52414d20",
          9192 => x"20202020",
          9193 => x"20202825",
          9194 => x"3038583a",
          9195 => x"25303858",
          9196 => x"292e0a00",
          9197 => x"20202020",
          9198 => x"53442043",
          9199 => x"41524420",
          9200 => x"20202844",
          9201 => x"65766963",
          9202 => x"6573203d",
          9203 => x"25303264",
          9204 => x"292e0a00",
          9205 => x"20202020",
          9206 => x"54494d45",
          9207 => x"52312020",
          9208 => x"20202854",
          9209 => x"696d6572",
          9210 => x"7320203d",
          9211 => x"25303264",
          9212 => x"292e0a00",
          9213 => x"20202020",
          9214 => x"494e5452",
          9215 => x"20435452",
          9216 => x"4c202843",
          9217 => x"68616e6e",
          9218 => x"656c733d",
          9219 => x"25303264",
          9220 => x"292e0a00",
          9221 => x"20202020",
          9222 => x"57495348",
          9223 => x"424f4e45",
          9224 => x"20425553",
          9225 => x"0a000000",
          9226 => x"20202020",
          9227 => x"57422049",
          9228 => x"32430a00",
          9229 => x"20202020",
          9230 => x"494f4354",
          9231 => x"4c0a0000",
          9232 => x"20202020",
          9233 => x"5053320a",
          9234 => x"00000000",
          9235 => x"20202020",
          9236 => x"5350490a",
          9237 => x"00000000",
          9238 => x"41646472",
          9239 => x"65737365",
          9240 => x"733a0a00",
          9241 => x"20202020",
          9242 => x"43505520",
          9243 => x"52657365",
          9244 => x"74205665",
          9245 => x"63746f72",
          9246 => x"20416464",
          9247 => x"72657373",
          9248 => x"203d2025",
          9249 => x"3038580a",
          9250 => x"00000000",
          9251 => x"20202020",
          9252 => x"43505520",
          9253 => x"4d656d6f",
          9254 => x"72792053",
          9255 => x"74617274",
          9256 => x"20416464",
          9257 => x"72657373",
          9258 => x"203d2025",
          9259 => x"3038580a",
          9260 => x"00000000",
          9261 => x"20202020",
          9262 => x"53746163",
          9263 => x"6b205374",
          9264 => x"61727420",
          9265 => x"41646472",
          9266 => x"65737320",
          9267 => x"20202020",
          9268 => x"203d2025",
          9269 => x"3038580a",
          9270 => x"00000000",
          9271 => x"4d697363",
          9272 => x"3a0a0000",
          9273 => x"20202020",
          9274 => x"5a505520",
          9275 => x"49642020",
          9276 => x"20202020",
          9277 => x"20202020",
          9278 => x"20202020",
          9279 => x"20202020",
          9280 => x"203d2025",
          9281 => x"3034580a",
          9282 => x"00000000",
          9283 => x"20202020",
          9284 => x"53797374",
          9285 => x"656d2043",
          9286 => x"6c6f636b",
          9287 => x"20467265",
          9288 => x"71202020",
          9289 => x"20202020",
          9290 => x"203d2025",
          9291 => x"642e2530",
          9292 => x"34644d48",
          9293 => x"7a0a0000",
          9294 => x"20202020",
          9295 => x"53445241",
          9296 => x"4d20436c",
          9297 => x"6f636b20",
          9298 => x"46726571",
          9299 => x"20202020",
          9300 => x"20202020",
          9301 => x"203d2025",
          9302 => x"642e2530",
          9303 => x"34644d48",
          9304 => x"7a0a0000",
          9305 => x"20202020",
          9306 => x"57697368",
          9307 => x"626f6e65",
          9308 => x"20534452",
          9309 => x"414d2043",
          9310 => x"6c6f636b",
          9311 => x"20467265",
          9312 => x"713d2025",
          9313 => x"642e2530",
          9314 => x"34644d48",
          9315 => x"7a0a0000",
          9316 => x"536d616c",
          9317 => x"6c000000",
          9318 => x"4d656469",
          9319 => x"756d0000",
          9320 => x"466c6578",
          9321 => x"00000000",
          9322 => x"45564f00",
          9323 => x"45564f6d",
          9324 => x"696e0000",
          9325 => x"556e6b6e",
          9326 => x"6f776e00",
          9327 => x"68697374",
          9328 => x"6f72792e",
          9329 => x"74787400",
          9330 => x"68697374",
          9331 => x"6f727900",
          9332 => x"68697374",
          9333 => x"00000000",
          9334 => x"21000000",
          9335 => x"25303464",
          9336 => x"20202573",
          9337 => x"0a000000",
          9338 => x"4661696c",
          9339 => x"65642074",
          9340 => x"6f207265",
          9341 => x"73657420",
          9342 => x"74686520",
          9343 => x"68697374",
          9344 => x"6f727920",
          9345 => x"66696c65",
          9346 => x"20746f20",
          9347 => x"454f462e",
          9348 => x"0a000000",
          9349 => x"43616e6e",
          9350 => x"6f74206f",
          9351 => x"70656e2f",
          9352 => x"63726561",
          9353 => x"74652068",
          9354 => x"6973746f",
          9355 => x"72792066",
          9356 => x"696c652c",
          9357 => x"20646973",
          9358 => x"61626c69",
          9359 => x"6e672e0a",
          9360 => x"00000000",
          9361 => x"000072f0",
          9362 => x"01000000",
          9363 => x"00000001",
          9364 => x"000072ec",
          9365 => x"01000000",
          9366 => x"00000002",
          9367 => x"000072e8",
          9368 => x"04000000",
          9369 => x"00000003",
          9370 => x"000072e4",
          9371 => x"04000000",
          9372 => x"00000004",
          9373 => x"000072e0",
          9374 => x"04000000",
          9375 => x"00000005",
          9376 => x"000072dc",
          9377 => x"04000000",
          9378 => x"00000006",
          9379 => x"000072d8",
          9380 => x"04000000",
          9381 => x"00000007",
          9382 => x"000072d4",
          9383 => x"03000000",
          9384 => x"00000008",
          9385 => x"000072d0",
          9386 => x"03000000",
          9387 => x"00000009",
          9388 => x"000072cc",
          9389 => x"03000000",
          9390 => x"0000000a",
          9391 => x"000072c8",
          9392 => x"03000000",
          9393 => x"0000000b",
          9394 => x"1b5b4400",
          9395 => x"1b5b4300",
          9396 => x"1b5b4200",
          9397 => x"1b5b4100",
          9398 => x"1b5b367e",
          9399 => x"1b5b357e",
          9400 => x"1b5b347e",
          9401 => x"1b5b337e",
          9402 => x"1b5b317e",
          9403 => x"0d000000",
          9404 => x"08000000",
          9405 => x"53440000",
          9406 => x"222a2b2c",
          9407 => x"3a3b3c3d",
          9408 => x"3e3f5b5d",
          9409 => x"7c7f0000",
          9410 => x"46415400",
          9411 => x"46415433",
          9412 => x"32000000",
          9413 => x"ebfe904d",
          9414 => x"53444f53",
          9415 => x"352e3000",
          9416 => x"4e4f204e",
          9417 => x"414d4520",
          9418 => x"20202046",
          9419 => x"41543332",
          9420 => x"20202000",
          9421 => x"4e4f204e",
          9422 => x"414d4520",
          9423 => x"20202046",
          9424 => x"41542020",
          9425 => x"20202000",
          9426 => x"000072f4",
          9427 => x"00000000",
          9428 => x"00000000",
          9429 => x"00000000",
          9430 => x"809a4541",
          9431 => x"8e418f80",
          9432 => x"45454549",
          9433 => x"49498e8f",
          9434 => x"9092924f",
          9435 => x"994f5555",
          9436 => x"59999a9b",
          9437 => x"9c9d9e9f",
          9438 => x"41494f55",
          9439 => x"a5a5a6a7",
          9440 => x"a8a9aaab",
          9441 => x"acadaeaf",
          9442 => x"b0b1b2b3",
          9443 => x"b4b5b6b7",
          9444 => x"b8b9babb",
          9445 => x"bcbdbebf",
          9446 => x"c0c1c2c3",
          9447 => x"c4c5c6c7",
          9448 => x"c8c9cacb",
          9449 => x"cccdcecf",
          9450 => x"d0d1d2d3",
          9451 => x"d4d5d6d7",
          9452 => x"d8d9dadb",
          9453 => x"dcdddedf",
          9454 => x"e0e1e2e3",
          9455 => x"e4e5e6e7",
          9456 => x"e8e9eaeb",
          9457 => x"ecedeeef",
          9458 => x"f0f1f2f3",
          9459 => x"f4f5f6f7",
          9460 => x"f8f9fafb",
          9461 => x"fcfdfeff",
          9462 => x"2b2e2c3b",
          9463 => x"3d5b5d2f",
          9464 => x"5c222a3a",
          9465 => x"3c3e3f7c",
          9466 => x"7f000000",
          9467 => x"00010004",
          9468 => x"00100040",
          9469 => x"01000200",
          9470 => x"00000000",
          9471 => x"00010002",
          9472 => x"00040008",
          9473 => x"00100020",
          9474 => x"00000000",
          9475 => x"64696e69",
          9476 => x"74000000",
          9477 => x"64696f63",
          9478 => x"746c0000",
          9479 => x"66696e69",
          9480 => x"74000000",
          9481 => x"666c6f61",
          9482 => x"64000000",
          9483 => x"66657865",
          9484 => x"63000000",
          9485 => x"6d636c65",
          9486 => x"61720000",
          9487 => x"6d636f70",
          9488 => x"79000000",
          9489 => x"6d646966",
          9490 => x"66000000",
          9491 => x"6d64756d",
          9492 => x"70000000",
          9493 => x"6d656200",
          9494 => x"6d656800",
          9495 => x"6d657700",
          9496 => x"68696400",
          9497 => x"68696500",
          9498 => x"68666400",
          9499 => x"68666500",
          9500 => x"63616c6c",
          9501 => x"00000000",
          9502 => x"6a6d7000",
          9503 => x"72657374",
          9504 => x"61727400",
          9505 => x"72657365",
          9506 => x"74000000",
          9507 => x"696e666f",
          9508 => x"00000000",
          9509 => x"74657374",
          9510 => x"00000000",
          9511 => x"74626173",
          9512 => x"69630000",
          9513 => x"6d626173",
          9514 => x"69630000",
          9515 => x"6b696c6f",
          9516 => x"00000000",
          9517 => x"4469736b",
          9518 => x"20457272",
          9519 => x"6f720a00",
          9520 => x"496e7465",
          9521 => x"726e616c",
          9522 => x"20657272",
          9523 => x"6f722e0a",
          9524 => x"00000000",
          9525 => x"4469736b",
          9526 => x"206e6f74",
          9527 => x"20726561",
          9528 => x"64792e0a",
          9529 => x"00000000",
          9530 => x"4e6f2066",
          9531 => x"696c6520",
          9532 => x"666f756e",
          9533 => x"642e0a00",
          9534 => x"4e6f2070",
          9535 => x"61746820",
          9536 => x"666f756e",
          9537 => x"642e0a00",
          9538 => x"496e7661",
          9539 => x"6c696420",
          9540 => x"66696c65",
          9541 => x"6e616d65",
          9542 => x"2e0a0000",
          9543 => x"41636365",
          9544 => x"73732064",
          9545 => x"656e6965",
          9546 => x"642e0a00",
          9547 => x"46696c65",
          9548 => x"20616c72",
          9549 => x"65616479",
          9550 => x"20657869",
          9551 => x"7374732e",
          9552 => x"0a000000",
          9553 => x"46696c65",
          9554 => x"2068616e",
          9555 => x"646c6520",
          9556 => x"696e7661",
          9557 => x"6c69642e",
          9558 => x"0a000000",
          9559 => x"53442069",
          9560 => x"73207772",
          9561 => x"69746520",
          9562 => x"70726f74",
          9563 => x"65637465",
          9564 => x"642e0a00",
          9565 => x"44726976",
          9566 => x"65206e75",
          9567 => x"6d626572",
          9568 => x"20697320",
          9569 => x"696e7661",
          9570 => x"6c69642e",
          9571 => x"0a000000",
          9572 => x"4469736b",
          9573 => x"206e6f74",
          9574 => x"20656e61",
          9575 => x"626c6564",
          9576 => x"2e0a0000",
          9577 => x"4e6f2063",
          9578 => x"6f6d7061",
          9579 => x"7469626c",
          9580 => x"65206669",
          9581 => x"6c657379",
          9582 => x"7374656d",
          9583 => x"20666f75",
          9584 => x"6e64206f",
          9585 => x"6e206469",
          9586 => x"736b2e0a",
          9587 => x"00000000",
          9588 => x"466f726d",
          9589 => x"61742061",
          9590 => x"626f7274",
          9591 => x"65642e0a",
          9592 => x"00000000",
          9593 => x"54696d65",
          9594 => x"6f75742c",
          9595 => x"206f7065",
          9596 => x"72617469",
          9597 => x"6f6e2063",
          9598 => x"616e6365",
          9599 => x"6c6c6564",
          9600 => x"2e0a0000",
          9601 => x"46696c65",
          9602 => x"20697320",
          9603 => x"6c6f636b",
          9604 => x"65642e0a",
          9605 => x"00000000",
          9606 => x"496e7375",
          9607 => x"66666963",
          9608 => x"69656e74",
          9609 => x"206d656d",
          9610 => x"6f72792e",
          9611 => x"0a000000",
          9612 => x"546f6f20",
          9613 => x"6d616e79",
          9614 => x"206f7065",
          9615 => x"6e206669",
          9616 => x"6c65732e",
          9617 => x"0a000000",
          9618 => x"50617261",
          9619 => x"6d657465",
          9620 => x"72732069",
          9621 => x"6e636f72",
          9622 => x"72656374",
          9623 => x"2e0a0000",
          9624 => x"53756363",
          9625 => x"6573732e",
          9626 => x"0a000000",
          9627 => x"556e6b6e",
          9628 => x"6f776e20",
          9629 => x"6572726f",
          9630 => x"722e0a00",
          9631 => x"0a256c75",
          9632 => x"20627974",
          9633 => x"65732025",
          9634 => x"73206174",
          9635 => x"20256c75",
          9636 => x"20627974",
          9637 => x"65732f73",
          9638 => x"65632e0a",
          9639 => x"00000000",
          9640 => x"72656164",
          9641 => x"00000000",
          9642 => x"25303858",
          9643 => x"00000000",
          9644 => x"3a202000",
          9645 => x"25303458",
          9646 => x"00000000",
          9647 => x"20202020",
          9648 => x"20202020",
          9649 => x"00000000",
          9650 => x"25303258",
          9651 => x"00000000",
          9652 => x"20200000",
          9653 => x"207c0000",
          9654 => x"7c0d0a00",
          9655 => x"7a4f5300",
          9656 => x"0a2a2a20",
          9657 => x"25732028",
          9658 => x"00000000",
          9659 => x"31372f30",
          9660 => x"342f3230",
          9661 => x"32300000",
          9662 => x"76312e30",
          9663 => x"31000000",
          9664 => x"205a5055",
          9665 => x"2c207265",
          9666 => x"76202530",
          9667 => x"32782920",
          9668 => x"25732025",
          9669 => x"73202a2a",
          9670 => x"0a0a0000",
          9671 => x"5a505520",
          9672 => x"496e7465",
          9673 => x"72727570",
          9674 => x"74204861",
          9675 => x"6e646c65",
          9676 => x"720a0000",
          9677 => x"54696d65",
          9678 => x"7220696e",
          9679 => x"74657272",
          9680 => x"7570740a",
          9681 => x"00000000",
          9682 => x"50533220",
          9683 => x"696e7465",
          9684 => x"72727570",
          9685 => x"740a0000",
          9686 => x"494f4354",
          9687 => x"4c205244",
          9688 => x"20696e74",
          9689 => x"65727275",
          9690 => x"70740a00",
          9691 => x"494f4354",
          9692 => x"4c205752",
          9693 => x"20696e74",
          9694 => x"65727275",
          9695 => x"70740a00",
          9696 => x"55415254",
          9697 => x"30205258",
          9698 => x"20696e74",
          9699 => x"65727275",
          9700 => x"70740a00",
          9701 => x"55415254",
          9702 => x"30205458",
          9703 => x"20696e74",
          9704 => x"65727275",
          9705 => x"70740a00",
          9706 => x"55415254",
          9707 => x"31205258",
          9708 => x"20696e74",
          9709 => x"65727275",
          9710 => x"70740a00",
          9711 => x"55415254",
          9712 => x"31205458",
          9713 => x"20696e74",
          9714 => x"65727275",
          9715 => x"70740a00",
          9716 => x"53657474",
          9717 => x"696e6720",
          9718 => x"75702074",
          9719 => x"696d6572",
          9720 => x"2e2e2e0a",
          9721 => x"00000000",
          9722 => x"456e6162",
          9723 => x"6c696e67",
          9724 => x"2074696d",
          9725 => x"65722e2e",
          9726 => x"2e0a0000",
          9727 => x"6175746f",
          9728 => x"65786563",
          9729 => x"2e626174",
          9730 => x"00000000",
          9731 => x"303a0000",
          9732 => x"4661696c",
          9733 => x"65642074",
          9734 => x"6f20696e",
          9735 => x"69746961",
          9736 => x"6c697365",
          9737 => x"20736420",
          9738 => x"63617264",
          9739 => x"20302c20",
          9740 => x"706c6561",
          9741 => x"73652069",
          9742 => x"6e697420",
          9743 => x"6d616e75",
          9744 => x"616c6c79",
          9745 => x"2e0a0000",
          9746 => x"2a200000",
          9747 => x"436c6561",
          9748 => x"72696e67",
          9749 => x"2e2e2e2e",
          9750 => x"00000000",
          9751 => x"436f7079",
          9752 => x"696e672e",
          9753 => x"2e2e0000",
          9754 => x"436f6d70",
          9755 => x"6172696e",
          9756 => x"672e2e2e",
          9757 => x"00000000",
          9758 => x"2530386c",
          9759 => x"78282530",
          9760 => x"3878292d",
          9761 => x"3e253038",
          9762 => x"6c782825",
          9763 => x"30387829",
          9764 => x"0a000000",
          9765 => x"44756d70",
          9766 => x"204d656d",
          9767 => x"6f72790a",
          9768 => x"00000000",
          9769 => x"0a436f6d",
          9770 => x"706c6574",
          9771 => x"652e0a00",
          9772 => x"25303858",
          9773 => x"20253032",
          9774 => x"582d0000",
          9775 => x"3f3f3f0a",
          9776 => x"00000000",
          9777 => x"25303858",
          9778 => x"20253034",
          9779 => x"582d0000",
          9780 => x"25303858",
          9781 => x"20253038",
          9782 => x"582d0000",
          9783 => x"45786563",
          9784 => x"7574696e",
          9785 => x"6720636f",
          9786 => x"64652040",
          9787 => x"20253038",
          9788 => x"78202e2e",
          9789 => x"2e0a0000",
          9790 => x"43616c6c",
          9791 => x"696e6720",
          9792 => x"636f6465",
          9793 => x"20402025",
          9794 => x"30387820",
          9795 => x"2e2e2e0a",
          9796 => x"00000000",
          9797 => x"43616c6c",
          9798 => x"20726574",
          9799 => x"75726e65",
          9800 => x"6420636f",
          9801 => x"64652028",
          9802 => x"2564292e",
          9803 => x"0a000000",
          9804 => x"52657374",
          9805 => x"61727469",
          9806 => x"6e672061",
          9807 => x"70706c69",
          9808 => x"63617469",
          9809 => x"6f6e2e2e",
          9810 => x"2e0a0000",
          9811 => x"436f6c64",
          9812 => x"20726562",
          9813 => x"6f6f7469",
          9814 => x"6e672e2e",
          9815 => x"2e0a0000",
          9816 => x"5a505500",
          9817 => x"62696e00",
          9818 => x"25643a5c",
          9819 => x"25735c25",
          9820 => x"732e2573",
          9821 => x"00000000",
          9822 => x"25643a5c",
          9823 => x"25735c25",
          9824 => x"73000000",
          9825 => x"25643a5c",
          9826 => x"25730000",
          9827 => x"42616420",
          9828 => x"636f6d6d",
          9829 => x"616e642e",
          9830 => x"0a000000",
          9831 => x"52756e6e",
          9832 => x"696e672e",
          9833 => x"2e2e0a00",
          9834 => x"456e6162",
          9835 => x"6c696e67",
          9836 => x"20696e74",
          9837 => x"65727275",
          9838 => x"7074732e",
          9839 => x"2e2e0a00",
          9840 => x"00000000",
          9841 => x"00000000",
          9842 => x"00007fff",
          9843 => x"00000000",
          9844 => x"00007fff",
          9845 => x"00010000",
          9846 => x"00007fff",
          9847 => x"00010000",
          9848 => x"00810000",
          9849 => x"01000000",
          9850 => x"017fffff",
          9851 => x"00000000",
          9852 => x"00000000",
          9853 => x"00007800",
          9854 => x"00000000",
          9855 => x"05f5e100",
          9856 => x"05f5e100",
          9857 => x"05f5e100",
          9858 => x"00000000",
          9859 => x"01010101",
          9860 => x"01010101",
          9861 => x"01011001",
          9862 => x"01000000",
          9863 => x"00000000",
          9864 => x"00000002",
          9865 => x"00000000",
          9866 => x"00007a20",
          9867 => x"00007a20",
          9868 => x"00007a20",
          9869 => x"00007a20",
          9870 => x"000071bc",
          9871 => x"00000000",
          9872 => x"00000000",
          9873 => x"00000000",
          9874 => x"00000000",
          9875 => x"00000000",
          9876 => x"00000000",
          9877 => x"00000000",
          9878 => x"00000000",
          9879 => x"00000000",
          9880 => x"00000000",
          9881 => x"00000000",
          9882 => x"00000000",
          9883 => x"00000000",
          9884 => x"00000000",
          9885 => x"00000000",
          9886 => x"00000000",
          9887 => x"00000000",
          9888 => x"00000000",
          9889 => x"00000000",
          9890 => x"00000000",
          9891 => x"00000000",
          9892 => x"00000000",
          9893 => x"00000000",
          9894 => x"000071c8",
          9895 => x"01000000",
          9896 => x"000071d0",
          9897 => x"01000000",
          9898 => x"000071d8",
          9899 => x"02000000",
          9900 => x"01000000",
          9901 => x"00000000",
          9902 => x"0000740c",
          9903 => x"01020100",
          9904 => x"00000000",
          9905 => x"00000000",
          9906 => x"00007414",
          9907 => x"01040100",
          9908 => x"00000000",
          9909 => x"00000000",
          9910 => x"0000741c",
          9911 => x"01140300",
          9912 => x"00000000",
          9913 => x"00000000",
          9914 => x"00007424",
          9915 => x"012b0300",
          9916 => x"00000000",
          9917 => x"00000000",
          9918 => x"0000742c",
          9919 => x"01300300",
          9920 => x"00000000",
          9921 => x"00000000",
          9922 => x"00007434",
          9923 => x"013c0400",
          9924 => x"00000000",
          9925 => x"00000000",
          9926 => x"0000743c",
          9927 => x"013d0400",
          9928 => x"00000000",
          9929 => x"00000000",
          9930 => x"00007444",
          9931 => x"013f0400",
          9932 => x"00000000",
          9933 => x"00000000",
          9934 => x"0000744c",
          9935 => x"01400400",
          9936 => x"00000000",
          9937 => x"00000000",
          9938 => x"00007454",
          9939 => x"01410400",
          9940 => x"00000000",
          9941 => x"00000000",
          9942 => x"00007458",
          9943 => x"01420400",
          9944 => x"00000000",
          9945 => x"00000000",
          9946 => x"0000745c",
          9947 => x"01430400",
          9948 => x"00000000",
          9949 => x"00000000",
          9950 => x"00007460",
          9951 => x"01500500",
          9952 => x"00000000",
          9953 => x"00000000",
          9954 => x"00007464",
          9955 => x"01510500",
          9956 => x"00000000",
          9957 => x"00000000",
          9958 => x"00007468",
          9959 => x"01540500",
          9960 => x"00000000",
          9961 => x"00000000",
          9962 => x"0000746c",
          9963 => x"01550500",
          9964 => x"00000000",
          9965 => x"00000000",
          9966 => x"00007470",
          9967 => x"01790700",
          9968 => x"00000000",
          9969 => x"00000000",
          9970 => x"00007478",
          9971 => x"01780700",
          9972 => x"00000000",
          9973 => x"00000000",
          9974 => x"0000747c",
          9975 => x"01820800",
          9976 => x"00000000",
          9977 => x"00000000",
          9978 => x"00007484",
          9979 => x"01830800",
          9980 => x"00000000",
          9981 => x"00000000",
          9982 => x"0000748c",
          9983 => x"01850800",
          9984 => x"00000000",
          9985 => x"00000000",
          9986 => x"00007494",
          9987 => x"01870800",
          9988 => x"00000000",
          9989 => x"00000000",
          9990 => x"0000749c",
          9991 => x"018c0900",
          9992 => x"00000000",
          9993 => x"00000000",
          9994 => x"000074a4",
          9995 => x"018d0900",
          9996 => x"00000000",
          9997 => x"00000000",
          9998 => x"000074ac",
          9999 => x"018e0900",
         10000 => x"00000000",
         10001 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

