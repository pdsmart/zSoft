-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"93",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"92",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"d3",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"e1",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"94",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"95",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"fc",
           386 => x"2d",
           387 => x"08",
           388 => x"04",
           389 => x"0c",
           390 => x"81",
           391 => x"83",
           392 => x"81",
           393 => x"b6",
           394 => x"fe",
           395 => x"80",
           396 => x"fe",
           397 => x"a5",
           398 => x"fc",
           399 => x"90",
           400 => x"fc",
           401 => x"2d",
           402 => x"08",
           403 => x"04",
           404 => x"0c",
           405 => x"81",
           406 => x"83",
           407 => x"81",
           408 => x"b6",
           409 => x"fe",
           410 => x"80",
           411 => x"fe",
           412 => x"fe",
           413 => x"fc",
           414 => x"90",
           415 => x"fc",
           416 => x"2d",
           417 => x"08",
           418 => x"04",
           419 => x"0c",
           420 => x"81",
           421 => x"83",
           422 => x"81",
           423 => x"b6",
           424 => x"fe",
           425 => x"80",
           426 => x"fe",
           427 => x"9f",
           428 => x"fc",
           429 => x"90",
           430 => x"fc",
           431 => x"2d",
           432 => x"08",
           433 => x"04",
           434 => x"0c",
           435 => x"81",
           436 => x"83",
           437 => x"81",
           438 => x"a6",
           439 => x"fe",
           440 => x"80",
           441 => x"fe",
           442 => x"f9",
           443 => x"fc",
           444 => x"90",
           445 => x"fc",
           446 => x"2d",
           447 => x"08",
           448 => x"04",
           449 => x"0c",
           450 => x"81",
           451 => x"83",
           452 => x"81",
           453 => x"81",
           454 => x"81",
           455 => x"83",
           456 => x"81",
           457 => x"81",
           458 => x"81",
           459 => x"83",
           460 => x"81",
           461 => x"81",
           462 => x"81",
           463 => x"83",
           464 => x"81",
           465 => x"81",
           466 => x"81",
           467 => x"83",
           468 => x"81",
           469 => x"81",
           470 => x"81",
           471 => x"83",
           472 => x"81",
           473 => x"81",
           474 => x"81",
           475 => x"83",
           476 => x"81",
           477 => x"81",
           478 => x"81",
           479 => x"83",
           480 => x"81",
           481 => x"81",
           482 => x"81",
           483 => x"83",
           484 => x"81",
           485 => x"81",
           486 => x"81",
           487 => x"83",
           488 => x"81",
           489 => x"81",
           490 => x"81",
           491 => x"83",
           492 => x"81",
           493 => x"81",
           494 => x"81",
           495 => x"83",
           496 => x"81",
           497 => x"81",
           498 => x"81",
           499 => x"83",
           500 => x"81",
           501 => x"81",
           502 => x"81",
           503 => x"83",
           504 => x"81",
           505 => x"81",
           506 => x"81",
           507 => x"83",
           508 => x"81",
           509 => x"81",
           510 => x"81",
           511 => x"83",
           512 => x"81",
           513 => x"81",
           514 => x"81",
           515 => x"83",
           516 => x"81",
           517 => x"81",
           518 => x"81",
           519 => x"83",
           520 => x"81",
           521 => x"81",
           522 => x"81",
           523 => x"83",
           524 => x"81",
           525 => x"81",
           526 => x"81",
           527 => x"83",
           528 => x"81",
           529 => x"81",
           530 => x"81",
           531 => x"83",
           532 => x"81",
           533 => x"81",
           534 => x"81",
           535 => x"83",
           536 => x"81",
           537 => x"81",
           538 => x"81",
           539 => x"83",
           540 => x"81",
           541 => x"81",
           542 => x"81",
           543 => x"83",
           544 => x"81",
           545 => x"81",
           546 => x"81",
           547 => x"83",
           548 => x"81",
           549 => x"81",
           550 => x"81",
           551 => x"83",
           552 => x"81",
           553 => x"81",
           554 => x"81",
           555 => x"83",
           556 => x"81",
           557 => x"81",
           558 => x"81",
           559 => x"83",
           560 => x"81",
           561 => x"80",
           562 => x"81",
           563 => x"83",
           564 => x"81",
           565 => x"80",
           566 => x"81",
           567 => x"83",
           568 => x"81",
           569 => x"80",
           570 => x"81",
           571 => x"83",
           572 => x"81",
           573 => x"9f",
           574 => x"fe",
           575 => x"80",
           576 => x"fe",
           577 => x"84",
           578 => x"fc",
           579 => x"90",
           580 => x"fc",
           581 => x"2d",
           582 => x"08",
           583 => x"04",
           584 => x"0c",
           585 => x"2d",
           586 => x"08",
           587 => x"04",
           588 => x"00",
           589 => x"10",
           590 => x"10",
           591 => x"10",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"53",
           597 => x"00",
           598 => x"06",
           599 => x"09",
           600 => x"05",
           601 => x"2b",
           602 => x"06",
           603 => x"04",
           604 => x"72",
           605 => x"05",
           606 => x"05",
           607 => x"72",
           608 => x"53",
           609 => x"51",
           610 => x"04",
           611 => x"70",
           612 => x"27",
           613 => x"71",
           614 => x"53",
           615 => x"0b",
           616 => x"8c",
           617 => x"e0",
           618 => x"81",
           619 => x"02",
           620 => x"0c",
           621 => x"80",
           622 => x"fc",
           623 => x"08",
           624 => x"fc",
           625 => x"08",
           626 => x"3f",
           627 => x"08",
           628 => x"f0",
           629 => x"3d",
           630 => x"fc",
           631 => x"fe",
           632 => x"81",
           633 => x"fd",
           634 => x"53",
           635 => x"08",
           636 => x"52",
           637 => x"08",
           638 => x"51",
           639 => x"81",
           640 => x"70",
           641 => x"0c",
           642 => x"0d",
           643 => x"0c",
           644 => x"fc",
           645 => x"fe",
           646 => x"3d",
           647 => x"81",
           648 => x"fc",
           649 => x"fe",
           650 => x"05",
           651 => x"b9",
           652 => x"fc",
           653 => x"08",
           654 => x"fc",
           655 => x"0c",
           656 => x"fe",
           657 => x"05",
           658 => x"fc",
           659 => x"08",
           660 => x"0b",
           661 => x"08",
           662 => x"81",
           663 => x"f4",
           664 => x"fe",
           665 => x"05",
           666 => x"fc",
           667 => x"08",
           668 => x"38",
           669 => x"08",
           670 => x"30",
           671 => x"08",
           672 => x"80",
           673 => x"fc",
           674 => x"0c",
           675 => x"08",
           676 => x"8a",
           677 => x"81",
           678 => x"f0",
           679 => x"fe",
           680 => x"05",
           681 => x"fc",
           682 => x"0c",
           683 => x"fe",
           684 => x"05",
           685 => x"fe",
           686 => x"05",
           687 => x"df",
           688 => x"f0",
           689 => x"fe",
           690 => x"05",
           691 => x"fe",
           692 => x"05",
           693 => x"90",
           694 => x"fc",
           695 => x"08",
           696 => x"fc",
           697 => x"0c",
           698 => x"08",
           699 => x"70",
           700 => x"0c",
           701 => x"0d",
           702 => x"0c",
           703 => x"fc",
           704 => x"fe",
           705 => x"3d",
           706 => x"81",
           707 => x"fc",
           708 => x"fe",
           709 => x"05",
           710 => x"99",
           711 => x"fc",
           712 => x"08",
           713 => x"fc",
           714 => x"0c",
           715 => x"fe",
           716 => x"05",
           717 => x"fc",
           718 => x"08",
           719 => x"38",
           720 => x"08",
           721 => x"30",
           722 => x"08",
           723 => x"81",
           724 => x"fc",
           725 => x"08",
           726 => x"fc",
           727 => x"08",
           728 => x"81",
           729 => x"70",
           730 => x"08",
           731 => x"54",
           732 => x"08",
           733 => x"80",
           734 => x"81",
           735 => x"f8",
           736 => x"81",
           737 => x"f8",
           738 => x"fe",
           739 => x"05",
           740 => x"fe",
           741 => x"87",
           742 => x"fe",
           743 => x"81",
           744 => x"02",
           745 => x"0c",
           746 => x"81",
           747 => x"fc",
           748 => x"0c",
           749 => x"fe",
           750 => x"05",
           751 => x"fc",
           752 => x"08",
           753 => x"08",
           754 => x"27",
           755 => x"fe",
           756 => x"05",
           757 => x"ae",
           758 => x"81",
           759 => x"8c",
           760 => x"a2",
           761 => x"fc",
           762 => x"08",
           763 => x"fc",
           764 => x"0c",
           765 => x"08",
           766 => x"10",
           767 => x"08",
           768 => x"ff",
           769 => x"fe",
           770 => x"05",
           771 => x"80",
           772 => x"fe",
           773 => x"05",
           774 => x"fc",
           775 => x"08",
           776 => x"81",
           777 => x"88",
           778 => x"fe",
           779 => x"05",
           780 => x"fe",
           781 => x"05",
           782 => x"fc",
           783 => x"08",
           784 => x"08",
           785 => x"07",
           786 => x"08",
           787 => x"81",
           788 => x"fc",
           789 => x"2a",
           790 => x"08",
           791 => x"81",
           792 => x"8c",
           793 => x"2a",
           794 => x"08",
           795 => x"ff",
           796 => x"fe",
           797 => x"05",
           798 => x"93",
           799 => x"fc",
           800 => x"08",
           801 => x"fc",
           802 => x"0c",
           803 => x"81",
           804 => x"f8",
           805 => x"81",
           806 => x"f4",
           807 => x"81",
           808 => x"f4",
           809 => x"fe",
           810 => x"3d",
           811 => x"fc",
           812 => x"3d",
           813 => x"79",
           814 => x"55",
           815 => x"27",
           816 => x"75",
           817 => x"51",
           818 => x"a9",
           819 => x"52",
           820 => x"98",
           821 => x"81",
           822 => x"74",
           823 => x"56",
           824 => x"52",
           825 => x"09",
           826 => x"38",
           827 => x"f0",
           828 => x"0d",
           829 => x"72",
           830 => x"54",
           831 => x"84",
           832 => x"72",
           833 => x"54",
           834 => x"84",
           835 => x"72",
           836 => x"54",
           837 => x"84",
           838 => x"72",
           839 => x"54",
           840 => x"84",
           841 => x"f0",
           842 => x"8f",
           843 => x"83",
           844 => x"38",
           845 => x"05",
           846 => x"70",
           847 => x"0c",
           848 => x"71",
           849 => x"38",
           850 => x"81",
           851 => x"0d",
           852 => x"02",
           853 => x"05",
           854 => x"53",
           855 => x"27",
           856 => x"83",
           857 => x"80",
           858 => x"ff",
           859 => x"ff",
           860 => x"73",
           861 => x"05",
           862 => x"12",
           863 => x"2e",
           864 => x"ef",
           865 => x"fe",
           866 => x"3d",
           867 => x"74",
           868 => x"07",
           869 => x"2b",
           870 => x"51",
           871 => x"a5",
           872 => x"70",
           873 => x"0c",
           874 => x"84",
           875 => x"72",
           876 => x"05",
           877 => x"71",
           878 => x"53",
           879 => x"52",
           880 => x"dd",
           881 => x"27",
           882 => x"71",
           883 => x"53",
           884 => x"52",
           885 => x"f2",
           886 => x"ff",
           887 => x"3d",
           888 => x"79",
           889 => x"83",
           890 => x"54",
           891 => x"c3",
           892 => x"08",
           893 => x"f7",
           894 => x"13",
           895 => x"84",
           896 => x"06",
           897 => x"53",
           898 => x"38",
           899 => x"74",
           900 => x"56",
           901 => x"70",
           902 => x"fb",
           903 => x"06",
           904 => x"82",
           905 => x"51",
           906 => x"54",
           907 => x"dc",
           908 => x"71",
           909 => x"53",
           910 => x"73",
           911 => x"55",
           912 => x"38",
           913 => x"f0",
           914 => x"0d",
           915 => x"0d",
           916 => x"83",
           917 => x"52",
           918 => x"71",
           919 => x"09",
           920 => x"ff",
           921 => x"f8",
           922 => x"80",
           923 => x"52",
           924 => x"38",
           925 => x"08",
           926 => x"fb",
           927 => x"06",
           928 => x"82",
           929 => x"51",
           930 => x"70",
           931 => x"38",
           932 => x"33",
           933 => x"2e",
           934 => x"12",
           935 => x"52",
           936 => x"71",
           937 => x"fe",
           938 => x"3d",
           939 => x"3d",
           940 => x"7c",
           941 => x"55",
           942 => x"2e",
           943 => x"71",
           944 => x"06",
           945 => x"2e",
           946 => x"ff",
           947 => x"ff",
           948 => x"71",
           949 => x"56",
           950 => x"2e",
           951 => x"a9",
           952 => x"2e",
           953 => x"70",
           954 => x"51",
           955 => x"80",
           956 => x"12",
           957 => x"15",
           958 => x"72",
           959 => x"81",
           960 => x"71",
           961 => x"56",
           962 => x"ff",
           963 => x"ff",
           964 => x"31",
           965 => x"70",
           966 => x"0c",
           967 => x"04",
           968 => x"55",
           969 => x"88",
           970 => x"74",
           971 => x"38",
           972 => x"52",
           973 => x"fc",
           974 => x"80",
           975 => x"74",
           976 => x"f7",
           977 => x"12",
           978 => x"84",
           979 => x"06",
           980 => x"70",
           981 => x"15",
           982 => x"55",
           983 => x"d0",
           984 => x"76",
           985 => x"38",
           986 => x"52",
           987 => x"80",
           988 => x"f0",
           989 => x"0d",
           990 => x"0d",
           991 => x"53",
           992 => x"52",
           993 => x"81",
           994 => x"81",
           995 => x"07",
           996 => x"52",
           997 => x"e8",
           998 => x"fe",
           999 => x"3d",
          1000 => x"3d",
          1001 => x"08",
          1002 => x"56",
          1003 => x"80",
          1004 => x"33",
          1005 => x"2e",
          1006 => x"86",
          1007 => x"52",
          1008 => x"53",
          1009 => x"13",
          1010 => x"33",
          1011 => x"06",
          1012 => x"70",
          1013 => x"38",
          1014 => x"80",
          1015 => x"74",
          1016 => x"81",
          1017 => x"70",
          1018 => x"81",
          1019 => x"80",
          1020 => x"05",
          1021 => x"76",
          1022 => x"70",
          1023 => x"0c",
          1024 => x"04",
          1025 => x"76",
          1026 => x"80",
          1027 => x"86",
          1028 => x"52",
          1029 => x"d8",
          1030 => x"f0",
          1031 => x"80",
          1032 => x"74",
          1033 => x"fe",
          1034 => x"3d",
          1035 => x"3d",
          1036 => x"11",
          1037 => x"52",
          1038 => x"70",
          1039 => x"98",
          1040 => x"33",
          1041 => x"82",
          1042 => x"26",
          1043 => x"84",
          1044 => x"83",
          1045 => x"26",
          1046 => x"85",
          1047 => x"84",
          1048 => x"26",
          1049 => x"86",
          1050 => x"85",
          1051 => x"26",
          1052 => x"88",
          1053 => x"86",
          1054 => x"e7",
          1055 => x"38",
          1056 => x"54",
          1057 => x"87",
          1058 => x"cc",
          1059 => x"87",
          1060 => x"0c",
          1061 => x"c0",
          1062 => x"82",
          1063 => x"c0",
          1064 => x"83",
          1065 => x"c0",
          1066 => x"84",
          1067 => x"c0",
          1068 => x"85",
          1069 => x"c0",
          1070 => x"86",
          1071 => x"c0",
          1072 => x"74",
          1073 => x"a4",
          1074 => x"c0",
          1075 => x"80",
          1076 => x"98",
          1077 => x"52",
          1078 => x"f0",
          1079 => x"0d",
          1080 => x"0d",
          1081 => x"c0",
          1082 => x"81",
          1083 => x"c0",
          1084 => x"5e",
          1085 => x"87",
          1086 => x"08",
          1087 => x"1c",
          1088 => x"98",
          1089 => x"79",
          1090 => x"87",
          1091 => x"08",
          1092 => x"1c",
          1093 => x"98",
          1094 => x"79",
          1095 => x"87",
          1096 => x"08",
          1097 => x"1c",
          1098 => x"98",
          1099 => x"7b",
          1100 => x"87",
          1101 => x"08",
          1102 => x"1c",
          1103 => x"0c",
          1104 => x"ff",
          1105 => x"83",
          1106 => x"58",
          1107 => x"57",
          1108 => x"56",
          1109 => x"55",
          1110 => x"54",
          1111 => x"53",
          1112 => x"ff",
          1113 => x"e2",
          1114 => x"9d",
          1115 => x"0d",
          1116 => x"0d",
          1117 => x"33",
          1118 => x"9f",
          1119 => x"52",
          1120 => x"81",
          1121 => x"83",
          1122 => x"fb",
          1123 => x"0b",
          1124 => x"e8",
          1125 => x"ff",
          1126 => x"56",
          1127 => x"84",
          1128 => x"2e",
          1129 => x"c0",
          1130 => x"70",
          1131 => x"2a",
          1132 => x"53",
          1133 => x"80",
          1134 => x"71",
          1135 => x"81",
          1136 => x"70",
          1137 => x"81",
          1138 => x"06",
          1139 => x"80",
          1140 => x"71",
          1141 => x"81",
          1142 => x"70",
          1143 => x"73",
          1144 => x"51",
          1145 => x"80",
          1146 => x"2e",
          1147 => x"c0",
          1148 => x"75",
          1149 => x"81",
          1150 => x"87",
          1151 => x"fb",
          1152 => x"9f",
          1153 => x"0b",
          1154 => x"33",
          1155 => x"06",
          1156 => x"87",
          1157 => x"51",
          1158 => x"86",
          1159 => x"94",
          1160 => x"08",
          1161 => x"70",
          1162 => x"54",
          1163 => x"2e",
          1164 => x"91",
          1165 => x"06",
          1166 => x"d7",
          1167 => x"32",
          1168 => x"51",
          1169 => x"2e",
          1170 => x"93",
          1171 => x"06",
          1172 => x"ff",
          1173 => x"81",
          1174 => x"87",
          1175 => x"52",
          1176 => x"86",
          1177 => x"94",
          1178 => x"72",
          1179 => x"0d",
          1180 => x"0d",
          1181 => x"74",
          1182 => x"ff",
          1183 => x"57",
          1184 => x"80",
          1185 => x"81",
          1186 => x"15",
          1187 => x"f9",
          1188 => x"81",
          1189 => x"57",
          1190 => x"c0",
          1191 => x"75",
          1192 => x"38",
          1193 => x"94",
          1194 => x"70",
          1195 => x"81",
          1196 => x"52",
          1197 => x"8c",
          1198 => x"2a",
          1199 => x"51",
          1200 => x"38",
          1201 => x"70",
          1202 => x"51",
          1203 => x"8d",
          1204 => x"2a",
          1205 => x"51",
          1206 => x"be",
          1207 => x"ff",
          1208 => x"c0",
          1209 => x"70",
          1210 => x"38",
          1211 => x"90",
          1212 => x"0c",
          1213 => x"33",
          1214 => x"06",
          1215 => x"70",
          1216 => x"76",
          1217 => x"0c",
          1218 => x"04",
          1219 => x"0b",
          1220 => x"e8",
          1221 => x"ff",
          1222 => x"87",
          1223 => x"51",
          1224 => x"86",
          1225 => x"94",
          1226 => x"08",
          1227 => x"70",
          1228 => x"51",
          1229 => x"2e",
          1230 => x"81",
          1231 => x"87",
          1232 => x"52",
          1233 => x"86",
          1234 => x"94",
          1235 => x"08",
          1236 => x"06",
          1237 => x"0c",
          1238 => x"0d",
          1239 => x"0d",
          1240 => x"f9",
          1241 => x"81",
          1242 => x"53",
          1243 => x"84",
          1244 => x"2e",
          1245 => x"c0",
          1246 => x"71",
          1247 => x"2a",
          1248 => x"51",
          1249 => x"52",
          1250 => x"a0",
          1251 => x"ff",
          1252 => x"c0",
          1253 => x"70",
          1254 => x"38",
          1255 => x"90",
          1256 => x"70",
          1257 => x"98",
          1258 => x"51",
          1259 => x"f0",
          1260 => x"0d",
          1261 => x"0d",
          1262 => x"80",
          1263 => x"2a",
          1264 => x"51",
          1265 => x"84",
          1266 => x"c0",
          1267 => x"81",
          1268 => x"87",
          1269 => x"08",
          1270 => x"0c",
          1271 => x"94",
          1272 => x"f4",
          1273 => x"9e",
          1274 => x"f9",
          1275 => x"c0",
          1276 => x"81",
          1277 => x"87",
          1278 => x"08",
          1279 => x"0c",
          1280 => x"ac",
          1281 => x"84",
          1282 => x"9e",
          1283 => x"fa",
          1284 => x"c0",
          1285 => x"81",
          1286 => x"87",
          1287 => x"08",
          1288 => x"0c",
          1289 => x"bc",
          1290 => x"94",
          1291 => x"9e",
          1292 => x"fa",
          1293 => x"c0",
          1294 => x"81",
          1295 => x"87",
          1296 => x"08",
          1297 => x"fa",
          1298 => x"c0",
          1299 => x"81",
          1300 => x"87",
          1301 => x"08",
          1302 => x"0c",
          1303 => x"8c",
          1304 => x"ac",
          1305 => x"81",
          1306 => x"80",
          1307 => x"9e",
          1308 => x"84",
          1309 => x"51",
          1310 => x"80",
          1311 => x"81",
          1312 => x"fa",
          1313 => x"0b",
          1314 => x"90",
          1315 => x"80",
          1316 => x"52",
          1317 => x"2e",
          1318 => x"52",
          1319 => x"b2",
          1320 => x"87",
          1321 => x"08",
          1322 => x"0a",
          1323 => x"52",
          1324 => x"83",
          1325 => x"71",
          1326 => x"34",
          1327 => x"c0",
          1328 => x"70",
          1329 => x"06",
          1330 => x"70",
          1331 => x"38",
          1332 => x"81",
          1333 => x"80",
          1334 => x"9e",
          1335 => x"a0",
          1336 => x"51",
          1337 => x"80",
          1338 => x"81",
          1339 => x"fa",
          1340 => x"0b",
          1341 => x"90",
          1342 => x"80",
          1343 => x"52",
          1344 => x"2e",
          1345 => x"52",
          1346 => x"b6",
          1347 => x"87",
          1348 => x"08",
          1349 => x"80",
          1350 => x"52",
          1351 => x"83",
          1352 => x"71",
          1353 => x"34",
          1354 => x"c0",
          1355 => x"70",
          1356 => x"06",
          1357 => x"70",
          1358 => x"38",
          1359 => x"81",
          1360 => x"80",
          1361 => x"9e",
          1362 => x"81",
          1363 => x"51",
          1364 => x"80",
          1365 => x"81",
          1366 => x"fa",
          1367 => x"0b",
          1368 => x"90",
          1369 => x"c0",
          1370 => x"52",
          1371 => x"2e",
          1372 => x"52",
          1373 => x"ba",
          1374 => x"87",
          1375 => x"08",
          1376 => x"06",
          1377 => x"70",
          1378 => x"38",
          1379 => x"81",
          1380 => x"87",
          1381 => x"08",
          1382 => x"06",
          1383 => x"51",
          1384 => x"81",
          1385 => x"80",
          1386 => x"9e",
          1387 => x"84",
          1388 => x"52",
          1389 => x"2e",
          1390 => x"52",
          1391 => x"bd",
          1392 => x"9e",
          1393 => x"83",
          1394 => x"84",
          1395 => x"51",
          1396 => x"be",
          1397 => x"87",
          1398 => x"08",
          1399 => x"51",
          1400 => x"80",
          1401 => x"81",
          1402 => x"fa",
          1403 => x"c0",
          1404 => x"70",
          1405 => x"51",
          1406 => x"c0",
          1407 => x"0d",
          1408 => x"0d",
          1409 => x"51",
          1410 => x"81",
          1411 => x"54",
          1412 => x"88",
          1413 => x"80",
          1414 => x"3f",
          1415 => x"51",
          1416 => x"81",
          1417 => x"54",
          1418 => x"93",
          1419 => x"8c",
          1420 => x"90",
          1421 => x"52",
          1422 => x"51",
          1423 => x"81",
          1424 => x"54",
          1425 => x"93",
          1426 => x"84",
          1427 => x"88",
          1428 => x"52",
          1429 => x"51",
          1430 => x"81",
          1431 => x"54",
          1432 => x"93",
          1433 => x"ec",
          1434 => x"f0",
          1435 => x"52",
          1436 => x"51",
          1437 => x"81",
          1438 => x"54",
          1439 => x"93",
          1440 => x"f4",
          1441 => x"f8",
          1442 => x"52",
          1443 => x"51",
          1444 => x"81",
          1445 => x"54",
          1446 => x"93",
          1447 => x"fc",
          1448 => x"80",
          1449 => x"52",
          1450 => x"51",
          1451 => x"81",
          1452 => x"54",
          1453 => x"8d",
          1454 => x"bc",
          1455 => x"e4",
          1456 => x"c5",
          1457 => x"bf",
          1458 => x"80",
          1459 => x"81",
          1460 => x"52",
          1461 => x"51",
          1462 => x"81",
          1463 => x"54",
          1464 => x"8d",
          1465 => x"be",
          1466 => x"e4",
          1467 => x"99",
          1468 => x"b1",
          1469 => x"80",
          1470 => x"81",
          1471 => x"88",
          1472 => x"fa",
          1473 => x"73",
          1474 => x"38",
          1475 => x"51",
          1476 => x"81",
          1477 => x"54",
          1478 => x"88",
          1479 => x"b8",
          1480 => x"3f",
          1481 => x"33",
          1482 => x"2e",
          1483 => x"e5",
          1484 => x"f1",
          1485 => x"ba",
          1486 => x"80",
          1487 => x"81",
          1488 => x"87",
          1489 => x"e5",
          1490 => x"d9",
          1491 => x"94",
          1492 => x"e5",
          1493 => x"b1",
          1494 => x"98",
          1495 => x"e6",
          1496 => x"a5",
          1497 => x"9c",
          1498 => x"e6",
          1499 => x"99",
          1500 => x"e0",
          1501 => x"3f",
          1502 => x"22",
          1503 => x"e8",
          1504 => x"3f",
          1505 => x"08",
          1506 => x"c0",
          1507 => x"e4",
          1508 => x"fe",
          1509 => x"84",
          1510 => x"71",
          1511 => x"81",
          1512 => x"52",
          1513 => x"51",
          1514 => x"81",
          1515 => x"54",
          1516 => x"a8",
          1517 => x"a8",
          1518 => x"84",
          1519 => x"51",
          1520 => x"81",
          1521 => x"bd",
          1522 => x"76",
          1523 => x"54",
          1524 => x"08",
          1525 => x"bc",
          1526 => x"3f",
          1527 => x"33",
          1528 => x"2e",
          1529 => x"fa",
          1530 => x"bd",
          1531 => x"75",
          1532 => x"3f",
          1533 => x"08",
          1534 => x"29",
          1535 => x"54",
          1536 => x"f0",
          1537 => x"e7",
          1538 => x"fd",
          1539 => x"e4",
          1540 => x"3f",
          1541 => x"04",
          1542 => x"02",
          1543 => x"ff",
          1544 => x"84",
          1545 => x"71",
          1546 => x"e1",
          1547 => x"71",
          1548 => x"e8",
          1549 => x"39",
          1550 => x"51",
          1551 => x"e8",
          1552 => x"39",
          1553 => x"51",
          1554 => x"e8",
          1555 => x"39",
          1556 => x"51",
          1557 => x"84",
          1558 => x"71",
          1559 => x"04",
          1560 => x"87",
          1561 => x"70",
          1562 => x"80",
          1563 => x"74",
          1564 => x"fa",
          1565 => x"0c",
          1566 => x"04",
          1567 => x"87",
          1568 => x"70",
          1569 => x"c4",
          1570 => x"72",
          1571 => x"70",
          1572 => x"08",
          1573 => x"fa",
          1574 => x"0c",
          1575 => x"0d",
          1576 => x"87",
          1577 => x"0c",
          1578 => x"c4",
          1579 => x"96",
          1580 => x"fe",
          1581 => x"ff",
          1582 => x"38",
          1583 => x"0b",
          1584 => x"0c",
          1585 => x"08",
          1586 => x"52",
          1587 => x"83",
          1588 => x"88",
          1589 => x"ff",
          1590 => x"53",
          1591 => x"f0",
          1592 => x"0d",
          1593 => x"0d",
          1594 => x"12",
          1595 => x"90",
          1596 => x"15",
          1597 => x"5e",
          1598 => x"59",
          1599 => x"77",
          1600 => x"75",
          1601 => x"08",
          1602 => x"71",
          1603 => x"31",
          1604 => x"80",
          1605 => x"84",
          1606 => x"8c",
          1607 => x"88",
          1608 => x"8c",
          1609 => x"88",
          1610 => x"90",
          1611 => x"94",
          1612 => x"94",
          1613 => x"90",
          1614 => x"39",
          1615 => x"73",
          1616 => x"74",
          1617 => x"77",
          1618 => x"0c",
          1619 => x"04",
          1620 => x"76",
          1621 => x"88",
          1622 => x"53",
          1623 => x"81",
          1624 => x"06",
          1625 => x"12",
          1626 => x"52",
          1627 => x"2e",
          1628 => x"94",
          1629 => x"08",
          1630 => x"0c",
          1631 => x"0c",
          1632 => x"0c",
          1633 => x"39",
          1634 => x"81",
          1635 => x"90",
          1636 => x"fa",
          1637 => x"14",
          1638 => x"fa",
          1639 => x"13",
          1640 => x"12",
          1641 => x"08",
          1642 => x"81",
          1643 => x"84",
          1644 => x"14",
          1645 => x"74",
          1646 => x"06",
          1647 => x"14",
          1648 => x"14",
          1649 => x"08",
          1650 => x"70",
          1651 => x"52",
          1652 => x"8c",
          1653 => x"15",
          1654 => x"13",
          1655 => x"12",
          1656 => x"fe",
          1657 => x"3d",
          1658 => x"3d",
          1659 => x"55",
          1660 => x"2e",
          1661 => x"9f",
          1662 => x"81",
          1663 => x"57",
          1664 => x"82",
          1665 => x"84",
          1666 => x"27",
          1667 => x"90",
          1668 => x"ed",
          1669 => x"ff",
          1670 => x"80",
          1671 => x"58",
          1672 => x"81",
          1673 => x"81",
          1674 => x"30",
          1675 => x"f0",
          1676 => x"25",
          1677 => x"08",
          1678 => x"70",
          1679 => x"25",
          1680 => x"58",
          1681 => x"56",
          1682 => x"74",
          1683 => x"06",
          1684 => x"88",
          1685 => x"75",
          1686 => x"39",
          1687 => x"fe",
          1688 => x"77",
          1689 => x"08",
          1690 => x"81",
          1691 => x"53",
          1692 => x"2e",
          1693 => x"73",
          1694 => x"8c",
          1695 => x"f0",
          1696 => x"08",
          1697 => x"72",
          1698 => x"75",
          1699 => x"88",
          1700 => x"8c",
          1701 => x"75",
          1702 => x"3f",
          1703 => x"fe",
          1704 => x"fc",
          1705 => x"fe",
          1706 => x"73",
          1707 => x"0c",
          1708 => x"04",
          1709 => x"73",
          1710 => x"2e",
          1711 => x"12",
          1712 => x"3f",
          1713 => x"04",
          1714 => x"02",
          1715 => x"53",
          1716 => x"09",
          1717 => x"38",
          1718 => x"3f",
          1719 => x"08",
          1720 => x"2e",
          1721 => x"72",
          1722 => x"8c",
          1723 => x"81",
          1724 => x"8f",
          1725 => x"84",
          1726 => x"80",
          1727 => x"72",
          1728 => x"84",
          1729 => x"fe",
          1730 => x"97",
          1731 => x"ff",
          1732 => x"81",
          1733 => x"54",
          1734 => x"3f",
          1735 => x"84",
          1736 => x"0d",
          1737 => x"0d",
          1738 => x"33",
          1739 => x"06",
          1740 => x"80",
          1741 => x"72",
          1742 => x"51",
          1743 => x"ff",
          1744 => x"39",
          1745 => x"04",
          1746 => x"77",
          1747 => x"08",
          1748 => x"84",
          1749 => x"73",
          1750 => x"ff",
          1751 => x"71",
          1752 => x"38",
          1753 => x"06",
          1754 => x"54",
          1755 => x"e7",
          1756 => x"ff",
          1757 => x"3d",
          1758 => x"3d",
          1759 => x"59",
          1760 => x"81",
          1761 => x"56",
          1762 => x"84",
          1763 => x"a5",
          1764 => x"06",
          1765 => x"80",
          1766 => x"81",
          1767 => x"58",
          1768 => x"b0",
          1769 => x"06",
          1770 => x"5a",
          1771 => x"ad",
          1772 => x"06",
          1773 => x"5a",
          1774 => x"05",
          1775 => x"75",
          1776 => x"81",
          1777 => x"77",
          1778 => x"08",
          1779 => x"05",
          1780 => x"5d",
          1781 => x"39",
          1782 => x"72",
          1783 => x"38",
          1784 => x"7b",
          1785 => x"05",
          1786 => x"70",
          1787 => x"33",
          1788 => x"39",
          1789 => x"32",
          1790 => x"72",
          1791 => x"78",
          1792 => x"70",
          1793 => x"07",
          1794 => x"07",
          1795 => x"51",
          1796 => x"80",
          1797 => x"79",
          1798 => x"70",
          1799 => x"33",
          1800 => x"80",
          1801 => x"38",
          1802 => x"e0",
          1803 => x"38",
          1804 => x"81",
          1805 => x"53",
          1806 => x"2e",
          1807 => x"73",
          1808 => x"a2",
          1809 => x"c3",
          1810 => x"38",
          1811 => x"24",
          1812 => x"80",
          1813 => x"8c",
          1814 => x"39",
          1815 => x"2e",
          1816 => x"81",
          1817 => x"80",
          1818 => x"80",
          1819 => x"d5",
          1820 => x"73",
          1821 => x"8e",
          1822 => x"39",
          1823 => x"2e",
          1824 => x"80",
          1825 => x"84",
          1826 => x"56",
          1827 => x"74",
          1828 => x"72",
          1829 => x"38",
          1830 => x"15",
          1831 => x"54",
          1832 => x"38",
          1833 => x"56",
          1834 => x"81",
          1835 => x"72",
          1836 => x"38",
          1837 => x"90",
          1838 => x"06",
          1839 => x"2e",
          1840 => x"51",
          1841 => x"74",
          1842 => x"53",
          1843 => x"fd",
          1844 => x"51",
          1845 => x"ef",
          1846 => x"19",
          1847 => x"53",
          1848 => x"39",
          1849 => x"39",
          1850 => x"39",
          1851 => x"39",
          1852 => x"39",
          1853 => x"d0",
          1854 => x"39",
          1855 => x"70",
          1856 => x"53",
          1857 => x"88",
          1858 => x"19",
          1859 => x"39",
          1860 => x"54",
          1861 => x"74",
          1862 => x"70",
          1863 => x"07",
          1864 => x"55",
          1865 => x"80",
          1866 => x"72",
          1867 => x"38",
          1868 => x"90",
          1869 => x"80",
          1870 => x"5e",
          1871 => x"74",
          1872 => x"3f",
          1873 => x"08",
          1874 => x"7c",
          1875 => x"54",
          1876 => x"81",
          1877 => x"55",
          1878 => x"92",
          1879 => x"53",
          1880 => x"2e",
          1881 => x"14",
          1882 => x"ff",
          1883 => x"14",
          1884 => x"70",
          1885 => x"34",
          1886 => x"30",
          1887 => x"9f",
          1888 => x"57",
          1889 => x"85",
          1890 => x"b1",
          1891 => x"2a",
          1892 => x"51",
          1893 => x"2e",
          1894 => x"3d",
          1895 => x"05",
          1896 => x"34",
          1897 => x"76",
          1898 => x"54",
          1899 => x"72",
          1900 => x"54",
          1901 => x"70",
          1902 => x"56",
          1903 => x"81",
          1904 => x"7b",
          1905 => x"73",
          1906 => x"3f",
          1907 => x"53",
          1908 => x"74",
          1909 => x"53",
          1910 => x"eb",
          1911 => x"77",
          1912 => x"53",
          1913 => x"14",
          1914 => x"54",
          1915 => x"3f",
          1916 => x"74",
          1917 => x"53",
          1918 => x"fb",
          1919 => x"51",
          1920 => x"ef",
          1921 => x"0d",
          1922 => x"0d",
          1923 => x"70",
          1924 => x"08",
          1925 => x"51",
          1926 => x"85",
          1927 => x"fe",
          1928 => x"81",
          1929 => x"85",
          1930 => x"52",
          1931 => x"ca",
          1932 => x"8c",
          1933 => x"73",
          1934 => x"81",
          1935 => x"84",
          1936 => x"fd",
          1937 => x"ff",
          1938 => x"81",
          1939 => x"87",
          1940 => x"53",
          1941 => x"fa",
          1942 => x"81",
          1943 => x"85",
          1944 => x"fb",
          1945 => x"79",
          1946 => x"08",
          1947 => x"57",
          1948 => x"71",
          1949 => x"e0",
          1950 => x"88",
          1951 => x"2d",
          1952 => x"08",
          1953 => x"53",
          1954 => x"80",
          1955 => x"8d",
          1956 => x"72",
          1957 => x"30",
          1958 => x"51",
          1959 => x"80",
          1960 => x"71",
          1961 => x"38",
          1962 => x"97",
          1963 => x"25",
          1964 => x"16",
          1965 => x"25",
          1966 => x"14",
          1967 => x"34",
          1968 => x"72",
          1969 => x"3f",
          1970 => x"73",
          1971 => x"72",
          1972 => x"f7",
          1973 => x"53",
          1974 => x"f0",
          1975 => x"0d",
          1976 => x"0d",
          1977 => x"08",
          1978 => x"88",
          1979 => x"76",
          1980 => x"ef",
          1981 => x"ff",
          1982 => x"3d",
          1983 => x"3d",
          1984 => x"5a",
          1985 => x"7a",
          1986 => x"08",
          1987 => x"53",
          1988 => x"09",
          1989 => x"38",
          1990 => x"0c",
          1991 => x"ad",
          1992 => x"06",
          1993 => x"76",
          1994 => x"0c",
          1995 => x"33",
          1996 => x"73",
          1997 => x"81",
          1998 => x"38",
          1999 => x"05",
          2000 => x"08",
          2001 => x"53",
          2002 => x"2e",
          2003 => x"57",
          2004 => x"2e",
          2005 => x"39",
          2006 => x"13",
          2007 => x"08",
          2008 => x"53",
          2009 => x"55",
          2010 => x"80",
          2011 => x"14",
          2012 => x"88",
          2013 => x"27",
          2014 => x"eb",
          2015 => x"53",
          2016 => x"89",
          2017 => x"38",
          2018 => x"55",
          2019 => x"8a",
          2020 => x"a0",
          2021 => x"c2",
          2022 => x"74",
          2023 => x"e0",
          2024 => x"ff",
          2025 => x"d0",
          2026 => x"ff",
          2027 => x"90",
          2028 => x"38",
          2029 => x"81",
          2030 => x"53",
          2031 => x"ca",
          2032 => x"27",
          2033 => x"77",
          2034 => x"08",
          2035 => x"0c",
          2036 => x"33",
          2037 => x"ff",
          2038 => x"80",
          2039 => x"74",
          2040 => x"79",
          2041 => x"74",
          2042 => x"0c",
          2043 => x"04",
          2044 => x"7a",
          2045 => x"80",
          2046 => x"58",
          2047 => x"33",
          2048 => x"a0",
          2049 => x"06",
          2050 => x"13",
          2051 => x"39",
          2052 => x"09",
          2053 => x"38",
          2054 => x"11",
          2055 => x"08",
          2056 => x"54",
          2057 => x"2e",
          2058 => x"80",
          2059 => x"08",
          2060 => x"0c",
          2061 => x"33",
          2062 => x"80",
          2063 => x"38",
          2064 => x"80",
          2065 => x"38",
          2066 => x"57",
          2067 => x"0c",
          2068 => x"33",
          2069 => x"39",
          2070 => x"74",
          2071 => x"38",
          2072 => x"80",
          2073 => x"89",
          2074 => x"38",
          2075 => x"d0",
          2076 => x"55",
          2077 => x"80",
          2078 => x"39",
          2079 => x"d9",
          2080 => x"80",
          2081 => x"27",
          2082 => x"80",
          2083 => x"89",
          2084 => x"70",
          2085 => x"55",
          2086 => x"70",
          2087 => x"55",
          2088 => x"27",
          2089 => x"14",
          2090 => x"06",
          2091 => x"74",
          2092 => x"73",
          2093 => x"38",
          2094 => x"14",
          2095 => x"05",
          2096 => x"08",
          2097 => x"54",
          2098 => x"39",
          2099 => x"84",
          2100 => x"55",
          2101 => x"81",
          2102 => x"fe",
          2103 => x"3d",
          2104 => x"3d",
          2105 => x"2b",
          2106 => x"79",
          2107 => x"98",
          2108 => x"13",
          2109 => x"51",
          2110 => x"51",
          2111 => x"81",
          2112 => x"33",
          2113 => x"74",
          2114 => x"81",
          2115 => x"08",
          2116 => x"05",
          2117 => x"71",
          2118 => x"52",
          2119 => x"09",
          2120 => x"38",
          2121 => x"81",
          2122 => x"85",
          2123 => x"fc",
          2124 => x"02",
          2125 => x"05",
          2126 => x"54",
          2127 => x"80",
          2128 => x"88",
          2129 => x"3f",
          2130 => x"fc",
          2131 => x"f2",
          2132 => x"33",
          2133 => x"71",
          2134 => x"81",
          2135 => x"de",
          2136 => x"f3",
          2137 => x"73",
          2138 => x"0d",
          2139 => x"0d",
          2140 => x"05",
          2141 => x"02",
          2142 => x"05",
          2143 => x"bc",
          2144 => x"29",
          2145 => x"05",
          2146 => x"59",
          2147 => x"59",
          2148 => x"86",
          2149 => x"f2",
          2150 => x"fb",
          2151 => x"84",
          2152 => x"e4",
          2153 => x"70",
          2154 => x"5a",
          2155 => x"81",
          2156 => x"75",
          2157 => x"bc",
          2158 => x"29",
          2159 => x"05",
          2160 => x"56",
          2161 => x"2e",
          2162 => x"53",
          2163 => x"51",
          2164 => x"81",
          2165 => x"81",
          2166 => x"81",
          2167 => x"74",
          2168 => x"55",
          2169 => x"87",
          2170 => x"81",
          2171 => x"77",
          2172 => x"38",
          2173 => x"08",
          2174 => x"2e",
          2175 => x"fb",
          2176 => x"74",
          2177 => x"3d",
          2178 => x"76",
          2179 => x"75",
          2180 => x"91",
          2181 => x"b8",
          2182 => x"51",
          2183 => x"3f",
          2184 => x"08",
          2185 => x"ee",
          2186 => x"0d",
          2187 => x"0d",
          2188 => x"52",
          2189 => x"08",
          2190 => x"87",
          2191 => x"f0",
          2192 => x"38",
          2193 => x"08",
          2194 => x"52",
          2195 => x"52",
          2196 => x"d5",
          2197 => x"f0",
          2198 => x"b8",
          2199 => x"d7",
          2200 => x"fe",
          2201 => x"80",
          2202 => x"f0",
          2203 => x"38",
          2204 => x"08",
          2205 => x"17",
          2206 => x"74",
          2207 => x"76",
          2208 => x"81",
          2209 => x"57",
          2210 => x"74",
          2211 => x"81",
          2212 => x"38",
          2213 => x"04",
          2214 => x"aa",
          2215 => x"3d",
          2216 => x"81",
          2217 => x"80",
          2218 => x"b8",
          2219 => x"d1",
          2220 => x"fe",
          2221 => x"91",
          2222 => x"81",
          2223 => x"54",
          2224 => x"52",
          2225 => x"52",
          2226 => x"dd",
          2227 => x"f0",
          2228 => x"a4",
          2229 => x"d6",
          2230 => x"fe",
          2231 => x"18",
          2232 => x"0b",
          2233 => x"08",
          2234 => x"81",
          2235 => x"ff",
          2236 => x"55",
          2237 => x"34",
          2238 => x"30",
          2239 => x"9f",
          2240 => x"55",
          2241 => x"85",
          2242 => x"ad",
          2243 => x"b8",
          2244 => x"08",
          2245 => x"d0",
          2246 => x"fe",
          2247 => x"2e",
          2248 => x"e8",
          2249 => x"fd",
          2250 => x"2e",
          2251 => x"99",
          2252 => x"79",
          2253 => x"3f",
          2254 => x"91",
          2255 => x"08",
          2256 => x"f0",
          2257 => x"80",
          2258 => x"fe",
          2259 => x"3d",
          2260 => x"3d",
          2261 => x"71",
          2262 => x"33",
          2263 => x"58",
          2264 => x"09",
          2265 => x"38",
          2266 => x"05",
          2267 => x"27",
          2268 => x"17",
          2269 => x"71",
          2270 => x"55",
          2271 => x"09",
          2272 => x"38",
          2273 => x"ea",
          2274 => x"73",
          2275 => x"fb",
          2276 => x"08",
          2277 => x"b5",
          2278 => x"f0",
          2279 => x"52",
          2280 => x"d6",
          2281 => x"fe",
          2282 => x"c4",
          2283 => x"33",
          2284 => x"2e",
          2285 => x"82",
          2286 => x"b4",
          2287 => x"3f",
          2288 => x"1a",
          2289 => x"fc",
          2290 => x"05",
          2291 => x"3f",
          2292 => x"08",
          2293 => x"38",
          2294 => x"52",
          2295 => x"b8",
          2296 => x"f0",
          2297 => x"06",
          2298 => x"38",
          2299 => x"39",
          2300 => x"81",
          2301 => x"54",
          2302 => x"ff",
          2303 => x"54",
          2304 => x"f0",
          2305 => x"0d",
          2306 => x"0d",
          2307 => x"02",
          2308 => x"c3",
          2309 => x"5a",
          2310 => x"3d",
          2311 => x"bc",
          2312 => x"fb",
          2313 => x"a3",
          2314 => x"b4",
          2315 => x"81",
          2316 => x"51",
          2317 => x"81",
          2318 => x"81",
          2319 => x"81",
          2320 => x"80",
          2321 => x"38",
          2322 => x"fa",
          2323 => x"81",
          2324 => x"51",
          2325 => x"81",
          2326 => x"80",
          2327 => x"81",
          2328 => x"f3",
          2329 => x"e3",
          2330 => x"b8",
          2331 => x"f8",
          2332 => x"70",
          2333 => x"f6",
          2334 => x"fe",
          2335 => x"81",
          2336 => x"74",
          2337 => x"06",
          2338 => x"81",
          2339 => x"51",
          2340 => x"81",
          2341 => x"55",
          2342 => x"fe",
          2343 => x"9a",
          2344 => x"f0",
          2345 => x"70",
          2346 => x"80",
          2347 => x"53",
          2348 => x"06",
          2349 => x"f9",
          2350 => x"ff",
          2351 => x"06",
          2352 => x"87",
          2353 => x"81",
          2354 => x"8f",
          2355 => x"8d",
          2356 => x"f0",
          2357 => x"70",
          2358 => x"59",
          2359 => x"ee",
          2360 => x"ff",
          2361 => x"94",
          2362 => x"2b",
          2363 => x"81",
          2364 => x"70",
          2365 => x"97",
          2366 => x"2c",
          2367 => x"29",
          2368 => x"05",
          2369 => x"70",
          2370 => x"51",
          2371 => x"51",
          2372 => x"81",
          2373 => x"2e",
          2374 => x"77",
          2375 => x"38",
          2376 => x"0a",
          2377 => x"0a",
          2378 => x"2c",
          2379 => x"75",
          2380 => x"38",
          2381 => x"52",
          2382 => x"a6",
          2383 => x"f0",
          2384 => x"06",
          2385 => x"2e",
          2386 => x"81",
          2387 => x"81",
          2388 => x"74",
          2389 => x"29",
          2390 => x"05",
          2391 => x"70",
          2392 => x"56",
          2393 => x"8a",
          2394 => x"76",
          2395 => x"77",
          2396 => x"3f",
          2397 => x"08",
          2398 => x"54",
          2399 => x"d3",
          2400 => x"75",
          2401 => x"ca",
          2402 => x"55",
          2403 => x"94",
          2404 => x"2b",
          2405 => x"81",
          2406 => x"70",
          2407 => x"98",
          2408 => x"11",
          2409 => x"81",
          2410 => x"33",
          2411 => x"51",
          2412 => x"55",
          2413 => x"09",
          2414 => x"92",
          2415 => x"d0",
          2416 => x"0c",
          2417 => x"ff",
          2418 => x"0b",
          2419 => x"34",
          2420 => x"81",
          2421 => x"75",
          2422 => x"34",
          2423 => x"34",
          2424 => x"7e",
          2425 => x"26",
          2426 => x"73",
          2427 => x"e1",
          2428 => x"73",
          2429 => x"ff",
          2430 => x"73",
          2431 => x"cb",
          2432 => x"98",
          2433 => x"75",
          2434 => x"74",
          2435 => x"98",
          2436 => x"73",
          2437 => x"38",
          2438 => x"73",
          2439 => x"34",
          2440 => x"0a",
          2441 => x"0a",
          2442 => x"2c",
          2443 => x"33",
          2444 => x"df",
          2445 => x"9c",
          2446 => x"56",
          2447 => x"ff",
          2448 => x"1a",
          2449 => x"33",
          2450 => x"ff",
          2451 => x"73",
          2452 => x"38",
          2453 => x"73",
          2454 => x"34",
          2455 => x"33",
          2456 => x"0a",
          2457 => x"0a",
          2458 => x"2c",
          2459 => x"33",
          2460 => x"56",
          2461 => x"a2",
          2462 => x"70",
          2463 => x"e8",
          2464 => x"81",
          2465 => x"81",
          2466 => x"70",
          2467 => x"ff",
          2468 => x"51",
          2469 => x"24",
          2470 => x"ff",
          2471 => x"98",
          2472 => x"2c",
          2473 => x"33",
          2474 => x"56",
          2475 => x"fc",
          2476 => x"51",
          2477 => x"74",
          2478 => x"29",
          2479 => x"05",
          2480 => x"81",
          2481 => x"56",
          2482 => x"75",
          2483 => x"fb",
          2484 => x"ff",
          2485 => x"81",
          2486 => x"55",
          2487 => x"fb",
          2488 => x"ff",
          2489 => x"05",
          2490 => x"ff",
          2491 => x"15",
          2492 => x"ff",
          2493 => x"51",
          2494 => x"81",
          2495 => x"70",
          2496 => x"98",
          2497 => x"98",
          2498 => x"56",
          2499 => x"25",
          2500 => x"1a",
          2501 => x"33",
          2502 => x"33",
          2503 => x"3f",
          2504 => x"0a",
          2505 => x"0a",
          2506 => x"2c",
          2507 => x"33",
          2508 => x"75",
          2509 => x"38",
          2510 => x"8c",
          2511 => x"9c",
          2512 => x"2b",
          2513 => x"81",
          2514 => x"57",
          2515 => x"74",
          2516 => x"f7",
          2517 => x"e6",
          2518 => x"81",
          2519 => x"81",
          2520 => x"70",
          2521 => x"ff",
          2522 => x"51",
          2523 => x"25",
          2524 => x"d7",
          2525 => x"98",
          2526 => x"54",
          2527 => x"8a",
          2528 => x"3f",
          2529 => x"52",
          2530 => x"c6",
          2531 => x"f0",
          2532 => x"06",
          2533 => x"38",
          2534 => x"33",
          2535 => x"2e",
          2536 => x"81",
          2537 => x"79",
          2538 => x"3f",
          2539 => x"80",
          2540 => x"b7",
          2541 => x"9c",
          2542 => x"80",
          2543 => x"38",
          2544 => x"84",
          2545 => x"9c",
          2546 => x"54",
          2547 => x"9c",
          2548 => x"ff",
          2549 => x"39",
          2550 => x"33",
          2551 => x"33",
          2552 => x"75",
          2553 => x"38",
          2554 => x"73",
          2555 => x"34",
          2556 => x"70",
          2557 => x"81",
          2558 => x"51",
          2559 => x"25",
          2560 => x"1a",
          2561 => x"33",
          2562 => x"33",
          2563 => x"3f",
          2564 => x"0a",
          2565 => x"0a",
          2566 => x"2c",
          2567 => x"33",
          2568 => x"75",
          2569 => x"38",
          2570 => x"9c",
          2571 => x"9c",
          2572 => x"2b",
          2573 => x"81",
          2574 => x"57",
          2575 => x"74",
          2576 => x"87",
          2577 => x"e4",
          2578 => x"81",
          2579 => x"81",
          2580 => x"70",
          2581 => x"ff",
          2582 => x"51",
          2583 => x"25",
          2584 => x"e7",
          2585 => x"9c",
          2586 => x"ff",
          2587 => x"98",
          2588 => x"54",
          2589 => x"f8",
          2590 => x"14",
          2591 => x"ff",
          2592 => x"1a",
          2593 => x"54",
          2594 => x"81",
          2595 => x"70",
          2596 => x"81",
          2597 => x"58",
          2598 => x"75",
          2599 => x"f8",
          2600 => x"ae",
          2601 => x"b0",
          2602 => x"80",
          2603 => x"74",
          2604 => x"3f",
          2605 => x"08",
          2606 => x"34",
          2607 => x"08",
          2608 => x"81",
          2609 => x"52",
          2610 => x"e6",
          2611 => x"81",
          2612 => x"84",
          2613 => x"e4",
          2614 => x"08",
          2615 => x"80",
          2616 => x"74",
          2617 => x"3f",
          2618 => x"08",
          2619 => x"34",
          2620 => x"08",
          2621 => x"81",
          2622 => x"52",
          2623 => x"b2",
          2624 => x"54",
          2625 => x"73",
          2626 => x"80",
          2627 => x"38",
          2628 => x"b9",
          2629 => x"39",
          2630 => x"09",
          2631 => x"38",
          2632 => x"08",
          2633 => x"2e",
          2634 => x"51",
          2635 => x"80",
          2636 => x"84",
          2637 => x"e4",
          2638 => x"08",
          2639 => x"80",
          2640 => x"74",
          2641 => x"3f",
          2642 => x"08",
          2643 => x"34",
          2644 => x"08",
          2645 => x"81",
          2646 => x"52",
          2647 => x"d2",
          2648 => x"54",
          2649 => x"06",
          2650 => x"73",
          2651 => x"80",
          2652 => x"38",
          2653 => x"d5",
          2654 => x"f0",
          2655 => x"98",
          2656 => x"f0",
          2657 => x"06",
          2658 => x"74",
          2659 => x"c6",
          2660 => x"ff",
          2661 => x"ff",
          2662 => x"79",
          2663 => x"3f",
          2664 => x"81",
          2665 => x"70",
          2666 => x"81",
          2667 => x"59",
          2668 => x"77",
          2669 => x"38",
          2670 => x"73",
          2671 => x"34",
          2672 => x"33",
          2673 => x"80",
          2674 => x"39",
          2675 => x"33",
          2676 => x"2e",
          2677 => x"88",
          2678 => x"3f",
          2679 => x"33",
          2680 => x"73",
          2681 => x"34",
          2682 => x"80",
          2683 => x"9c",
          2684 => x"81",
          2685 => x"79",
          2686 => x"0c",
          2687 => x"04",
          2688 => x"02",
          2689 => x"51",
          2690 => x"72",
          2691 => x"81",
          2692 => x"33",
          2693 => x"fe",
          2694 => x"3d",
          2695 => x"3d",
          2696 => x"05",
          2697 => x"05",
          2698 => x"56",
          2699 => x"72",
          2700 => x"e0",
          2701 => x"2b",
          2702 => x"8c",
          2703 => x"88",
          2704 => x"2e",
          2705 => x"88",
          2706 => x"0c",
          2707 => x"8c",
          2708 => x"71",
          2709 => x"87",
          2710 => x"0c",
          2711 => x"08",
          2712 => x"51",
          2713 => x"2e",
          2714 => x"c0",
          2715 => x"51",
          2716 => x"71",
          2717 => x"80",
          2718 => x"92",
          2719 => x"98",
          2720 => x"70",
          2721 => x"38",
          2722 => x"d8",
          2723 => x"fb",
          2724 => x"51",
          2725 => x"f0",
          2726 => x"0d",
          2727 => x"0d",
          2728 => x"02",
          2729 => x"05",
          2730 => x"58",
          2731 => x"52",
          2732 => x"3f",
          2733 => x"08",
          2734 => x"54",
          2735 => x"be",
          2736 => x"75",
          2737 => x"c0",
          2738 => x"87",
          2739 => x"12",
          2740 => x"84",
          2741 => x"40",
          2742 => x"85",
          2743 => x"98",
          2744 => x"7d",
          2745 => x"0c",
          2746 => x"85",
          2747 => x"06",
          2748 => x"71",
          2749 => x"38",
          2750 => x"71",
          2751 => x"05",
          2752 => x"19",
          2753 => x"a2",
          2754 => x"71",
          2755 => x"38",
          2756 => x"83",
          2757 => x"38",
          2758 => x"8a",
          2759 => x"98",
          2760 => x"71",
          2761 => x"c0",
          2762 => x"52",
          2763 => x"87",
          2764 => x"80",
          2765 => x"81",
          2766 => x"c0",
          2767 => x"53",
          2768 => x"82",
          2769 => x"71",
          2770 => x"1a",
          2771 => x"84",
          2772 => x"19",
          2773 => x"06",
          2774 => x"79",
          2775 => x"38",
          2776 => x"80",
          2777 => x"87",
          2778 => x"26",
          2779 => x"73",
          2780 => x"06",
          2781 => x"2e",
          2782 => x"52",
          2783 => x"81",
          2784 => x"8f",
          2785 => x"f3",
          2786 => x"62",
          2787 => x"05",
          2788 => x"57",
          2789 => x"83",
          2790 => x"52",
          2791 => x"3f",
          2792 => x"08",
          2793 => x"54",
          2794 => x"2e",
          2795 => x"81",
          2796 => x"74",
          2797 => x"c0",
          2798 => x"87",
          2799 => x"12",
          2800 => x"84",
          2801 => x"5f",
          2802 => x"0b",
          2803 => x"8c",
          2804 => x"0c",
          2805 => x"80",
          2806 => x"70",
          2807 => x"81",
          2808 => x"54",
          2809 => x"8c",
          2810 => x"81",
          2811 => x"7c",
          2812 => x"58",
          2813 => x"70",
          2814 => x"52",
          2815 => x"8a",
          2816 => x"98",
          2817 => x"71",
          2818 => x"c0",
          2819 => x"52",
          2820 => x"87",
          2821 => x"80",
          2822 => x"81",
          2823 => x"c0",
          2824 => x"53",
          2825 => x"82",
          2826 => x"71",
          2827 => x"19",
          2828 => x"81",
          2829 => x"ff",
          2830 => x"19",
          2831 => x"78",
          2832 => x"38",
          2833 => x"80",
          2834 => x"87",
          2835 => x"26",
          2836 => x"73",
          2837 => x"06",
          2838 => x"2e",
          2839 => x"52",
          2840 => x"81",
          2841 => x"8f",
          2842 => x"fa",
          2843 => x"02",
          2844 => x"05",
          2845 => x"05",
          2846 => x"71",
          2847 => x"57",
          2848 => x"81",
          2849 => x"81",
          2850 => x"54",
          2851 => x"38",
          2852 => x"c0",
          2853 => x"81",
          2854 => x"2e",
          2855 => x"71",
          2856 => x"38",
          2857 => x"87",
          2858 => x"11",
          2859 => x"80",
          2860 => x"80",
          2861 => x"83",
          2862 => x"38",
          2863 => x"72",
          2864 => x"2a",
          2865 => x"51",
          2866 => x"80",
          2867 => x"87",
          2868 => x"08",
          2869 => x"38",
          2870 => x"8c",
          2871 => x"96",
          2872 => x"0c",
          2873 => x"8c",
          2874 => x"08",
          2875 => x"51",
          2876 => x"38",
          2877 => x"56",
          2878 => x"80",
          2879 => x"85",
          2880 => x"77",
          2881 => x"83",
          2882 => x"75",
          2883 => x"fe",
          2884 => x"3d",
          2885 => x"3d",
          2886 => x"11",
          2887 => x"71",
          2888 => x"81",
          2889 => x"53",
          2890 => x"0d",
          2891 => x"0d",
          2892 => x"33",
          2893 => x"71",
          2894 => x"88",
          2895 => x"14",
          2896 => x"07",
          2897 => x"33",
          2898 => x"fe",
          2899 => x"53",
          2900 => x"52",
          2901 => x"04",
          2902 => x"73",
          2903 => x"92",
          2904 => x"52",
          2905 => x"81",
          2906 => x"70",
          2907 => x"70",
          2908 => x"3d",
          2909 => x"3d",
          2910 => x"52",
          2911 => x"70",
          2912 => x"34",
          2913 => x"51",
          2914 => x"81",
          2915 => x"70",
          2916 => x"70",
          2917 => x"05",
          2918 => x"88",
          2919 => x"72",
          2920 => x"0d",
          2921 => x"0d",
          2922 => x"54",
          2923 => x"80",
          2924 => x"71",
          2925 => x"53",
          2926 => x"81",
          2927 => x"ff",
          2928 => x"39",
          2929 => x"04",
          2930 => x"75",
          2931 => x"52",
          2932 => x"70",
          2933 => x"34",
          2934 => x"70",
          2935 => x"3d",
          2936 => x"3d",
          2937 => x"79",
          2938 => x"74",
          2939 => x"56",
          2940 => x"81",
          2941 => x"71",
          2942 => x"16",
          2943 => x"52",
          2944 => x"86",
          2945 => x"2e",
          2946 => x"81",
          2947 => x"86",
          2948 => x"fe",
          2949 => x"76",
          2950 => x"39",
          2951 => x"8a",
          2952 => x"51",
          2953 => x"71",
          2954 => x"33",
          2955 => x"0c",
          2956 => x"04",
          2957 => x"fe",
          2958 => x"80",
          2959 => x"f0",
          2960 => x"3d",
          2961 => x"80",
          2962 => x"33",
          2963 => x"7a",
          2964 => x"38",
          2965 => x"16",
          2966 => x"16",
          2967 => x"17",
          2968 => x"fa",
          2969 => x"fe",
          2970 => x"2e",
          2971 => x"b7",
          2972 => x"f0",
          2973 => x"34",
          2974 => x"70",
          2975 => x"31",
          2976 => x"59",
          2977 => x"77",
          2978 => x"82",
          2979 => x"74",
          2980 => x"81",
          2981 => x"81",
          2982 => x"53",
          2983 => x"16",
          2984 => x"e3",
          2985 => x"81",
          2986 => x"fe",
          2987 => x"3d",
          2988 => x"3d",
          2989 => x"56",
          2990 => x"74",
          2991 => x"2e",
          2992 => x"51",
          2993 => x"81",
          2994 => x"57",
          2995 => x"08",
          2996 => x"54",
          2997 => x"16",
          2998 => x"33",
          2999 => x"3f",
          3000 => x"08",
          3001 => x"38",
          3002 => x"57",
          3003 => x"0c",
          3004 => x"f0",
          3005 => x"0d",
          3006 => x"0d",
          3007 => x"57",
          3008 => x"81",
          3009 => x"58",
          3010 => x"08",
          3011 => x"76",
          3012 => x"83",
          3013 => x"06",
          3014 => x"84",
          3015 => x"78",
          3016 => x"81",
          3017 => x"38",
          3018 => x"81",
          3019 => x"52",
          3020 => x"52",
          3021 => x"3f",
          3022 => x"52",
          3023 => x"51",
          3024 => x"84",
          3025 => x"d2",
          3026 => x"fc",
          3027 => x"8a",
          3028 => x"52",
          3029 => x"51",
          3030 => x"90",
          3031 => x"84",
          3032 => x"fc",
          3033 => x"17",
          3034 => x"a0",
          3035 => x"86",
          3036 => x"08",
          3037 => x"b0",
          3038 => x"55",
          3039 => x"81",
          3040 => x"f8",
          3041 => x"84",
          3042 => x"53",
          3043 => x"17",
          3044 => x"d7",
          3045 => x"f0",
          3046 => x"83",
          3047 => x"77",
          3048 => x"0c",
          3049 => x"04",
          3050 => x"77",
          3051 => x"12",
          3052 => x"55",
          3053 => x"56",
          3054 => x"8d",
          3055 => x"22",
          3056 => x"ac",
          3057 => x"57",
          3058 => x"fe",
          3059 => x"3d",
          3060 => x"3d",
          3061 => x"70",
          3062 => x"57",
          3063 => x"81",
          3064 => x"98",
          3065 => x"81",
          3066 => x"74",
          3067 => x"72",
          3068 => x"f5",
          3069 => x"24",
          3070 => x"81",
          3071 => x"81",
          3072 => x"83",
          3073 => x"38",
          3074 => x"76",
          3075 => x"70",
          3076 => x"16",
          3077 => x"74",
          3078 => x"96",
          3079 => x"f0",
          3080 => x"38",
          3081 => x"06",
          3082 => x"33",
          3083 => x"89",
          3084 => x"08",
          3085 => x"54",
          3086 => x"fc",
          3087 => x"fe",
          3088 => x"fe",
          3089 => x"ff",
          3090 => x"11",
          3091 => x"2b",
          3092 => x"81",
          3093 => x"2a",
          3094 => x"51",
          3095 => x"e2",
          3096 => x"ff",
          3097 => x"da",
          3098 => x"2a",
          3099 => x"05",
          3100 => x"fc",
          3101 => x"fe",
          3102 => x"c6",
          3103 => x"83",
          3104 => x"05",
          3105 => x"f9",
          3106 => x"fe",
          3107 => x"ff",
          3108 => x"ae",
          3109 => x"2a",
          3110 => x"05",
          3111 => x"fc",
          3112 => x"fe",
          3113 => x"38",
          3114 => x"83",
          3115 => x"05",
          3116 => x"f8",
          3117 => x"fe",
          3118 => x"0a",
          3119 => x"39",
          3120 => x"81",
          3121 => x"89",
          3122 => x"f8",
          3123 => x"7c",
          3124 => x"56",
          3125 => x"77",
          3126 => x"38",
          3127 => x"08",
          3128 => x"38",
          3129 => x"72",
          3130 => x"9d",
          3131 => x"24",
          3132 => x"81",
          3133 => x"82",
          3134 => x"83",
          3135 => x"38",
          3136 => x"76",
          3137 => x"70",
          3138 => x"18",
          3139 => x"76",
          3140 => x"9e",
          3141 => x"f0",
          3142 => x"fe",
          3143 => x"d9",
          3144 => x"ff",
          3145 => x"05",
          3146 => x"81",
          3147 => x"54",
          3148 => x"80",
          3149 => x"77",
          3150 => x"f0",
          3151 => x"8f",
          3152 => x"51",
          3153 => x"34",
          3154 => x"17",
          3155 => x"2a",
          3156 => x"05",
          3157 => x"fa",
          3158 => x"fe",
          3159 => x"81",
          3160 => x"81",
          3161 => x"83",
          3162 => x"b4",
          3163 => x"2a",
          3164 => x"8f",
          3165 => x"2a",
          3166 => x"f0",
          3167 => x"06",
          3168 => x"72",
          3169 => x"ec",
          3170 => x"2a",
          3171 => x"05",
          3172 => x"fa",
          3173 => x"fe",
          3174 => x"81",
          3175 => x"80",
          3176 => x"83",
          3177 => x"52",
          3178 => x"fe",
          3179 => x"b4",
          3180 => x"a4",
          3181 => x"76",
          3182 => x"17",
          3183 => x"75",
          3184 => x"3f",
          3185 => x"08",
          3186 => x"f0",
          3187 => x"77",
          3188 => x"77",
          3189 => x"fc",
          3190 => x"b4",
          3191 => x"51",
          3192 => x"c9",
          3193 => x"f0",
          3194 => x"06",
          3195 => x"72",
          3196 => x"3f",
          3197 => x"17",
          3198 => x"fe",
          3199 => x"3d",
          3200 => x"3d",
          3201 => x"7e",
          3202 => x"56",
          3203 => x"75",
          3204 => x"74",
          3205 => x"27",
          3206 => x"80",
          3207 => x"ff",
          3208 => x"75",
          3209 => x"3f",
          3210 => x"08",
          3211 => x"f0",
          3212 => x"38",
          3213 => x"54",
          3214 => x"81",
          3215 => x"39",
          3216 => x"08",
          3217 => x"39",
          3218 => x"51",
          3219 => x"81",
          3220 => x"58",
          3221 => x"08",
          3222 => x"c7",
          3223 => x"f0",
          3224 => x"d2",
          3225 => x"f0",
          3226 => x"cf",
          3227 => x"74",
          3228 => x"fc",
          3229 => x"fe",
          3230 => x"38",
          3231 => x"fe",
          3232 => x"08",
          3233 => x"74",
          3234 => x"38",
          3235 => x"17",
          3236 => x"33",
          3237 => x"73",
          3238 => x"77",
          3239 => x"26",
          3240 => x"80",
          3241 => x"fe",
          3242 => x"3d",
          3243 => x"3d",
          3244 => x"71",
          3245 => x"5b",
          3246 => x"8c",
          3247 => x"77",
          3248 => x"38",
          3249 => x"78",
          3250 => x"81",
          3251 => x"79",
          3252 => x"f9",
          3253 => x"55",
          3254 => x"f0",
          3255 => x"e0",
          3256 => x"f0",
          3257 => x"fe",
          3258 => x"2e",
          3259 => x"98",
          3260 => x"fe",
          3261 => x"82",
          3262 => x"58",
          3263 => x"70",
          3264 => x"80",
          3265 => x"38",
          3266 => x"09",
          3267 => x"e2",
          3268 => x"56",
          3269 => x"76",
          3270 => x"82",
          3271 => x"7a",
          3272 => x"3f",
          3273 => x"fe",
          3274 => x"2e",
          3275 => x"86",
          3276 => x"f0",
          3277 => x"fe",
          3278 => x"70",
          3279 => x"07",
          3280 => x"7c",
          3281 => x"f0",
          3282 => x"51",
          3283 => x"81",
          3284 => x"fe",
          3285 => x"2e",
          3286 => x"17",
          3287 => x"74",
          3288 => x"73",
          3289 => x"27",
          3290 => x"58",
          3291 => x"80",
          3292 => x"56",
          3293 => x"98",
          3294 => x"26",
          3295 => x"56",
          3296 => x"81",
          3297 => x"52",
          3298 => x"c6",
          3299 => x"f0",
          3300 => x"b8",
          3301 => x"81",
          3302 => x"81",
          3303 => x"06",
          3304 => x"fe",
          3305 => x"81",
          3306 => x"09",
          3307 => x"72",
          3308 => x"70",
          3309 => x"51",
          3310 => x"80",
          3311 => x"78",
          3312 => x"06",
          3313 => x"73",
          3314 => x"39",
          3315 => x"52",
          3316 => x"f7",
          3317 => x"f0",
          3318 => x"f0",
          3319 => x"81",
          3320 => x"07",
          3321 => x"55",
          3322 => x"2e",
          3323 => x"80",
          3324 => x"75",
          3325 => x"76",
          3326 => x"3f",
          3327 => x"08",
          3328 => x"38",
          3329 => x"0c",
          3330 => x"fe",
          3331 => x"08",
          3332 => x"74",
          3333 => x"ff",
          3334 => x"0c",
          3335 => x"81",
          3336 => x"84",
          3337 => x"39",
          3338 => x"81",
          3339 => x"8c",
          3340 => x"8c",
          3341 => x"f0",
          3342 => x"39",
          3343 => x"55",
          3344 => x"f0",
          3345 => x"0d",
          3346 => x"0d",
          3347 => x"55",
          3348 => x"81",
          3349 => x"58",
          3350 => x"fe",
          3351 => x"d8",
          3352 => x"74",
          3353 => x"3f",
          3354 => x"08",
          3355 => x"08",
          3356 => x"59",
          3357 => x"77",
          3358 => x"70",
          3359 => x"c8",
          3360 => x"84",
          3361 => x"56",
          3362 => x"58",
          3363 => x"97",
          3364 => x"75",
          3365 => x"52",
          3366 => x"51",
          3367 => x"81",
          3368 => x"80",
          3369 => x"8a",
          3370 => x"32",
          3371 => x"72",
          3372 => x"2a",
          3373 => x"56",
          3374 => x"f0",
          3375 => x"0d",
          3376 => x"0d",
          3377 => x"08",
          3378 => x"74",
          3379 => x"26",
          3380 => x"74",
          3381 => x"72",
          3382 => x"74",
          3383 => x"88",
          3384 => x"73",
          3385 => x"33",
          3386 => x"27",
          3387 => x"16",
          3388 => x"9b",
          3389 => x"2a",
          3390 => x"88",
          3391 => x"58",
          3392 => x"80",
          3393 => x"16",
          3394 => x"0c",
          3395 => x"8a",
          3396 => x"89",
          3397 => x"72",
          3398 => x"38",
          3399 => x"51",
          3400 => x"81",
          3401 => x"54",
          3402 => x"08",
          3403 => x"38",
          3404 => x"fe",
          3405 => x"8b",
          3406 => x"08",
          3407 => x"08",
          3408 => x"82",
          3409 => x"74",
          3410 => x"cb",
          3411 => x"75",
          3412 => x"3f",
          3413 => x"08",
          3414 => x"73",
          3415 => x"98",
          3416 => x"82",
          3417 => x"2e",
          3418 => x"39",
          3419 => x"39",
          3420 => x"13",
          3421 => x"74",
          3422 => x"16",
          3423 => x"18",
          3424 => x"77",
          3425 => x"0c",
          3426 => x"04",
          3427 => x"7a",
          3428 => x"12",
          3429 => x"59",
          3430 => x"80",
          3431 => x"86",
          3432 => x"98",
          3433 => x"14",
          3434 => x"55",
          3435 => x"81",
          3436 => x"83",
          3437 => x"77",
          3438 => x"81",
          3439 => x"0c",
          3440 => x"55",
          3441 => x"76",
          3442 => x"17",
          3443 => x"74",
          3444 => x"9b",
          3445 => x"39",
          3446 => x"ff",
          3447 => x"2a",
          3448 => x"81",
          3449 => x"52",
          3450 => x"e6",
          3451 => x"f0",
          3452 => x"55",
          3453 => x"fe",
          3454 => x"80",
          3455 => x"55",
          3456 => x"08",
          3457 => x"f4",
          3458 => x"08",
          3459 => x"08",
          3460 => x"38",
          3461 => x"77",
          3462 => x"84",
          3463 => x"39",
          3464 => x"52",
          3465 => x"86",
          3466 => x"f0",
          3467 => x"55",
          3468 => x"08",
          3469 => x"c4",
          3470 => x"81",
          3471 => x"81",
          3472 => x"81",
          3473 => x"f0",
          3474 => x"b0",
          3475 => x"f0",
          3476 => x"51",
          3477 => x"81",
          3478 => x"a0",
          3479 => x"15",
          3480 => x"75",
          3481 => x"3f",
          3482 => x"08",
          3483 => x"76",
          3484 => x"77",
          3485 => x"9c",
          3486 => x"55",
          3487 => x"f0",
          3488 => x"0d",
          3489 => x"0d",
          3490 => x"08",
          3491 => x"80",
          3492 => x"fc",
          3493 => x"fe",
          3494 => x"81",
          3495 => x"80",
          3496 => x"fe",
          3497 => x"98",
          3498 => x"78",
          3499 => x"3f",
          3500 => x"08",
          3501 => x"f0",
          3502 => x"38",
          3503 => x"08",
          3504 => x"70",
          3505 => x"58",
          3506 => x"2e",
          3507 => x"83",
          3508 => x"81",
          3509 => x"55",
          3510 => x"81",
          3511 => x"07",
          3512 => x"2e",
          3513 => x"16",
          3514 => x"2e",
          3515 => x"88",
          3516 => x"81",
          3517 => x"56",
          3518 => x"51",
          3519 => x"81",
          3520 => x"54",
          3521 => x"08",
          3522 => x"9b",
          3523 => x"2e",
          3524 => x"83",
          3525 => x"73",
          3526 => x"0c",
          3527 => x"04",
          3528 => x"76",
          3529 => x"54",
          3530 => x"81",
          3531 => x"83",
          3532 => x"76",
          3533 => x"53",
          3534 => x"2e",
          3535 => x"90",
          3536 => x"51",
          3537 => x"81",
          3538 => x"90",
          3539 => x"53",
          3540 => x"f0",
          3541 => x"0d",
          3542 => x"0d",
          3543 => x"83",
          3544 => x"54",
          3545 => x"55",
          3546 => x"3f",
          3547 => x"51",
          3548 => x"2e",
          3549 => x"8b",
          3550 => x"2a",
          3551 => x"51",
          3552 => x"86",
          3553 => x"f7",
          3554 => x"7d",
          3555 => x"75",
          3556 => x"98",
          3557 => x"2e",
          3558 => x"98",
          3559 => x"78",
          3560 => x"3f",
          3561 => x"08",
          3562 => x"f0",
          3563 => x"38",
          3564 => x"70",
          3565 => x"73",
          3566 => x"58",
          3567 => x"8b",
          3568 => x"bf",
          3569 => x"ff",
          3570 => x"53",
          3571 => x"34",
          3572 => x"08",
          3573 => x"e5",
          3574 => x"81",
          3575 => x"2e",
          3576 => x"70",
          3577 => x"57",
          3578 => x"9e",
          3579 => x"2e",
          3580 => x"fe",
          3581 => x"df",
          3582 => x"72",
          3583 => x"81",
          3584 => x"76",
          3585 => x"2e",
          3586 => x"52",
          3587 => x"fc",
          3588 => x"f0",
          3589 => x"fe",
          3590 => x"38",
          3591 => x"fe",
          3592 => x"39",
          3593 => x"16",
          3594 => x"fe",
          3595 => x"3d",
          3596 => x"3d",
          3597 => x"08",
          3598 => x"52",
          3599 => x"c5",
          3600 => x"f0",
          3601 => x"fe",
          3602 => x"38",
          3603 => x"52",
          3604 => x"de",
          3605 => x"f0",
          3606 => x"fe",
          3607 => x"38",
          3608 => x"fe",
          3609 => x"9c",
          3610 => x"ea",
          3611 => x"53",
          3612 => x"9c",
          3613 => x"ea",
          3614 => x"0b",
          3615 => x"74",
          3616 => x"0c",
          3617 => x"04",
          3618 => x"75",
          3619 => x"12",
          3620 => x"53",
          3621 => x"9a",
          3622 => x"f0",
          3623 => x"9c",
          3624 => x"e5",
          3625 => x"0b",
          3626 => x"85",
          3627 => x"fa",
          3628 => x"7a",
          3629 => x"0b",
          3630 => x"98",
          3631 => x"2e",
          3632 => x"80",
          3633 => x"55",
          3634 => x"17",
          3635 => x"33",
          3636 => x"51",
          3637 => x"2e",
          3638 => x"85",
          3639 => x"06",
          3640 => x"e5",
          3641 => x"2e",
          3642 => x"8b",
          3643 => x"70",
          3644 => x"34",
          3645 => x"71",
          3646 => x"05",
          3647 => x"15",
          3648 => x"27",
          3649 => x"15",
          3650 => x"80",
          3651 => x"34",
          3652 => x"52",
          3653 => x"88",
          3654 => x"17",
          3655 => x"52",
          3656 => x"3f",
          3657 => x"08",
          3658 => x"12",
          3659 => x"3f",
          3660 => x"08",
          3661 => x"98",
          3662 => x"da",
          3663 => x"f0",
          3664 => x"23",
          3665 => x"04",
          3666 => x"7f",
          3667 => x"5b",
          3668 => x"33",
          3669 => x"73",
          3670 => x"38",
          3671 => x"80",
          3672 => x"38",
          3673 => x"8c",
          3674 => x"08",
          3675 => x"aa",
          3676 => x"41",
          3677 => x"33",
          3678 => x"73",
          3679 => x"81",
          3680 => x"81",
          3681 => x"dc",
          3682 => x"70",
          3683 => x"07",
          3684 => x"73",
          3685 => x"88",
          3686 => x"70",
          3687 => x"73",
          3688 => x"38",
          3689 => x"ab",
          3690 => x"52",
          3691 => x"91",
          3692 => x"f0",
          3693 => x"98",
          3694 => x"61",
          3695 => x"5a",
          3696 => x"a0",
          3697 => x"e7",
          3698 => x"70",
          3699 => x"79",
          3700 => x"73",
          3701 => x"81",
          3702 => x"38",
          3703 => x"33",
          3704 => x"ae",
          3705 => x"70",
          3706 => x"82",
          3707 => x"51",
          3708 => x"54",
          3709 => x"79",
          3710 => x"74",
          3711 => x"57",
          3712 => x"af",
          3713 => x"70",
          3714 => x"51",
          3715 => x"dc",
          3716 => x"73",
          3717 => x"38",
          3718 => x"82",
          3719 => x"19",
          3720 => x"54",
          3721 => x"82",
          3722 => x"54",
          3723 => x"78",
          3724 => x"81",
          3725 => x"54",
          3726 => x"81",
          3727 => x"af",
          3728 => x"77",
          3729 => x"70",
          3730 => x"25",
          3731 => x"07",
          3732 => x"51",
          3733 => x"2e",
          3734 => x"39",
          3735 => x"80",
          3736 => x"33",
          3737 => x"73",
          3738 => x"81",
          3739 => x"81",
          3740 => x"dc",
          3741 => x"70",
          3742 => x"07",
          3743 => x"73",
          3744 => x"b5",
          3745 => x"2e",
          3746 => x"83",
          3747 => x"76",
          3748 => x"07",
          3749 => x"2e",
          3750 => x"8b",
          3751 => x"77",
          3752 => x"30",
          3753 => x"71",
          3754 => x"53",
          3755 => x"55",
          3756 => x"38",
          3757 => x"5c",
          3758 => x"75",
          3759 => x"73",
          3760 => x"38",
          3761 => x"06",
          3762 => x"11",
          3763 => x"75",
          3764 => x"3f",
          3765 => x"08",
          3766 => x"38",
          3767 => x"33",
          3768 => x"54",
          3769 => x"e6",
          3770 => x"fe",
          3771 => x"2e",
          3772 => x"ff",
          3773 => x"74",
          3774 => x"38",
          3775 => x"75",
          3776 => x"17",
          3777 => x"57",
          3778 => x"a7",
          3779 => x"81",
          3780 => x"e5",
          3781 => x"fe",
          3782 => x"38",
          3783 => x"54",
          3784 => x"89",
          3785 => x"70",
          3786 => x"57",
          3787 => x"54",
          3788 => x"81",
          3789 => x"f7",
          3790 => x"7e",
          3791 => x"2e",
          3792 => x"33",
          3793 => x"e5",
          3794 => x"06",
          3795 => x"7a",
          3796 => x"a0",
          3797 => x"38",
          3798 => x"55",
          3799 => x"84",
          3800 => x"39",
          3801 => x"8b",
          3802 => x"7b",
          3803 => x"7a",
          3804 => x"3f",
          3805 => x"08",
          3806 => x"f0",
          3807 => x"38",
          3808 => x"52",
          3809 => x"aa",
          3810 => x"f0",
          3811 => x"fe",
          3812 => x"c2",
          3813 => x"08",
          3814 => x"55",
          3815 => x"ff",
          3816 => x"15",
          3817 => x"54",
          3818 => x"34",
          3819 => x"70",
          3820 => x"81",
          3821 => x"58",
          3822 => x"8b",
          3823 => x"74",
          3824 => x"3f",
          3825 => x"08",
          3826 => x"38",
          3827 => x"51",
          3828 => x"ff",
          3829 => x"ab",
          3830 => x"55",
          3831 => x"bb",
          3832 => x"2e",
          3833 => x"80",
          3834 => x"85",
          3835 => x"06",
          3836 => x"58",
          3837 => x"80",
          3838 => x"75",
          3839 => x"73",
          3840 => x"b5",
          3841 => x"0b",
          3842 => x"80",
          3843 => x"39",
          3844 => x"54",
          3845 => x"85",
          3846 => x"75",
          3847 => x"81",
          3848 => x"73",
          3849 => x"1b",
          3850 => x"2a",
          3851 => x"51",
          3852 => x"80",
          3853 => x"90",
          3854 => x"ff",
          3855 => x"05",
          3856 => x"f5",
          3857 => x"fe",
          3858 => x"1c",
          3859 => x"39",
          3860 => x"f0",
          3861 => x"0d",
          3862 => x"0d",
          3863 => x"7b",
          3864 => x"73",
          3865 => x"55",
          3866 => x"2e",
          3867 => x"75",
          3868 => x"57",
          3869 => x"26",
          3870 => x"ba",
          3871 => x"70",
          3872 => x"ba",
          3873 => x"06",
          3874 => x"73",
          3875 => x"70",
          3876 => x"51",
          3877 => x"89",
          3878 => x"82",
          3879 => x"ff",
          3880 => x"56",
          3881 => x"2e",
          3882 => x"80",
          3883 => x"cc",
          3884 => x"08",
          3885 => x"76",
          3886 => x"58",
          3887 => x"81",
          3888 => x"ff",
          3889 => x"53",
          3890 => x"26",
          3891 => x"13",
          3892 => x"06",
          3893 => x"9f",
          3894 => x"99",
          3895 => x"e0",
          3896 => x"ff",
          3897 => x"72",
          3898 => x"2a",
          3899 => x"72",
          3900 => x"06",
          3901 => x"ff",
          3902 => x"30",
          3903 => x"70",
          3904 => x"07",
          3905 => x"9f",
          3906 => x"54",
          3907 => x"80",
          3908 => x"81",
          3909 => x"59",
          3910 => x"25",
          3911 => x"8b",
          3912 => x"24",
          3913 => x"76",
          3914 => x"78",
          3915 => x"81",
          3916 => x"51",
          3917 => x"f0",
          3918 => x"0d",
          3919 => x"0d",
          3920 => x"0b",
          3921 => x"ff",
          3922 => x"0c",
          3923 => x"51",
          3924 => x"84",
          3925 => x"f0",
          3926 => x"38",
          3927 => x"51",
          3928 => x"81",
          3929 => x"83",
          3930 => x"54",
          3931 => x"82",
          3932 => x"09",
          3933 => x"e3",
          3934 => x"b4",
          3935 => x"57",
          3936 => x"2e",
          3937 => x"83",
          3938 => x"74",
          3939 => x"70",
          3940 => x"25",
          3941 => x"51",
          3942 => x"38",
          3943 => x"2e",
          3944 => x"b5",
          3945 => x"81",
          3946 => x"80",
          3947 => x"e0",
          3948 => x"fe",
          3949 => x"81",
          3950 => x"80",
          3951 => x"85",
          3952 => x"90",
          3953 => x"16",
          3954 => x"3f",
          3955 => x"08",
          3956 => x"f0",
          3957 => x"83",
          3958 => x"74",
          3959 => x"0c",
          3960 => x"04",
          3961 => x"61",
          3962 => x"80",
          3963 => x"58",
          3964 => x"0c",
          3965 => x"e1",
          3966 => x"f0",
          3967 => x"56",
          3968 => x"fe",
          3969 => x"86",
          3970 => x"fe",
          3971 => x"29",
          3972 => x"05",
          3973 => x"53",
          3974 => x"80",
          3975 => x"38",
          3976 => x"76",
          3977 => x"74",
          3978 => x"72",
          3979 => x"38",
          3980 => x"51",
          3981 => x"81",
          3982 => x"81",
          3983 => x"81",
          3984 => x"72",
          3985 => x"80",
          3986 => x"38",
          3987 => x"70",
          3988 => x"53",
          3989 => x"86",
          3990 => x"a7",
          3991 => x"34",
          3992 => x"34",
          3993 => x"14",
          3994 => x"b2",
          3995 => x"f0",
          3996 => x"06",
          3997 => x"54",
          3998 => x"72",
          3999 => x"76",
          4000 => x"38",
          4001 => x"70",
          4002 => x"53",
          4003 => x"85",
          4004 => x"70",
          4005 => x"5b",
          4006 => x"81",
          4007 => x"81",
          4008 => x"76",
          4009 => x"81",
          4010 => x"38",
          4011 => x"56",
          4012 => x"83",
          4013 => x"70",
          4014 => x"80",
          4015 => x"83",
          4016 => x"dc",
          4017 => x"fe",
          4018 => x"76",
          4019 => x"05",
          4020 => x"16",
          4021 => x"56",
          4022 => x"d7",
          4023 => x"8d",
          4024 => x"72",
          4025 => x"54",
          4026 => x"57",
          4027 => x"95",
          4028 => x"73",
          4029 => x"3f",
          4030 => x"08",
          4031 => x"57",
          4032 => x"89",
          4033 => x"56",
          4034 => x"d7",
          4035 => x"76",
          4036 => x"f1",
          4037 => x"76",
          4038 => x"e9",
          4039 => x"51",
          4040 => x"81",
          4041 => x"83",
          4042 => x"53",
          4043 => x"2e",
          4044 => x"84",
          4045 => x"ca",
          4046 => x"da",
          4047 => x"f0",
          4048 => x"ff",
          4049 => x"8d",
          4050 => x"14",
          4051 => x"3f",
          4052 => x"08",
          4053 => x"15",
          4054 => x"14",
          4055 => x"34",
          4056 => x"33",
          4057 => x"81",
          4058 => x"54",
          4059 => x"72",
          4060 => x"91",
          4061 => x"ff",
          4062 => x"29",
          4063 => x"33",
          4064 => x"72",
          4065 => x"72",
          4066 => x"38",
          4067 => x"06",
          4068 => x"2e",
          4069 => x"56",
          4070 => x"80",
          4071 => x"da",
          4072 => x"fe",
          4073 => x"81",
          4074 => x"88",
          4075 => x"8f",
          4076 => x"56",
          4077 => x"38",
          4078 => x"51",
          4079 => x"81",
          4080 => x"83",
          4081 => x"55",
          4082 => x"80",
          4083 => x"da",
          4084 => x"fe",
          4085 => x"80",
          4086 => x"da",
          4087 => x"fe",
          4088 => x"ff",
          4089 => x"8d",
          4090 => x"2e",
          4091 => x"88",
          4092 => x"14",
          4093 => x"05",
          4094 => x"75",
          4095 => x"38",
          4096 => x"52",
          4097 => x"51",
          4098 => x"3f",
          4099 => x"08",
          4100 => x"f0",
          4101 => x"82",
          4102 => x"fe",
          4103 => x"ff",
          4104 => x"26",
          4105 => x"57",
          4106 => x"f5",
          4107 => x"82",
          4108 => x"f5",
          4109 => x"81",
          4110 => x"8d",
          4111 => x"2e",
          4112 => x"82",
          4113 => x"16",
          4114 => x"16",
          4115 => x"70",
          4116 => x"7a",
          4117 => x"0c",
          4118 => x"83",
          4119 => x"06",
          4120 => x"de",
          4121 => x"ae",
          4122 => x"f0",
          4123 => x"ff",
          4124 => x"56",
          4125 => x"38",
          4126 => x"38",
          4127 => x"51",
          4128 => x"81",
          4129 => x"a8",
          4130 => x"82",
          4131 => x"39",
          4132 => x"80",
          4133 => x"38",
          4134 => x"15",
          4135 => x"53",
          4136 => x"8d",
          4137 => x"15",
          4138 => x"76",
          4139 => x"51",
          4140 => x"13",
          4141 => x"8d",
          4142 => x"15",
          4143 => x"c5",
          4144 => x"90",
          4145 => x"0b",
          4146 => x"ff",
          4147 => x"15",
          4148 => x"2e",
          4149 => x"81",
          4150 => x"e4",
          4151 => x"b6",
          4152 => x"f0",
          4153 => x"ff",
          4154 => x"81",
          4155 => x"06",
          4156 => x"81",
          4157 => x"51",
          4158 => x"81",
          4159 => x"80",
          4160 => x"fe",
          4161 => x"15",
          4162 => x"14",
          4163 => x"3f",
          4164 => x"08",
          4165 => x"06",
          4166 => x"d4",
          4167 => x"81",
          4168 => x"38",
          4169 => x"d8",
          4170 => x"fe",
          4171 => x"8b",
          4172 => x"2e",
          4173 => x"b3",
          4174 => x"14",
          4175 => x"3f",
          4176 => x"08",
          4177 => x"e4",
          4178 => x"81",
          4179 => x"84",
          4180 => x"d7",
          4181 => x"fe",
          4182 => x"15",
          4183 => x"14",
          4184 => x"3f",
          4185 => x"08",
          4186 => x"76",
          4187 => x"ff",
          4188 => x"05",
          4189 => x"ff",
          4190 => x"86",
          4191 => x"0b",
          4192 => x"80",
          4193 => x"fe",
          4194 => x"3d",
          4195 => x"3d",
          4196 => x"89",
          4197 => x"2e",
          4198 => x"08",
          4199 => x"2e",
          4200 => x"33",
          4201 => x"2e",
          4202 => x"13",
          4203 => x"22",
          4204 => x"76",
          4205 => x"06",
          4206 => x"13",
          4207 => x"c0",
          4208 => x"f0",
          4209 => x"52",
          4210 => x"71",
          4211 => x"55",
          4212 => x"53",
          4213 => x"0c",
          4214 => x"fe",
          4215 => x"3d",
          4216 => x"3d",
          4217 => x"05",
          4218 => x"89",
          4219 => x"52",
          4220 => x"3f",
          4221 => x"0b",
          4222 => x"08",
          4223 => x"81",
          4224 => x"84",
          4225 => x"a0",
          4226 => x"55",
          4227 => x"2e",
          4228 => x"74",
          4229 => x"73",
          4230 => x"38",
          4231 => x"78",
          4232 => x"54",
          4233 => x"92",
          4234 => x"89",
          4235 => x"84",
          4236 => x"b0",
          4237 => x"f0",
          4238 => x"81",
          4239 => x"88",
          4240 => x"eb",
          4241 => x"02",
          4242 => x"e7",
          4243 => x"59",
          4244 => x"80",
          4245 => x"38",
          4246 => x"70",
          4247 => x"d0",
          4248 => x"3d",
          4249 => x"58",
          4250 => x"81",
          4251 => x"55",
          4252 => x"08",
          4253 => x"7a",
          4254 => x"8c",
          4255 => x"56",
          4256 => x"81",
          4257 => x"55",
          4258 => x"08",
          4259 => x"80",
          4260 => x"70",
          4261 => x"57",
          4262 => x"83",
          4263 => x"77",
          4264 => x"73",
          4265 => x"ab",
          4266 => x"2e",
          4267 => x"84",
          4268 => x"06",
          4269 => x"51",
          4270 => x"81",
          4271 => x"55",
          4272 => x"b2",
          4273 => x"06",
          4274 => x"b8",
          4275 => x"2a",
          4276 => x"51",
          4277 => x"2e",
          4278 => x"55",
          4279 => x"77",
          4280 => x"74",
          4281 => x"77",
          4282 => x"81",
          4283 => x"73",
          4284 => x"af",
          4285 => x"7a",
          4286 => x"3f",
          4287 => x"08",
          4288 => x"b2",
          4289 => x"8e",
          4290 => x"ea",
          4291 => x"a0",
          4292 => x"34",
          4293 => x"52",
          4294 => x"bd",
          4295 => x"62",
          4296 => x"d4",
          4297 => x"54",
          4298 => x"15",
          4299 => x"2e",
          4300 => x"7a",
          4301 => x"51",
          4302 => x"75",
          4303 => x"d4",
          4304 => x"be",
          4305 => x"f0",
          4306 => x"fe",
          4307 => x"ca",
          4308 => x"74",
          4309 => x"02",
          4310 => x"70",
          4311 => x"81",
          4312 => x"56",
          4313 => x"86",
          4314 => x"82",
          4315 => x"81",
          4316 => x"06",
          4317 => x"80",
          4318 => x"75",
          4319 => x"73",
          4320 => x"38",
          4321 => x"92",
          4322 => x"7a",
          4323 => x"3f",
          4324 => x"08",
          4325 => x"8c",
          4326 => x"55",
          4327 => x"08",
          4328 => x"77",
          4329 => x"81",
          4330 => x"73",
          4331 => x"38",
          4332 => x"07",
          4333 => x"11",
          4334 => x"0c",
          4335 => x"0c",
          4336 => x"52",
          4337 => x"3f",
          4338 => x"08",
          4339 => x"08",
          4340 => x"63",
          4341 => x"5a",
          4342 => x"81",
          4343 => x"81",
          4344 => x"8c",
          4345 => x"7a",
          4346 => x"17",
          4347 => x"23",
          4348 => x"34",
          4349 => x"1a",
          4350 => x"9c",
          4351 => x"0b",
          4352 => x"77",
          4353 => x"81",
          4354 => x"73",
          4355 => x"8d",
          4356 => x"f0",
          4357 => x"81",
          4358 => x"fe",
          4359 => x"1a",
          4360 => x"22",
          4361 => x"7b",
          4362 => x"a8",
          4363 => x"78",
          4364 => x"3f",
          4365 => x"08",
          4366 => x"f0",
          4367 => x"83",
          4368 => x"81",
          4369 => x"ff",
          4370 => x"06",
          4371 => x"55",
          4372 => x"56",
          4373 => x"76",
          4374 => x"51",
          4375 => x"27",
          4376 => x"70",
          4377 => x"5a",
          4378 => x"76",
          4379 => x"74",
          4380 => x"83",
          4381 => x"73",
          4382 => x"38",
          4383 => x"51",
          4384 => x"81",
          4385 => x"85",
          4386 => x"8e",
          4387 => x"2a",
          4388 => x"08",
          4389 => x"0c",
          4390 => x"79",
          4391 => x"73",
          4392 => x"0c",
          4393 => x"04",
          4394 => x"60",
          4395 => x"40",
          4396 => x"80",
          4397 => x"3d",
          4398 => x"78",
          4399 => x"3f",
          4400 => x"08",
          4401 => x"f0",
          4402 => x"91",
          4403 => x"74",
          4404 => x"38",
          4405 => x"c4",
          4406 => x"33",
          4407 => x"87",
          4408 => x"2e",
          4409 => x"95",
          4410 => x"91",
          4411 => x"56",
          4412 => x"81",
          4413 => x"34",
          4414 => x"a0",
          4415 => x"08",
          4416 => x"31",
          4417 => x"27",
          4418 => x"5c",
          4419 => x"82",
          4420 => x"19",
          4421 => x"ff",
          4422 => x"74",
          4423 => x"7e",
          4424 => x"ff",
          4425 => x"2a",
          4426 => x"79",
          4427 => x"87",
          4428 => x"08",
          4429 => x"98",
          4430 => x"78",
          4431 => x"3f",
          4432 => x"08",
          4433 => x"27",
          4434 => x"74",
          4435 => x"a3",
          4436 => x"1a",
          4437 => x"08",
          4438 => x"d4",
          4439 => x"fe",
          4440 => x"2e",
          4441 => x"81",
          4442 => x"1a",
          4443 => x"59",
          4444 => x"2e",
          4445 => x"77",
          4446 => x"11",
          4447 => x"55",
          4448 => x"85",
          4449 => x"31",
          4450 => x"76",
          4451 => x"81",
          4452 => x"ca",
          4453 => x"fe",
          4454 => x"d7",
          4455 => x"11",
          4456 => x"74",
          4457 => x"38",
          4458 => x"77",
          4459 => x"78",
          4460 => x"84",
          4461 => x"16",
          4462 => x"08",
          4463 => x"2b",
          4464 => x"cf",
          4465 => x"89",
          4466 => x"39",
          4467 => x"0c",
          4468 => x"83",
          4469 => x"80",
          4470 => x"55",
          4471 => x"83",
          4472 => x"9c",
          4473 => x"7e",
          4474 => x"3f",
          4475 => x"08",
          4476 => x"75",
          4477 => x"08",
          4478 => x"1f",
          4479 => x"7c",
          4480 => x"3f",
          4481 => x"7e",
          4482 => x"0c",
          4483 => x"1b",
          4484 => x"1c",
          4485 => x"fd",
          4486 => x"56",
          4487 => x"f0",
          4488 => x"0d",
          4489 => x"0d",
          4490 => x"64",
          4491 => x"58",
          4492 => x"90",
          4493 => x"52",
          4494 => x"d2",
          4495 => x"f0",
          4496 => x"fe",
          4497 => x"38",
          4498 => x"55",
          4499 => x"86",
          4500 => x"83",
          4501 => x"18",
          4502 => x"2a",
          4503 => x"51",
          4504 => x"56",
          4505 => x"83",
          4506 => x"39",
          4507 => x"19",
          4508 => x"83",
          4509 => x"0b",
          4510 => x"81",
          4511 => x"39",
          4512 => x"7c",
          4513 => x"74",
          4514 => x"38",
          4515 => x"7b",
          4516 => x"ec",
          4517 => x"08",
          4518 => x"06",
          4519 => x"81",
          4520 => x"8a",
          4521 => x"05",
          4522 => x"06",
          4523 => x"bf",
          4524 => x"38",
          4525 => x"55",
          4526 => x"7a",
          4527 => x"98",
          4528 => x"77",
          4529 => x"3f",
          4530 => x"08",
          4531 => x"f0",
          4532 => x"82",
          4533 => x"81",
          4534 => x"38",
          4535 => x"ff",
          4536 => x"98",
          4537 => x"18",
          4538 => x"74",
          4539 => x"7e",
          4540 => x"08",
          4541 => x"2e",
          4542 => x"8d",
          4543 => x"ce",
          4544 => x"fe",
          4545 => x"ee",
          4546 => x"08",
          4547 => x"d1",
          4548 => x"fe",
          4549 => x"2e",
          4550 => x"81",
          4551 => x"1b",
          4552 => x"5a",
          4553 => x"2e",
          4554 => x"78",
          4555 => x"11",
          4556 => x"55",
          4557 => x"85",
          4558 => x"31",
          4559 => x"76",
          4560 => x"81",
          4561 => x"c8",
          4562 => x"fe",
          4563 => x"a6",
          4564 => x"11",
          4565 => x"56",
          4566 => x"27",
          4567 => x"80",
          4568 => x"08",
          4569 => x"2b",
          4570 => x"b4",
          4571 => x"b5",
          4572 => x"80",
          4573 => x"34",
          4574 => x"56",
          4575 => x"8c",
          4576 => x"19",
          4577 => x"38",
          4578 => x"b6",
          4579 => x"f0",
          4580 => x"38",
          4581 => x"12",
          4582 => x"9c",
          4583 => x"18",
          4584 => x"06",
          4585 => x"31",
          4586 => x"76",
          4587 => x"7b",
          4588 => x"08",
          4589 => x"cd",
          4590 => x"fe",
          4591 => x"b6",
          4592 => x"7c",
          4593 => x"08",
          4594 => x"1f",
          4595 => x"cb",
          4596 => x"55",
          4597 => x"16",
          4598 => x"31",
          4599 => x"7f",
          4600 => x"94",
          4601 => x"70",
          4602 => x"8c",
          4603 => x"58",
          4604 => x"76",
          4605 => x"75",
          4606 => x"19",
          4607 => x"39",
          4608 => x"80",
          4609 => x"74",
          4610 => x"80",
          4611 => x"fe",
          4612 => x"3d",
          4613 => x"3d",
          4614 => x"3d",
          4615 => x"70",
          4616 => x"ea",
          4617 => x"f0",
          4618 => x"fe",
          4619 => x"fb",
          4620 => x"33",
          4621 => x"70",
          4622 => x"55",
          4623 => x"2e",
          4624 => x"a0",
          4625 => x"78",
          4626 => x"3f",
          4627 => x"08",
          4628 => x"f0",
          4629 => x"38",
          4630 => x"8b",
          4631 => x"07",
          4632 => x"8b",
          4633 => x"16",
          4634 => x"52",
          4635 => x"dd",
          4636 => x"16",
          4637 => x"15",
          4638 => x"3f",
          4639 => x"0a",
          4640 => x"51",
          4641 => x"76",
          4642 => x"51",
          4643 => x"78",
          4644 => x"83",
          4645 => x"51",
          4646 => x"81",
          4647 => x"90",
          4648 => x"bf",
          4649 => x"73",
          4650 => x"76",
          4651 => x"0c",
          4652 => x"04",
          4653 => x"76",
          4654 => x"fe",
          4655 => x"fe",
          4656 => x"81",
          4657 => x"9c",
          4658 => x"fc",
          4659 => x"51",
          4660 => x"81",
          4661 => x"53",
          4662 => x"08",
          4663 => x"fe",
          4664 => x"0c",
          4665 => x"f0",
          4666 => x"0d",
          4667 => x"0d",
          4668 => x"e6",
          4669 => x"52",
          4670 => x"fe",
          4671 => x"8b",
          4672 => x"f0",
          4673 => x"b4",
          4674 => x"71",
          4675 => x"0c",
          4676 => x"04",
          4677 => x"80",
          4678 => x"d0",
          4679 => x"3d",
          4680 => x"3f",
          4681 => x"08",
          4682 => x"f0",
          4683 => x"38",
          4684 => x"52",
          4685 => x"05",
          4686 => x"3f",
          4687 => x"08",
          4688 => x"f0",
          4689 => x"02",
          4690 => x"33",
          4691 => x"55",
          4692 => x"25",
          4693 => x"7a",
          4694 => x"54",
          4695 => x"a2",
          4696 => x"84",
          4697 => x"06",
          4698 => x"73",
          4699 => x"38",
          4700 => x"70",
          4701 => x"a8",
          4702 => x"f0",
          4703 => x"0c",
          4704 => x"fe",
          4705 => x"2e",
          4706 => x"83",
          4707 => x"74",
          4708 => x"0c",
          4709 => x"04",
          4710 => x"6f",
          4711 => x"80",
          4712 => x"53",
          4713 => x"b8",
          4714 => x"3d",
          4715 => x"3f",
          4716 => x"08",
          4717 => x"f0",
          4718 => x"38",
          4719 => x"7c",
          4720 => x"47",
          4721 => x"54",
          4722 => x"81",
          4723 => x"52",
          4724 => x"52",
          4725 => x"3f",
          4726 => x"08",
          4727 => x"f0",
          4728 => x"38",
          4729 => x"51",
          4730 => x"81",
          4731 => x"57",
          4732 => x"08",
          4733 => x"69",
          4734 => x"da",
          4735 => x"fe",
          4736 => x"76",
          4737 => x"d5",
          4738 => x"fe",
          4739 => x"81",
          4740 => x"82",
          4741 => x"52",
          4742 => x"eb",
          4743 => x"f0",
          4744 => x"fe",
          4745 => x"38",
          4746 => x"51",
          4747 => x"73",
          4748 => x"08",
          4749 => x"76",
          4750 => x"d6",
          4751 => x"fe",
          4752 => x"81",
          4753 => x"80",
          4754 => x"76",
          4755 => x"81",
          4756 => x"82",
          4757 => x"39",
          4758 => x"38",
          4759 => x"bc",
          4760 => x"51",
          4761 => x"76",
          4762 => x"11",
          4763 => x"51",
          4764 => x"73",
          4765 => x"38",
          4766 => x"55",
          4767 => x"16",
          4768 => x"56",
          4769 => x"38",
          4770 => x"73",
          4771 => x"90",
          4772 => x"2e",
          4773 => x"16",
          4774 => x"ff",
          4775 => x"ff",
          4776 => x"58",
          4777 => x"74",
          4778 => x"75",
          4779 => x"18",
          4780 => x"58",
          4781 => x"fe",
          4782 => x"7b",
          4783 => x"06",
          4784 => x"18",
          4785 => x"58",
          4786 => x"80",
          4787 => x"b4",
          4788 => x"29",
          4789 => x"05",
          4790 => x"33",
          4791 => x"56",
          4792 => x"2e",
          4793 => x"16",
          4794 => x"33",
          4795 => x"73",
          4796 => x"16",
          4797 => x"26",
          4798 => x"55",
          4799 => x"91",
          4800 => x"54",
          4801 => x"70",
          4802 => x"34",
          4803 => x"ec",
          4804 => x"70",
          4805 => x"34",
          4806 => x"09",
          4807 => x"38",
          4808 => x"39",
          4809 => x"19",
          4810 => x"33",
          4811 => x"05",
          4812 => x"78",
          4813 => x"80",
          4814 => x"81",
          4815 => x"9e",
          4816 => x"f7",
          4817 => x"7d",
          4818 => x"05",
          4819 => x"57",
          4820 => x"3f",
          4821 => x"08",
          4822 => x"f0",
          4823 => x"38",
          4824 => x"53",
          4825 => x"38",
          4826 => x"54",
          4827 => x"92",
          4828 => x"33",
          4829 => x"70",
          4830 => x"54",
          4831 => x"38",
          4832 => x"15",
          4833 => x"70",
          4834 => x"58",
          4835 => x"82",
          4836 => x"8a",
          4837 => x"89",
          4838 => x"53",
          4839 => x"b7",
          4840 => x"ff",
          4841 => x"fc",
          4842 => x"fe",
          4843 => x"15",
          4844 => x"53",
          4845 => x"fb",
          4846 => x"fe",
          4847 => x"26",
          4848 => x"30",
          4849 => x"70",
          4850 => x"77",
          4851 => x"18",
          4852 => x"51",
          4853 => x"88",
          4854 => x"73",
          4855 => x"52",
          4856 => x"ca",
          4857 => x"f0",
          4858 => x"fe",
          4859 => x"2e",
          4860 => x"81",
          4861 => x"ff",
          4862 => x"38",
          4863 => x"08",
          4864 => x"73",
          4865 => x"73",
          4866 => x"9c",
          4867 => x"27",
          4868 => x"75",
          4869 => x"16",
          4870 => x"17",
          4871 => x"33",
          4872 => x"70",
          4873 => x"55",
          4874 => x"80",
          4875 => x"73",
          4876 => x"cc",
          4877 => x"fe",
          4878 => x"81",
          4879 => x"94",
          4880 => x"f0",
          4881 => x"39",
          4882 => x"51",
          4883 => x"81",
          4884 => x"54",
          4885 => x"be",
          4886 => x"27",
          4887 => x"53",
          4888 => x"08",
          4889 => x"73",
          4890 => x"ff",
          4891 => x"15",
          4892 => x"16",
          4893 => x"ff",
          4894 => x"80",
          4895 => x"73",
          4896 => x"c6",
          4897 => x"fe",
          4898 => x"38",
          4899 => x"16",
          4900 => x"80",
          4901 => x"0b",
          4902 => x"81",
          4903 => x"75",
          4904 => x"fe",
          4905 => x"58",
          4906 => x"54",
          4907 => x"74",
          4908 => x"73",
          4909 => x"90",
          4910 => x"c0",
          4911 => x"90",
          4912 => x"83",
          4913 => x"72",
          4914 => x"38",
          4915 => x"08",
          4916 => x"77",
          4917 => x"80",
          4918 => x"fe",
          4919 => x"3d",
          4920 => x"3d",
          4921 => x"89",
          4922 => x"2e",
          4923 => x"80",
          4924 => x"fc",
          4925 => x"3d",
          4926 => x"e1",
          4927 => x"fe",
          4928 => x"81",
          4929 => x"80",
          4930 => x"76",
          4931 => x"75",
          4932 => x"3f",
          4933 => x"08",
          4934 => x"f0",
          4935 => x"38",
          4936 => x"70",
          4937 => x"57",
          4938 => x"a2",
          4939 => x"33",
          4940 => x"70",
          4941 => x"55",
          4942 => x"2e",
          4943 => x"16",
          4944 => x"51",
          4945 => x"81",
          4946 => x"88",
          4947 => x"54",
          4948 => x"84",
          4949 => x"52",
          4950 => x"e5",
          4951 => x"f0",
          4952 => x"84",
          4953 => x"06",
          4954 => x"55",
          4955 => x"80",
          4956 => x"80",
          4957 => x"54",
          4958 => x"f0",
          4959 => x"0d",
          4960 => x"0d",
          4961 => x"fc",
          4962 => x"52",
          4963 => x"3f",
          4964 => x"08",
          4965 => x"fe",
          4966 => x"0c",
          4967 => x"04",
          4968 => x"77",
          4969 => x"fc",
          4970 => x"53",
          4971 => x"de",
          4972 => x"f0",
          4973 => x"fe",
          4974 => x"df",
          4975 => x"38",
          4976 => x"08",
          4977 => x"cd",
          4978 => x"fe",
          4979 => x"80",
          4980 => x"fe",
          4981 => x"73",
          4982 => x"3f",
          4983 => x"08",
          4984 => x"f0",
          4985 => x"09",
          4986 => x"38",
          4987 => x"39",
          4988 => x"08",
          4989 => x"52",
          4990 => x"b3",
          4991 => x"73",
          4992 => x"3f",
          4993 => x"08",
          4994 => x"30",
          4995 => x"9f",
          4996 => x"fe",
          4997 => x"51",
          4998 => x"72",
          4999 => x"0c",
          5000 => x"04",
          5001 => x"65",
          5002 => x"89",
          5003 => x"96",
          5004 => x"df",
          5005 => x"fe",
          5006 => x"81",
          5007 => x"b2",
          5008 => x"75",
          5009 => x"3f",
          5010 => x"08",
          5011 => x"f0",
          5012 => x"02",
          5013 => x"33",
          5014 => x"55",
          5015 => x"25",
          5016 => x"55",
          5017 => x"80",
          5018 => x"76",
          5019 => x"d4",
          5020 => x"81",
          5021 => x"94",
          5022 => x"f0",
          5023 => x"65",
          5024 => x"53",
          5025 => x"05",
          5026 => x"51",
          5027 => x"81",
          5028 => x"5b",
          5029 => x"08",
          5030 => x"7c",
          5031 => x"08",
          5032 => x"fe",
          5033 => x"08",
          5034 => x"55",
          5035 => x"91",
          5036 => x"0c",
          5037 => x"81",
          5038 => x"39",
          5039 => x"c7",
          5040 => x"f0",
          5041 => x"55",
          5042 => x"2e",
          5043 => x"bf",
          5044 => x"5f",
          5045 => x"92",
          5046 => x"51",
          5047 => x"81",
          5048 => x"ff",
          5049 => x"81",
          5050 => x"81",
          5051 => x"81",
          5052 => x"30",
          5053 => x"f0",
          5054 => x"25",
          5055 => x"19",
          5056 => x"5a",
          5057 => x"08",
          5058 => x"38",
          5059 => x"a4",
          5060 => x"fe",
          5061 => x"58",
          5062 => x"77",
          5063 => x"7d",
          5064 => x"bf",
          5065 => x"fe",
          5066 => x"81",
          5067 => x"80",
          5068 => x"70",
          5069 => x"ff",
          5070 => x"56",
          5071 => x"2e",
          5072 => x"9e",
          5073 => x"51",
          5074 => x"3f",
          5075 => x"08",
          5076 => x"06",
          5077 => x"80",
          5078 => x"19",
          5079 => x"54",
          5080 => x"14",
          5081 => x"c5",
          5082 => x"f0",
          5083 => x"06",
          5084 => x"80",
          5085 => x"19",
          5086 => x"54",
          5087 => x"06",
          5088 => x"79",
          5089 => x"78",
          5090 => x"79",
          5091 => x"84",
          5092 => x"07",
          5093 => x"84",
          5094 => x"81",
          5095 => x"92",
          5096 => x"f9",
          5097 => x"8a",
          5098 => x"53",
          5099 => x"e3",
          5100 => x"fe",
          5101 => x"81",
          5102 => x"81",
          5103 => x"17",
          5104 => x"81",
          5105 => x"17",
          5106 => x"2a",
          5107 => x"51",
          5108 => x"55",
          5109 => x"81",
          5110 => x"17",
          5111 => x"8c",
          5112 => x"81",
          5113 => x"9b",
          5114 => x"f0",
          5115 => x"17",
          5116 => x"51",
          5117 => x"81",
          5118 => x"74",
          5119 => x"56",
          5120 => x"98",
          5121 => x"76",
          5122 => x"c6",
          5123 => x"f0",
          5124 => x"09",
          5125 => x"38",
          5126 => x"fe",
          5127 => x"2e",
          5128 => x"85",
          5129 => x"a3",
          5130 => x"38",
          5131 => x"fe",
          5132 => x"15",
          5133 => x"38",
          5134 => x"53",
          5135 => x"08",
          5136 => x"c3",
          5137 => x"fe",
          5138 => x"94",
          5139 => x"18",
          5140 => x"33",
          5141 => x"54",
          5142 => x"34",
          5143 => x"85",
          5144 => x"18",
          5145 => x"74",
          5146 => x"0c",
          5147 => x"04",
          5148 => x"82",
          5149 => x"ff",
          5150 => x"a1",
          5151 => x"e4",
          5152 => x"f0",
          5153 => x"fe",
          5154 => x"f5",
          5155 => x"a1",
          5156 => x"95",
          5157 => x"58",
          5158 => x"81",
          5159 => x"55",
          5160 => x"08",
          5161 => x"02",
          5162 => x"33",
          5163 => x"70",
          5164 => x"55",
          5165 => x"73",
          5166 => x"75",
          5167 => x"80",
          5168 => x"bd",
          5169 => x"d6",
          5170 => x"81",
          5171 => x"87",
          5172 => x"ad",
          5173 => x"78",
          5174 => x"3f",
          5175 => x"08",
          5176 => x"70",
          5177 => x"55",
          5178 => x"2e",
          5179 => x"78",
          5180 => x"f0",
          5181 => x"08",
          5182 => x"38",
          5183 => x"fe",
          5184 => x"76",
          5185 => x"70",
          5186 => x"b5",
          5187 => x"f0",
          5188 => x"fe",
          5189 => x"e9",
          5190 => x"f0",
          5191 => x"51",
          5192 => x"81",
          5193 => x"55",
          5194 => x"08",
          5195 => x"55",
          5196 => x"81",
          5197 => x"84",
          5198 => x"81",
          5199 => x"80",
          5200 => x"51",
          5201 => x"81",
          5202 => x"81",
          5203 => x"30",
          5204 => x"f0",
          5205 => x"25",
          5206 => x"75",
          5207 => x"38",
          5208 => x"8f",
          5209 => x"75",
          5210 => x"c1",
          5211 => x"fe",
          5212 => x"74",
          5213 => x"51",
          5214 => x"3f",
          5215 => x"08",
          5216 => x"fe",
          5217 => x"3d",
          5218 => x"3d",
          5219 => x"99",
          5220 => x"52",
          5221 => x"d8",
          5222 => x"fe",
          5223 => x"81",
          5224 => x"82",
          5225 => x"5e",
          5226 => x"3d",
          5227 => x"cf",
          5228 => x"fe",
          5229 => x"81",
          5230 => x"86",
          5231 => x"82",
          5232 => x"fe",
          5233 => x"2e",
          5234 => x"82",
          5235 => x"80",
          5236 => x"70",
          5237 => x"06",
          5238 => x"54",
          5239 => x"38",
          5240 => x"52",
          5241 => x"52",
          5242 => x"3f",
          5243 => x"08",
          5244 => x"81",
          5245 => x"83",
          5246 => x"81",
          5247 => x"81",
          5248 => x"06",
          5249 => x"54",
          5250 => x"08",
          5251 => x"81",
          5252 => x"81",
          5253 => x"39",
          5254 => x"38",
          5255 => x"08",
          5256 => x"c4",
          5257 => x"fe",
          5258 => x"81",
          5259 => x"81",
          5260 => x"53",
          5261 => x"19",
          5262 => x"8c",
          5263 => x"ae",
          5264 => x"34",
          5265 => x"0b",
          5266 => x"82",
          5267 => x"52",
          5268 => x"51",
          5269 => x"3f",
          5270 => x"b4",
          5271 => x"c9",
          5272 => x"53",
          5273 => x"53",
          5274 => x"51",
          5275 => x"3f",
          5276 => x"0b",
          5277 => x"34",
          5278 => x"80",
          5279 => x"51",
          5280 => x"78",
          5281 => x"83",
          5282 => x"51",
          5283 => x"81",
          5284 => x"54",
          5285 => x"08",
          5286 => x"88",
          5287 => x"64",
          5288 => x"ff",
          5289 => x"75",
          5290 => x"78",
          5291 => x"3f",
          5292 => x"0b",
          5293 => x"78",
          5294 => x"83",
          5295 => x"51",
          5296 => x"3f",
          5297 => x"08",
          5298 => x"80",
          5299 => x"76",
          5300 => x"ae",
          5301 => x"fe",
          5302 => x"3d",
          5303 => x"3d",
          5304 => x"84",
          5305 => x"f1",
          5306 => x"a8",
          5307 => x"05",
          5308 => x"51",
          5309 => x"81",
          5310 => x"55",
          5311 => x"08",
          5312 => x"78",
          5313 => x"08",
          5314 => x"70",
          5315 => x"b8",
          5316 => x"f0",
          5317 => x"fe",
          5318 => x"b9",
          5319 => x"9b",
          5320 => x"a0",
          5321 => x"55",
          5322 => x"38",
          5323 => x"3d",
          5324 => x"3d",
          5325 => x"51",
          5326 => x"3f",
          5327 => x"52",
          5328 => x"52",
          5329 => x"dd",
          5330 => x"08",
          5331 => x"cb",
          5332 => x"fe",
          5333 => x"81",
          5334 => x"95",
          5335 => x"2e",
          5336 => x"88",
          5337 => x"3d",
          5338 => x"38",
          5339 => x"e5",
          5340 => x"f0",
          5341 => x"09",
          5342 => x"b8",
          5343 => x"c9",
          5344 => x"fe",
          5345 => x"81",
          5346 => x"81",
          5347 => x"56",
          5348 => x"3d",
          5349 => x"52",
          5350 => x"ff",
          5351 => x"02",
          5352 => x"8b",
          5353 => x"16",
          5354 => x"2a",
          5355 => x"51",
          5356 => x"89",
          5357 => x"07",
          5358 => x"17",
          5359 => x"81",
          5360 => x"34",
          5361 => x"70",
          5362 => x"81",
          5363 => x"55",
          5364 => x"80",
          5365 => x"64",
          5366 => x"38",
          5367 => x"51",
          5368 => x"81",
          5369 => x"52",
          5370 => x"b7",
          5371 => x"55",
          5372 => x"08",
          5373 => x"dd",
          5374 => x"f0",
          5375 => x"51",
          5376 => x"3f",
          5377 => x"08",
          5378 => x"11",
          5379 => x"81",
          5380 => x"80",
          5381 => x"16",
          5382 => x"ae",
          5383 => x"06",
          5384 => x"53",
          5385 => x"51",
          5386 => x"78",
          5387 => x"83",
          5388 => x"39",
          5389 => x"08",
          5390 => x"51",
          5391 => x"81",
          5392 => x"55",
          5393 => x"08",
          5394 => x"51",
          5395 => x"3f",
          5396 => x"08",
          5397 => x"fe",
          5398 => x"3d",
          5399 => x"3d",
          5400 => x"db",
          5401 => x"84",
          5402 => x"05",
          5403 => x"82",
          5404 => x"d0",
          5405 => x"3d",
          5406 => x"3f",
          5407 => x"08",
          5408 => x"f0",
          5409 => x"38",
          5410 => x"52",
          5411 => x"05",
          5412 => x"3f",
          5413 => x"08",
          5414 => x"f0",
          5415 => x"02",
          5416 => x"33",
          5417 => x"54",
          5418 => x"aa",
          5419 => x"06",
          5420 => x"8b",
          5421 => x"06",
          5422 => x"07",
          5423 => x"56",
          5424 => x"34",
          5425 => x"0b",
          5426 => x"78",
          5427 => x"a9",
          5428 => x"f0",
          5429 => x"81",
          5430 => x"95",
          5431 => x"ef",
          5432 => x"56",
          5433 => x"3d",
          5434 => x"94",
          5435 => x"f4",
          5436 => x"f0",
          5437 => x"fe",
          5438 => x"cb",
          5439 => x"63",
          5440 => x"d4",
          5441 => x"c0",
          5442 => x"f0",
          5443 => x"fe",
          5444 => x"38",
          5445 => x"05",
          5446 => x"06",
          5447 => x"73",
          5448 => x"16",
          5449 => x"22",
          5450 => x"07",
          5451 => x"1f",
          5452 => x"c2",
          5453 => x"81",
          5454 => x"34",
          5455 => x"b3",
          5456 => x"fe",
          5457 => x"74",
          5458 => x"0c",
          5459 => x"04",
          5460 => x"69",
          5461 => x"80",
          5462 => x"d0",
          5463 => x"3d",
          5464 => x"3f",
          5465 => x"08",
          5466 => x"08",
          5467 => x"fe",
          5468 => x"80",
          5469 => x"57",
          5470 => x"81",
          5471 => x"70",
          5472 => x"55",
          5473 => x"80",
          5474 => x"5d",
          5475 => x"52",
          5476 => x"52",
          5477 => x"a9",
          5478 => x"f0",
          5479 => x"fe",
          5480 => x"d1",
          5481 => x"73",
          5482 => x"3f",
          5483 => x"08",
          5484 => x"f0",
          5485 => x"81",
          5486 => x"81",
          5487 => x"65",
          5488 => x"78",
          5489 => x"7b",
          5490 => x"55",
          5491 => x"34",
          5492 => x"8a",
          5493 => x"38",
          5494 => x"1a",
          5495 => x"34",
          5496 => x"9e",
          5497 => x"70",
          5498 => x"51",
          5499 => x"a0",
          5500 => x"8e",
          5501 => x"2e",
          5502 => x"86",
          5503 => x"34",
          5504 => x"30",
          5505 => x"80",
          5506 => x"7a",
          5507 => x"c1",
          5508 => x"2e",
          5509 => x"a0",
          5510 => x"51",
          5511 => x"3f",
          5512 => x"08",
          5513 => x"f0",
          5514 => x"7b",
          5515 => x"55",
          5516 => x"73",
          5517 => x"38",
          5518 => x"73",
          5519 => x"38",
          5520 => x"15",
          5521 => x"ff",
          5522 => x"81",
          5523 => x"7b",
          5524 => x"fe",
          5525 => x"3d",
          5526 => x"3d",
          5527 => x"9c",
          5528 => x"05",
          5529 => x"51",
          5530 => x"81",
          5531 => x"81",
          5532 => x"56",
          5533 => x"f0",
          5534 => x"38",
          5535 => x"52",
          5536 => x"52",
          5537 => x"c0",
          5538 => x"70",
          5539 => x"ff",
          5540 => x"55",
          5541 => x"27",
          5542 => x"78",
          5543 => x"ff",
          5544 => x"05",
          5545 => x"55",
          5546 => x"3f",
          5547 => x"08",
          5548 => x"38",
          5549 => x"70",
          5550 => x"ff",
          5551 => x"81",
          5552 => x"80",
          5553 => x"74",
          5554 => x"07",
          5555 => x"4e",
          5556 => x"81",
          5557 => x"55",
          5558 => x"70",
          5559 => x"06",
          5560 => x"99",
          5561 => x"e0",
          5562 => x"ff",
          5563 => x"54",
          5564 => x"27",
          5565 => x"ea",
          5566 => x"55",
          5567 => x"a3",
          5568 => x"81",
          5569 => x"ff",
          5570 => x"81",
          5571 => x"93",
          5572 => x"75",
          5573 => x"76",
          5574 => x"38",
          5575 => x"77",
          5576 => x"86",
          5577 => x"39",
          5578 => x"27",
          5579 => x"88",
          5580 => x"78",
          5581 => x"5a",
          5582 => x"57",
          5583 => x"81",
          5584 => x"81",
          5585 => x"33",
          5586 => x"06",
          5587 => x"57",
          5588 => x"fe",
          5589 => x"3d",
          5590 => x"55",
          5591 => x"2e",
          5592 => x"76",
          5593 => x"38",
          5594 => x"55",
          5595 => x"33",
          5596 => x"a0",
          5597 => x"06",
          5598 => x"17",
          5599 => x"38",
          5600 => x"43",
          5601 => x"3d",
          5602 => x"ff",
          5603 => x"81",
          5604 => x"54",
          5605 => x"08",
          5606 => x"81",
          5607 => x"ff",
          5608 => x"81",
          5609 => x"54",
          5610 => x"08",
          5611 => x"80",
          5612 => x"54",
          5613 => x"80",
          5614 => x"fe",
          5615 => x"2e",
          5616 => x"80",
          5617 => x"54",
          5618 => x"80",
          5619 => x"52",
          5620 => x"bd",
          5621 => x"fe",
          5622 => x"81",
          5623 => x"b1",
          5624 => x"81",
          5625 => x"52",
          5626 => x"ab",
          5627 => x"54",
          5628 => x"15",
          5629 => x"78",
          5630 => x"ff",
          5631 => x"79",
          5632 => x"83",
          5633 => x"51",
          5634 => x"3f",
          5635 => x"08",
          5636 => x"74",
          5637 => x"0c",
          5638 => x"04",
          5639 => x"60",
          5640 => x"05",
          5641 => x"33",
          5642 => x"05",
          5643 => x"40",
          5644 => x"da",
          5645 => x"f0",
          5646 => x"fe",
          5647 => x"bd",
          5648 => x"33",
          5649 => x"b5",
          5650 => x"2e",
          5651 => x"1a",
          5652 => x"90",
          5653 => x"33",
          5654 => x"70",
          5655 => x"55",
          5656 => x"38",
          5657 => x"97",
          5658 => x"82",
          5659 => x"58",
          5660 => x"7e",
          5661 => x"70",
          5662 => x"55",
          5663 => x"56",
          5664 => x"a7",
          5665 => x"7d",
          5666 => x"70",
          5667 => x"2a",
          5668 => x"08",
          5669 => x"08",
          5670 => x"5d",
          5671 => x"77",
          5672 => x"98",
          5673 => x"26",
          5674 => x"57",
          5675 => x"59",
          5676 => x"52",
          5677 => x"ae",
          5678 => x"15",
          5679 => x"98",
          5680 => x"26",
          5681 => x"55",
          5682 => x"08",
          5683 => x"99",
          5684 => x"f0",
          5685 => x"ff",
          5686 => x"fe",
          5687 => x"38",
          5688 => x"75",
          5689 => x"81",
          5690 => x"93",
          5691 => x"80",
          5692 => x"2e",
          5693 => x"ff",
          5694 => x"58",
          5695 => x"7d",
          5696 => x"38",
          5697 => x"55",
          5698 => x"b4",
          5699 => x"56",
          5700 => x"09",
          5701 => x"38",
          5702 => x"53",
          5703 => x"51",
          5704 => x"3f",
          5705 => x"08",
          5706 => x"f0",
          5707 => x"38",
          5708 => x"ff",
          5709 => x"5c",
          5710 => x"84",
          5711 => x"5c",
          5712 => x"12",
          5713 => x"80",
          5714 => x"78",
          5715 => x"7c",
          5716 => x"90",
          5717 => x"c0",
          5718 => x"90",
          5719 => x"15",
          5720 => x"90",
          5721 => x"54",
          5722 => x"91",
          5723 => x"31",
          5724 => x"84",
          5725 => x"07",
          5726 => x"16",
          5727 => x"73",
          5728 => x"0c",
          5729 => x"04",
          5730 => x"6b",
          5731 => x"05",
          5732 => x"33",
          5733 => x"5a",
          5734 => x"bd",
          5735 => x"80",
          5736 => x"f0",
          5737 => x"f8",
          5738 => x"f0",
          5739 => x"81",
          5740 => x"70",
          5741 => x"74",
          5742 => x"38",
          5743 => x"81",
          5744 => x"81",
          5745 => x"81",
          5746 => x"ff",
          5747 => x"81",
          5748 => x"81",
          5749 => x"81",
          5750 => x"83",
          5751 => x"c0",
          5752 => x"2a",
          5753 => x"51",
          5754 => x"74",
          5755 => x"99",
          5756 => x"53",
          5757 => x"51",
          5758 => x"3f",
          5759 => x"08",
          5760 => x"55",
          5761 => x"92",
          5762 => x"80",
          5763 => x"38",
          5764 => x"06",
          5765 => x"2e",
          5766 => x"48",
          5767 => x"87",
          5768 => x"79",
          5769 => x"78",
          5770 => x"26",
          5771 => x"19",
          5772 => x"74",
          5773 => x"38",
          5774 => x"e4",
          5775 => x"2a",
          5776 => x"70",
          5777 => x"59",
          5778 => x"7a",
          5779 => x"56",
          5780 => x"80",
          5781 => x"51",
          5782 => x"74",
          5783 => x"99",
          5784 => x"53",
          5785 => x"51",
          5786 => x"3f",
          5787 => x"fe",
          5788 => x"ac",
          5789 => x"2a",
          5790 => x"81",
          5791 => x"43",
          5792 => x"83",
          5793 => x"66",
          5794 => x"60",
          5795 => x"90",
          5796 => x"31",
          5797 => x"80",
          5798 => x"8a",
          5799 => x"56",
          5800 => x"26",
          5801 => x"77",
          5802 => x"81",
          5803 => x"74",
          5804 => x"38",
          5805 => x"55",
          5806 => x"83",
          5807 => x"81",
          5808 => x"80",
          5809 => x"38",
          5810 => x"55",
          5811 => x"5e",
          5812 => x"89",
          5813 => x"5a",
          5814 => x"09",
          5815 => x"e1",
          5816 => x"38",
          5817 => x"57",
          5818 => x"ed",
          5819 => x"5a",
          5820 => x"9d",
          5821 => x"26",
          5822 => x"ed",
          5823 => x"10",
          5824 => x"22",
          5825 => x"74",
          5826 => x"38",
          5827 => x"ee",
          5828 => x"66",
          5829 => x"93",
          5830 => x"f0",
          5831 => x"84",
          5832 => x"89",
          5833 => x"a0",
          5834 => x"81",
          5835 => x"fc",
          5836 => x"56",
          5837 => x"f0",
          5838 => x"80",
          5839 => x"d3",
          5840 => x"38",
          5841 => x"57",
          5842 => x"ec",
          5843 => x"5a",
          5844 => x"9d",
          5845 => x"26",
          5846 => x"ec",
          5847 => x"10",
          5848 => x"22",
          5849 => x"74",
          5850 => x"38",
          5851 => x"ee",
          5852 => x"66",
          5853 => x"b3",
          5854 => x"f0",
          5855 => x"05",
          5856 => x"f0",
          5857 => x"26",
          5858 => x"0b",
          5859 => x"08",
          5860 => x"f0",
          5861 => x"11",
          5862 => x"05",
          5863 => x"83",
          5864 => x"2a",
          5865 => x"a0",
          5866 => x"7d",
          5867 => x"69",
          5868 => x"05",
          5869 => x"72",
          5870 => x"5c",
          5871 => x"59",
          5872 => x"2e",
          5873 => x"89",
          5874 => x"60",
          5875 => x"84",
          5876 => x"5d",
          5877 => x"18",
          5878 => x"68",
          5879 => x"74",
          5880 => x"af",
          5881 => x"31",
          5882 => x"53",
          5883 => x"52",
          5884 => x"b7",
          5885 => x"f0",
          5886 => x"83",
          5887 => x"06",
          5888 => x"fe",
          5889 => x"ff",
          5890 => x"dd",
          5891 => x"83",
          5892 => x"2a",
          5893 => x"be",
          5894 => x"39",
          5895 => x"09",
          5896 => x"c5",
          5897 => x"f5",
          5898 => x"f0",
          5899 => x"38",
          5900 => x"79",
          5901 => x"80",
          5902 => x"38",
          5903 => x"96",
          5904 => x"06",
          5905 => x"2e",
          5906 => x"5e",
          5907 => x"81",
          5908 => x"9f",
          5909 => x"38",
          5910 => x"38",
          5911 => x"81",
          5912 => x"fc",
          5913 => x"ab",
          5914 => x"7d",
          5915 => x"81",
          5916 => x"7d",
          5917 => x"78",
          5918 => x"74",
          5919 => x"8e",
          5920 => x"9c",
          5921 => x"53",
          5922 => x"51",
          5923 => x"3f",
          5924 => x"eb",
          5925 => x"51",
          5926 => x"3f",
          5927 => x"8b",
          5928 => x"a1",
          5929 => x"8d",
          5930 => x"83",
          5931 => x"52",
          5932 => x"ff",
          5933 => x"81",
          5934 => x"34",
          5935 => x"70",
          5936 => x"2a",
          5937 => x"54",
          5938 => x"1b",
          5939 => x"88",
          5940 => x"74",
          5941 => x"26",
          5942 => x"83",
          5943 => x"52",
          5944 => x"ff",
          5945 => x"8a",
          5946 => x"a0",
          5947 => x"a1",
          5948 => x"0b",
          5949 => x"bf",
          5950 => x"51",
          5951 => x"3f",
          5952 => x"9a",
          5953 => x"a0",
          5954 => x"52",
          5955 => x"ff",
          5956 => x"7d",
          5957 => x"81",
          5958 => x"38",
          5959 => x"0a",
          5960 => x"1b",
          5961 => x"ce",
          5962 => x"a4",
          5963 => x"a0",
          5964 => x"52",
          5965 => x"ff",
          5966 => x"81",
          5967 => x"51",
          5968 => x"3f",
          5969 => x"1b",
          5970 => x"8c",
          5971 => x"0b",
          5972 => x"34",
          5973 => x"c2",
          5974 => x"53",
          5975 => x"52",
          5976 => x"51",
          5977 => x"88",
          5978 => x"a7",
          5979 => x"a0",
          5980 => x"83",
          5981 => x"52",
          5982 => x"ff",
          5983 => x"ff",
          5984 => x"1c",
          5985 => x"a6",
          5986 => x"53",
          5987 => x"52",
          5988 => x"ff",
          5989 => x"82",
          5990 => x"83",
          5991 => x"52",
          5992 => x"b4",
          5993 => x"60",
          5994 => x"7e",
          5995 => x"d7",
          5996 => x"81",
          5997 => x"83",
          5998 => x"83",
          5999 => x"06",
          6000 => x"75",
          6001 => x"05",
          6002 => x"7e",
          6003 => x"b7",
          6004 => x"53",
          6005 => x"51",
          6006 => x"3f",
          6007 => x"a4",
          6008 => x"51",
          6009 => x"3f",
          6010 => x"e4",
          6011 => x"e4",
          6012 => x"9f",
          6013 => x"18",
          6014 => x"1b",
          6015 => x"f6",
          6016 => x"83",
          6017 => x"ff",
          6018 => x"82",
          6019 => x"78",
          6020 => x"c4",
          6021 => x"60",
          6022 => x"7a",
          6023 => x"ff",
          6024 => x"75",
          6025 => x"53",
          6026 => x"51",
          6027 => x"3f",
          6028 => x"52",
          6029 => x"9f",
          6030 => x"56",
          6031 => x"83",
          6032 => x"06",
          6033 => x"52",
          6034 => x"9e",
          6035 => x"52",
          6036 => x"ff",
          6037 => x"f0",
          6038 => x"1b",
          6039 => x"87",
          6040 => x"55",
          6041 => x"83",
          6042 => x"74",
          6043 => x"ff",
          6044 => x"7c",
          6045 => x"74",
          6046 => x"38",
          6047 => x"54",
          6048 => x"52",
          6049 => x"99",
          6050 => x"fe",
          6051 => x"87",
          6052 => x"53",
          6053 => x"08",
          6054 => x"ff",
          6055 => x"76",
          6056 => x"31",
          6057 => x"cd",
          6058 => x"58",
          6059 => x"ff",
          6060 => x"55",
          6061 => x"83",
          6062 => x"61",
          6063 => x"26",
          6064 => x"57",
          6065 => x"53",
          6066 => x"51",
          6067 => x"3f",
          6068 => x"08",
          6069 => x"76",
          6070 => x"31",
          6071 => x"db",
          6072 => x"7d",
          6073 => x"38",
          6074 => x"83",
          6075 => x"8a",
          6076 => x"7d",
          6077 => x"38",
          6078 => x"81",
          6079 => x"80",
          6080 => x"80",
          6081 => x"7a",
          6082 => x"bc",
          6083 => x"d5",
          6084 => x"ff",
          6085 => x"83",
          6086 => x"77",
          6087 => x"0b",
          6088 => x"81",
          6089 => x"34",
          6090 => x"34",
          6091 => x"34",
          6092 => x"56",
          6093 => x"52",
          6094 => x"d4",
          6095 => x"0b",
          6096 => x"81",
          6097 => x"82",
          6098 => x"56",
          6099 => x"34",
          6100 => x"08",
          6101 => x"60",
          6102 => x"1b",
          6103 => x"96",
          6104 => x"83",
          6105 => x"ff",
          6106 => x"81",
          6107 => x"7a",
          6108 => x"ff",
          6109 => x"81",
          6110 => x"f0",
          6111 => x"80",
          6112 => x"7e",
          6113 => x"e3",
          6114 => x"81",
          6115 => x"90",
          6116 => x"8e",
          6117 => x"81",
          6118 => x"81",
          6119 => x"56",
          6120 => x"f0",
          6121 => x"0d",
          6122 => x"0d",
          6123 => x"59",
          6124 => x"ff",
          6125 => x"57",
          6126 => x"b4",
          6127 => x"f8",
          6128 => x"81",
          6129 => x"52",
          6130 => x"dc",
          6131 => x"2e",
          6132 => x"9c",
          6133 => x"33",
          6134 => x"2e",
          6135 => x"76",
          6136 => x"58",
          6137 => x"57",
          6138 => x"09",
          6139 => x"38",
          6140 => x"78",
          6141 => x"38",
          6142 => x"81",
          6143 => x"8d",
          6144 => x"f7",
          6145 => x"02",
          6146 => x"05",
          6147 => x"77",
          6148 => x"81",
          6149 => x"8d",
          6150 => x"e7",
          6151 => x"08",
          6152 => x"24",
          6153 => x"17",
          6154 => x"8c",
          6155 => x"77",
          6156 => x"16",
          6157 => x"25",
          6158 => x"3d",
          6159 => x"75",
          6160 => x"52",
          6161 => x"cb",
          6162 => x"76",
          6163 => x"70",
          6164 => x"2a",
          6165 => x"51",
          6166 => x"84",
          6167 => x"19",
          6168 => x"8b",
          6169 => x"f9",
          6170 => x"84",
          6171 => x"56",
          6172 => x"a7",
          6173 => x"fc",
          6174 => x"53",
          6175 => x"75",
          6176 => x"a1",
          6177 => x"f0",
          6178 => x"84",
          6179 => x"2e",
          6180 => x"87",
          6181 => x"08",
          6182 => x"ff",
          6183 => x"fe",
          6184 => x"3d",
          6185 => x"3d",
          6186 => x"80",
          6187 => x"52",
          6188 => x"9a",
          6189 => x"74",
          6190 => x"0d",
          6191 => x"0d",
          6192 => x"05",
          6193 => x"86",
          6194 => x"54",
          6195 => x"73",
          6196 => x"fe",
          6197 => x"51",
          6198 => x"98",
          6199 => x"f8",
          6200 => x"70",
          6201 => x"56",
          6202 => x"2e",
          6203 => x"8c",
          6204 => x"79",
          6205 => x"33",
          6206 => x"39",
          6207 => x"73",
          6208 => x"81",
          6209 => x"81",
          6210 => x"39",
          6211 => x"90",
          6212 => x"e0",
          6213 => x"52",
          6214 => x"b1",
          6215 => x"f0",
          6216 => x"f0",
          6217 => x"53",
          6218 => x"58",
          6219 => x"3f",
          6220 => x"08",
          6221 => x"16",
          6222 => x"81",
          6223 => x"38",
          6224 => x"81",
          6225 => x"54",
          6226 => x"c2",
          6227 => x"73",
          6228 => x"0c",
          6229 => x"04",
          6230 => x"73",
          6231 => x"26",
          6232 => x"71",
          6233 => x"e2",
          6234 => x"71",
          6235 => x"ee",
          6236 => x"80",
          6237 => x"c4",
          6238 => x"39",
          6239 => x"51",
          6240 => x"81",
          6241 => x"80",
          6242 => x"ee",
          6243 => x"e4",
          6244 => x"8c",
          6245 => x"39",
          6246 => x"51",
          6247 => x"81",
          6248 => x"80",
          6249 => x"ef",
          6250 => x"c8",
          6251 => x"e0",
          6252 => x"39",
          6253 => x"51",
          6254 => x"f0",
          6255 => x"39",
          6256 => x"51",
          6257 => x"f0",
          6258 => x"39",
          6259 => x"51",
          6260 => x"f1",
          6261 => x"39",
          6262 => x"51",
          6263 => x"f1",
          6264 => x"39",
          6265 => x"51",
          6266 => x"f1",
          6267 => x"39",
          6268 => x"51",
          6269 => x"3f",
          6270 => x"04",
          6271 => x"77",
          6272 => x"74",
          6273 => x"8a",
          6274 => x"75",
          6275 => x"51",
          6276 => x"e8",
          6277 => x"fe",
          6278 => x"81",
          6279 => x"52",
          6280 => x"cf",
          6281 => x"fe",
          6282 => x"79",
          6283 => x"81",
          6284 => x"fe",
          6285 => x"87",
          6286 => x"ec",
          6287 => x"02",
          6288 => x"e3",
          6289 => x"57",
          6290 => x"30",
          6291 => x"73",
          6292 => x"59",
          6293 => x"77",
          6294 => x"83",
          6295 => x"74",
          6296 => x"81",
          6297 => x"55",
          6298 => x"81",
          6299 => x"53",
          6300 => x"3d",
          6301 => x"ff",
          6302 => x"81",
          6303 => x"57",
          6304 => x"08",
          6305 => x"fe",
          6306 => x"c0",
          6307 => x"81",
          6308 => x"59",
          6309 => x"05",
          6310 => x"53",
          6311 => x"51",
          6312 => x"81",
          6313 => x"57",
          6314 => x"08",
          6315 => x"55",
          6316 => x"89",
          6317 => x"75",
          6318 => x"d8",
          6319 => x"d8",
          6320 => x"f0",
          6321 => x"70",
          6322 => x"25",
          6323 => x"9f",
          6324 => x"51",
          6325 => x"74",
          6326 => x"38",
          6327 => x"53",
          6328 => x"88",
          6329 => x"51",
          6330 => x"76",
          6331 => x"fe",
          6332 => x"3d",
          6333 => x"3d",
          6334 => x"84",
          6335 => x"33",
          6336 => x"57",
          6337 => x"52",
          6338 => x"af",
          6339 => x"f0",
          6340 => x"75",
          6341 => x"38",
          6342 => x"98",
          6343 => x"60",
          6344 => x"81",
          6345 => x"7e",
          6346 => x"77",
          6347 => x"f0",
          6348 => x"39",
          6349 => x"81",
          6350 => x"89",
          6351 => x"f3",
          6352 => x"61",
          6353 => x"05",
          6354 => x"33",
          6355 => x"68",
          6356 => x"5c",
          6357 => x"7a",
          6358 => x"ac",
          6359 => x"a9",
          6360 => x"b4",
          6361 => x"bd",
          6362 => x"74",
          6363 => x"fc",
          6364 => x"2e",
          6365 => x"a0",
          6366 => x"80",
          6367 => x"18",
          6368 => x"27",
          6369 => x"22",
          6370 => x"b8",
          6371 => x"f9",
          6372 => x"81",
          6373 => x"fe",
          6374 => x"82",
          6375 => x"c3",
          6376 => x"53",
          6377 => x"8e",
          6378 => x"52",
          6379 => x"51",
          6380 => x"3f",
          6381 => x"f2",
          6382 => x"ee",
          6383 => x"15",
          6384 => x"74",
          6385 => x"7a",
          6386 => x"72",
          6387 => x"f2",
          6388 => x"f4",
          6389 => x"39",
          6390 => x"51",
          6391 => x"3f",
          6392 => x"a0",
          6393 => x"e0",
          6394 => x"39",
          6395 => x"51",
          6396 => x"3f",
          6397 => x"79",
          6398 => x"74",
          6399 => x"55",
          6400 => x"72",
          6401 => x"38",
          6402 => x"53",
          6403 => x"83",
          6404 => x"75",
          6405 => x"81",
          6406 => x"53",
          6407 => x"8b",
          6408 => x"fe",
          6409 => x"73",
          6410 => x"a0",
          6411 => x"98",
          6412 => x"55",
          6413 => x"f2",
          6414 => x"ed",
          6415 => x"18",
          6416 => x"58",
          6417 => x"3f",
          6418 => x"08",
          6419 => x"98",
          6420 => x"76",
          6421 => x"81",
          6422 => x"fe",
          6423 => x"81",
          6424 => x"98",
          6425 => x"2c",
          6426 => x"70",
          6427 => x"32",
          6428 => x"72",
          6429 => x"07",
          6430 => x"58",
          6431 => x"57",
          6432 => x"d7",
          6433 => x"2e",
          6434 => x"85",
          6435 => x"8c",
          6436 => x"53",
          6437 => x"fd",
          6438 => x"53",
          6439 => x"f0",
          6440 => x"0d",
          6441 => x"0d",
          6442 => x"33",
          6443 => x"53",
          6444 => x"52",
          6445 => x"d1",
          6446 => x"a0",
          6447 => x"e6",
          6448 => x"f2",
          6449 => x"f3",
          6450 => x"fa",
          6451 => x"81",
          6452 => x"fe",
          6453 => x"74",
          6454 => x"38",
          6455 => x"3f",
          6456 => x"04",
          6457 => x"87",
          6458 => x"08",
          6459 => x"b1",
          6460 => x"fe",
          6461 => x"81",
          6462 => x"fe",
          6463 => x"80",
          6464 => x"ed",
          6465 => x"2a",
          6466 => x"51",
          6467 => x"2e",
          6468 => x"51",
          6469 => x"3f",
          6470 => x"51",
          6471 => x"3f",
          6472 => x"d8",
          6473 => x"82",
          6474 => x"06",
          6475 => x"80",
          6476 => x"81",
          6477 => x"b9",
          6478 => x"d4",
          6479 => x"b1",
          6480 => x"fe",
          6481 => x"72",
          6482 => x"81",
          6483 => x"71",
          6484 => x"38",
          6485 => x"d8",
          6486 => x"f3",
          6487 => x"da",
          6488 => x"51",
          6489 => x"3f",
          6490 => x"70",
          6491 => x"52",
          6492 => x"95",
          6493 => x"fe",
          6494 => x"81",
          6495 => x"fe",
          6496 => x"80",
          6497 => x"e9",
          6498 => x"2a",
          6499 => x"51",
          6500 => x"2e",
          6501 => x"51",
          6502 => x"3f",
          6503 => x"51",
          6504 => x"3f",
          6505 => x"d7",
          6506 => x"86",
          6507 => x"06",
          6508 => x"80",
          6509 => x"81",
          6510 => x"b5",
          6511 => x"a0",
          6512 => x"ad",
          6513 => x"fe",
          6514 => x"72",
          6515 => x"81",
          6516 => x"71",
          6517 => x"38",
          6518 => x"d7",
          6519 => x"f4",
          6520 => x"d9",
          6521 => x"51",
          6522 => x"3f",
          6523 => x"70",
          6524 => x"52",
          6525 => x"95",
          6526 => x"fe",
          6527 => x"81",
          6528 => x"fe",
          6529 => x"80",
          6530 => x"e5",
          6531 => x"99",
          6532 => x"0d",
          6533 => x"0d",
          6534 => x"05",
          6535 => x"70",
          6536 => x"80",
          6537 => x"fe",
          6538 => x"81",
          6539 => x"54",
          6540 => x"81",
          6541 => x"88",
          6542 => x"88",
          6543 => x"83",
          6544 => x"f0",
          6545 => x"81",
          6546 => x"07",
          6547 => x"71",
          6548 => x"54",
          6549 => x"dc",
          6550 => x"dc",
          6551 => x"81",
          6552 => x"06",
          6553 => x"96",
          6554 => x"52",
          6555 => x"b9",
          6556 => x"f0",
          6557 => x"8c",
          6558 => x"f0",
          6559 => x"e9",
          6560 => x"39",
          6561 => x"51",
          6562 => x"82",
          6563 => x"dc",
          6564 => x"dc",
          6565 => x"82",
          6566 => x"06",
          6567 => x"52",
          6568 => x"fa",
          6569 => x"0b",
          6570 => x"0c",
          6571 => x"04",
          6572 => x"80",
          6573 => x"96",
          6574 => x"5d",
          6575 => x"51",
          6576 => x"3f",
          6577 => x"08",
          6578 => x"59",
          6579 => x"09",
          6580 => x"38",
          6581 => x"52",
          6582 => x"52",
          6583 => x"bf",
          6584 => x"78",
          6585 => x"b4",
          6586 => x"f6",
          6587 => x"f0",
          6588 => x"88",
          6589 => x"9c",
          6590 => x"39",
          6591 => x"5d",
          6592 => x"51",
          6593 => x"3f",
          6594 => x"46",
          6595 => x"52",
          6596 => x"81",
          6597 => x"ff",
          6598 => x"f3",
          6599 => x"fe",
          6600 => x"2b",
          6601 => x"51",
          6602 => x"c1",
          6603 => x"38",
          6604 => x"24",
          6605 => x"78",
          6606 => x"c0",
          6607 => x"24",
          6608 => x"82",
          6609 => x"38",
          6610 => x"8a",
          6611 => x"2e",
          6612 => x"8f",
          6613 => x"84",
          6614 => x"38",
          6615 => x"82",
          6616 => x"96",
          6617 => x"2e",
          6618 => x"78",
          6619 => x"38",
          6620 => x"83",
          6621 => x"bc",
          6622 => x"38",
          6623 => x"78",
          6624 => x"d7",
          6625 => x"c0",
          6626 => x"38",
          6627 => x"78",
          6628 => x"8d",
          6629 => x"80",
          6630 => x"38",
          6631 => x"2e",
          6632 => x"78",
          6633 => x"92",
          6634 => x"c2",
          6635 => x"38",
          6636 => x"2e",
          6637 => x"8e",
          6638 => x"80",
          6639 => x"e9",
          6640 => x"d4",
          6641 => x"38",
          6642 => x"78",
          6643 => x"8e",
          6644 => x"81",
          6645 => x"38",
          6646 => x"2e",
          6647 => x"78",
          6648 => x"8d",
          6649 => x"92",
          6650 => x"83",
          6651 => x"38",
          6652 => x"2e",
          6653 => x"8e",
          6654 => x"3d",
          6655 => x"53",
          6656 => x"51",
          6657 => x"3f",
          6658 => x"08",
          6659 => x"f5",
          6660 => x"e5",
          6661 => x"fe",
          6662 => x"ff",
          6663 => x"fe",
          6664 => x"81",
          6665 => x"80",
          6666 => x"81",
          6667 => x"38",
          6668 => x"80",
          6669 => x"52",
          6670 => x"05",
          6671 => x"83",
          6672 => x"fe",
          6673 => x"ff",
          6674 => x"8e",
          6675 => x"e8",
          6676 => x"d1",
          6677 => x"fd",
          6678 => x"f5",
          6679 => x"b9",
          6680 => x"ff",
          6681 => x"ff",
          6682 => x"fe",
          6683 => x"81",
          6684 => x"80",
          6685 => x"38",
          6686 => x"52",
          6687 => x"05",
          6688 => x"87",
          6689 => x"fe",
          6690 => x"81",
          6691 => x"8c",
          6692 => x"3d",
          6693 => x"53",
          6694 => x"51",
          6695 => x"3f",
          6696 => x"08",
          6697 => x"38",
          6698 => x"fc",
          6699 => x"3d",
          6700 => x"53",
          6701 => x"51",
          6702 => x"3f",
          6703 => x"08",
          6704 => x"fe",
          6705 => x"63",
          6706 => x"98",
          6707 => x"fe",
          6708 => x"02",
          6709 => x"33",
          6710 => x"63",
          6711 => x"82",
          6712 => x"51",
          6713 => x"3f",
          6714 => x"08",
          6715 => x"81",
          6716 => x"fe",
          6717 => x"81",
          6718 => x"39",
          6719 => x"84",
          6720 => x"cd",
          6721 => x"fe",
          6722 => x"3d",
          6723 => x"52",
          6724 => x"f0",
          6725 => x"81",
          6726 => x"52",
          6727 => x"9b",
          6728 => x"39",
          6729 => x"84",
          6730 => x"cc",
          6731 => x"fe",
          6732 => x"3d",
          6733 => x"52",
          6734 => x"c8",
          6735 => x"f0",
          6736 => x"ff",
          6737 => x"5a",
          6738 => x"3f",
          6739 => x"08",
          6740 => x"84",
          6741 => x"fe",
          6742 => x"81",
          6743 => x"81",
          6744 => x"80",
          6745 => x"81",
          6746 => x"81",
          6747 => x"78",
          6748 => x"7a",
          6749 => x"3f",
          6750 => x"08",
          6751 => x"80",
          6752 => x"f0",
          6753 => x"d0",
          6754 => x"39",
          6755 => x"80",
          6756 => x"84",
          6757 => x"ea",
          6758 => x"fe",
          6759 => x"2e",
          6760 => x"b4",
          6761 => x"11",
          6762 => x"05",
          6763 => x"ce",
          6764 => x"f0",
          6765 => x"fa",
          6766 => x"3d",
          6767 => x"53",
          6768 => x"51",
          6769 => x"3f",
          6770 => x"08",
          6771 => x"fe",
          6772 => x"81",
          6773 => x"fe",
          6774 => x"63",
          6775 => x"79",
          6776 => x"f2",
          6777 => x"78",
          6778 => x"05",
          6779 => x"7a",
          6780 => x"81",
          6781 => x"3d",
          6782 => x"53",
          6783 => x"51",
          6784 => x"3f",
          6785 => x"08",
          6786 => x"f4",
          6787 => x"fe",
          6788 => x"ff",
          6789 => x"fe",
          6790 => x"81",
          6791 => x"80",
          6792 => x"38",
          6793 => x"f8",
          6794 => x"84",
          6795 => x"e9",
          6796 => x"fe",
          6797 => x"2e",
          6798 => x"81",
          6799 => x"fe",
          6800 => x"63",
          6801 => x"27",
          6802 => x"61",
          6803 => x"81",
          6804 => x"79",
          6805 => x"05",
          6806 => x"b4",
          6807 => x"11",
          6808 => x"05",
          6809 => x"96",
          6810 => x"f0",
          6811 => x"f9",
          6812 => x"3d",
          6813 => x"53",
          6814 => x"51",
          6815 => x"3f",
          6816 => x"08",
          6817 => x"f8",
          6818 => x"fe",
          6819 => x"ff",
          6820 => x"fe",
          6821 => x"81",
          6822 => x"80",
          6823 => x"38",
          6824 => x"51",
          6825 => x"3f",
          6826 => x"63",
          6827 => x"61",
          6828 => x"33",
          6829 => x"78",
          6830 => x"38",
          6831 => x"54",
          6832 => x"79",
          6833 => x"c8",
          6834 => x"bd",
          6835 => x"62",
          6836 => x"5a",
          6837 => x"f5",
          6838 => x"bd",
          6839 => x"ff",
          6840 => x"ff",
          6841 => x"fe",
          6842 => x"81",
          6843 => x"80",
          6844 => x"fa",
          6845 => x"78",
          6846 => x"38",
          6847 => x"08",
          6848 => x"39",
          6849 => x"33",
          6850 => x"2e",
          6851 => x"f9",
          6852 => x"bc",
          6853 => x"b6",
          6854 => x"80",
          6855 => x"81",
          6856 => x"44",
          6857 => x"fa",
          6858 => x"78",
          6859 => x"38",
          6860 => x"08",
          6861 => x"81",
          6862 => x"59",
          6863 => x"88",
          6864 => x"8c",
          6865 => x"39",
          6866 => x"08",
          6867 => x"44",
          6868 => x"fc",
          6869 => x"84",
          6870 => x"e7",
          6871 => x"fe",
          6872 => x"de",
          6873 => x"b4",
          6874 => x"80",
          6875 => x"81",
          6876 => x"43",
          6877 => x"81",
          6878 => x"59",
          6879 => x"88",
          6880 => x"f8",
          6881 => x"39",
          6882 => x"33",
          6883 => x"2e",
          6884 => x"fa",
          6885 => x"aa",
          6886 => x"b7",
          6887 => x"80",
          6888 => x"81",
          6889 => x"43",
          6890 => x"fa",
          6891 => x"78",
          6892 => x"38",
          6893 => x"08",
          6894 => x"81",
          6895 => x"88",
          6896 => x"3d",
          6897 => x"53",
          6898 => x"51",
          6899 => x"3f",
          6900 => x"08",
          6901 => x"38",
          6902 => x"5c",
          6903 => x"83",
          6904 => x"7a",
          6905 => x"30",
          6906 => x"9f",
          6907 => x"06",
          6908 => x"5a",
          6909 => x"88",
          6910 => x"2e",
          6911 => x"42",
          6912 => x"51",
          6913 => x"3f",
          6914 => x"54",
          6915 => x"52",
          6916 => x"ab",
          6917 => x"f4",
          6918 => x"89",
          6919 => x"39",
          6920 => x"80",
          6921 => x"84",
          6922 => x"e5",
          6923 => x"fe",
          6924 => x"2e",
          6925 => x"b4",
          6926 => x"11",
          6927 => x"05",
          6928 => x"ba",
          6929 => x"f0",
          6930 => x"a5",
          6931 => x"02",
          6932 => x"33",
          6933 => x"81",
          6934 => x"3d",
          6935 => x"53",
          6936 => x"51",
          6937 => x"3f",
          6938 => x"08",
          6939 => x"90",
          6940 => x"33",
          6941 => x"f7",
          6942 => x"e3",
          6943 => x"f8",
          6944 => x"fe",
          6945 => x"79",
          6946 => x"59",
          6947 => x"f4",
          6948 => x"79",
          6949 => x"b4",
          6950 => x"11",
          6951 => x"05",
          6952 => x"da",
          6953 => x"f0",
          6954 => x"91",
          6955 => x"02",
          6956 => x"33",
          6957 => x"81",
          6958 => x"b5",
          6959 => x"8c",
          6960 => x"e1",
          6961 => x"39",
          6962 => x"f4",
          6963 => x"84",
          6964 => x"e6",
          6965 => x"fe",
          6966 => x"2e",
          6967 => x"b4",
          6968 => x"11",
          6969 => x"05",
          6970 => x"84",
          6971 => x"f0",
          6972 => x"a6",
          6973 => x"02",
          6974 => x"79",
          6975 => x"5b",
          6976 => x"b4",
          6977 => x"11",
          6978 => x"05",
          6979 => x"e0",
          6980 => x"f0",
          6981 => x"f3",
          6982 => x"70",
          6983 => x"81",
          6984 => x"fe",
          6985 => x"80",
          6986 => x"51",
          6987 => x"3f",
          6988 => x"33",
          6989 => x"2e",
          6990 => x"78",
          6991 => x"38",
          6992 => x"41",
          6993 => x"3d",
          6994 => x"53",
          6995 => x"51",
          6996 => x"3f",
          6997 => x"08",
          6998 => x"38",
          6999 => x"be",
          7000 => x"70",
          7001 => x"23",
          7002 => x"ae",
          7003 => x"8c",
          7004 => x"b1",
          7005 => x"39",
          7006 => x"f4",
          7007 => x"84",
          7008 => x"e4",
          7009 => x"fe",
          7010 => x"2e",
          7011 => x"b4",
          7012 => x"11",
          7013 => x"05",
          7014 => x"d4",
          7015 => x"f0",
          7016 => x"a1",
          7017 => x"71",
          7018 => x"84",
          7019 => x"3d",
          7020 => x"53",
          7021 => x"51",
          7022 => x"3f",
          7023 => x"08",
          7024 => x"bc",
          7025 => x"08",
          7026 => x"f7",
          7027 => x"e0",
          7028 => x"f8",
          7029 => x"fe",
          7030 => x"79",
          7031 => x"59",
          7032 => x"f2",
          7033 => x"79",
          7034 => x"b4",
          7035 => x"11",
          7036 => x"05",
          7037 => x"f8",
          7038 => x"f0",
          7039 => x"8d",
          7040 => x"71",
          7041 => x"84",
          7042 => x"b9",
          7043 => x"8c",
          7044 => x"91",
          7045 => x"39",
          7046 => x"51",
          7047 => x"3f",
          7048 => x"d4",
          7049 => x"d8",
          7050 => x"c4",
          7051 => x"f5",
          7052 => x"fe",
          7053 => x"f1",
          7054 => x"f7",
          7055 => x"d9",
          7056 => x"80",
          7057 => x"c0",
          7058 => x"84",
          7059 => x"87",
          7060 => x"0c",
          7061 => x"81",
          7062 => x"fe",
          7063 => x"8c",
          7064 => x"87",
          7065 => x"0c",
          7066 => x"0b",
          7067 => x"94",
          7068 => x"39",
          7069 => x"80",
          7070 => x"84",
          7071 => x"e0",
          7072 => x"fe",
          7073 => x"2e",
          7074 => x"63",
          7075 => x"84",
          7076 => x"f5",
          7077 => x"78",
          7078 => x"ff",
          7079 => x"ff",
          7080 => x"fe",
          7081 => x"81",
          7082 => x"80",
          7083 => x"38",
          7084 => x"f8",
          7085 => x"de",
          7086 => x"59",
          7087 => x"fe",
          7088 => x"2e",
          7089 => x"81",
          7090 => x"52",
          7091 => x"51",
          7092 => x"3f",
          7093 => x"81",
          7094 => x"fe",
          7095 => x"fe",
          7096 => x"f0",
          7097 => x"f8",
          7098 => x"d8",
          7099 => x"59",
          7100 => x"fe",
          7101 => x"f0",
          7102 => x"45",
          7103 => x"78",
          7104 => x"fc",
          7105 => x"06",
          7106 => x"2e",
          7107 => x"b4",
          7108 => x"05",
          7109 => x"8a",
          7110 => x"f0",
          7111 => x"5c",
          7112 => x"b2",
          7113 => x"24",
          7114 => x"81",
          7115 => x"80",
          7116 => x"83",
          7117 => x"80",
          7118 => x"f9",
          7119 => x"55",
          7120 => x"54",
          7121 => x"f9",
          7122 => x"3d",
          7123 => x"51",
          7124 => x"3f",
          7125 => x"f9",
          7126 => x"3d",
          7127 => x"51",
          7128 => x"3f",
          7129 => x"55",
          7130 => x"54",
          7131 => x"f9",
          7132 => x"3d",
          7133 => x"51",
          7134 => x"3f",
          7135 => x"54",
          7136 => x"f9",
          7137 => x"3d",
          7138 => x"51",
          7139 => x"3f",
          7140 => x"58",
          7141 => x"57",
          7142 => x"55",
          7143 => x"80",
          7144 => x"80",
          7145 => x"3d",
          7146 => x"51",
          7147 => x"81",
          7148 => x"81",
          7149 => x"09",
          7150 => x"72",
          7151 => x"51",
          7152 => x"80",
          7153 => x"26",
          7154 => x"5a",
          7155 => x"59",
          7156 => x"8d",
          7157 => x"70",
          7158 => x"5d",
          7159 => x"c0",
          7160 => x"32",
          7161 => x"07",
          7162 => x"38",
          7163 => x"09",
          7164 => x"8c",
          7165 => x"b4",
          7166 => x"8d",
          7167 => x"39",
          7168 => x"80",
          7169 => x"b8",
          7170 => x"94",
          7171 => x"54",
          7172 => x"80",
          7173 => x"fe",
          7174 => x"81",
          7175 => x"90",
          7176 => x"55",
          7177 => x"80",
          7178 => x"fe",
          7179 => x"72",
          7180 => x"08",
          7181 => x"87",
          7182 => x"70",
          7183 => x"87",
          7184 => x"72",
          7185 => x"e3",
          7186 => x"f0",
          7187 => x"75",
          7188 => x"87",
          7189 => x"73",
          7190 => x"cf",
          7191 => x"fe",
          7192 => x"75",
          7193 => x"83",
          7194 => x"94",
          7195 => x"80",
          7196 => x"c0",
          7197 => x"a3",
          7198 => x"ff",
          7199 => x"8c",
          7200 => x"88",
          7201 => x"ad",
          7202 => x"95",
          7203 => x"c4",
          7204 => x"91",
          7205 => x"d0",
          7206 => x"89",
          7207 => x"e4",
          7208 => x"b7",
          7209 => x"e7",
          7210 => x"84",
          7211 => x"00",
          7212 => x"ff",
          7213 => x"ff",
          7214 => x"ff",
          7215 => x"00",
          7216 => x"32",
          7217 => x"38",
          7218 => x"3e",
          7219 => x"44",
          7220 => x"4a",
          7221 => x"f6",
          7222 => x"d2",
          7223 => x"75",
          7224 => x"b5",
          7225 => x"d8",
          7226 => x"65",
          7227 => x"cb",
          7228 => x"cb",
          7229 => x"a2",
          7230 => x"18",
          7231 => x"a3",
          7232 => x"cc",
          7233 => x"ea",
          7234 => x"6e",
          7235 => x"75",
          7236 => x"7c",
          7237 => x"83",
          7238 => x"8a",
          7239 => x"91",
          7240 => x"98",
          7241 => x"9f",
          7242 => x"a6",
          7243 => x"ad",
          7244 => x"b4",
          7245 => x"ba",
          7246 => x"c0",
          7247 => x"c6",
          7248 => x"cc",
          7249 => x"d2",
          7250 => x"d8",
          7251 => x"de",
          7252 => x"e4",
          7253 => x"25",
          7254 => x"64",
          7255 => x"3a",
          7256 => x"25",
          7257 => x"64",
          7258 => x"00",
          7259 => x"20",
          7260 => x"66",
          7261 => x"72",
          7262 => x"6f",
          7263 => x"00",
          7264 => x"72",
          7265 => x"53",
          7266 => x"63",
          7267 => x"69",
          7268 => x"00",
          7269 => x"65",
          7270 => x"65",
          7271 => x"6d",
          7272 => x"6d",
          7273 => x"65",
          7274 => x"00",
          7275 => x"20",
          7276 => x"53",
          7277 => x"4d",
          7278 => x"25",
          7279 => x"3a",
          7280 => x"58",
          7281 => x"00",
          7282 => x"20",
          7283 => x"41",
          7284 => x"20",
          7285 => x"25",
          7286 => x"3a",
          7287 => x"58",
          7288 => x"00",
          7289 => x"20",
          7290 => x"4e",
          7291 => x"41",
          7292 => x"25",
          7293 => x"3a",
          7294 => x"58",
          7295 => x"00",
          7296 => x"20",
          7297 => x"4d",
          7298 => x"20",
          7299 => x"25",
          7300 => x"3a",
          7301 => x"58",
          7302 => x"00",
          7303 => x"20",
          7304 => x"20",
          7305 => x"20",
          7306 => x"25",
          7307 => x"3a",
          7308 => x"58",
          7309 => x"00",
          7310 => x"20",
          7311 => x"43",
          7312 => x"20",
          7313 => x"44",
          7314 => x"63",
          7315 => x"3d",
          7316 => x"64",
          7317 => x"00",
          7318 => x"20",
          7319 => x"45",
          7320 => x"20",
          7321 => x"54",
          7322 => x"72",
          7323 => x"3d",
          7324 => x"64",
          7325 => x"00",
          7326 => x"20",
          7327 => x"52",
          7328 => x"52",
          7329 => x"43",
          7330 => x"6e",
          7331 => x"3d",
          7332 => x"64",
          7333 => x"00",
          7334 => x"20",
          7335 => x"48",
          7336 => x"45",
          7337 => x"53",
          7338 => x"00",
          7339 => x"20",
          7340 => x"49",
          7341 => x"00",
          7342 => x"20",
          7343 => x"54",
          7344 => x"00",
          7345 => x"20",
          7346 => x"0a",
          7347 => x"00",
          7348 => x"20",
          7349 => x"0a",
          7350 => x"00",
          7351 => x"72",
          7352 => x"65",
          7353 => x"00",
          7354 => x"20",
          7355 => x"20",
          7356 => x"65",
          7357 => x"65",
          7358 => x"72",
          7359 => x"64",
          7360 => x"73",
          7361 => x"25",
          7362 => x"0a",
          7363 => x"00",
          7364 => x"20",
          7365 => x"20",
          7366 => x"6f",
          7367 => x"53",
          7368 => x"74",
          7369 => x"64",
          7370 => x"73",
          7371 => x"25",
          7372 => x"0a",
          7373 => x"00",
          7374 => x"20",
          7375 => x"63",
          7376 => x"74",
          7377 => x"20",
          7378 => x"72",
          7379 => x"20",
          7380 => x"20",
          7381 => x"25",
          7382 => x"0a",
          7383 => x"00",
          7384 => x"63",
          7385 => x"00",
          7386 => x"20",
          7387 => x"20",
          7388 => x"20",
          7389 => x"20",
          7390 => x"20",
          7391 => x"20",
          7392 => x"20",
          7393 => x"25",
          7394 => x"0a",
          7395 => x"00",
          7396 => x"20",
          7397 => x"74",
          7398 => x"43",
          7399 => x"6b",
          7400 => x"65",
          7401 => x"20",
          7402 => x"20",
          7403 => x"25",
          7404 => x"30",
          7405 => x"48",
          7406 => x"00",
          7407 => x"20",
          7408 => x"41",
          7409 => x"6c",
          7410 => x"20",
          7411 => x"71",
          7412 => x"20",
          7413 => x"20",
          7414 => x"25",
          7415 => x"30",
          7416 => x"48",
          7417 => x"00",
          7418 => x"20",
          7419 => x"68",
          7420 => x"65",
          7421 => x"52",
          7422 => x"43",
          7423 => x"6b",
          7424 => x"65",
          7425 => x"25",
          7426 => x"30",
          7427 => x"48",
          7428 => x"00",
          7429 => x"6c",
          7430 => x"00",
          7431 => x"69",
          7432 => x"00",
          7433 => x"78",
          7434 => x"00",
          7435 => x"00",
          7436 => x"6d",
          7437 => x"00",
          7438 => x"6e",
          7439 => x"00",
          7440 => x"74",
          7441 => x"2e",
          7442 => x"00",
          7443 => x"74",
          7444 => x"00",
          7445 => x"74",
          7446 => x"00",
          7447 => x"00",
          7448 => x"64",
          7449 => x"73",
          7450 => x"00",
          7451 => x"6c",
          7452 => x"74",
          7453 => x"65",
          7454 => x"20",
          7455 => x"20",
          7456 => x"74",
          7457 => x"20",
          7458 => x"65",
          7459 => x"20",
          7460 => x"2e",
          7461 => x"00",
          7462 => x"6e",
          7463 => x"6f",
          7464 => x"2f",
          7465 => x"61",
          7466 => x"68",
          7467 => x"6f",
          7468 => x"66",
          7469 => x"2c",
          7470 => x"73",
          7471 => x"69",
          7472 => x"0a",
          7473 => x"00",
          7474 => x"74",
          7475 => x"00",
          7476 => x"01",
          7477 => x"70",
          7478 => x"00",
          7479 => x"02",
          7480 => x"6c",
          7481 => x"00",
          7482 => x"03",
          7483 => x"68",
          7484 => x"00",
          7485 => x"04",
          7486 => x"64",
          7487 => x"00",
          7488 => x"05",
          7489 => x"60",
          7490 => x"00",
          7491 => x"06",
          7492 => x"5c",
          7493 => x"00",
          7494 => x"07",
          7495 => x"58",
          7496 => x"00",
          7497 => x"08",
          7498 => x"54",
          7499 => x"00",
          7500 => x"09",
          7501 => x"50",
          7502 => x"00",
          7503 => x"0a",
          7504 => x"4c",
          7505 => x"00",
          7506 => x"0b",
          7507 => x"00",
          7508 => x"00",
          7509 => x"00",
          7510 => x"00",
          7511 => x"7e",
          7512 => x"7e",
          7513 => x"7e",
          7514 => x"7e",
          7515 => x"7e",
          7516 => x"00",
          7517 => x"00",
          7518 => x"00",
          7519 => x"2c",
          7520 => x"3d",
          7521 => x"5d",
          7522 => x"00",
          7523 => x"00",
          7524 => x"33",
          7525 => x"00",
          7526 => x"4d",
          7527 => x"53",
          7528 => x"00",
          7529 => x"4e",
          7530 => x"20",
          7531 => x"46",
          7532 => x"32",
          7533 => x"00",
          7534 => x"4e",
          7535 => x"20",
          7536 => x"46",
          7537 => x"20",
          7538 => x"00",
          7539 => x"78",
          7540 => x"00",
          7541 => x"00",
          7542 => x"00",
          7543 => x"41",
          7544 => x"80",
          7545 => x"49",
          7546 => x"8f",
          7547 => x"4f",
          7548 => x"55",
          7549 => x"9b",
          7550 => x"9f",
          7551 => x"55",
          7552 => x"a7",
          7553 => x"ab",
          7554 => x"af",
          7555 => x"b3",
          7556 => x"b7",
          7557 => x"bb",
          7558 => x"bf",
          7559 => x"c3",
          7560 => x"c7",
          7561 => x"cb",
          7562 => x"cf",
          7563 => x"d3",
          7564 => x"d7",
          7565 => x"db",
          7566 => x"df",
          7567 => x"e3",
          7568 => x"e7",
          7569 => x"eb",
          7570 => x"ef",
          7571 => x"f3",
          7572 => x"f7",
          7573 => x"fb",
          7574 => x"ff",
          7575 => x"3b",
          7576 => x"2f",
          7577 => x"3a",
          7578 => x"7c",
          7579 => x"00",
          7580 => x"04",
          7581 => x"40",
          7582 => x"00",
          7583 => x"00",
          7584 => x"02",
          7585 => x"08",
          7586 => x"20",
          7587 => x"00",
          7588 => x"69",
          7589 => x"00",
          7590 => x"63",
          7591 => x"00",
          7592 => x"69",
          7593 => x"00",
          7594 => x"61",
          7595 => x"00",
          7596 => x"65",
          7597 => x"00",
          7598 => x"65",
          7599 => x"00",
          7600 => x"70",
          7601 => x"00",
          7602 => x"66",
          7603 => x"00",
          7604 => x"6d",
          7605 => x"00",
          7606 => x"00",
          7607 => x"00",
          7608 => x"00",
          7609 => x"00",
          7610 => x"00",
          7611 => x"00",
          7612 => x"00",
          7613 => x"6c",
          7614 => x"00",
          7615 => x"00",
          7616 => x"74",
          7617 => x"00",
          7618 => x"65",
          7619 => x"00",
          7620 => x"6f",
          7621 => x"00",
          7622 => x"74",
          7623 => x"00",
          7624 => x"73",
          7625 => x"00",
          7626 => x"73",
          7627 => x"00",
          7628 => x"6f",
          7629 => x"00",
          7630 => x"6b",
          7631 => x"72",
          7632 => x"00",
          7633 => x"65",
          7634 => x"6c",
          7635 => x"72",
          7636 => x"0a",
          7637 => x"00",
          7638 => x"6b",
          7639 => x"74",
          7640 => x"61",
          7641 => x"0a",
          7642 => x"00",
          7643 => x"66",
          7644 => x"20",
          7645 => x"6e",
          7646 => x"00",
          7647 => x"70",
          7648 => x"20",
          7649 => x"6e",
          7650 => x"00",
          7651 => x"61",
          7652 => x"20",
          7653 => x"65",
          7654 => x"65",
          7655 => x"00",
          7656 => x"65",
          7657 => x"64",
          7658 => x"65",
          7659 => x"00",
          7660 => x"65",
          7661 => x"72",
          7662 => x"79",
          7663 => x"69",
          7664 => x"2e",
          7665 => x"00",
          7666 => x"65",
          7667 => x"6e",
          7668 => x"20",
          7669 => x"61",
          7670 => x"2e",
          7671 => x"00",
          7672 => x"69",
          7673 => x"72",
          7674 => x"20",
          7675 => x"74",
          7676 => x"65",
          7677 => x"00",
          7678 => x"76",
          7679 => x"75",
          7680 => x"72",
          7681 => x"20",
          7682 => x"61",
          7683 => x"2e",
          7684 => x"00",
          7685 => x"6b",
          7686 => x"74",
          7687 => x"61",
          7688 => x"64",
          7689 => x"00",
          7690 => x"63",
          7691 => x"61",
          7692 => x"6c",
          7693 => x"69",
          7694 => x"79",
          7695 => x"6d",
          7696 => x"75",
          7697 => x"6f",
          7698 => x"69",
          7699 => x"0a",
          7700 => x"00",
          7701 => x"6d",
          7702 => x"61",
          7703 => x"74",
          7704 => x"0a",
          7705 => x"00",
          7706 => x"65",
          7707 => x"2c",
          7708 => x"65",
          7709 => x"69",
          7710 => x"63",
          7711 => x"65",
          7712 => x"64",
          7713 => x"00",
          7714 => x"65",
          7715 => x"20",
          7716 => x"6b",
          7717 => x"0a",
          7718 => x"00",
          7719 => x"75",
          7720 => x"63",
          7721 => x"74",
          7722 => x"6d",
          7723 => x"2e",
          7724 => x"00",
          7725 => x"20",
          7726 => x"79",
          7727 => x"65",
          7728 => x"69",
          7729 => x"2e",
          7730 => x"00",
          7731 => x"61",
          7732 => x"65",
          7733 => x"69",
          7734 => x"72",
          7735 => x"74",
          7736 => x"00",
          7737 => x"63",
          7738 => x"2e",
          7739 => x"00",
          7740 => x"6e",
          7741 => x"20",
          7742 => x"6f",
          7743 => x"00",
          7744 => x"75",
          7745 => x"74",
          7746 => x"25",
          7747 => x"74",
          7748 => x"75",
          7749 => x"74",
          7750 => x"73",
          7751 => x"0a",
          7752 => x"00",
          7753 => x"64",
          7754 => x"00",
          7755 => x"58",
          7756 => x"00",
          7757 => x"00",
          7758 => x"58",
          7759 => x"00",
          7760 => x"20",
          7761 => x"20",
          7762 => x"00",
          7763 => x"58",
          7764 => x"00",
          7765 => x"00",
          7766 => x"00",
          7767 => x"00",
          7768 => x"54",
          7769 => x"00",
          7770 => x"20",
          7771 => x"28",
          7772 => x"00",
          7773 => x"30",
          7774 => x"30",
          7775 => x"00",
          7776 => x"35",
          7777 => x"00",
          7778 => x"55",
          7779 => x"65",
          7780 => x"30",
          7781 => x"20",
          7782 => x"25",
          7783 => x"2a",
          7784 => x"00",
          7785 => x"54",
          7786 => x"6e",
          7787 => x"72",
          7788 => x"20",
          7789 => x"64",
          7790 => x"0a",
          7791 => x"00",
          7792 => x"65",
          7793 => x"6e",
          7794 => x"72",
          7795 => x"0a",
          7796 => x"00",
          7797 => x"20",
          7798 => x"65",
          7799 => x"70",
          7800 => x"00",
          7801 => x"54",
          7802 => x"44",
          7803 => x"74",
          7804 => x"75",
          7805 => x"00",
          7806 => x"54",
          7807 => x"52",
          7808 => x"74",
          7809 => x"75",
          7810 => x"00",
          7811 => x"54",
          7812 => x"58",
          7813 => x"74",
          7814 => x"75",
          7815 => x"00",
          7816 => x"54",
          7817 => x"58",
          7818 => x"74",
          7819 => x"75",
          7820 => x"00",
          7821 => x"54",
          7822 => x"58",
          7823 => x"74",
          7824 => x"75",
          7825 => x"00",
          7826 => x"54",
          7827 => x"58",
          7828 => x"74",
          7829 => x"75",
          7830 => x"00",
          7831 => x"74",
          7832 => x"20",
          7833 => x"74",
          7834 => x"72",
          7835 => x"0a",
          7836 => x"00",
          7837 => x"62",
          7838 => x"67",
          7839 => x"6d",
          7840 => x"2e",
          7841 => x"00",
          7842 => x"6f",
          7843 => x"63",
          7844 => x"74",
          7845 => x"00",
          7846 => x"00",
          7847 => x"6c",
          7848 => x"74",
          7849 => x"6e",
          7850 => x"61",
          7851 => x"65",
          7852 => x"20",
          7853 => x"64",
          7854 => x"20",
          7855 => x"61",
          7856 => x"69",
          7857 => x"20",
          7858 => x"75",
          7859 => x"79",
          7860 => x"00",
          7861 => x"00",
          7862 => x"20",
          7863 => x"6b",
          7864 => x"21",
          7865 => x"00",
          7866 => x"74",
          7867 => x"69",
          7868 => x"2e",
          7869 => x"00",
          7870 => x"6c",
          7871 => x"74",
          7872 => x"6e",
          7873 => x"61",
          7874 => x"65",
          7875 => x"00",
          7876 => x"25",
          7877 => x"00",
          7878 => x"00",
          7879 => x"61",
          7880 => x"67",
          7881 => x"2e",
          7882 => x"00",
          7883 => x"79",
          7884 => x"2e",
          7885 => x"00",
          7886 => x"70",
          7887 => x"6e",
          7888 => x"2e",
          7889 => x"00",
          7890 => x"6c",
          7891 => x"30",
          7892 => x"2d",
          7893 => x"38",
          7894 => x"25",
          7895 => x"29",
          7896 => x"00",
          7897 => x"70",
          7898 => x"6d",
          7899 => x"0a",
          7900 => x"00",
          7901 => x"6d",
          7902 => x"74",
          7903 => x"00",
          7904 => x"58",
          7905 => x"32",
          7906 => x"00",
          7907 => x"0a",
          7908 => x"00",
          7909 => x"58",
          7910 => x"34",
          7911 => x"00",
          7912 => x"58",
          7913 => x"38",
          7914 => x"00",
          7915 => x"61",
          7916 => x"6e",
          7917 => x"6e",
          7918 => x"72",
          7919 => x"73",
          7920 => x"00",
          7921 => x"62",
          7922 => x"67",
          7923 => x"74",
          7924 => x"75",
          7925 => x"0a",
          7926 => x"00",
          7927 => x"61",
          7928 => x"64",
          7929 => x"72",
          7930 => x"69",
          7931 => x"00",
          7932 => x"62",
          7933 => x"67",
          7934 => x"72",
          7935 => x"69",
          7936 => x"00",
          7937 => x"63",
          7938 => x"6e",
          7939 => x"6f",
          7940 => x"40",
          7941 => x"38",
          7942 => x"2e",
          7943 => x"00",
          7944 => x"6c",
          7945 => x"20",
          7946 => x"65",
          7947 => x"25",
          7948 => x"20",
          7949 => x"0a",
          7950 => x"00",
          7951 => x"6c",
          7952 => x"74",
          7953 => x"65",
          7954 => x"6f",
          7955 => x"28",
          7956 => x"2e",
          7957 => x"00",
          7958 => x"74",
          7959 => x"69",
          7960 => x"61",
          7961 => x"69",
          7962 => x"69",
          7963 => x"2e",
          7964 => x"00",
          7965 => x"64",
          7966 => x"62",
          7967 => x"69",
          7968 => x"2e",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"5c",
          7973 => x"25",
          7974 => x"73",
          7975 => x"00",
          7976 => x"5c",
          7977 => x"25",
          7978 => x"00",
          7979 => x"5c",
          7980 => x"00",
          7981 => x"20",
          7982 => x"6d",
          7983 => x"2e",
          7984 => x"00",
          7985 => x"6e",
          7986 => x"2e",
          7987 => x"00",
          7988 => x"62",
          7989 => x"67",
          7990 => x"74",
          7991 => x"75",
          7992 => x"2e",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"ff",
          7997 => x"00",
          7998 => x"ff",
          7999 => x"00",
          8000 => x"ff",
          8001 => x"00",
          8002 => x"00",
          8003 => x"00",
          8004 => x"ff",
          8005 => x"00",
          8006 => x"00",
          8007 => x"00",
          8008 => x"00",
          8009 => x"00",
          8010 => x"00",
          8011 => x"00",
          8012 => x"00",
          8013 => x"01",
          8014 => x"01",
          8015 => x"01",
          8016 => x"00",
          8017 => x"00",
          8018 => x"02",
          8019 => x"00",
          8020 => x"48",
          8021 => x"48",
          8022 => x"48",
          8023 => x"48",
          8024 => x"40",
          8025 => x"00",
          8026 => x"00",
          8027 => x"00",
          8028 => x"00",
          8029 => x"00",
          8030 => x"00",
          8031 => x"00",
          8032 => x"00",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"4c",
          8049 => x"00",
          8050 => x"54",
          8051 => x"00",
          8052 => x"5c",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"90",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"98",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"a0",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"a8",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"b0",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"b8",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"c0",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"c8",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"d0",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"d8",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"dc",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"e0",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"e4",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"e8",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"ec",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"f0",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"f4",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"fc",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"08",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"10",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"18",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"20",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"28",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"30",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"92",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"81",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a3",
           270 => x"0b",
           271 => x"0b",
           272 => x"c1",
           273 => x"0b",
           274 => x"0b",
           275 => x"df",
           276 => x"0b",
           277 => x"0b",
           278 => x"fd",
           279 => x"0b",
           280 => x"0b",
           281 => x"9b",
           282 => x"0b",
           283 => x"0b",
           284 => x"b9",
           285 => x"0b",
           286 => x"0b",
           287 => x"d7",
           288 => x"0b",
           289 => x"0b",
           290 => x"f5",
           291 => x"0b",
           292 => x"0b",
           293 => x"93",
           294 => x"0b",
           295 => x"0b",
           296 => x"b3",
           297 => x"0b",
           298 => x"0b",
           299 => x"d3",
           300 => x"0b",
           301 => x"0b",
           302 => x"f3",
           303 => x"0b",
           304 => x"0b",
           305 => x"93",
           306 => x"0b",
           307 => x"0b",
           308 => x"b3",
           309 => x"0b",
           310 => x"0b",
           311 => x"d3",
           312 => x"0b",
           313 => x"0b",
           314 => x"f3",
           315 => x"0b",
           316 => x"0b",
           317 => x"93",
           318 => x"0b",
           319 => x"0b",
           320 => x"b3",
           321 => x"0b",
           322 => x"0b",
           323 => x"d3",
           324 => x"0b",
           325 => x"0b",
           326 => x"f3",
           327 => x"0b",
           328 => x"0b",
           329 => x"93",
           330 => x"0b",
           331 => x"0b",
           332 => x"b3",
           333 => x"0b",
           334 => x"0b",
           335 => x"d3",
           336 => x"0b",
           337 => x"0b",
           338 => x"f3",
           339 => x"0b",
           340 => x"0b",
           341 => x"91",
           342 => x"0b",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"fe",
           386 => x"ff",
           387 => x"fc",
           388 => x"90",
           389 => x"fc",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"81",
           395 => x"83",
           396 => x"81",
           397 => x"b6",
           398 => x"fe",
           399 => x"80",
           400 => x"fe",
           401 => x"e3",
           402 => x"fc",
           403 => x"90",
           404 => x"fc",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"81",
           410 => x"83",
           411 => x"81",
           412 => x"bd",
           413 => x"fe",
           414 => x"80",
           415 => x"fe",
           416 => x"f0",
           417 => x"fc",
           418 => x"90",
           419 => x"fc",
           420 => x"2d",
           421 => x"08",
           422 => x"04",
           423 => x"0c",
           424 => x"81",
           425 => x"83",
           426 => x"81",
           427 => x"bc",
           428 => x"fe",
           429 => x"80",
           430 => x"fe",
           431 => x"c3",
           432 => x"fc",
           433 => x"90",
           434 => x"fc",
           435 => x"2d",
           436 => x"08",
           437 => x"04",
           438 => x"0c",
           439 => x"81",
           440 => x"83",
           441 => x"81",
           442 => x"9e",
           443 => x"fe",
           444 => x"80",
           445 => x"fe",
           446 => x"ae",
           447 => x"fc",
           448 => x"90",
           449 => x"fc",
           450 => x"2d",
           451 => x"08",
           452 => x"04",
           453 => x"0c",
           454 => x"2d",
           455 => x"08",
           456 => x"04",
           457 => x"0c",
           458 => x"2d",
           459 => x"08",
           460 => x"04",
           461 => x"0c",
           462 => x"2d",
           463 => x"08",
           464 => x"04",
           465 => x"0c",
           466 => x"2d",
           467 => x"08",
           468 => x"04",
           469 => x"0c",
           470 => x"2d",
           471 => x"08",
           472 => x"04",
           473 => x"0c",
           474 => x"2d",
           475 => x"08",
           476 => x"04",
           477 => x"0c",
           478 => x"2d",
           479 => x"08",
           480 => x"04",
           481 => x"0c",
           482 => x"2d",
           483 => x"08",
           484 => x"04",
           485 => x"0c",
           486 => x"2d",
           487 => x"08",
           488 => x"04",
           489 => x"0c",
           490 => x"2d",
           491 => x"08",
           492 => x"04",
           493 => x"0c",
           494 => x"2d",
           495 => x"08",
           496 => x"04",
           497 => x"0c",
           498 => x"2d",
           499 => x"08",
           500 => x"04",
           501 => x"0c",
           502 => x"2d",
           503 => x"08",
           504 => x"04",
           505 => x"0c",
           506 => x"2d",
           507 => x"08",
           508 => x"04",
           509 => x"0c",
           510 => x"2d",
           511 => x"08",
           512 => x"04",
           513 => x"0c",
           514 => x"2d",
           515 => x"08",
           516 => x"04",
           517 => x"0c",
           518 => x"2d",
           519 => x"08",
           520 => x"04",
           521 => x"0c",
           522 => x"2d",
           523 => x"08",
           524 => x"04",
           525 => x"0c",
           526 => x"2d",
           527 => x"08",
           528 => x"04",
           529 => x"0c",
           530 => x"2d",
           531 => x"08",
           532 => x"04",
           533 => x"0c",
           534 => x"2d",
           535 => x"08",
           536 => x"04",
           537 => x"0c",
           538 => x"2d",
           539 => x"08",
           540 => x"04",
           541 => x"0c",
           542 => x"2d",
           543 => x"08",
           544 => x"04",
           545 => x"0c",
           546 => x"2d",
           547 => x"08",
           548 => x"04",
           549 => x"0c",
           550 => x"2d",
           551 => x"08",
           552 => x"04",
           553 => x"0c",
           554 => x"2d",
           555 => x"08",
           556 => x"04",
           557 => x"0c",
           558 => x"2d",
           559 => x"08",
           560 => x"04",
           561 => x"0c",
           562 => x"2d",
           563 => x"08",
           564 => x"04",
           565 => x"0c",
           566 => x"2d",
           567 => x"08",
           568 => x"04",
           569 => x"0c",
           570 => x"2d",
           571 => x"08",
           572 => x"04",
           573 => x"0c",
           574 => x"81",
           575 => x"83",
           576 => x"81",
           577 => x"a0",
           578 => x"fe",
           579 => x"80",
           580 => x"fe",
           581 => x"f1",
           582 => x"fc",
           583 => x"90",
           584 => x"fc",
           585 => x"d8",
           586 => x"fc",
           587 => x"90",
           588 => x"00",
           589 => x"10",
           590 => x"10",
           591 => x"10",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"00",
           598 => x"ff",
           599 => x"06",
           600 => x"83",
           601 => x"10",
           602 => x"fc",
           603 => x"51",
           604 => x"80",
           605 => x"ff",
           606 => x"06",
           607 => x"52",
           608 => x"0a",
           609 => x"38",
           610 => x"51",
           611 => x"f0",
           612 => x"b0",
           613 => x"80",
           614 => x"05",
           615 => x"0b",
           616 => x"04",
           617 => x"81",
           618 => x"00",
           619 => x"08",
           620 => x"fc",
           621 => x"0d",
           622 => x"fe",
           623 => x"05",
           624 => x"fe",
           625 => x"05",
           626 => x"d4",
           627 => x"f0",
           628 => x"fe",
           629 => x"85",
           630 => x"fe",
           631 => x"81",
           632 => x"02",
           633 => x"0c",
           634 => x"81",
           635 => x"fc",
           636 => x"08",
           637 => x"fc",
           638 => x"08",
           639 => x"3f",
           640 => x"08",
           641 => x"f0",
           642 => x"3d",
           643 => x"fc",
           644 => x"fe",
           645 => x"81",
           646 => x"f9",
           647 => x"0b",
           648 => x"08",
           649 => x"81",
           650 => x"88",
           651 => x"25",
           652 => x"fe",
           653 => x"05",
           654 => x"fe",
           655 => x"05",
           656 => x"81",
           657 => x"f4",
           658 => x"fe",
           659 => x"05",
           660 => x"81",
           661 => x"fc",
           662 => x"0c",
           663 => x"08",
           664 => x"81",
           665 => x"fc",
           666 => x"fe",
           667 => x"05",
           668 => x"b9",
           669 => x"fc",
           670 => x"08",
           671 => x"fc",
           672 => x"0c",
           673 => x"fe",
           674 => x"05",
           675 => x"fc",
           676 => x"08",
           677 => x"0b",
           678 => x"08",
           679 => x"81",
           680 => x"f0",
           681 => x"fe",
           682 => x"05",
           683 => x"81",
           684 => x"8c",
           685 => x"81",
           686 => x"88",
           687 => x"81",
           688 => x"fe",
           689 => x"81",
           690 => x"f8",
           691 => x"81",
           692 => x"fc",
           693 => x"2e",
           694 => x"fe",
           695 => x"05",
           696 => x"fe",
           697 => x"05",
           698 => x"fc",
           699 => x"08",
           700 => x"f0",
           701 => x"3d",
           702 => x"fc",
           703 => x"fe",
           704 => x"81",
           705 => x"fb",
           706 => x"0b",
           707 => x"08",
           708 => x"81",
           709 => x"88",
           710 => x"25",
           711 => x"fe",
           712 => x"05",
           713 => x"fe",
           714 => x"05",
           715 => x"81",
           716 => x"fc",
           717 => x"fe",
           718 => x"05",
           719 => x"90",
           720 => x"fc",
           721 => x"08",
           722 => x"fc",
           723 => x"0c",
           724 => x"fe",
           725 => x"05",
           726 => x"fe",
           727 => x"05",
           728 => x"3f",
           729 => x"08",
           730 => x"fc",
           731 => x"0c",
           732 => x"fc",
           733 => x"08",
           734 => x"38",
           735 => x"08",
           736 => x"30",
           737 => x"08",
           738 => x"81",
           739 => x"f8",
           740 => x"81",
           741 => x"54",
           742 => x"81",
           743 => x"04",
           744 => x"08",
           745 => x"fc",
           746 => x"0d",
           747 => x"fe",
           748 => x"05",
           749 => x"81",
           750 => x"f8",
           751 => x"fe",
           752 => x"05",
           753 => x"fc",
           754 => x"08",
           755 => x"81",
           756 => x"fc",
           757 => x"2e",
           758 => x"0b",
           759 => x"08",
           760 => x"24",
           761 => x"fe",
           762 => x"05",
           763 => x"fe",
           764 => x"05",
           765 => x"fc",
           766 => x"08",
           767 => x"fc",
           768 => x"0c",
           769 => x"81",
           770 => x"fc",
           771 => x"2e",
           772 => x"81",
           773 => x"8c",
           774 => x"fe",
           775 => x"05",
           776 => x"38",
           777 => x"08",
           778 => x"81",
           779 => x"8c",
           780 => x"81",
           781 => x"88",
           782 => x"fe",
           783 => x"05",
           784 => x"fc",
           785 => x"08",
           786 => x"fc",
           787 => x"0c",
           788 => x"08",
           789 => x"81",
           790 => x"fc",
           791 => x"0c",
           792 => x"08",
           793 => x"81",
           794 => x"fc",
           795 => x"0c",
           796 => x"81",
           797 => x"90",
           798 => x"2e",
           799 => x"fe",
           800 => x"05",
           801 => x"fe",
           802 => x"05",
           803 => x"39",
           804 => x"08",
           805 => x"70",
           806 => x"08",
           807 => x"51",
           808 => x"08",
           809 => x"81",
           810 => x"85",
           811 => x"fe",
           812 => x"fc",
           813 => x"70",
           814 => x"55",
           815 => x"72",
           816 => x"72",
           817 => x"06",
           818 => x"2e",
           819 => x"12",
           820 => x"2e",
           821 => x"70",
           822 => x"33",
           823 => x"05",
           824 => x"12",
           825 => x"2e",
           826 => x"ea",
           827 => x"fe",
           828 => x"3d",
           829 => x"51",
           830 => x"05",
           831 => x"70",
           832 => x"0c",
           833 => x"05",
           834 => x"70",
           835 => x"0c",
           836 => x"05",
           837 => x"70",
           838 => x"0c",
           839 => x"05",
           840 => x"70",
           841 => x"0c",
           842 => x"71",
           843 => x"38",
           844 => x"95",
           845 => x"84",
           846 => x"71",
           847 => x"53",
           848 => x"52",
           849 => x"ed",
           850 => x"ff",
           851 => x"3d",
           852 => x"71",
           853 => x"9f",
           854 => x"55",
           855 => x"72",
           856 => x"74",
           857 => x"70",
           858 => x"38",
           859 => x"71",
           860 => x"38",
           861 => x"81",
           862 => x"ff",
           863 => x"ff",
           864 => x"06",
           865 => x"81",
           866 => x"86",
           867 => x"74",
           868 => x"75",
           869 => x"90",
           870 => x"54",
           871 => x"27",
           872 => x"71",
           873 => x"53",
           874 => x"70",
           875 => x"0c",
           876 => x"84",
           877 => x"72",
           878 => x"05",
           879 => x"12",
           880 => x"26",
           881 => x"72",
           882 => x"72",
           883 => x"05",
           884 => x"12",
           885 => x"26",
           886 => x"53",
           887 => x"fc",
           888 => x"70",
           889 => x"07",
           890 => x"54",
           891 => x"80",
           892 => x"70",
           893 => x"70",
           894 => x"ff",
           895 => x"f8",
           896 => x"80",
           897 => x"53",
           898 => x"a6",
           899 => x"72",
           900 => x"05",
           901 => x"08",
           902 => x"f7",
           903 => x"13",
           904 => x"84",
           905 => x"06",
           906 => x"53",
           907 => x"2e",
           908 => x"52",
           909 => x"05",
           910 => x"70",
           911 => x"05",
           912 => x"f0",
           913 => x"fe",
           914 => x"3d",
           915 => x"3d",
           916 => x"71",
           917 => x"55",
           918 => x"38",
           919 => x"70",
           920 => x"fd",
           921 => x"70",
           922 => x"81",
           923 => x"51",
           924 => x"9d",
           925 => x"70",
           926 => x"f7",
           927 => x"12",
           928 => x"84",
           929 => x"06",
           930 => x"53",
           931 => x"e5",
           932 => x"71",
           933 => x"80",
           934 => x"81",
           935 => x"52",
           936 => x"38",
           937 => x"81",
           938 => x"85",
           939 => x"fa",
           940 => x"7a",
           941 => x"55",
           942 => x"80",
           943 => x"38",
           944 => x"83",
           945 => x"80",
           946 => x"38",
           947 => x"72",
           948 => x"38",
           949 => x"33",
           950 => x"71",
           951 => x"06",
           952 => x"80",
           953 => x"38",
           954 => x"06",
           955 => x"2e",
           956 => x"81",
           957 => x"ff",
           958 => x"52",
           959 => x"09",
           960 => x"38",
           961 => x"33",
           962 => x"81",
           963 => x"81",
           964 => x"71",
           965 => x"52",
           966 => x"f0",
           967 => x"0d",
           968 => x"57",
           969 => x"27",
           970 => x"08",
           971 => x"88",
           972 => x"55",
           973 => x"39",
           974 => x"72",
           975 => x"38",
           976 => x"09",
           977 => x"ff",
           978 => x"f8",
           979 => x"80",
           980 => x"51",
           981 => x"84",
           982 => x"57",
           983 => x"27",
           984 => x"08",
           985 => x"d0",
           986 => x"55",
           987 => x"39",
           988 => x"fe",
           989 => x"3d",
           990 => x"3d",
           991 => x"83",
           992 => x"2b",
           993 => x"3f",
           994 => x"08",
           995 => x"72",
           996 => x"54",
           997 => x"25",
           998 => x"81",
           999 => x"84",
          1000 => x"fb",
          1001 => x"70",
          1002 => x"53",
          1003 => x"2e",
          1004 => x"71",
          1005 => x"a0",
          1006 => x"06",
          1007 => x"12",
          1008 => x"71",
          1009 => x"81",
          1010 => x"73",
          1011 => x"ff",
          1012 => x"55",
          1013 => x"83",
          1014 => x"70",
          1015 => x"38",
          1016 => x"73",
          1017 => x"51",
          1018 => x"09",
          1019 => x"38",
          1020 => x"81",
          1021 => x"72",
          1022 => x"51",
          1023 => x"f0",
          1024 => x"0d",
          1025 => x"0d",
          1026 => x"08",
          1027 => x"38",
          1028 => x"05",
          1029 => x"9f",
          1030 => x"fe",
          1031 => x"38",
          1032 => x"39",
          1033 => x"81",
          1034 => x"86",
          1035 => x"fc",
          1036 => x"82",
          1037 => x"05",
          1038 => x"52",
          1039 => x"81",
          1040 => x"13",
          1041 => x"51",
          1042 => x"9e",
          1043 => x"38",
          1044 => x"51",
          1045 => x"97",
          1046 => x"38",
          1047 => x"51",
          1048 => x"bb",
          1049 => x"38",
          1050 => x"51",
          1051 => x"bb",
          1052 => x"38",
          1053 => x"55",
          1054 => x"87",
          1055 => x"d9",
          1056 => x"22",
          1057 => x"73",
          1058 => x"80",
          1059 => x"0b",
          1060 => x"9c",
          1061 => x"87",
          1062 => x"0c",
          1063 => x"87",
          1064 => x"0c",
          1065 => x"87",
          1066 => x"0c",
          1067 => x"87",
          1068 => x"0c",
          1069 => x"87",
          1070 => x"0c",
          1071 => x"87",
          1072 => x"0c",
          1073 => x"98",
          1074 => x"87",
          1075 => x"0c",
          1076 => x"c0",
          1077 => x"80",
          1078 => x"fe",
          1079 => x"3d",
          1080 => x"3d",
          1081 => x"87",
          1082 => x"5d",
          1083 => x"87",
          1084 => x"08",
          1085 => x"23",
          1086 => x"b8",
          1087 => x"82",
          1088 => x"c0",
          1089 => x"5a",
          1090 => x"34",
          1091 => x"b0",
          1092 => x"84",
          1093 => x"c0",
          1094 => x"5a",
          1095 => x"34",
          1096 => x"a8",
          1097 => x"86",
          1098 => x"c0",
          1099 => x"5c",
          1100 => x"23",
          1101 => x"a0",
          1102 => x"8a",
          1103 => x"7d",
          1104 => x"ff",
          1105 => x"7b",
          1106 => x"06",
          1107 => x"33",
          1108 => x"33",
          1109 => x"33",
          1110 => x"33",
          1111 => x"33",
          1112 => x"ff",
          1113 => x"81",
          1114 => x"99",
          1115 => x"3d",
          1116 => x"3d",
          1117 => x"05",
          1118 => x"70",
          1119 => x"52",
          1120 => x"0b",
          1121 => x"34",
          1122 => x"04",
          1123 => x"77",
          1124 => x"f9",
          1125 => x"81",
          1126 => x"55",
          1127 => x"94",
          1128 => x"80",
          1129 => x"87",
          1130 => x"51",
          1131 => x"96",
          1132 => x"06",
          1133 => x"70",
          1134 => x"38",
          1135 => x"70",
          1136 => x"51",
          1137 => x"72",
          1138 => x"81",
          1139 => x"70",
          1140 => x"38",
          1141 => x"70",
          1142 => x"51",
          1143 => x"38",
          1144 => x"06",
          1145 => x"94",
          1146 => x"80",
          1147 => x"87",
          1148 => x"52",
          1149 => x"75",
          1150 => x"0c",
          1151 => x"04",
          1152 => x"02",
          1153 => x"0b",
          1154 => x"e8",
          1155 => x"ff",
          1156 => x"56",
          1157 => x"84",
          1158 => x"2e",
          1159 => x"c0",
          1160 => x"70",
          1161 => x"2a",
          1162 => x"53",
          1163 => x"80",
          1164 => x"71",
          1165 => x"81",
          1166 => x"70",
          1167 => x"81",
          1168 => x"06",
          1169 => x"80",
          1170 => x"71",
          1171 => x"81",
          1172 => x"70",
          1173 => x"73",
          1174 => x"51",
          1175 => x"80",
          1176 => x"2e",
          1177 => x"c0",
          1178 => x"75",
          1179 => x"3d",
          1180 => x"3d",
          1181 => x"80",
          1182 => x"81",
          1183 => x"53",
          1184 => x"2e",
          1185 => x"71",
          1186 => x"81",
          1187 => x"81",
          1188 => x"70",
          1189 => x"59",
          1190 => x"87",
          1191 => x"51",
          1192 => x"86",
          1193 => x"94",
          1194 => x"08",
          1195 => x"70",
          1196 => x"54",
          1197 => x"2e",
          1198 => x"91",
          1199 => x"06",
          1200 => x"d7",
          1201 => x"32",
          1202 => x"51",
          1203 => x"2e",
          1204 => x"93",
          1205 => x"06",
          1206 => x"ff",
          1207 => x"81",
          1208 => x"87",
          1209 => x"52",
          1210 => x"86",
          1211 => x"94",
          1212 => x"72",
          1213 => x"74",
          1214 => x"ff",
          1215 => x"57",
          1216 => x"38",
          1217 => x"f0",
          1218 => x"0d",
          1219 => x"0d",
          1220 => x"f9",
          1221 => x"81",
          1222 => x"52",
          1223 => x"84",
          1224 => x"2e",
          1225 => x"c0",
          1226 => x"70",
          1227 => x"2a",
          1228 => x"51",
          1229 => x"80",
          1230 => x"71",
          1231 => x"51",
          1232 => x"80",
          1233 => x"2e",
          1234 => x"c0",
          1235 => x"71",
          1236 => x"ff",
          1237 => x"f0",
          1238 => x"3d",
          1239 => x"3d",
          1240 => x"81",
          1241 => x"70",
          1242 => x"52",
          1243 => x"94",
          1244 => x"80",
          1245 => x"87",
          1246 => x"52",
          1247 => x"82",
          1248 => x"06",
          1249 => x"ff",
          1250 => x"2e",
          1251 => x"81",
          1252 => x"87",
          1253 => x"52",
          1254 => x"86",
          1255 => x"94",
          1256 => x"08",
          1257 => x"70",
          1258 => x"53",
          1259 => x"fe",
          1260 => x"3d",
          1261 => x"3d",
          1262 => x"9e",
          1263 => x"9c",
          1264 => x"51",
          1265 => x"2e",
          1266 => x"87",
          1267 => x"08",
          1268 => x"0c",
          1269 => x"a8",
          1270 => x"f0",
          1271 => x"9e",
          1272 => x"f9",
          1273 => x"c0",
          1274 => x"81",
          1275 => x"87",
          1276 => x"08",
          1277 => x"0c",
          1278 => x"a0",
          1279 => x"80",
          1280 => x"9e",
          1281 => x"fa",
          1282 => x"c0",
          1283 => x"81",
          1284 => x"87",
          1285 => x"08",
          1286 => x"0c",
          1287 => x"b8",
          1288 => x"90",
          1289 => x"9e",
          1290 => x"fa",
          1291 => x"c0",
          1292 => x"81",
          1293 => x"87",
          1294 => x"08",
          1295 => x"0c",
          1296 => x"80",
          1297 => x"81",
          1298 => x"87",
          1299 => x"08",
          1300 => x"0c",
          1301 => x"88",
          1302 => x"a8",
          1303 => x"9e",
          1304 => x"fa",
          1305 => x"0b",
          1306 => x"34",
          1307 => x"c0",
          1308 => x"70",
          1309 => x"06",
          1310 => x"70",
          1311 => x"38",
          1312 => x"81",
          1313 => x"80",
          1314 => x"9e",
          1315 => x"88",
          1316 => x"51",
          1317 => x"80",
          1318 => x"81",
          1319 => x"fa",
          1320 => x"0b",
          1321 => x"90",
          1322 => x"80",
          1323 => x"52",
          1324 => x"2e",
          1325 => x"52",
          1326 => x"b3",
          1327 => x"87",
          1328 => x"08",
          1329 => x"80",
          1330 => x"52",
          1331 => x"83",
          1332 => x"71",
          1333 => x"34",
          1334 => x"c0",
          1335 => x"70",
          1336 => x"06",
          1337 => x"70",
          1338 => x"38",
          1339 => x"81",
          1340 => x"80",
          1341 => x"9e",
          1342 => x"90",
          1343 => x"51",
          1344 => x"80",
          1345 => x"81",
          1346 => x"fa",
          1347 => x"0b",
          1348 => x"90",
          1349 => x"80",
          1350 => x"52",
          1351 => x"2e",
          1352 => x"52",
          1353 => x"b7",
          1354 => x"87",
          1355 => x"08",
          1356 => x"80",
          1357 => x"52",
          1358 => x"83",
          1359 => x"71",
          1360 => x"34",
          1361 => x"c0",
          1362 => x"70",
          1363 => x"06",
          1364 => x"70",
          1365 => x"38",
          1366 => x"81",
          1367 => x"80",
          1368 => x"9e",
          1369 => x"80",
          1370 => x"51",
          1371 => x"80",
          1372 => x"81",
          1373 => x"fa",
          1374 => x"0b",
          1375 => x"90",
          1376 => x"80",
          1377 => x"52",
          1378 => x"83",
          1379 => x"71",
          1380 => x"34",
          1381 => x"90",
          1382 => x"80",
          1383 => x"2a",
          1384 => x"70",
          1385 => x"34",
          1386 => x"c0",
          1387 => x"70",
          1388 => x"51",
          1389 => x"80",
          1390 => x"81",
          1391 => x"fa",
          1392 => x"c0",
          1393 => x"70",
          1394 => x"70",
          1395 => x"51",
          1396 => x"fa",
          1397 => x"0b",
          1398 => x"90",
          1399 => x"06",
          1400 => x"70",
          1401 => x"38",
          1402 => x"81",
          1403 => x"87",
          1404 => x"08",
          1405 => x"51",
          1406 => x"fa",
          1407 => x"3d",
          1408 => x"3d",
          1409 => x"ec",
          1410 => x"3f",
          1411 => x"33",
          1412 => x"2e",
          1413 => x"e3",
          1414 => x"8a",
          1415 => x"94",
          1416 => x"3f",
          1417 => x"33",
          1418 => x"2e",
          1419 => x"fa",
          1420 => x"fa",
          1421 => x"54",
          1422 => x"ac",
          1423 => x"3f",
          1424 => x"33",
          1425 => x"2e",
          1426 => x"fa",
          1427 => x"fa",
          1428 => x"54",
          1429 => x"c8",
          1430 => x"3f",
          1431 => x"33",
          1432 => x"2e",
          1433 => x"f9",
          1434 => x"f9",
          1435 => x"54",
          1436 => x"e4",
          1437 => x"3f",
          1438 => x"33",
          1439 => x"2e",
          1440 => x"f9",
          1441 => x"f9",
          1442 => x"54",
          1443 => x"80",
          1444 => x"3f",
          1445 => x"33",
          1446 => x"2e",
          1447 => x"f9",
          1448 => x"fa",
          1449 => x"54",
          1450 => x"9c",
          1451 => x"3f",
          1452 => x"33",
          1453 => x"2e",
          1454 => x"fa",
          1455 => x"81",
          1456 => x"8e",
          1457 => x"fa",
          1458 => x"73",
          1459 => x"38",
          1460 => x"33",
          1461 => x"d8",
          1462 => x"3f",
          1463 => x"33",
          1464 => x"2e",
          1465 => x"fa",
          1466 => x"81",
          1467 => x"8e",
          1468 => x"fa",
          1469 => x"73",
          1470 => x"38",
          1471 => x"51",
          1472 => x"81",
          1473 => x"54",
          1474 => x"88",
          1475 => x"ac",
          1476 => x"3f",
          1477 => x"33",
          1478 => x"2e",
          1479 => x"e5",
          1480 => x"82",
          1481 => x"b9",
          1482 => x"80",
          1483 => x"81",
          1484 => x"87",
          1485 => x"fa",
          1486 => x"73",
          1487 => x"38",
          1488 => x"51",
          1489 => x"81",
          1490 => x"87",
          1491 => x"fa",
          1492 => x"81",
          1493 => x"8d",
          1494 => x"fa",
          1495 => x"81",
          1496 => x"8d",
          1497 => x"fa",
          1498 => x"81",
          1499 => x"8d",
          1500 => x"e6",
          1501 => x"ae",
          1502 => x"a0",
          1503 => x"e6",
          1504 => x"86",
          1505 => x"a4",
          1506 => x"84",
          1507 => x"51",
          1508 => x"81",
          1509 => x"bd",
          1510 => x"76",
          1511 => x"54",
          1512 => x"08",
          1513 => x"90",
          1514 => x"3f",
          1515 => x"33",
          1516 => x"2e",
          1517 => x"fa",
          1518 => x"bd",
          1519 => x"75",
          1520 => x"3f",
          1521 => x"08",
          1522 => x"29",
          1523 => x"54",
          1524 => x"f0",
          1525 => x"e7",
          1526 => x"ae",
          1527 => x"b2",
          1528 => x"80",
          1529 => x"81",
          1530 => x"56",
          1531 => x"52",
          1532 => x"b8",
          1533 => x"f0",
          1534 => x"c0",
          1535 => x"31",
          1536 => x"fe",
          1537 => x"81",
          1538 => x"8b",
          1539 => x"f5",
          1540 => x"92",
          1541 => x"0d",
          1542 => x"0d",
          1543 => x"33",
          1544 => x"71",
          1545 => x"38",
          1546 => x"81",
          1547 => x"52",
          1548 => x"81",
          1549 => x"9d",
          1550 => x"9c",
          1551 => x"81",
          1552 => x"91",
          1553 => x"ac",
          1554 => x"81",
          1555 => x"85",
          1556 => x"b8",
          1557 => x"3f",
          1558 => x"04",
          1559 => x"0c",
          1560 => x"0d",
          1561 => x"84",
          1562 => x"52",
          1563 => x"70",
          1564 => x"81",
          1565 => x"72",
          1566 => x"0d",
          1567 => x"0d",
          1568 => x"84",
          1569 => x"fa",
          1570 => x"80",
          1571 => x"09",
          1572 => x"c4",
          1573 => x"81",
          1574 => x"73",
          1575 => x"3d",
          1576 => x"0b",
          1577 => x"84",
          1578 => x"fa",
          1579 => x"c0",
          1580 => x"04",
          1581 => x"81",
          1582 => x"89",
          1583 => x"b0",
          1584 => x"80",
          1585 => x"80",
          1586 => x"52",
          1587 => x"70",
          1588 => x"26",
          1589 => x"81",
          1590 => x"71",
          1591 => x"fe",
          1592 => x"3d",
          1593 => x"3d",
          1594 => x"84",
          1595 => x"12",
          1596 => x"94",
          1597 => x"16",
          1598 => x"54",
          1599 => x"70",
          1600 => x"38",
          1601 => x"14",
          1602 => x"81",
          1603 => x"76",
          1604 => x"0c",
          1605 => x"75",
          1606 => x"72",
          1607 => x"71",
          1608 => x"70",
          1609 => x"70",
          1610 => x"73",
          1611 => x"74",
          1612 => x"70",
          1613 => x"70",
          1614 => x"8c",
          1615 => x"0c",
          1616 => x"0c",
          1617 => x"0c",
          1618 => x"f0",
          1619 => x"0d",
          1620 => x"0d",
          1621 => x"08",
          1622 => x"56",
          1623 => x"08",
          1624 => x"81",
          1625 => x"84",
          1626 => x"13",
          1627 => x"73",
          1628 => x"06",
          1629 => x"13",
          1630 => x"13",
          1631 => x"13",
          1632 => x"15",
          1633 => x"9f",
          1634 => x"0c",
          1635 => x"08",
          1636 => x"81",
          1637 => x"94",
          1638 => x"81",
          1639 => x"90",
          1640 => x"94",
          1641 => x"73",
          1642 => x"09",
          1643 => x"38",
          1644 => x"70",
          1645 => x"70",
          1646 => x"81",
          1647 => x"84",
          1648 => x"84",
          1649 => x"14",
          1650 => x"08",
          1651 => x"0c",
          1652 => x"0c",
          1653 => x"88",
          1654 => x"88",
          1655 => x"8c",
          1656 => x"81",
          1657 => x"86",
          1658 => x"f9",
          1659 => x"70",
          1660 => x"80",
          1661 => x"38",
          1662 => x"06",
          1663 => x"08",
          1664 => x"08",
          1665 => x"38",
          1666 => x"77",
          1667 => x"38",
          1668 => x"56",
          1669 => x"ff",
          1670 => x"80",
          1671 => x"52",
          1672 => x"3f",
          1673 => x"08",
          1674 => x"08",
          1675 => x"fe",
          1676 => x"80",
          1677 => x"f0",
          1678 => x"30",
          1679 => x"80",
          1680 => x"53",
          1681 => x"54",
          1682 => x"72",
          1683 => x"81",
          1684 => x"38",
          1685 => x"52",
          1686 => x"c8",
          1687 => x"81",
          1688 => x"0c",
          1689 => x"f0",
          1690 => x"0c",
          1691 => x"08",
          1692 => x"82",
          1693 => x"75",
          1694 => x"38",
          1695 => x"53",
          1696 => x"13",
          1697 => x"0c",
          1698 => x"0c",
          1699 => x"0c",
          1700 => x"76",
          1701 => x"53",
          1702 => x"b5",
          1703 => x"81",
          1704 => x"51",
          1705 => x"81",
          1706 => x"54",
          1707 => x"f0",
          1708 => x"0d",
          1709 => x"0d",
          1710 => x"80",
          1711 => x"f0",
          1712 => x"8d",
          1713 => x"0d",
          1714 => x"0d",
          1715 => x"33",
          1716 => x"2e",
          1717 => x"85",
          1718 => x"ed",
          1719 => x"8c",
          1720 => x"80",
          1721 => x"72",
          1722 => x"ff",
          1723 => x"05",
          1724 => x"0c",
          1725 => x"ff",
          1726 => x"71",
          1727 => x"38",
          1728 => x"2d",
          1729 => x"04",
          1730 => x"02",
          1731 => x"81",
          1732 => x"76",
          1733 => x"0c",
          1734 => x"ad",
          1735 => x"ff",
          1736 => x"3d",
          1737 => x"3d",
          1738 => x"73",
          1739 => x"ff",
          1740 => x"71",
          1741 => x"38",
          1742 => x"06",
          1743 => x"54",
          1744 => x"e7",
          1745 => x"0d",
          1746 => x"0d",
          1747 => x"84",
          1748 => x"ff",
          1749 => x"54",
          1750 => x"81",
          1751 => x"53",
          1752 => x"8e",
          1753 => x"ff",
          1754 => x"14",
          1755 => x"3f",
          1756 => x"81",
          1757 => x"86",
          1758 => x"ec",
          1759 => x"68",
          1760 => x"70",
          1761 => x"33",
          1762 => x"2e",
          1763 => x"75",
          1764 => x"81",
          1765 => x"38",
          1766 => x"70",
          1767 => x"33",
          1768 => x"75",
          1769 => x"81",
          1770 => x"81",
          1771 => x"75",
          1772 => x"81",
          1773 => x"82",
          1774 => x"81",
          1775 => x"56",
          1776 => x"09",
          1777 => x"38",
          1778 => x"71",
          1779 => x"81",
          1780 => x"59",
          1781 => x"9d",
          1782 => x"53",
          1783 => x"95",
          1784 => x"29",
          1785 => x"76",
          1786 => x"79",
          1787 => x"5b",
          1788 => x"e5",
          1789 => x"ec",
          1790 => x"70",
          1791 => x"25",
          1792 => x"32",
          1793 => x"72",
          1794 => x"73",
          1795 => x"58",
          1796 => x"73",
          1797 => x"38",
          1798 => x"79",
          1799 => x"5b",
          1800 => x"75",
          1801 => x"de",
          1802 => x"80",
          1803 => x"89",
          1804 => x"70",
          1805 => x"55",
          1806 => x"cf",
          1807 => x"38",
          1808 => x"24",
          1809 => x"80",
          1810 => x"8e",
          1811 => x"c3",
          1812 => x"73",
          1813 => x"81",
          1814 => x"99",
          1815 => x"c4",
          1816 => x"38",
          1817 => x"73",
          1818 => x"81",
          1819 => x"80",
          1820 => x"38",
          1821 => x"2e",
          1822 => x"f9",
          1823 => x"d8",
          1824 => x"38",
          1825 => x"77",
          1826 => x"08",
          1827 => x"80",
          1828 => x"55",
          1829 => x"8d",
          1830 => x"70",
          1831 => x"51",
          1832 => x"f5",
          1833 => x"2a",
          1834 => x"74",
          1835 => x"53",
          1836 => x"8f",
          1837 => x"fc",
          1838 => x"81",
          1839 => x"80",
          1840 => x"73",
          1841 => x"3f",
          1842 => x"56",
          1843 => x"27",
          1844 => x"a0",
          1845 => x"3f",
          1846 => x"84",
          1847 => x"33",
          1848 => x"93",
          1849 => x"95",
          1850 => x"91",
          1851 => x"8d",
          1852 => x"89",
          1853 => x"fb",
          1854 => x"86",
          1855 => x"2a",
          1856 => x"51",
          1857 => x"2e",
          1858 => x"84",
          1859 => x"86",
          1860 => x"78",
          1861 => x"08",
          1862 => x"32",
          1863 => x"72",
          1864 => x"51",
          1865 => x"74",
          1866 => x"38",
          1867 => x"88",
          1868 => x"7a",
          1869 => x"55",
          1870 => x"3d",
          1871 => x"52",
          1872 => x"9b",
          1873 => x"f0",
          1874 => x"06",
          1875 => x"52",
          1876 => x"3f",
          1877 => x"08",
          1878 => x"27",
          1879 => x"14",
          1880 => x"f8",
          1881 => x"87",
          1882 => x"81",
          1883 => x"b0",
          1884 => x"7d",
          1885 => x"5f",
          1886 => x"75",
          1887 => x"07",
          1888 => x"54",
          1889 => x"26",
          1890 => x"ff",
          1891 => x"84",
          1892 => x"06",
          1893 => x"80",
          1894 => x"96",
          1895 => x"e0",
          1896 => x"73",
          1897 => x"57",
          1898 => x"06",
          1899 => x"54",
          1900 => x"a0",
          1901 => x"2a",
          1902 => x"54",
          1903 => x"38",
          1904 => x"76",
          1905 => x"38",
          1906 => x"fd",
          1907 => x"06",
          1908 => x"38",
          1909 => x"56",
          1910 => x"26",
          1911 => x"3d",
          1912 => x"05",
          1913 => x"ff",
          1914 => x"53",
          1915 => x"d9",
          1916 => x"38",
          1917 => x"56",
          1918 => x"27",
          1919 => x"a0",
          1920 => x"3f",
          1921 => x"3d",
          1922 => x"3d",
          1923 => x"70",
          1924 => x"52",
          1925 => x"73",
          1926 => x"3f",
          1927 => x"04",
          1928 => x"74",
          1929 => x"0c",
          1930 => x"05",
          1931 => x"fa",
          1932 => x"ff",
          1933 => x"80",
          1934 => x"0b",
          1935 => x"0c",
          1936 => x"04",
          1937 => x"81",
          1938 => x"76",
          1939 => x"0c",
          1940 => x"05",
          1941 => x"53",
          1942 => x"72",
          1943 => x"0c",
          1944 => x"04",
          1945 => x"77",
          1946 => x"88",
          1947 => x"54",
          1948 => x"54",
          1949 => x"80",
          1950 => x"ff",
          1951 => x"71",
          1952 => x"f0",
          1953 => x"06",
          1954 => x"2e",
          1955 => x"72",
          1956 => x"38",
          1957 => x"70",
          1958 => x"25",
          1959 => x"73",
          1960 => x"38",
          1961 => x"86",
          1962 => x"54",
          1963 => x"73",
          1964 => x"ff",
          1965 => x"72",
          1966 => x"74",
          1967 => x"72",
          1968 => x"54",
          1969 => x"81",
          1970 => x"39",
          1971 => x"80",
          1972 => x"51",
          1973 => x"81",
          1974 => x"fe",
          1975 => x"3d",
          1976 => x"3d",
          1977 => x"88",
          1978 => x"ff",
          1979 => x"53",
          1980 => x"fe",
          1981 => x"81",
          1982 => x"84",
          1983 => x"f8",
          1984 => x"7c",
          1985 => x"70",
          1986 => x"75",
          1987 => x"55",
          1988 => x"2e",
          1989 => x"87",
          1990 => x"76",
          1991 => x"73",
          1992 => x"81",
          1993 => x"81",
          1994 => x"77",
          1995 => x"70",
          1996 => x"58",
          1997 => x"09",
          1998 => x"c2",
          1999 => x"81",
          2000 => x"75",
          2001 => x"55",
          2002 => x"e2",
          2003 => x"90",
          2004 => x"f8",
          2005 => x"8f",
          2006 => x"81",
          2007 => x"75",
          2008 => x"55",
          2009 => x"81",
          2010 => x"27",
          2011 => x"d0",
          2012 => x"55",
          2013 => x"73",
          2014 => x"80",
          2015 => x"14",
          2016 => x"72",
          2017 => x"e0",
          2018 => x"80",
          2019 => x"39",
          2020 => x"55",
          2021 => x"80",
          2022 => x"e0",
          2023 => x"38",
          2024 => x"81",
          2025 => x"53",
          2026 => x"81",
          2027 => x"53",
          2028 => x"8e",
          2029 => x"70",
          2030 => x"55",
          2031 => x"27",
          2032 => x"77",
          2033 => x"74",
          2034 => x"76",
          2035 => x"77",
          2036 => x"70",
          2037 => x"55",
          2038 => x"77",
          2039 => x"38",
          2040 => x"74",
          2041 => x"55",
          2042 => x"f0",
          2043 => x"0d",
          2044 => x"0d",
          2045 => x"56",
          2046 => x"0c",
          2047 => x"70",
          2048 => x"73",
          2049 => x"81",
          2050 => x"81",
          2051 => x"ed",
          2052 => x"2e",
          2053 => x"8e",
          2054 => x"08",
          2055 => x"76",
          2056 => x"56",
          2057 => x"b0",
          2058 => x"06",
          2059 => x"75",
          2060 => x"76",
          2061 => x"70",
          2062 => x"73",
          2063 => x"8b",
          2064 => x"73",
          2065 => x"85",
          2066 => x"82",
          2067 => x"76",
          2068 => x"70",
          2069 => x"ac",
          2070 => x"a0",
          2071 => x"fa",
          2072 => x"53",
          2073 => x"57",
          2074 => x"98",
          2075 => x"39",
          2076 => x"80",
          2077 => x"26",
          2078 => x"86",
          2079 => x"80",
          2080 => x"57",
          2081 => x"74",
          2082 => x"38",
          2083 => x"27",
          2084 => x"14",
          2085 => x"06",
          2086 => x"14",
          2087 => x"06",
          2088 => x"74",
          2089 => x"f9",
          2090 => x"ff",
          2091 => x"89",
          2092 => x"38",
          2093 => x"c5",
          2094 => x"29",
          2095 => x"81",
          2096 => x"76",
          2097 => x"56",
          2098 => x"ba",
          2099 => x"2e",
          2100 => x"30",
          2101 => x"0c",
          2102 => x"81",
          2103 => x"8a",
          2104 => x"fd",
          2105 => x"98",
          2106 => x"2c",
          2107 => x"70",
          2108 => x"10",
          2109 => x"2b",
          2110 => x"54",
          2111 => x"0b",
          2112 => x"12",
          2113 => x"71",
          2114 => x"38",
          2115 => x"11",
          2116 => x"84",
          2117 => x"33",
          2118 => x"52",
          2119 => x"2e",
          2120 => x"83",
          2121 => x"72",
          2122 => x"0c",
          2123 => x"04",
          2124 => x"78",
          2125 => x"9f",
          2126 => x"33",
          2127 => x"71",
          2128 => x"38",
          2129 => x"81",
          2130 => x"f2",
          2131 => x"51",
          2132 => x"72",
          2133 => x"52",
          2134 => x"71",
          2135 => x"52",
          2136 => x"51",
          2137 => x"73",
          2138 => x"3d",
          2139 => x"3d",
          2140 => x"84",
          2141 => x"33",
          2142 => x"bb",
          2143 => x"fb",
          2144 => x"84",
          2145 => x"e4",
          2146 => x"51",
          2147 => x"58",
          2148 => x"2e",
          2149 => x"51",
          2150 => x"81",
          2151 => x"70",
          2152 => x"fa",
          2153 => x"19",
          2154 => x"56",
          2155 => x"3f",
          2156 => x"08",
          2157 => x"fb",
          2158 => x"84",
          2159 => x"e4",
          2160 => x"51",
          2161 => x"80",
          2162 => x"75",
          2163 => x"74",
          2164 => x"3f",
          2165 => x"33",
          2166 => x"74",
          2167 => x"34",
          2168 => x"06",
          2169 => x"27",
          2170 => x"0b",
          2171 => x"34",
          2172 => x"b6",
          2173 => x"b8",
          2174 => x"80",
          2175 => x"81",
          2176 => x"55",
          2177 => x"8c",
          2178 => x"54",
          2179 => x"52",
          2180 => x"c8",
          2181 => x"fb",
          2182 => x"8a",
          2183 => x"9e",
          2184 => x"b8",
          2185 => x"cb",
          2186 => x"3d",
          2187 => x"3d",
          2188 => x"80",
          2189 => x"b8",
          2190 => x"d2",
          2191 => x"fe",
          2192 => x"d1",
          2193 => x"b8",
          2194 => x"f8",
          2195 => x"70",
          2196 => x"fa",
          2197 => x"fe",
          2198 => x"2e",
          2199 => x"51",
          2200 => x"81",
          2201 => x"55",
          2202 => x"fe",
          2203 => x"9c",
          2204 => x"f0",
          2205 => x"70",
          2206 => x"80",
          2207 => x"53",
          2208 => x"17",
          2209 => x"52",
          2210 => x"3f",
          2211 => x"09",
          2212 => x"b1",
          2213 => x"0d",
          2214 => x"0d",
          2215 => x"ad",
          2216 => x"5a",
          2217 => x"58",
          2218 => x"fb",
          2219 => x"80",
          2220 => x"81",
          2221 => x"81",
          2222 => x"0b",
          2223 => x"08",
          2224 => x"f8",
          2225 => x"70",
          2226 => x"f9",
          2227 => x"fe",
          2228 => x"2e",
          2229 => x"51",
          2230 => x"81",
          2231 => x"81",
          2232 => x"80",
          2233 => x"f0",
          2234 => x"38",
          2235 => x"08",
          2236 => x"17",
          2237 => x"74",
          2238 => x"70",
          2239 => x"07",
          2240 => x"55",
          2241 => x"2e",
          2242 => x"ff",
          2243 => x"fb",
          2244 => x"11",
          2245 => x"80",
          2246 => x"81",
          2247 => x"80",
          2248 => x"81",
          2249 => x"ef",
          2250 => x"77",
          2251 => x"06",
          2252 => x"52",
          2253 => x"a7",
          2254 => x"d6",
          2255 => x"3d",
          2256 => x"fe",
          2257 => x"34",
          2258 => x"81",
          2259 => x"a9",
          2260 => x"f6",
          2261 => x"7e",
          2262 => x"72",
          2263 => x"5a",
          2264 => x"2e",
          2265 => x"a2",
          2266 => x"78",
          2267 => x"76",
          2268 => x"81",
          2269 => x"70",
          2270 => x"58",
          2271 => x"2e",
          2272 => x"86",
          2273 => x"26",
          2274 => x"54",
          2275 => x"81",
          2276 => x"70",
          2277 => x"d5",
          2278 => x"fe",
          2279 => x"79",
          2280 => x"51",
          2281 => x"81",
          2282 => x"80",
          2283 => x"15",
          2284 => x"81",
          2285 => x"74",
          2286 => x"38",
          2287 => x"ee",
          2288 => x"81",
          2289 => x"3d",
          2290 => x"f8",
          2291 => x"af",
          2292 => x"f0",
          2293 => x"99",
          2294 => x"78",
          2295 => x"fd",
          2296 => x"fe",
          2297 => x"ff",
          2298 => x"85",
          2299 => x"91",
          2300 => x"70",
          2301 => x"51",
          2302 => x"27",
          2303 => x"80",
          2304 => x"fe",
          2305 => x"3d",
          2306 => x"3d",
          2307 => x"08",
          2308 => x"81",
          2309 => x"5f",
          2310 => x"af",
          2311 => x"fb",
          2312 => x"81",
          2313 => x"81",
          2314 => x"fb",
          2315 => x"73",
          2316 => x"a8",
          2317 => x"3f",
          2318 => x"08",
          2319 => x"0c",
          2320 => x"08",
          2321 => x"fe",
          2322 => x"81",
          2323 => x"52",
          2324 => x"08",
          2325 => x"3f",
          2326 => x"08",
          2327 => x"38",
          2328 => x"51",
          2329 => x"80",
          2330 => x"fb",
          2331 => x"80",
          2332 => x"3d",
          2333 => x"80",
          2334 => x"81",
          2335 => x"56",
          2336 => x"08",
          2337 => x"81",
          2338 => x"38",
          2339 => x"08",
          2340 => x"3f",
          2341 => x"08",
          2342 => x"81",
          2343 => x"25",
          2344 => x"fe",
          2345 => x"05",
          2346 => x"55",
          2347 => x"80",
          2348 => x"ff",
          2349 => x"51",
          2350 => x"74",
          2351 => x"81",
          2352 => x"38",
          2353 => x"0b",
          2354 => x"34",
          2355 => x"dd",
          2356 => x"fe",
          2357 => x"2b",
          2358 => x"51",
          2359 => x"2e",
          2360 => x"81",
          2361 => x"ff",
          2362 => x"98",
          2363 => x"2c",
          2364 => x"33",
          2365 => x"70",
          2366 => x"98",
          2367 => x"84",
          2368 => x"c8",
          2369 => x"15",
          2370 => x"51",
          2371 => x"59",
          2372 => x"58",
          2373 => x"78",
          2374 => x"38",
          2375 => x"b4",
          2376 => x"80",
          2377 => x"ff",
          2378 => x"98",
          2379 => x"80",
          2380 => x"ce",
          2381 => x"74",
          2382 => x"f7",
          2383 => x"fe",
          2384 => x"ff",
          2385 => x"80",
          2386 => x"74",
          2387 => x"34",
          2388 => x"39",
          2389 => x"0a",
          2390 => x"0a",
          2391 => x"2c",
          2392 => x"06",
          2393 => x"73",
          2394 => x"38",
          2395 => x"52",
          2396 => x"ef",
          2397 => x"f0",
          2398 => x"06",
          2399 => x"38",
          2400 => x"56",
          2401 => x"80",
          2402 => x"1c",
          2403 => x"ff",
          2404 => x"98",
          2405 => x"2c",
          2406 => x"33",
          2407 => x"70",
          2408 => x"10",
          2409 => x"2b",
          2410 => x"11",
          2411 => x"51",
          2412 => x"51",
          2413 => x"2e",
          2414 => x"fe",
          2415 => x"e9",
          2416 => x"7d",
          2417 => x"81",
          2418 => x"80",
          2419 => x"90",
          2420 => x"75",
          2421 => x"34",
          2422 => x"90",
          2423 => x"3d",
          2424 => x"0c",
          2425 => x"8b",
          2426 => x"38",
          2427 => x"81",
          2428 => x"54",
          2429 => x"81",
          2430 => x"54",
          2431 => x"fd",
          2432 => x"ff",
          2433 => x"73",
          2434 => x"38",
          2435 => x"70",
          2436 => x"55",
          2437 => x"9e",
          2438 => x"54",
          2439 => x"15",
          2440 => x"80",
          2441 => x"ff",
          2442 => x"98",
          2443 => x"9c",
          2444 => x"55",
          2445 => x"ff",
          2446 => x"11",
          2447 => x"81",
          2448 => x"73",
          2449 => x"3d",
          2450 => x"81",
          2451 => x"54",
          2452 => x"89",
          2453 => x"54",
          2454 => x"98",
          2455 => x"9c",
          2456 => x"80",
          2457 => x"ff",
          2458 => x"98",
          2459 => x"98",
          2460 => x"56",
          2461 => x"25",
          2462 => x"1a",
          2463 => x"54",
          2464 => x"74",
          2465 => x"29",
          2466 => x"05",
          2467 => x"81",
          2468 => x"56",
          2469 => x"75",
          2470 => x"81",
          2471 => x"70",
          2472 => x"98",
          2473 => x"98",
          2474 => x"56",
          2475 => x"25",
          2476 => x"88",
          2477 => x"3f",
          2478 => x"0a",
          2479 => x"0a",
          2480 => x"2c",
          2481 => x"33",
          2482 => x"73",
          2483 => x"38",
          2484 => x"81",
          2485 => x"70",
          2486 => x"55",
          2487 => x"2e",
          2488 => x"81",
          2489 => x"ff",
          2490 => x"81",
          2491 => x"ff",
          2492 => x"81",
          2493 => x"88",
          2494 => x"3f",
          2495 => x"33",
          2496 => x"70",
          2497 => x"ff",
          2498 => x"51",
          2499 => x"74",
          2500 => x"74",
          2501 => x"14",
          2502 => x"73",
          2503 => x"a9",
          2504 => x"80",
          2505 => x"80",
          2506 => x"98",
          2507 => x"98",
          2508 => x"55",
          2509 => x"db",
          2510 => x"e7",
          2511 => x"ff",
          2512 => x"98",
          2513 => x"2c",
          2514 => x"33",
          2515 => x"57",
          2516 => x"fa",
          2517 => x"51",
          2518 => x"74",
          2519 => x"29",
          2520 => x"05",
          2521 => x"81",
          2522 => x"58",
          2523 => x"75",
          2524 => x"fa",
          2525 => x"ff",
          2526 => x"05",
          2527 => x"34",
          2528 => x"c5",
          2529 => x"98",
          2530 => x"f7",
          2531 => x"fe",
          2532 => x"ff",
          2533 => x"98",
          2534 => x"98",
          2535 => x"80",
          2536 => x"38",
          2537 => x"52",
          2538 => x"c2",
          2539 => x"39",
          2540 => x"84",
          2541 => x"ff",
          2542 => x"73",
          2543 => x"8c",
          2544 => x"e6",
          2545 => x"ff",
          2546 => x"05",
          2547 => x"ff",
          2548 => x"81",
          2549 => x"e3",
          2550 => x"9c",
          2551 => x"98",
          2552 => x"73",
          2553 => x"e4",
          2554 => x"54",
          2555 => x"98",
          2556 => x"2b",
          2557 => x"75",
          2558 => x"56",
          2559 => x"74",
          2560 => x"74",
          2561 => x"14",
          2562 => x"73",
          2563 => x"b9",
          2564 => x"80",
          2565 => x"80",
          2566 => x"98",
          2567 => x"98",
          2568 => x"55",
          2569 => x"db",
          2570 => x"e5",
          2571 => x"ff",
          2572 => x"98",
          2573 => x"2c",
          2574 => x"33",
          2575 => x"57",
          2576 => x"f9",
          2577 => x"51",
          2578 => x"74",
          2579 => x"29",
          2580 => x"05",
          2581 => x"81",
          2582 => x"58",
          2583 => x"75",
          2584 => x"f8",
          2585 => x"ff",
          2586 => x"81",
          2587 => x"ff",
          2588 => x"56",
          2589 => x"27",
          2590 => x"81",
          2591 => x"81",
          2592 => x"74",
          2593 => x"52",
          2594 => x"3f",
          2595 => x"33",
          2596 => x"06",
          2597 => x"33",
          2598 => x"75",
          2599 => x"38",
          2600 => x"7a",
          2601 => x"fb",
          2602 => x"74",
          2603 => x"38",
          2604 => x"9a",
          2605 => x"f0",
          2606 => x"98",
          2607 => x"f0",
          2608 => x"06",
          2609 => x"74",
          2610 => x"c7",
          2611 => x"5b",
          2612 => x"7a",
          2613 => x"fa",
          2614 => x"11",
          2615 => x"74",
          2616 => x"38",
          2617 => x"e6",
          2618 => x"f0",
          2619 => x"98",
          2620 => x"f0",
          2621 => x"06",
          2622 => x"74",
          2623 => x"c7",
          2624 => x"1b",
          2625 => x"39",
          2626 => x"74",
          2627 => x"bc",
          2628 => x"ca",
          2629 => x"e2",
          2630 => x"2e",
          2631 => x"93",
          2632 => x"e4",
          2633 => x"80",
          2634 => x"74",
          2635 => x"3f",
          2636 => x"7a",
          2637 => x"fa",
          2638 => x"11",
          2639 => x"74",
          2640 => x"38",
          2641 => x"86",
          2642 => x"f0",
          2643 => x"98",
          2644 => x"f0",
          2645 => x"06",
          2646 => x"74",
          2647 => x"c6",
          2648 => x"1b",
          2649 => x"ff",
          2650 => x"39",
          2651 => x"74",
          2652 => x"d8",
          2653 => x"c9",
          2654 => x"fe",
          2655 => x"ff",
          2656 => x"fe",
          2657 => x"ff",
          2658 => x"53",
          2659 => x"51",
          2660 => x"81",
          2661 => x"81",
          2662 => x"52",
          2663 => x"90",
          2664 => x"39",
          2665 => x"33",
          2666 => x"06",
          2667 => x"33",
          2668 => x"74",
          2669 => x"94",
          2670 => x"54",
          2671 => x"9c",
          2672 => x"70",
          2673 => x"e2",
          2674 => x"80",
          2675 => x"9c",
          2676 => x"80",
          2677 => x"38",
          2678 => x"ed",
          2679 => x"9c",
          2680 => x"54",
          2681 => x"9c",
          2682 => x"39",
          2683 => x"ff",
          2684 => x"0b",
          2685 => x"34",
          2686 => x"f0",
          2687 => x"0d",
          2688 => x"0d",
          2689 => x"33",
          2690 => x"70",
          2691 => x"38",
          2692 => x"11",
          2693 => x"81",
          2694 => x"83",
          2695 => x"fc",
          2696 => x"9b",
          2697 => x"84",
          2698 => x"33",
          2699 => x"51",
          2700 => x"80",
          2701 => x"84",
          2702 => x"92",
          2703 => x"51",
          2704 => x"80",
          2705 => x"81",
          2706 => x"72",
          2707 => x"92",
          2708 => x"81",
          2709 => x"0b",
          2710 => x"8c",
          2711 => x"71",
          2712 => x"06",
          2713 => x"80",
          2714 => x"87",
          2715 => x"08",
          2716 => x"38",
          2717 => x"80",
          2718 => x"71",
          2719 => x"c0",
          2720 => x"51",
          2721 => x"87",
          2722 => x"fb",
          2723 => x"81",
          2724 => x"33",
          2725 => x"fe",
          2726 => x"3d",
          2727 => x"3d",
          2728 => x"64",
          2729 => x"bf",
          2730 => x"40",
          2731 => x"74",
          2732 => x"cd",
          2733 => x"f0",
          2734 => x"7a",
          2735 => x"81",
          2736 => x"72",
          2737 => x"87",
          2738 => x"11",
          2739 => x"8c",
          2740 => x"92",
          2741 => x"5a",
          2742 => x"58",
          2743 => x"c0",
          2744 => x"76",
          2745 => x"76",
          2746 => x"70",
          2747 => x"81",
          2748 => x"54",
          2749 => x"8e",
          2750 => x"52",
          2751 => x"81",
          2752 => x"81",
          2753 => x"74",
          2754 => x"53",
          2755 => x"83",
          2756 => x"78",
          2757 => x"8f",
          2758 => x"2e",
          2759 => x"c0",
          2760 => x"52",
          2761 => x"87",
          2762 => x"08",
          2763 => x"2e",
          2764 => x"84",
          2765 => x"38",
          2766 => x"87",
          2767 => x"15",
          2768 => x"70",
          2769 => x"52",
          2770 => x"ff",
          2771 => x"39",
          2772 => x"81",
          2773 => x"ff",
          2774 => x"57",
          2775 => x"90",
          2776 => x"80",
          2777 => x"71",
          2778 => x"78",
          2779 => x"38",
          2780 => x"80",
          2781 => x"80",
          2782 => x"81",
          2783 => x"72",
          2784 => x"0c",
          2785 => x"04",
          2786 => x"60",
          2787 => x"8c",
          2788 => x"33",
          2789 => x"5b",
          2790 => x"74",
          2791 => x"e1",
          2792 => x"f0",
          2793 => x"79",
          2794 => x"78",
          2795 => x"06",
          2796 => x"77",
          2797 => x"87",
          2798 => x"11",
          2799 => x"8c",
          2800 => x"92",
          2801 => x"59",
          2802 => x"85",
          2803 => x"98",
          2804 => x"7d",
          2805 => x"0c",
          2806 => x"08",
          2807 => x"70",
          2808 => x"53",
          2809 => x"2e",
          2810 => x"70",
          2811 => x"33",
          2812 => x"18",
          2813 => x"2a",
          2814 => x"51",
          2815 => x"2e",
          2816 => x"c0",
          2817 => x"52",
          2818 => x"87",
          2819 => x"08",
          2820 => x"2e",
          2821 => x"84",
          2822 => x"38",
          2823 => x"87",
          2824 => x"15",
          2825 => x"70",
          2826 => x"52",
          2827 => x"ff",
          2828 => x"39",
          2829 => x"81",
          2830 => x"80",
          2831 => x"52",
          2832 => x"90",
          2833 => x"80",
          2834 => x"71",
          2835 => x"7a",
          2836 => x"38",
          2837 => x"80",
          2838 => x"80",
          2839 => x"81",
          2840 => x"72",
          2841 => x"0c",
          2842 => x"04",
          2843 => x"7a",
          2844 => x"a3",
          2845 => x"88",
          2846 => x"33",
          2847 => x"56",
          2848 => x"3f",
          2849 => x"08",
          2850 => x"83",
          2851 => x"fe",
          2852 => x"87",
          2853 => x"0c",
          2854 => x"76",
          2855 => x"38",
          2856 => x"93",
          2857 => x"2b",
          2858 => x"8c",
          2859 => x"71",
          2860 => x"38",
          2861 => x"71",
          2862 => x"c6",
          2863 => x"39",
          2864 => x"81",
          2865 => x"06",
          2866 => x"71",
          2867 => x"38",
          2868 => x"8c",
          2869 => x"e8",
          2870 => x"98",
          2871 => x"71",
          2872 => x"73",
          2873 => x"92",
          2874 => x"72",
          2875 => x"06",
          2876 => x"f7",
          2877 => x"80",
          2878 => x"88",
          2879 => x"0c",
          2880 => x"80",
          2881 => x"56",
          2882 => x"56",
          2883 => x"81",
          2884 => x"88",
          2885 => x"fe",
          2886 => x"81",
          2887 => x"33",
          2888 => x"07",
          2889 => x"0c",
          2890 => x"3d",
          2891 => x"3d",
          2892 => x"11",
          2893 => x"33",
          2894 => x"71",
          2895 => x"81",
          2896 => x"72",
          2897 => x"75",
          2898 => x"81",
          2899 => x"52",
          2900 => x"54",
          2901 => x"0d",
          2902 => x"0d",
          2903 => x"05",
          2904 => x"52",
          2905 => x"70",
          2906 => x"34",
          2907 => x"51",
          2908 => x"83",
          2909 => x"ff",
          2910 => x"75",
          2911 => x"72",
          2912 => x"54",
          2913 => x"2a",
          2914 => x"70",
          2915 => x"34",
          2916 => x"51",
          2917 => x"81",
          2918 => x"70",
          2919 => x"70",
          2920 => x"3d",
          2921 => x"3d",
          2922 => x"77",
          2923 => x"70",
          2924 => x"38",
          2925 => x"05",
          2926 => x"70",
          2927 => x"34",
          2928 => x"eb",
          2929 => x"0d",
          2930 => x"0d",
          2931 => x"54",
          2932 => x"72",
          2933 => x"54",
          2934 => x"51",
          2935 => x"84",
          2936 => x"fc",
          2937 => x"77",
          2938 => x"53",
          2939 => x"05",
          2940 => x"70",
          2941 => x"33",
          2942 => x"ff",
          2943 => x"52",
          2944 => x"2e",
          2945 => x"80",
          2946 => x"71",
          2947 => x"0c",
          2948 => x"04",
          2949 => x"74",
          2950 => x"89",
          2951 => x"2e",
          2952 => x"11",
          2953 => x"52",
          2954 => x"70",
          2955 => x"f0",
          2956 => x"0d",
          2957 => x"81",
          2958 => x"04",
          2959 => x"fe",
          2960 => x"f7",
          2961 => x"56",
          2962 => x"17",
          2963 => x"74",
          2964 => x"d6",
          2965 => x"b0",
          2966 => x"b4",
          2967 => x"81",
          2968 => x"59",
          2969 => x"81",
          2970 => x"7a",
          2971 => x"06",
          2972 => x"fe",
          2973 => x"17",
          2974 => x"08",
          2975 => x"08",
          2976 => x"08",
          2977 => x"74",
          2978 => x"38",
          2979 => x"55",
          2980 => x"09",
          2981 => x"38",
          2982 => x"18",
          2983 => x"81",
          2984 => x"f9",
          2985 => x"39",
          2986 => x"81",
          2987 => x"8b",
          2988 => x"fa",
          2989 => x"7a",
          2990 => x"57",
          2991 => x"08",
          2992 => x"75",
          2993 => x"3f",
          2994 => x"08",
          2995 => x"f0",
          2996 => x"81",
          2997 => x"b4",
          2998 => x"16",
          2999 => x"be",
          3000 => x"f0",
          3001 => x"85",
          3002 => x"81",
          3003 => x"17",
          3004 => x"fe",
          3005 => x"3d",
          3006 => x"3d",
          3007 => x"52",
          3008 => x"3f",
          3009 => x"08",
          3010 => x"f0",
          3011 => x"38",
          3012 => x"74",
          3013 => x"81",
          3014 => x"38",
          3015 => x"59",
          3016 => x"09",
          3017 => x"e3",
          3018 => x"53",
          3019 => x"08",
          3020 => x"70",
          3021 => x"91",
          3022 => x"d5",
          3023 => x"17",
          3024 => x"3f",
          3025 => x"a4",
          3026 => x"51",
          3027 => x"86",
          3028 => x"f2",
          3029 => x"17",
          3030 => x"3f",
          3031 => x"52",
          3032 => x"51",
          3033 => x"8c",
          3034 => x"84",
          3035 => x"fc",
          3036 => x"17",
          3037 => x"70",
          3038 => x"79",
          3039 => x"52",
          3040 => x"51",
          3041 => x"77",
          3042 => x"80",
          3043 => x"81",
          3044 => x"f9",
          3045 => x"fe",
          3046 => x"2e",
          3047 => x"58",
          3048 => x"f0",
          3049 => x"0d",
          3050 => x"0d",
          3051 => x"98",
          3052 => x"05",
          3053 => x"80",
          3054 => x"27",
          3055 => x"14",
          3056 => x"29",
          3057 => x"05",
          3058 => x"81",
          3059 => x"87",
          3060 => x"f9",
          3061 => x"7a",
          3062 => x"54",
          3063 => x"27",
          3064 => x"76",
          3065 => x"27",
          3066 => x"ff",
          3067 => x"58",
          3068 => x"80",
          3069 => x"82",
          3070 => x"72",
          3071 => x"38",
          3072 => x"72",
          3073 => x"8e",
          3074 => x"39",
          3075 => x"17",
          3076 => x"a4",
          3077 => x"53",
          3078 => x"fd",
          3079 => x"fe",
          3080 => x"9f",
          3081 => x"ff",
          3082 => x"11",
          3083 => x"70",
          3084 => x"18",
          3085 => x"76",
          3086 => x"53",
          3087 => x"81",
          3088 => x"80",
          3089 => x"83",
          3090 => x"b4",
          3091 => x"88",
          3092 => x"79",
          3093 => x"84",
          3094 => x"58",
          3095 => x"80",
          3096 => x"9f",
          3097 => x"80",
          3098 => x"88",
          3099 => x"08",
          3100 => x"51",
          3101 => x"81",
          3102 => x"80",
          3103 => x"10",
          3104 => x"74",
          3105 => x"51",
          3106 => x"81",
          3107 => x"83",
          3108 => x"58",
          3109 => x"87",
          3110 => x"08",
          3111 => x"51",
          3112 => x"81",
          3113 => x"9b",
          3114 => x"2b",
          3115 => x"74",
          3116 => x"51",
          3117 => x"81",
          3118 => x"f0",
          3119 => x"83",
          3120 => x"77",
          3121 => x"0c",
          3122 => x"04",
          3123 => x"7a",
          3124 => x"58",
          3125 => x"81",
          3126 => x"9e",
          3127 => x"17",
          3128 => x"96",
          3129 => x"53",
          3130 => x"81",
          3131 => x"79",
          3132 => x"72",
          3133 => x"38",
          3134 => x"72",
          3135 => x"b8",
          3136 => x"39",
          3137 => x"17",
          3138 => x"a4",
          3139 => x"53",
          3140 => x"fb",
          3141 => x"fe",
          3142 => x"81",
          3143 => x"81",
          3144 => x"83",
          3145 => x"b4",
          3146 => x"78",
          3147 => x"56",
          3148 => x"76",
          3149 => x"38",
          3150 => x"9f",
          3151 => x"33",
          3152 => x"07",
          3153 => x"74",
          3154 => x"83",
          3155 => x"89",
          3156 => x"08",
          3157 => x"51",
          3158 => x"81",
          3159 => x"59",
          3160 => x"08",
          3161 => x"74",
          3162 => x"16",
          3163 => x"84",
          3164 => x"76",
          3165 => x"88",
          3166 => x"81",
          3167 => x"8f",
          3168 => x"53",
          3169 => x"80",
          3170 => x"88",
          3171 => x"08",
          3172 => x"51",
          3173 => x"81",
          3174 => x"59",
          3175 => x"08",
          3176 => x"77",
          3177 => x"06",
          3178 => x"83",
          3179 => x"05",
          3180 => x"f7",
          3181 => x"39",
          3182 => x"a4",
          3183 => x"52",
          3184 => x"ef",
          3185 => x"f0",
          3186 => x"fe",
          3187 => x"38",
          3188 => x"06",
          3189 => x"83",
          3190 => x"18",
          3191 => x"54",
          3192 => x"f6",
          3193 => x"fe",
          3194 => x"0a",
          3195 => x"52",
          3196 => x"83",
          3197 => x"83",
          3198 => x"81",
          3199 => x"8a",
          3200 => x"f8",
          3201 => x"7c",
          3202 => x"59",
          3203 => x"81",
          3204 => x"38",
          3205 => x"08",
          3206 => x"73",
          3207 => x"38",
          3208 => x"52",
          3209 => x"a4",
          3210 => x"f0",
          3211 => x"fe",
          3212 => x"f2",
          3213 => x"82",
          3214 => x"39",
          3215 => x"e6",
          3216 => x"f0",
          3217 => x"de",
          3218 => x"78",
          3219 => x"3f",
          3220 => x"08",
          3221 => x"f0",
          3222 => x"80",
          3223 => x"fe",
          3224 => x"2e",
          3225 => x"fe",
          3226 => x"2e",
          3227 => x"53",
          3228 => x"51",
          3229 => x"81",
          3230 => x"c5",
          3231 => x"08",
          3232 => x"18",
          3233 => x"57",
          3234 => x"90",
          3235 => x"90",
          3236 => x"16",
          3237 => x"54",
          3238 => x"34",
          3239 => x"78",
          3240 => x"38",
          3241 => x"81",
          3242 => x"8a",
          3243 => x"f6",
          3244 => x"7e",
          3245 => x"5b",
          3246 => x"38",
          3247 => x"58",
          3248 => x"88",
          3249 => x"08",
          3250 => x"38",
          3251 => x"39",
          3252 => x"51",
          3253 => x"81",
          3254 => x"fe",
          3255 => x"82",
          3256 => x"fe",
          3257 => x"81",
          3258 => x"ff",
          3259 => x"38",
          3260 => x"81",
          3261 => x"26",
          3262 => x"79",
          3263 => x"08",
          3264 => x"73",
          3265 => x"b9",
          3266 => x"2e",
          3267 => x"80",
          3268 => x"1a",
          3269 => x"08",
          3270 => x"38",
          3271 => x"52",
          3272 => x"af",
          3273 => x"81",
          3274 => x"81",
          3275 => x"06",
          3276 => x"fe",
          3277 => x"81",
          3278 => x"09",
          3279 => x"72",
          3280 => x"70",
          3281 => x"fe",
          3282 => x"51",
          3283 => x"73",
          3284 => x"81",
          3285 => x"80",
          3286 => x"8c",
          3287 => x"81",
          3288 => x"38",
          3289 => x"08",
          3290 => x"73",
          3291 => x"75",
          3292 => x"77",
          3293 => x"56",
          3294 => x"76",
          3295 => x"82",
          3296 => x"26",
          3297 => x"75",
          3298 => x"f8",
          3299 => x"fe",
          3300 => x"2e",
          3301 => x"59",
          3302 => x"08",
          3303 => x"81",
          3304 => x"81",
          3305 => x"59",
          3306 => x"08",
          3307 => x"70",
          3308 => x"25",
          3309 => x"51",
          3310 => x"73",
          3311 => x"75",
          3312 => x"81",
          3313 => x"38",
          3314 => x"f5",
          3315 => x"75",
          3316 => x"f9",
          3317 => x"fe",
          3318 => x"fe",
          3319 => x"70",
          3320 => x"08",
          3321 => x"51",
          3322 => x"80",
          3323 => x"73",
          3324 => x"38",
          3325 => x"52",
          3326 => x"d0",
          3327 => x"f0",
          3328 => x"a5",
          3329 => x"18",
          3330 => x"08",
          3331 => x"18",
          3332 => x"74",
          3333 => x"38",
          3334 => x"18",
          3335 => x"33",
          3336 => x"73",
          3337 => x"97",
          3338 => x"74",
          3339 => x"38",
          3340 => x"55",
          3341 => x"fe",
          3342 => x"85",
          3343 => x"75",
          3344 => x"fe",
          3345 => x"3d",
          3346 => x"3d",
          3347 => x"52",
          3348 => x"3f",
          3349 => x"08",
          3350 => x"81",
          3351 => x"80",
          3352 => x"52",
          3353 => x"c1",
          3354 => x"f0",
          3355 => x"f0",
          3356 => x"0c",
          3357 => x"53",
          3358 => x"15",
          3359 => x"f2",
          3360 => x"56",
          3361 => x"16",
          3362 => x"22",
          3363 => x"27",
          3364 => x"54",
          3365 => x"76",
          3366 => x"33",
          3367 => x"3f",
          3368 => x"08",
          3369 => x"38",
          3370 => x"76",
          3371 => x"70",
          3372 => x"9f",
          3373 => x"56",
          3374 => x"fe",
          3375 => x"3d",
          3376 => x"3d",
          3377 => x"71",
          3378 => x"57",
          3379 => x"0a",
          3380 => x"38",
          3381 => x"53",
          3382 => x"38",
          3383 => x"0c",
          3384 => x"54",
          3385 => x"75",
          3386 => x"73",
          3387 => x"a8",
          3388 => x"73",
          3389 => x"85",
          3390 => x"0b",
          3391 => x"5a",
          3392 => x"27",
          3393 => x"a8",
          3394 => x"18",
          3395 => x"39",
          3396 => x"70",
          3397 => x"58",
          3398 => x"b2",
          3399 => x"76",
          3400 => x"3f",
          3401 => x"08",
          3402 => x"f0",
          3403 => x"bd",
          3404 => x"81",
          3405 => x"27",
          3406 => x"16",
          3407 => x"f0",
          3408 => x"38",
          3409 => x"39",
          3410 => x"55",
          3411 => x"52",
          3412 => x"d5",
          3413 => x"f0",
          3414 => x"0c",
          3415 => x"0c",
          3416 => x"53",
          3417 => x"80",
          3418 => x"85",
          3419 => x"94",
          3420 => x"2a",
          3421 => x"0c",
          3422 => x"06",
          3423 => x"9c",
          3424 => x"58",
          3425 => x"f0",
          3426 => x"0d",
          3427 => x"0d",
          3428 => x"90",
          3429 => x"05",
          3430 => x"f0",
          3431 => x"27",
          3432 => x"0b",
          3433 => x"98",
          3434 => x"84",
          3435 => x"2e",
          3436 => x"76",
          3437 => x"58",
          3438 => x"38",
          3439 => x"15",
          3440 => x"08",
          3441 => x"38",
          3442 => x"88",
          3443 => x"53",
          3444 => x"81",
          3445 => x"c0",
          3446 => x"22",
          3447 => x"89",
          3448 => x"72",
          3449 => x"74",
          3450 => x"f3",
          3451 => x"fe",
          3452 => x"82",
          3453 => x"81",
          3454 => x"27",
          3455 => x"81",
          3456 => x"f0",
          3457 => x"80",
          3458 => x"16",
          3459 => x"f0",
          3460 => x"ca",
          3461 => x"38",
          3462 => x"0c",
          3463 => x"dd",
          3464 => x"08",
          3465 => x"f9",
          3466 => x"fe",
          3467 => x"87",
          3468 => x"f0",
          3469 => x"80",
          3470 => x"55",
          3471 => x"08",
          3472 => x"38",
          3473 => x"fe",
          3474 => x"2e",
          3475 => x"fe",
          3476 => x"75",
          3477 => x"3f",
          3478 => x"08",
          3479 => x"94",
          3480 => x"52",
          3481 => x"c1",
          3482 => x"f0",
          3483 => x"0c",
          3484 => x"0c",
          3485 => x"05",
          3486 => x"80",
          3487 => x"fe",
          3488 => x"3d",
          3489 => x"3d",
          3490 => x"71",
          3491 => x"57",
          3492 => x"51",
          3493 => x"81",
          3494 => x"54",
          3495 => x"08",
          3496 => x"81",
          3497 => x"56",
          3498 => x"52",
          3499 => x"83",
          3500 => x"f0",
          3501 => x"fe",
          3502 => x"d2",
          3503 => x"f0",
          3504 => x"08",
          3505 => x"54",
          3506 => x"e5",
          3507 => x"06",
          3508 => x"58",
          3509 => x"08",
          3510 => x"38",
          3511 => x"75",
          3512 => x"80",
          3513 => x"81",
          3514 => x"7a",
          3515 => x"06",
          3516 => x"39",
          3517 => x"08",
          3518 => x"76",
          3519 => x"3f",
          3520 => x"08",
          3521 => x"f0",
          3522 => x"ff",
          3523 => x"84",
          3524 => x"06",
          3525 => x"54",
          3526 => x"f0",
          3527 => x"0d",
          3528 => x"0d",
          3529 => x"52",
          3530 => x"3f",
          3531 => x"08",
          3532 => x"06",
          3533 => x"51",
          3534 => x"83",
          3535 => x"06",
          3536 => x"14",
          3537 => x"3f",
          3538 => x"08",
          3539 => x"07",
          3540 => x"fe",
          3541 => x"3d",
          3542 => x"3d",
          3543 => x"70",
          3544 => x"06",
          3545 => x"53",
          3546 => x"ed",
          3547 => x"33",
          3548 => x"83",
          3549 => x"06",
          3550 => x"90",
          3551 => x"15",
          3552 => x"3f",
          3553 => x"04",
          3554 => x"7b",
          3555 => x"84",
          3556 => x"58",
          3557 => x"80",
          3558 => x"38",
          3559 => x"52",
          3560 => x"8f",
          3561 => x"f0",
          3562 => x"fe",
          3563 => x"f5",
          3564 => x"08",
          3565 => x"53",
          3566 => x"84",
          3567 => x"39",
          3568 => x"70",
          3569 => x"81",
          3570 => x"51",
          3571 => x"16",
          3572 => x"f0",
          3573 => x"81",
          3574 => x"38",
          3575 => x"ae",
          3576 => x"81",
          3577 => x"54",
          3578 => x"2e",
          3579 => x"8f",
          3580 => x"81",
          3581 => x"76",
          3582 => x"54",
          3583 => x"09",
          3584 => x"38",
          3585 => x"7a",
          3586 => x"80",
          3587 => x"fa",
          3588 => x"fe",
          3589 => x"81",
          3590 => x"89",
          3591 => x"08",
          3592 => x"86",
          3593 => x"98",
          3594 => x"81",
          3595 => x"8b",
          3596 => x"fb",
          3597 => x"70",
          3598 => x"81",
          3599 => x"fc",
          3600 => x"fe",
          3601 => x"81",
          3602 => x"b4",
          3603 => x"08",
          3604 => x"ec",
          3605 => x"fe",
          3606 => x"81",
          3607 => x"a0",
          3608 => x"81",
          3609 => x"52",
          3610 => x"51",
          3611 => x"8b",
          3612 => x"52",
          3613 => x"51",
          3614 => x"81",
          3615 => x"34",
          3616 => x"f0",
          3617 => x"0d",
          3618 => x"0d",
          3619 => x"98",
          3620 => x"70",
          3621 => x"ec",
          3622 => x"fe",
          3623 => x"38",
          3624 => x"53",
          3625 => x"81",
          3626 => x"34",
          3627 => x"04",
          3628 => x"78",
          3629 => x"80",
          3630 => x"34",
          3631 => x"80",
          3632 => x"38",
          3633 => x"18",
          3634 => x"9c",
          3635 => x"70",
          3636 => x"56",
          3637 => x"a0",
          3638 => x"71",
          3639 => x"81",
          3640 => x"81",
          3641 => x"89",
          3642 => x"06",
          3643 => x"73",
          3644 => x"55",
          3645 => x"55",
          3646 => x"81",
          3647 => x"81",
          3648 => x"74",
          3649 => x"75",
          3650 => x"52",
          3651 => x"13",
          3652 => x"08",
          3653 => x"33",
          3654 => x"9c",
          3655 => x"11",
          3656 => x"8a",
          3657 => x"f0",
          3658 => x"96",
          3659 => x"e7",
          3660 => x"f0",
          3661 => x"23",
          3662 => x"e7",
          3663 => x"fe",
          3664 => x"17",
          3665 => x"0d",
          3666 => x"0d",
          3667 => x"5e",
          3668 => x"70",
          3669 => x"55",
          3670 => x"83",
          3671 => x"73",
          3672 => x"91",
          3673 => x"2e",
          3674 => x"1d",
          3675 => x"0c",
          3676 => x"15",
          3677 => x"70",
          3678 => x"56",
          3679 => x"09",
          3680 => x"38",
          3681 => x"80",
          3682 => x"30",
          3683 => x"78",
          3684 => x"54",
          3685 => x"73",
          3686 => x"60",
          3687 => x"54",
          3688 => x"96",
          3689 => x"0b",
          3690 => x"80",
          3691 => x"f6",
          3692 => x"fe",
          3693 => x"85",
          3694 => x"3d",
          3695 => x"5c",
          3696 => x"53",
          3697 => x"51",
          3698 => x"80",
          3699 => x"88",
          3700 => x"5c",
          3701 => x"09",
          3702 => x"d4",
          3703 => x"70",
          3704 => x"71",
          3705 => x"30",
          3706 => x"73",
          3707 => x"51",
          3708 => x"57",
          3709 => x"38",
          3710 => x"75",
          3711 => x"17",
          3712 => x"75",
          3713 => x"30",
          3714 => x"51",
          3715 => x"80",
          3716 => x"38",
          3717 => x"87",
          3718 => x"26",
          3719 => x"77",
          3720 => x"a4",
          3721 => x"27",
          3722 => x"a0",
          3723 => x"39",
          3724 => x"33",
          3725 => x"57",
          3726 => x"27",
          3727 => x"75",
          3728 => x"30",
          3729 => x"32",
          3730 => x"80",
          3731 => x"25",
          3732 => x"56",
          3733 => x"80",
          3734 => x"84",
          3735 => x"58",
          3736 => x"70",
          3737 => x"55",
          3738 => x"09",
          3739 => x"38",
          3740 => x"80",
          3741 => x"30",
          3742 => x"77",
          3743 => x"54",
          3744 => x"81",
          3745 => x"ae",
          3746 => x"06",
          3747 => x"54",
          3748 => x"74",
          3749 => x"80",
          3750 => x"7b",
          3751 => x"30",
          3752 => x"70",
          3753 => x"25",
          3754 => x"07",
          3755 => x"51",
          3756 => x"a7",
          3757 => x"8b",
          3758 => x"39",
          3759 => x"54",
          3760 => x"8c",
          3761 => x"ff",
          3762 => x"dc",
          3763 => x"54",
          3764 => x"e1",
          3765 => x"f0",
          3766 => x"b2",
          3767 => x"70",
          3768 => x"71",
          3769 => x"54",
          3770 => x"81",
          3771 => x"80",
          3772 => x"38",
          3773 => x"76",
          3774 => x"df",
          3775 => x"54",
          3776 => x"81",
          3777 => x"55",
          3778 => x"34",
          3779 => x"52",
          3780 => x"51",
          3781 => x"81",
          3782 => x"bf",
          3783 => x"16",
          3784 => x"26",
          3785 => x"16",
          3786 => x"06",
          3787 => x"17",
          3788 => x"34",
          3789 => x"fd",
          3790 => x"19",
          3791 => x"80",
          3792 => x"79",
          3793 => x"81",
          3794 => x"81",
          3795 => x"85",
          3796 => x"54",
          3797 => x"8f",
          3798 => x"86",
          3799 => x"39",
          3800 => x"f3",
          3801 => x"73",
          3802 => x"80",
          3803 => x"52",
          3804 => x"ce",
          3805 => x"f0",
          3806 => x"fe",
          3807 => x"d7",
          3808 => x"08",
          3809 => x"e6",
          3810 => x"fe",
          3811 => x"81",
          3812 => x"80",
          3813 => x"1b",
          3814 => x"55",
          3815 => x"2e",
          3816 => x"8b",
          3817 => x"06",
          3818 => x"1c",
          3819 => x"33",
          3820 => x"70",
          3821 => x"55",
          3822 => x"38",
          3823 => x"52",
          3824 => x"9f",
          3825 => x"f0",
          3826 => x"8b",
          3827 => x"7a",
          3828 => x"3f",
          3829 => x"75",
          3830 => x"57",
          3831 => x"2e",
          3832 => x"84",
          3833 => x"06",
          3834 => x"75",
          3835 => x"81",
          3836 => x"2a",
          3837 => x"73",
          3838 => x"38",
          3839 => x"54",
          3840 => x"fb",
          3841 => x"80",
          3842 => x"34",
          3843 => x"c1",
          3844 => x"06",
          3845 => x"38",
          3846 => x"39",
          3847 => x"70",
          3848 => x"54",
          3849 => x"86",
          3850 => x"84",
          3851 => x"06",
          3852 => x"73",
          3853 => x"38",
          3854 => x"83",
          3855 => x"b4",
          3856 => x"51",
          3857 => x"81",
          3858 => x"88",
          3859 => x"ea",
          3860 => x"fe",
          3861 => x"3d",
          3862 => x"3d",
          3863 => x"ff",
          3864 => x"71",
          3865 => x"5c",
          3866 => x"80",
          3867 => x"38",
          3868 => x"05",
          3869 => x"a0",
          3870 => x"71",
          3871 => x"38",
          3872 => x"71",
          3873 => x"81",
          3874 => x"38",
          3875 => x"11",
          3876 => x"06",
          3877 => x"70",
          3878 => x"38",
          3879 => x"81",
          3880 => x"05",
          3881 => x"76",
          3882 => x"38",
          3883 => x"eb",
          3884 => x"77",
          3885 => x"57",
          3886 => x"05",
          3887 => x"70",
          3888 => x"33",
          3889 => x"53",
          3890 => x"99",
          3891 => x"e0",
          3892 => x"ff",
          3893 => x"ff",
          3894 => x"70",
          3895 => x"38",
          3896 => x"81",
          3897 => x"51",
          3898 => x"9f",
          3899 => x"72",
          3900 => x"81",
          3901 => x"70",
          3902 => x"72",
          3903 => x"32",
          3904 => x"72",
          3905 => x"73",
          3906 => x"53",
          3907 => x"70",
          3908 => x"38",
          3909 => x"19",
          3910 => x"75",
          3911 => x"38",
          3912 => x"83",
          3913 => x"74",
          3914 => x"59",
          3915 => x"39",
          3916 => x"33",
          3917 => x"fe",
          3918 => x"3d",
          3919 => x"3d",
          3920 => x"80",
          3921 => x"34",
          3922 => x"17",
          3923 => x"75",
          3924 => x"3f",
          3925 => x"fe",
          3926 => x"80",
          3927 => x"16",
          3928 => x"3f",
          3929 => x"08",
          3930 => x"06",
          3931 => x"73",
          3932 => x"2e",
          3933 => x"80",
          3934 => x"0b",
          3935 => x"56",
          3936 => x"e9",
          3937 => x"06",
          3938 => x"57",
          3939 => x"32",
          3940 => x"80",
          3941 => x"51",
          3942 => x"8a",
          3943 => x"e8",
          3944 => x"06",
          3945 => x"53",
          3946 => x"52",
          3947 => x"51",
          3948 => x"81",
          3949 => x"55",
          3950 => x"08",
          3951 => x"38",
          3952 => x"eb",
          3953 => x"86",
          3954 => x"97",
          3955 => x"f0",
          3956 => x"fe",
          3957 => x"2e",
          3958 => x"55",
          3959 => x"f0",
          3960 => x"0d",
          3961 => x"0d",
          3962 => x"05",
          3963 => x"33",
          3964 => x"75",
          3965 => x"fc",
          3966 => x"fe",
          3967 => x"8b",
          3968 => x"81",
          3969 => x"24",
          3970 => x"81",
          3971 => x"84",
          3972 => x"a0",
          3973 => x"55",
          3974 => x"73",
          3975 => x"e6",
          3976 => x"0c",
          3977 => x"06",
          3978 => x"57",
          3979 => x"ae",
          3980 => x"33",
          3981 => x"3f",
          3982 => x"08",
          3983 => x"70",
          3984 => x"55",
          3985 => x"76",
          3986 => x"b8",
          3987 => x"2a",
          3988 => x"51",
          3989 => x"72",
          3990 => x"86",
          3991 => x"74",
          3992 => x"15",
          3993 => x"81",
          3994 => x"d7",
          3995 => x"fe",
          3996 => x"ff",
          3997 => x"06",
          3998 => x"56",
          3999 => x"38",
          4000 => x"8f",
          4001 => x"2a",
          4002 => x"51",
          4003 => x"72",
          4004 => x"80",
          4005 => x"52",
          4006 => x"3f",
          4007 => x"08",
          4008 => x"57",
          4009 => x"09",
          4010 => x"e2",
          4011 => x"74",
          4012 => x"56",
          4013 => x"33",
          4014 => x"72",
          4015 => x"38",
          4016 => x"51",
          4017 => x"81",
          4018 => x"57",
          4019 => x"84",
          4020 => x"ff",
          4021 => x"56",
          4022 => x"25",
          4023 => x"0b",
          4024 => x"56",
          4025 => x"05",
          4026 => x"83",
          4027 => x"2e",
          4028 => x"52",
          4029 => x"c6",
          4030 => x"f0",
          4031 => x"06",
          4032 => x"27",
          4033 => x"16",
          4034 => x"27",
          4035 => x"56",
          4036 => x"84",
          4037 => x"56",
          4038 => x"84",
          4039 => x"14",
          4040 => x"3f",
          4041 => x"08",
          4042 => x"06",
          4043 => x"80",
          4044 => x"06",
          4045 => x"80",
          4046 => x"db",
          4047 => x"fe",
          4048 => x"ff",
          4049 => x"77",
          4050 => x"d8",
          4051 => x"de",
          4052 => x"f0",
          4053 => x"9c",
          4054 => x"c4",
          4055 => x"15",
          4056 => x"14",
          4057 => x"70",
          4058 => x"51",
          4059 => x"56",
          4060 => x"84",
          4061 => x"81",
          4062 => x"71",
          4063 => x"16",
          4064 => x"53",
          4065 => x"23",
          4066 => x"8b",
          4067 => x"73",
          4068 => x"80",
          4069 => x"8d",
          4070 => x"39",
          4071 => x"51",
          4072 => x"81",
          4073 => x"53",
          4074 => x"08",
          4075 => x"72",
          4076 => x"8d",
          4077 => x"ce",
          4078 => x"14",
          4079 => x"3f",
          4080 => x"08",
          4081 => x"06",
          4082 => x"38",
          4083 => x"51",
          4084 => x"81",
          4085 => x"55",
          4086 => x"51",
          4087 => x"81",
          4088 => x"83",
          4089 => x"53",
          4090 => x"80",
          4091 => x"38",
          4092 => x"78",
          4093 => x"2a",
          4094 => x"78",
          4095 => x"86",
          4096 => x"22",
          4097 => x"31",
          4098 => x"a0",
          4099 => x"f0",
          4100 => x"fe",
          4101 => x"2e",
          4102 => x"81",
          4103 => x"80",
          4104 => x"f5",
          4105 => x"83",
          4106 => x"ff",
          4107 => x"38",
          4108 => x"9f",
          4109 => x"38",
          4110 => x"39",
          4111 => x"80",
          4112 => x"38",
          4113 => x"98",
          4114 => x"a0",
          4115 => x"1c",
          4116 => x"0c",
          4117 => x"17",
          4118 => x"76",
          4119 => x"81",
          4120 => x"80",
          4121 => x"d9",
          4122 => x"fe",
          4123 => x"ff",
          4124 => x"8d",
          4125 => x"8e",
          4126 => x"8a",
          4127 => x"14",
          4128 => x"3f",
          4129 => x"08",
          4130 => x"74",
          4131 => x"a2",
          4132 => x"79",
          4133 => x"ee",
          4134 => x"a8",
          4135 => x"15",
          4136 => x"2e",
          4137 => x"10",
          4138 => x"2a",
          4139 => x"05",
          4140 => x"ff",
          4141 => x"53",
          4142 => x"9c",
          4143 => x"81",
          4144 => x"0b",
          4145 => x"ff",
          4146 => x"0c",
          4147 => x"84",
          4148 => x"83",
          4149 => x"06",
          4150 => x"80",
          4151 => x"d8",
          4152 => x"fe",
          4153 => x"ff",
          4154 => x"72",
          4155 => x"81",
          4156 => x"38",
          4157 => x"73",
          4158 => x"3f",
          4159 => x"08",
          4160 => x"81",
          4161 => x"84",
          4162 => x"b2",
          4163 => x"87",
          4164 => x"f0",
          4165 => x"ff",
          4166 => x"82",
          4167 => x"09",
          4168 => x"c8",
          4169 => x"51",
          4170 => x"81",
          4171 => x"84",
          4172 => x"d2",
          4173 => x"06",
          4174 => x"98",
          4175 => x"ee",
          4176 => x"f0",
          4177 => x"85",
          4178 => x"09",
          4179 => x"38",
          4180 => x"51",
          4181 => x"81",
          4182 => x"90",
          4183 => x"a0",
          4184 => x"ca",
          4185 => x"f0",
          4186 => x"0c",
          4187 => x"81",
          4188 => x"81",
          4189 => x"81",
          4190 => x"72",
          4191 => x"80",
          4192 => x"0c",
          4193 => x"81",
          4194 => x"90",
          4195 => x"fb",
          4196 => x"54",
          4197 => x"80",
          4198 => x"73",
          4199 => x"80",
          4200 => x"72",
          4201 => x"80",
          4202 => x"86",
          4203 => x"15",
          4204 => x"71",
          4205 => x"81",
          4206 => x"81",
          4207 => x"d0",
          4208 => x"fe",
          4209 => x"06",
          4210 => x"38",
          4211 => x"54",
          4212 => x"80",
          4213 => x"71",
          4214 => x"81",
          4215 => x"87",
          4216 => x"fa",
          4217 => x"ab",
          4218 => x"58",
          4219 => x"05",
          4220 => x"e6",
          4221 => x"80",
          4222 => x"f0",
          4223 => x"38",
          4224 => x"08",
          4225 => x"ff",
          4226 => x"08",
          4227 => x"80",
          4228 => x"80",
          4229 => x"54",
          4230 => x"84",
          4231 => x"34",
          4232 => x"75",
          4233 => x"2e",
          4234 => x"53",
          4235 => x"53",
          4236 => x"f7",
          4237 => x"fe",
          4238 => x"73",
          4239 => x"0c",
          4240 => x"04",
          4241 => x"67",
          4242 => x"80",
          4243 => x"59",
          4244 => x"78",
          4245 => x"c8",
          4246 => x"06",
          4247 => x"3d",
          4248 => x"99",
          4249 => x"52",
          4250 => x"3f",
          4251 => x"08",
          4252 => x"f0",
          4253 => x"38",
          4254 => x"52",
          4255 => x"52",
          4256 => x"3f",
          4257 => x"08",
          4258 => x"f0",
          4259 => x"02",
          4260 => x"33",
          4261 => x"55",
          4262 => x"25",
          4263 => x"55",
          4264 => x"54",
          4265 => x"81",
          4266 => x"80",
          4267 => x"74",
          4268 => x"81",
          4269 => x"75",
          4270 => x"3f",
          4271 => x"08",
          4272 => x"02",
          4273 => x"91",
          4274 => x"81",
          4275 => x"82",
          4276 => x"06",
          4277 => x"80",
          4278 => x"88",
          4279 => x"39",
          4280 => x"58",
          4281 => x"38",
          4282 => x"70",
          4283 => x"54",
          4284 => x"81",
          4285 => x"52",
          4286 => x"a5",
          4287 => x"f0",
          4288 => x"88",
          4289 => x"62",
          4290 => x"d4",
          4291 => x"54",
          4292 => x"15",
          4293 => x"62",
          4294 => x"e8",
          4295 => x"52",
          4296 => x"51",
          4297 => x"7a",
          4298 => x"83",
          4299 => x"80",
          4300 => x"38",
          4301 => x"08",
          4302 => x"53",
          4303 => x"3d",
          4304 => x"dd",
          4305 => x"fe",
          4306 => x"81",
          4307 => x"82",
          4308 => x"39",
          4309 => x"38",
          4310 => x"33",
          4311 => x"70",
          4312 => x"55",
          4313 => x"2e",
          4314 => x"55",
          4315 => x"77",
          4316 => x"81",
          4317 => x"73",
          4318 => x"38",
          4319 => x"54",
          4320 => x"a0",
          4321 => x"82",
          4322 => x"52",
          4323 => x"a3",
          4324 => x"f0",
          4325 => x"18",
          4326 => x"55",
          4327 => x"f0",
          4328 => x"38",
          4329 => x"70",
          4330 => x"54",
          4331 => x"86",
          4332 => x"c0",
          4333 => x"b0",
          4334 => x"1b",
          4335 => x"1b",
          4336 => x"70",
          4337 => x"d9",
          4338 => x"f0",
          4339 => x"f0",
          4340 => x"0c",
          4341 => x"52",
          4342 => x"3f",
          4343 => x"08",
          4344 => x"08",
          4345 => x"77",
          4346 => x"86",
          4347 => x"1a",
          4348 => x"1a",
          4349 => x"91",
          4350 => x"0b",
          4351 => x"80",
          4352 => x"0c",
          4353 => x"70",
          4354 => x"54",
          4355 => x"81",
          4356 => x"fe",
          4357 => x"2e",
          4358 => x"81",
          4359 => x"94",
          4360 => x"17",
          4361 => x"2b",
          4362 => x"57",
          4363 => x"52",
          4364 => x"9f",
          4365 => x"f0",
          4366 => x"fe",
          4367 => x"26",
          4368 => x"55",
          4369 => x"08",
          4370 => x"81",
          4371 => x"79",
          4372 => x"31",
          4373 => x"70",
          4374 => x"25",
          4375 => x"76",
          4376 => x"81",
          4377 => x"55",
          4378 => x"38",
          4379 => x"0c",
          4380 => x"75",
          4381 => x"54",
          4382 => x"a2",
          4383 => x"7a",
          4384 => x"3f",
          4385 => x"08",
          4386 => x"55",
          4387 => x"89",
          4388 => x"f0",
          4389 => x"1a",
          4390 => x"80",
          4391 => x"54",
          4392 => x"f0",
          4393 => x"0d",
          4394 => x"0d",
          4395 => x"64",
          4396 => x"59",
          4397 => x"90",
          4398 => x"52",
          4399 => x"cf",
          4400 => x"f0",
          4401 => x"fe",
          4402 => x"38",
          4403 => x"55",
          4404 => x"86",
          4405 => x"82",
          4406 => x"19",
          4407 => x"55",
          4408 => x"80",
          4409 => x"38",
          4410 => x"0b",
          4411 => x"82",
          4412 => x"39",
          4413 => x"1a",
          4414 => x"82",
          4415 => x"19",
          4416 => x"08",
          4417 => x"7c",
          4418 => x"74",
          4419 => x"2e",
          4420 => x"94",
          4421 => x"83",
          4422 => x"56",
          4423 => x"38",
          4424 => x"22",
          4425 => x"89",
          4426 => x"55",
          4427 => x"75",
          4428 => x"19",
          4429 => x"39",
          4430 => x"52",
          4431 => x"93",
          4432 => x"f0",
          4433 => x"75",
          4434 => x"38",
          4435 => x"ff",
          4436 => x"98",
          4437 => x"19",
          4438 => x"51",
          4439 => x"81",
          4440 => x"80",
          4441 => x"38",
          4442 => x"08",
          4443 => x"2a",
          4444 => x"80",
          4445 => x"38",
          4446 => x"8a",
          4447 => x"5c",
          4448 => x"27",
          4449 => x"7a",
          4450 => x"54",
          4451 => x"52",
          4452 => x"51",
          4453 => x"81",
          4454 => x"fe",
          4455 => x"83",
          4456 => x"56",
          4457 => x"9f",
          4458 => x"08",
          4459 => x"74",
          4460 => x"38",
          4461 => x"b4",
          4462 => x"16",
          4463 => x"89",
          4464 => x"51",
          4465 => x"77",
          4466 => x"b9",
          4467 => x"1a",
          4468 => x"08",
          4469 => x"84",
          4470 => x"57",
          4471 => x"27",
          4472 => x"56",
          4473 => x"52",
          4474 => x"c7",
          4475 => x"f0",
          4476 => x"38",
          4477 => x"19",
          4478 => x"06",
          4479 => x"52",
          4480 => x"a2",
          4481 => x"31",
          4482 => x"7f",
          4483 => x"94",
          4484 => x"94",
          4485 => x"5c",
          4486 => x"80",
          4487 => x"fe",
          4488 => x"3d",
          4489 => x"3d",
          4490 => x"65",
          4491 => x"5d",
          4492 => x"0c",
          4493 => x"05",
          4494 => x"f6",
          4495 => x"fe",
          4496 => x"81",
          4497 => x"8a",
          4498 => x"33",
          4499 => x"2e",
          4500 => x"56",
          4501 => x"90",
          4502 => x"81",
          4503 => x"06",
          4504 => x"87",
          4505 => x"2e",
          4506 => x"95",
          4507 => x"91",
          4508 => x"56",
          4509 => x"81",
          4510 => x"34",
          4511 => x"8e",
          4512 => x"08",
          4513 => x"56",
          4514 => x"84",
          4515 => x"5c",
          4516 => x"82",
          4517 => x"18",
          4518 => x"ff",
          4519 => x"74",
          4520 => x"7e",
          4521 => x"ff",
          4522 => x"2a",
          4523 => x"7a",
          4524 => x"8c",
          4525 => x"08",
          4526 => x"38",
          4527 => x"39",
          4528 => x"52",
          4529 => x"e7",
          4530 => x"f0",
          4531 => x"fe",
          4532 => x"2e",
          4533 => x"74",
          4534 => x"91",
          4535 => x"2e",
          4536 => x"74",
          4537 => x"88",
          4538 => x"38",
          4539 => x"0c",
          4540 => x"15",
          4541 => x"08",
          4542 => x"06",
          4543 => x"51",
          4544 => x"81",
          4545 => x"fe",
          4546 => x"18",
          4547 => x"51",
          4548 => x"81",
          4549 => x"80",
          4550 => x"38",
          4551 => x"08",
          4552 => x"2a",
          4553 => x"80",
          4554 => x"38",
          4555 => x"8a",
          4556 => x"5b",
          4557 => x"27",
          4558 => x"7b",
          4559 => x"54",
          4560 => x"52",
          4561 => x"51",
          4562 => x"81",
          4563 => x"fe",
          4564 => x"b0",
          4565 => x"31",
          4566 => x"79",
          4567 => x"84",
          4568 => x"16",
          4569 => x"89",
          4570 => x"52",
          4571 => x"cc",
          4572 => x"55",
          4573 => x"16",
          4574 => x"2b",
          4575 => x"39",
          4576 => x"94",
          4577 => x"93",
          4578 => x"cd",
          4579 => x"fe",
          4580 => x"e3",
          4581 => x"b0",
          4582 => x"76",
          4583 => x"94",
          4584 => x"ff",
          4585 => x"71",
          4586 => x"7b",
          4587 => x"38",
          4588 => x"18",
          4589 => x"51",
          4590 => x"81",
          4591 => x"fd",
          4592 => x"53",
          4593 => x"18",
          4594 => x"06",
          4595 => x"51",
          4596 => x"7e",
          4597 => x"83",
          4598 => x"76",
          4599 => x"17",
          4600 => x"1e",
          4601 => x"18",
          4602 => x"0c",
          4603 => x"58",
          4604 => x"74",
          4605 => x"38",
          4606 => x"8c",
          4607 => x"90",
          4608 => x"33",
          4609 => x"55",
          4610 => x"34",
          4611 => x"81",
          4612 => x"90",
          4613 => x"f8",
          4614 => x"8b",
          4615 => x"53",
          4616 => x"f2",
          4617 => x"fe",
          4618 => x"81",
          4619 => x"80",
          4620 => x"16",
          4621 => x"2a",
          4622 => x"51",
          4623 => x"80",
          4624 => x"38",
          4625 => x"52",
          4626 => x"e7",
          4627 => x"f0",
          4628 => x"fe",
          4629 => x"d4",
          4630 => x"08",
          4631 => x"a0",
          4632 => x"73",
          4633 => x"88",
          4634 => x"74",
          4635 => x"51",
          4636 => x"8c",
          4637 => x"9c",
          4638 => x"fb",
          4639 => x"b2",
          4640 => x"15",
          4641 => x"3f",
          4642 => x"15",
          4643 => x"3f",
          4644 => x"0b",
          4645 => x"78",
          4646 => x"3f",
          4647 => x"08",
          4648 => x"81",
          4649 => x"57",
          4650 => x"34",
          4651 => x"f0",
          4652 => x"0d",
          4653 => x"0d",
          4654 => x"54",
          4655 => x"81",
          4656 => x"53",
          4657 => x"08",
          4658 => x"3d",
          4659 => x"73",
          4660 => x"3f",
          4661 => x"08",
          4662 => x"f0",
          4663 => x"81",
          4664 => x"74",
          4665 => x"fe",
          4666 => x"3d",
          4667 => x"3d",
          4668 => x"51",
          4669 => x"8b",
          4670 => x"81",
          4671 => x"24",
          4672 => x"fe",
          4673 => x"ff",
          4674 => x"52",
          4675 => x"f0",
          4676 => x"0d",
          4677 => x"0d",
          4678 => x"3d",
          4679 => x"94",
          4680 => x"c1",
          4681 => x"f0",
          4682 => x"fe",
          4683 => x"e0",
          4684 => x"63",
          4685 => x"d4",
          4686 => x"8d",
          4687 => x"f0",
          4688 => x"fe",
          4689 => x"38",
          4690 => x"05",
          4691 => x"2b",
          4692 => x"80",
          4693 => x"76",
          4694 => x"0c",
          4695 => x"02",
          4696 => x"70",
          4697 => x"81",
          4698 => x"56",
          4699 => x"9e",
          4700 => x"53",
          4701 => x"db",
          4702 => x"fe",
          4703 => x"15",
          4704 => x"81",
          4705 => x"84",
          4706 => x"06",
          4707 => x"55",
          4708 => x"f0",
          4709 => x"0d",
          4710 => x"0d",
          4711 => x"5b",
          4712 => x"80",
          4713 => x"ff",
          4714 => x"9f",
          4715 => x"b5",
          4716 => x"f0",
          4717 => x"fe",
          4718 => x"fc",
          4719 => x"7a",
          4720 => x"08",
          4721 => x"64",
          4722 => x"2e",
          4723 => x"a0",
          4724 => x"70",
          4725 => x"ea",
          4726 => x"f0",
          4727 => x"fe",
          4728 => x"d4",
          4729 => x"7b",
          4730 => x"3f",
          4731 => x"08",
          4732 => x"f0",
          4733 => x"38",
          4734 => x"51",
          4735 => x"81",
          4736 => x"45",
          4737 => x"51",
          4738 => x"81",
          4739 => x"57",
          4740 => x"08",
          4741 => x"80",
          4742 => x"da",
          4743 => x"fe",
          4744 => x"81",
          4745 => x"a4",
          4746 => x"7b",
          4747 => x"3f",
          4748 => x"f0",
          4749 => x"38",
          4750 => x"51",
          4751 => x"81",
          4752 => x"57",
          4753 => x"08",
          4754 => x"38",
          4755 => x"09",
          4756 => x"38",
          4757 => x"e0",
          4758 => x"dc",
          4759 => x"ff",
          4760 => x"74",
          4761 => x"3f",
          4762 => x"78",
          4763 => x"33",
          4764 => x"56",
          4765 => x"91",
          4766 => x"05",
          4767 => x"81",
          4768 => x"56",
          4769 => x"f5",
          4770 => x"54",
          4771 => x"81",
          4772 => x"80",
          4773 => x"78",
          4774 => x"55",
          4775 => x"11",
          4776 => x"18",
          4777 => x"58",
          4778 => x"34",
          4779 => x"ff",
          4780 => x"55",
          4781 => x"34",
          4782 => x"77",
          4783 => x"81",
          4784 => x"ff",
          4785 => x"55",
          4786 => x"34",
          4787 => x"ff",
          4788 => x"84",
          4789 => x"cc",
          4790 => x"70",
          4791 => x"56",
          4792 => x"76",
          4793 => x"81",
          4794 => x"70",
          4795 => x"56",
          4796 => x"82",
          4797 => x"78",
          4798 => x"80",
          4799 => x"27",
          4800 => x"19",
          4801 => x"7a",
          4802 => x"5c",
          4803 => x"55",
          4804 => x"7a",
          4805 => x"5c",
          4806 => x"2e",
          4807 => x"85",
          4808 => x"94",
          4809 => x"81",
          4810 => x"73",
          4811 => x"81",
          4812 => x"7a",
          4813 => x"38",
          4814 => x"76",
          4815 => x"0c",
          4816 => x"04",
          4817 => x"7b",
          4818 => x"fc",
          4819 => x"53",
          4820 => x"bb",
          4821 => x"f0",
          4822 => x"fe",
          4823 => x"fa",
          4824 => x"33",
          4825 => x"f2",
          4826 => x"08",
          4827 => x"27",
          4828 => x"15",
          4829 => x"2a",
          4830 => x"51",
          4831 => x"83",
          4832 => x"94",
          4833 => x"80",
          4834 => x"0c",
          4835 => x"2e",
          4836 => x"79",
          4837 => x"70",
          4838 => x"51",
          4839 => x"2e",
          4840 => x"52",
          4841 => x"fe",
          4842 => x"81",
          4843 => x"ff",
          4844 => x"70",
          4845 => x"fe",
          4846 => x"81",
          4847 => x"73",
          4848 => x"76",
          4849 => x"06",
          4850 => x"0c",
          4851 => x"98",
          4852 => x"58",
          4853 => x"39",
          4854 => x"54",
          4855 => x"73",
          4856 => x"cd",
          4857 => x"fe",
          4858 => x"81",
          4859 => x"81",
          4860 => x"38",
          4861 => x"08",
          4862 => x"9b",
          4863 => x"f0",
          4864 => x"0c",
          4865 => x"0c",
          4866 => x"81",
          4867 => x"76",
          4868 => x"38",
          4869 => x"94",
          4870 => x"94",
          4871 => x"16",
          4872 => x"2a",
          4873 => x"51",
          4874 => x"72",
          4875 => x"38",
          4876 => x"51",
          4877 => x"81",
          4878 => x"54",
          4879 => x"08",
          4880 => x"fe",
          4881 => x"a7",
          4882 => x"74",
          4883 => x"3f",
          4884 => x"08",
          4885 => x"2e",
          4886 => x"74",
          4887 => x"79",
          4888 => x"14",
          4889 => x"38",
          4890 => x"0c",
          4891 => x"94",
          4892 => x"94",
          4893 => x"83",
          4894 => x"72",
          4895 => x"38",
          4896 => x"51",
          4897 => x"81",
          4898 => x"94",
          4899 => x"91",
          4900 => x"53",
          4901 => x"81",
          4902 => x"34",
          4903 => x"39",
          4904 => x"81",
          4905 => x"05",
          4906 => x"08",
          4907 => x"08",
          4908 => x"38",
          4909 => x"0c",
          4910 => x"80",
          4911 => x"72",
          4912 => x"73",
          4913 => x"53",
          4914 => x"8c",
          4915 => x"16",
          4916 => x"38",
          4917 => x"0c",
          4918 => x"81",
          4919 => x"8b",
          4920 => x"f9",
          4921 => x"56",
          4922 => x"80",
          4923 => x"38",
          4924 => x"3d",
          4925 => x"8a",
          4926 => x"51",
          4927 => x"81",
          4928 => x"55",
          4929 => x"08",
          4930 => x"77",
          4931 => x"52",
          4932 => x"b5",
          4933 => x"f0",
          4934 => x"fe",
          4935 => x"c3",
          4936 => x"33",
          4937 => x"55",
          4938 => x"24",
          4939 => x"16",
          4940 => x"2a",
          4941 => x"51",
          4942 => x"80",
          4943 => x"9c",
          4944 => x"77",
          4945 => x"3f",
          4946 => x"08",
          4947 => x"77",
          4948 => x"22",
          4949 => x"74",
          4950 => x"ce",
          4951 => x"fe",
          4952 => x"74",
          4953 => x"81",
          4954 => x"85",
          4955 => x"74",
          4956 => x"38",
          4957 => x"74",
          4958 => x"fe",
          4959 => x"3d",
          4960 => x"3d",
          4961 => x"3d",
          4962 => x"70",
          4963 => x"ff",
          4964 => x"f0",
          4965 => x"81",
          4966 => x"73",
          4967 => x"0d",
          4968 => x"0d",
          4969 => x"3d",
          4970 => x"71",
          4971 => x"e7",
          4972 => x"fe",
          4973 => x"81",
          4974 => x"80",
          4975 => x"93",
          4976 => x"f0",
          4977 => x"51",
          4978 => x"81",
          4979 => x"53",
          4980 => x"81",
          4981 => x"52",
          4982 => x"ac",
          4983 => x"f0",
          4984 => x"fe",
          4985 => x"2e",
          4986 => x"85",
          4987 => x"87",
          4988 => x"f0",
          4989 => x"74",
          4990 => x"d5",
          4991 => x"52",
          4992 => x"89",
          4993 => x"f0",
          4994 => x"70",
          4995 => x"07",
          4996 => x"81",
          4997 => x"06",
          4998 => x"54",
          4999 => x"f0",
          5000 => x"0d",
          5001 => x"0d",
          5002 => x"53",
          5003 => x"53",
          5004 => x"56",
          5005 => x"81",
          5006 => x"55",
          5007 => x"08",
          5008 => x"52",
          5009 => x"81",
          5010 => x"f0",
          5011 => x"fe",
          5012 => x"38",
          5013 => x"05",
          5014 => x"2b",
          5015 => x"80",
          5016 => x"86",
          5017 => x"76",
          5018 => x"38",
          5019 => x"51",
          5020 => x"74",
          5021 => x"0c",
          5022 => x"04",
          5023 => x"63",
          5024 => x"80",
          5025 => x"ec",
          5026 => x"3d",
          5027 => x"3f",
          5028 => x"08",
          5029 => x"f0",
          5030 => x"38",
          5031 => x"73",
          5032 => x"08",
          5033 => x"13",
          5034 => x"58",
          5035 => x"26",
          5036 => x"7c",
          5037 => x"39",
          5038 => x"cc",
          5039 => x"81",
          5040 => x"fe",
          5041 => x"33",
          5042 => x"81",
          5043 => x"06",
          5044 => x"75",
          5045 => x"52",
          5046 => x"05",
          5047 => x"3f",
          5048 => x"08",
          5049 => x"38",
          5050 => x"08",
          5051 => x"38",
          5052 => x"08",
          5053 => x"fe",
          5054 => x"80",
          5055 => x"81",
          5056 => x"59",
          5057 => x"14",
          5058 => x"ca",
          5059 => x"39",
          5060 => x"81",
          5061 => x"57",
          5062 => x"38",
          5063 => x"18",
          5064 => x"ff",
          5065 => x"81",
          5066 => x"5b",
          5067 => x"08",
          5068 => x"7c",
          5069 => x"12",
          5070 => x"52",
          5071 => x"82",
          5072 => x"06",
          5073 => x"14",
          5074 => x"cb",
          5075 => x"f0",
          5076 => x"ff",
          5077 => x"70",
          5078 => x"82",
          5079 => x"51",
          5080 => x"b4",
          5081 => x"bb",
          5082 => x"fe",
          5083 => x"0a",
          5084 => x"70",
          5085 => x"84",
          5086 => x"51",
          5087 => x"ff",
          5088 => x"56",
          5089 => x"38",
          5090 => x"7c",
          5091 => x"0c",
          5092 => x"81",
          5093 => x"74",
          5094 => x"7a",
          5095 => x"0c",
          5096 => x"04",
          5097 => x"79",
          5098 => x"05",
          5099 => x"57",
          5100 => x"81",
          5101 => x"56",
          5102 => x"08",
          5103 => x"91",
          5104 => x"75",
          5105 => x"90",
          5106 => x"81",
          5107 => x"06",
          5108 => x"87",
          5109 => x"2e",
          5110 => x"94",
          5111 => x"73",
          5112 => x"27",
          5113 => x"73",
          5114 => x"fe",
          5115 => x"88",
          5116 => x"76",
          5117 => x"3f",
          5118 => x"08",
          5119 => x"0c",
          5120 => x"39",
          5121 => x"52",
          5122 => x"bf",
          5123 => x"fe",
          5124 => x"2e",
          5125 => x"83",
          5126 => x"81",
          5127 => x"81",
          5128 => x"06",
          5129 => x"56",
          5130 => x"a0",
          5131 => x"81",
          5132 => x"98",
          5133 => x"94",
          5134 => x"08",
          5135 => x"f0",
          5136 => x"51",
          5137 => x"81",
          5138 => x"56",
          5139 => x"8c",
          5140 => x"17",
          5141 => x"07",
          5142 => x"18",
          5143 => x"2e",
          5144 => x"91",
          5145 => x"55",
          5146 => x"f0",
          5147 => x"0d",
          5148 => x"0d",
          5149 => x"3d",
          5150 => x"52",
          5151 => x"da",
          5152 => x"fe",
          5153 => x"81",
          5154 => x"81",
          5155 => x"45",
          5156 => x"52",
          5157 => x"52",
          5158 => x"3f",
          5159 => x"08",
          5160 => x"f0",
          5161 => x"38",
          5162 => x"05",
          5163 => x"2a",
          5164 => x"51",
          5165 => x"55",
          5166 => x"38",
          5167 => x"54",
          5168 => x"81",
          5169 => x"80",
          5170 => x"70",
          5171 => x"54",
          5172 => x"81",
          5173 => x"52",
          5174 => x"c5",
          5175 => x"f0",
          5176 => x"2a",
          5177 => x"51",
          5178 => x"80",
          5179 => x"38",
          5180 => x"fe",
          5181 => x"15",
          5182 => x"86",
          5183 => x"81",
          5184 => x"5c",
          5185 => x"3d",
          5186 => x"c7",
          5187 => x"fe",
          5188 => x"81",
          5189 => x"80",
          5190 => x"fe",
          5191 => x"73",
          5192 => x"3f",
          5193 => x"08",
          5194 => x"f0",
          5195 => x"87",
          5196 => x"39",
          5197 => x"08",
          5198 => x"38",
          5199 => x"08",
          5200 => x"77",
          5201 => x"3f",
          5202 => x"08",
          5203 => x"08",
          5204 => x"fe",
          5205 => x"80",
          5206 => x"55",
          5207 => x"94",
          5208 => x"2e",
          5209 => x"53",
          5210 => x"51",
          5211 => x"81",
          5212 => x"55",
          5213 => x"78",
          5214 => x"fe",
          5215 => x"f0",
          5216 => x"81",
          5217 => x"a0",
          5218 => x"e9",
          5219 => x"53",
          5220 => x"05",
          5221 => x"51",
          5222 => x"81",
          5223 => x"54",
          5224 => x"08",
          5225 => x"78",
          5226 => x"8e",
          5227 => x"58",
          5228 => x"81",
          5229 => x"54",
          5230 => x"08",
          5231 => x"54",
          5232 => x"81",
          5233 => x"84",
          5234 => x"06",
          5235 => x"02",
          5236 => x"33",
          5237 => x"81",
          5238 => x"86",
          5239 => x"f6",
          5240 => x"74",
          5241 => x"70",
          5242 => x"c3",
          5243 => x"f0",
          5244 => x"56",
          5245 => x"08",
          5246 => x"54",
          5247 => x"08",
          5248 => x"81",
          5249 => x"82",
          5250 => x"f0",
          5251 => x"09",
          5252 => x"38",
          5253 => x"b4",
          5254 => x"b0",
          5255 => x"f0",
          5256 => x"51",
          5257 => x"81",
          5258 => x"54",
          5259 => x"08",
          5260 => x"8b",
          5261 => x"b4",
          5262 => x"b7",
          5263 => x"54",
          5264 => x"15",
          5265 => x"90",
          5266 => x"34",
          5267 => x"0a",
          5268 => x"19",
          5269 => x"9f",
          5270 => x"78",
          5271 => x"51",
          5272 => x"a0",
          5273 => x"11",
          5274 => x"05",
          5275 => x"b6",
          5276 => x"ae",
          5277 => x"15",
          5278 => x"78",
          5279 => x"53",
          5280 => x"3f",
          5281 => x"0b",
          5282 => x"77",
          5283 => x"3f",
          5284 => x"08",
          5285 => x"f0",
          5286 => x"82",
          5287 => x"52",
          5288 => x"51",
          5289 => x"3f",
          5290 => x"52",
          5291 => x"aa",
          5292 => x"90",
          5293 => x"34",
          5294 => x"0b",
          5295 => x"78",
          5296 => x"b6",
          5297 => x"f0",
          5298 => x"39",
          5299 => x"52",
          5300 => x"be",
          5301 => x"81",
          5302 => x"99",
          5303 => x"da",
          5304 => x"3d",
          5305 => x"d2",
          5306 => x"53",
          5307 => x"84",
          5308 => x"3d",
          5309 => x"3f",
          5310 => x"08",
          5311 => x"f0",
          5312 => x"38",
          5313 => x"3d",
          5314 => x"3d",
          5315 => x"cc",
          5316 => x"fe",
          5317 => x"81",
          5318 => x"82",
          5319 => x"81",
          5320 => x"81",
          5321 => x"86",
          5322 => x"aa",
          5323 => x"a4",
          5324 => x"a8",
          5325 => x"05",
          5326 => x"ea",
          5327 => x"77",
          5328 => x"70",
          5329 => x"b4",
          5330 => x"3d",
          5331 => x"51",
          5332 => x"81",
          5333 => x"55",
          5334 => x"08",
          5335 => x"6f",
          5336 => x"06",
          5337 => x"a2",
          5338 => x"92",
          5339 => x"81",
          5340 => x"fe",
          5341 => x"2e",
          5342 => x"81",
          5343 => x"51",
          5344 => x"81",
          5345 => x"55",
          5346 => x"08",
          5347 => x"68",
          5348 => x"a8",
          5349 => x"05",
          5350 => x"51",
          5351 => x"3f",
          5352 => x"33",
          5353 => x"8b",
          5354 => x"84",
          5355 => x"06",
          5356 => x"73",
          5357 => x"a0",
          5358 => x"8b",
          5359 => x"54",
          5360 => x"15",
          5361 => x"33",
          5362 => x"70",
          5363 => x"55",
          5364 => x"2e",
          5365 => x"6e",
          5366 => x"df",
          5367 => x"78",
          5368 => x"3f",
          5369 => x"08",
          5370 => x"ff",
          5371 => x"82",
          5372 => x"f0",
          5373 => x"80",
          5374 => x"fe",
          5375 => x"78",
          5376 => x"af",
          5377 => x"f0",
          5378 => x"d4",
          5379 => x"55",
          5380 => x"08",
          5381 => x"81",
          5382 => x"73",
          5383 => x"81",
          5384 => x"63",
          5385 => x"76",
          5386 => x"3f",
          5387 => x"0b",
          5388 => x"87",
          5389 => x"f0",
          5390 => x"77",
          5391 => x"3f",
          5392 => x"08",
          5393 => x"f0",
          5394 => x"78",
          5395 => x"aa",
          5396 => x"f0",
          5397 => x"81",
          5398 => x"a8",
          5399 => x"ed",
          5400 => x"80",
          5401 => x"02",
          5402 => x"df",
          5403 => x"57",
          5404 => x"3d",
          5405 => x"96",
          5406 => x"e9",
          5407 => x"f0",
          5408 => x"fe",
          5409 => x"cf",
          5410 => x"65",
          5411 => x"d4",
          5412 => x"b5",
          5413 => x"f0",
          5414 => x"fe",
          5415 => x"38",
          5416 => x"05",
          5417 => x"06",
          5418 => x"73",
          5419 => x"a7",
          5420 => x"09",
          5421 => x"71",
          5422 => x"06",
          5423 => x"55",
          5424 => x"15",
          5425 => x"81",
          5426 => x"34",
          5427 => x"b4",
          5428 => x"fe",
          5429 => x"74",
          5430 => x"0c",
          5431 => x"04",
          5432 => x"64",
          5433 => x"93",
          5434 => x"52",
          5435 => x"d1",
          5436 => x"fe",
          5437 => x"81",
          5438 => x"80",
          5439 => x"58",
          5440 => x"3d",
          5441 => x"c8",
          5442 => x"fe",
          5443 => x"81",
          5444 => x"b4",
          5445 => x"c7",
          5446 => x"a0",
          5447 => x"55",
          5448 => x"84",
          5449 => x"17",
          5450 => x"2b",
          5451 => x"96",
          5452 => x"b0",
          5453 => x"54",
          5454 => x"15",
          5455 => x"ff",
          5456 => x"81",
          5457 => x"55",
          5458 => x"f0",
          5459 => x"0d",
          5460 => x"0d",
          5461 => x"5a",
          5462 => x"3d",
          5463 => x"99",
          5464 => x"81",
          5465 => x"f0",
          5466 => x"f0",
          5467 => x"81",
          5468 => x"07",
          5469 => x"55",
          5470 => x"2e",
          5471 => x"81",
          5472 => x"55",
          5473 => x"2e",
          5474 => x"7b",
          5475 => x"80",
          5476 => x"70",
          5477 => x"be",
          5478 => x"fe",
          5479 => x"81",
          5480 => x"80",
          5481 => x"52",
          5482 => x"dc",
          5483 => x"f0",
          5484 => x"fe",
          5485 => x"38",
          5486 => x"08",
          5487 => x"08",
          5488 => x"56",
          5489 => x"19",
          5490 => x"59",
          5491 => x"74",
          5492 => x"56",
          5493 => x"ec",
          5494 => x"75",
          5495 => x"74",
          5496 => x"2e",
          5497 => x"16",
          5498 => x"33",
          5499 => x"73",
          5500 => x"38",
          5501 => x"84",
          5502 => x"06",
          5503 => x"7a",
          5504 => x"76",
          5505 => x"07",
          5506 => x"54",
          5507 => x"80",
          5508 => x"80",
          5509 => x"7b",
          5510 => x"53",
          5511 => x"93",
          5512 => x"f0",
          5513 => x"fe",
          5514 => x"38",
          5515 => x"55",
          5516 => x"56",
          5517 => x"8b",
          5518 => x"56",
          5519 => x"83",
          5520 => x"75",
          5521 => x"51",
          5522 => x"3f",
          5523 => x"08",
          5524 => x"81",
          5525 => x"98",
          5526 => x"e6",
          5527 => x"53",
          5528 => x"b8",
          5529 => x"3d",
          5530 => x"3f",
          5531 => x"08",
          5532 => x"08",
          5533 => x"fe",
          5534 => x"98",
          5535 => x"a0",
          5536 => x"70",
          5537 => x"ae",
          5538 => x"6d",
          5539 => x"81",
          5540 => x"57",
          5541 => x"74",
          5542 => x"38",
          5543 => x"81",
          5544 => x"81",
          5545 => x"52",
          5546 => x"89",
          5547 => x"f0",
          5548 => x"a5",
          5549 => x"33",
          5550 => x"54",
          5551 => x"3f",
          5552 => x"08",
          5553 => x"38",
          5554 => x"76",
          5555 => x"05",
          5556 => x"39",
          5557 => x"08",
          5558 => x"15",
          5559 => x"ff",
          5560 => x"73",
          5561 => x"38",
          5562 => x"83",
          5563 => x"56",
          5564 => x"75",
          5565 => x"81",
          5566 => x"33",
          5567 => x"2e",
          5568 => x"52",
          5569 => x"51",
          5570 => x"3f",
          5571 => x"08",
          5572 => x"ff",
          5573 => x"38",
          5574 => x"88",
          5575 => x"8a",
          5576 => x"38",
          5577 => x"ec",
          5578 => x"75",
          5579 => x"74",
          5580 => x"73",
          5581 => x"05",
          5582 => x"17",
          5583 => x"70",
          5584 => x"34",
          5585 => x"70",
          5586 => x"ff",
          5587 => x"55",
          5588 => x"26",
          5589 => x"8b",
          5590 => x"86",
          5591 => x"e5",
          5592 => x"38",
          5593 => x"99",
          5594 => x"05",
          5595 => x"70",
          5596 => x"73",
          5597 => x"81",
          5598 => x"ff",
          5599 => x"ed",
          5600 => x"80",
          5601 => x"91",
          5602 => x"55",
          5603 => x"3f",
          5604 => x"08",
          5605 => x"f0",
          5606 => x"38",
          5607 => x"51",
          5608 => x"3f",
          5609 => x"08",
          5610 => x"f0",
          5611 => x"76",
          5612 => x"67",
          5613 => x"34",
          5614 => x"81",
          5615 => x"84",
          5616 => x"06",
          5617 => x"80",
          5618 => x"2e",
          5619 => x"81",
          5620 => x"ff",
          5621 => x"81",
          5622 => x"54",
          5623 => x"08",
          5624 => x"53",
          5625 => x"08",
          5626 => x"ff",
          5627 => x"67",
          5628 => x"8b",
          5629 => x"53",
          5630 => x"51",
          5631 => x"3f",
          5632 => x"0b",
          5633 => x"79",
          5634 => x"ee",
          5635 => x"f0",
          5636 => x"55",
          5637 => x"f0",
          5638 => x"0d",
          5639 => x"0d",
          5640 => x"88",
          5641 => x"05",
          5642 => x"fc",
          5643 => x"54",
          5644 => x"d2",
          5645 => x"fe",
          5646 => x"81",
          5647 => x"82",
          5648 => x"1a",
          5649 => x"82",
          5650 => x"80",
          5651 => x"8c",
          5652 => x"78",
          5653 => x"1a",
          5654 => x"2a",
          5655 => x"51",
          5656 => x"90",
          5657 => x"82",
          5658 => x"58",
          5659 => x"81",
          5660 => x"39",
          5661 => x"22",
          5662 => x"70",
          5663 => x"56",
          5664 => x"e2",
          5665 => x"14",
          5666 => x"30",
          5667 => x"9f",
          5668 => x"f0",
          5669 => x"19",
          5670 => x"5a",
          5671 => x"81",
          5672 => x"38",
          5673 => x"77",
          5674 => x"82",
          5675 => x"56",
          5676 => x"74",
          5677 => x"ff",
          5678 => x"81",
          5679 => x"55",
          5680 => x"75",
          5681 => x"82",
          5682 => x"f0",
          5683 => x"ff",
          5684 => x"fe",
          5685 => x"2e",
          5686 => x"81",
          5687 => x"8e",
          5688 => x"56",
          5689 => x"09",
          5690 => x"38",
          5691 => x"59",
          5692 => x"77",
          5693 => x"06",
          5694 => x"87",
          5695 => x"39",
          5696 => x"ba",
          5697 => x"55",
          5698 => x"2e",
          5699 => x"15",
          5700 => x"2e",
          5701 => x"83",
          5702 => x"75",
          5703 => x"7e",
          5704 => x"a8",
          5705 => x"f0",
          5706 => x"fe",
          5707 => x"ce",
          5708 => x"16",
          5709 => x"56",
          5710 => x"38",
          5711 => x"19",
          5712 => x"8c",
          5713 => x"7d",
          5714 => x"38",
          5715 => x"0c",
          5716 => x"0c",
          5717 => x"80",
          5718 => x"73",
          5719 => x"98",
          5720 => x"05",
          5721 => x"57",
          5722 => x"26",
          5723 => x"7b",
          5724 => x"0c",
          5725 => x"81",
          5726 => x"84",
          5727 => x"54",
          5728 => x"f0",
          5729 => x"0d",
          5730 => x"0d",
          5731 => x"88",
          5732 => x"05",
          5733 => x"54",
          5734 => x"c5",
          5735 => x"56",
          5736 => x"fe",
          5737 => x"8b",
          5738 => x"fe",
          5739 => x"29",
          5740 => x"05",
          5741 => x"55",
          5742 => x"84",
          5743 => x"34",
          5744 => x"08",
          5745 => x"5f",
          5746 => x"51",
          5747 => x"3f",
          5748 => x"08",
          5749 => x"70",
          5750 => x"57",
          5751 => x"8b",
          5752 => x"82",
          5753 => x"06",
          5754 => x"56",
          5755 => x"38",
          5756 => x"05",
          5757 => x"7e",
          5758 => x"f0",
          5759 => x"f0",
          5760 => x"67",
          5761 => x"2e",
          5762 => x"82",
          5763 => x"8b",
          5764 => x"75",
          5765 => x"80",
          5766 => x"81",
          5767 => x"2e",
          5768 => x"80",
          5769 => x"38",
          5770 => x"0a",
          5771 => x"ff",
          5772 => x"55",
          5773 => x"86",
          5774 => x"8a",
          5775 => x"89",
          5776 => x"2a",
          5777 => x"77",
          5778 => x"59",
          5779 => x"81",
          5780 => x"70",
          5781 => x"07",
          5782 => x"56",
          5783 => x"38",
          5784 => x"05",
          5785 => x"7e",
          5786 => x"80",
          5787 => x"81",
          5788 => x"8a",
          5789 => x"83",
          5790 => x"06",
          5791 => x"08",
          5792 => x"74",
          5793 => x"41",
          5794 => x"56",
          5795 => x"8a",
          5796 => x"61",
          5797 => x"55",
          5798 => x"27",
          5799 => x"93",
          5800 => x"80",
          5801 => x"38",
          5802 => x"70",
          5803 => x"43",
          5804 => x"95",
          5805 => x"06",
          5806 => x"2e",
          5807 => x"77",
          5808 => x"74",
          5809 => x"83",
          5810 => x"06",
          5811 => x"82",
          5812 => x"2e",
          5813 => x"78",
          5814 => x"2e",
          5815 => x"80",
          5816 => x"ae",
          5817 => x"2a",
          5818 => x"81",
          5819 => x"56",
          5820 => x"2e",
          5821 => x"77",
          5822 => x"81",
          5823 => x"79",
          5824 => x"70",
          5825 => x"5a",
          5826 => x"86",
          5827 => x"27",
          5828 => x"52",
          5829 => x"dd",
          5830 => x"fe",
          5831 => x"29",
          5832 => x"70",
          5833 => x"55",
          5834 => x"0b",
          5835 => x"08",
          5836 => x"05",
          5837 => x"ff",
          5838 => x"27",
          5839 => x"88",
          5840 => x"ae",
          5841 => x"2a",
          5842 => x"81",
          5843 => x"56",
          5844 => x"2e",
          5845 => x"77",
          5846 => x"81",
          5847 => x"79",
          5848 => x"70",
          5849 => x"5a",
          5850 => x"86",
          5851 => x"27",
          5852 => x"52",
          5853 => x"dc",
          5854 => x"fe",
          5855 => x"84",
          5856 => x"fe",
          5857 => x"f5",
          5858 => x"81",
          5859 => x"f0",
          5860 => x"fe",
          5861 => x"71",
          5862 => x"83",
          5863 => x"5e",
          5864 => x"89",
          5865 => x"5c",
          5866 => x"1c",
          5867 => x"05",
          5868 => x"ff",
          5869 => x"70",
          5870 => x"31",
          5871 => x"57",
          5872 => x"83",
          5873 => x"06",
          5874 => x"1c",
          5875 => x"5c",
          5876 => x"1d",
          5877 => x"29",
          5878 => x"31",
          5879 => x"55",
          5880 => x"87",
          5881 => x"7c",
          5882 => x"7a",
          5883 => x"31",
          5884 => x"db",
          5885 => x"fe",
          5886 => x"7d",
          5887 => x"81",
          5888 => x"81",
          5889 => x"83",
          5890 => x"80",
          5891 => x"87",
          5892 => x"81",
          5893 => x"fd",
          5894 => x"f8",
          5895 => x"2e",
          5896 => x"80",
          5897 => x"ff",
          5898 => x"fe",
          5899 => x"a0",
          5900 => x"38",
          5901 => x"74",
          5902 => x"86",
          5903 => x"fd",
          5904 => x"81",
          5905 => x"80",
          5906 => x"83",
          5907 => x"39",
          5908 => x"08",
          5909 => x"92",
          5910 => x"b8",
          5911 => x"59",
          5912 => x"27",
          5913 => x"86",
          5914 => x"55",
          5915 => x"09",
          5916 => x"38",
          5917 => x"f5",
          5918 => x"38",
          5919 => x"55",
          5920 => x"86",
          5921 => x"80",
          5922 => x"7a",
          5923 => x"b9",
          5924 => x"81",
          5925 => x"7a",
          5926 => x"8a",
          5927 => x"52",
          5928 => x"ff",
          5929 => x"79",
          5930 => x"7b",
          5931 => x"06",
          5932 => x"51",
          5933 => x"3f",
          5934 => x"1c",
          5935 => x"32",
          5936 => x"96",
          5937 => x"06",
          5938 => x"91",
          5939 => x"a1",
          5940 => x"55",
          5941 => x"ff",
          5942 => x"74",
          5943 => x"06",
          5944 => x"51",
          5945 => x"3f",
          5946 => x"52",
          5947 => x"ff",
          5948 => x"f8",
          5949 => x"34",
          5950 => x"1b",
          5951 => x"d9",
          5952 => x"52",
          5953 => x"ff",
          5954 => x"60",
          5955 => x"51",
          5956 => x"3f",
          5957 => x"09",
          5958 => x"cb",
          5959 => x"b2",
          5960 => x"c3",
          5961 => x"a0",
          5962 => x"52",
          5963 => x"ff",
          5964 => x"82",
          5965 => x"51",
          5966 => x"3f",
          5967 => x"1b",
          5968 => x"95",
          5969 => x"b2",
          5970 => x"a0",
          5971 => x"80",
          5972 => x"1c",
          5973 => x"80",
          5974 => x"93",
          5975 => x"a4",
          5976 => x"1b",
          5977 => x"82",
          5978 => x"52",
          5979 => x"ff",
          5980 => x"7c",
          5981 => x"06",
          5982 => x"51",
          5983 => x"3f",
          5984 => x"a4",
          5985 => x"0b",
          5986 => x"93",
          5987 => x"b8",
          5988 => x"51",
          5989 => x"3f",
          5990 => x"52",
          5991 => x"70",
          5992 => x"9f",
          5993 => x"54",
          5994 => x"52",
          5995 => x"9b",
          5996 => x"56",
          5997 => x"08",
          5998 => x"7d",
          5999 => x"81",
          6000 => x"38",
          6001 => x"86",
          6002 => x"52",
          6003 => x"9b",
          6004 => x"80",
          6005 => x"7a",
          6006 => x"ed",
          6007 => x"85",
          6008 => x"7a",
          6009 => x"8f",
          6010 => x"85",
          6011 => x"83",
          6012 => x"ff",
          6013 => x"ff",
          6014 => x"e8",
          6015 => x"9e",
          6016 => x"52",
          6017 => x"51",
          6018 => x"3f",
          6019 => x"52",
          6020 => x"9e",
          6021 => x"54",
          6022 => x"53",
          6023 => x"51",
          6024 => x"3f",
          6025 => x"16",
          6026 => x"7e",
          6027 => x"d8",
          6028 => x"80",
          6029 => x"ff",
          6030 => x"7f",
          6031 => x"7d",
          6032 => x"81",
          6033 => x"f8",
          6034 => x"ff",
          6035 => x"ff",
          6036 => x"51",
          6037 => x"3f",
          6038 => x"88",
          6039 => x"39",
          6040 => x"f8",
          6041 => x"2e",
          6042 => x"55",
          6043 => x"51",
          6044 => x"3f",
          6045 => x"57",
          6046 => x"83",
          6047 => x"76",
          6048 => x"7a",
          6049 => x"ff",
          6050 => x"81",
          6051 => x"82",
          6052 => x"80",
          6053 => x"f0",
          6054 => x"51",
          6055 => x"3f",
          6056 => x"78",
          6057 => x"74",
          6058 => x"18",
          6059 => x"2e",
          6060 => x"79",
          6061 => x"2e",
          6062 => x"55",
          6063 => x"62",
          6064 => x"74",
          6065 => x"75",
          6066 => x"7e",
          6067 => x"b8",
          6068 => x"f0",
          6069 => x"38",
          6070 => x"78",
          6071 => x"74",
          6072 => x"56",
          6073 => x"93",
          6074 => x"66",
          6075 => x"26",
          6076 => x"56",
          6077 => x"83",
          6078 => x"64",
          6079 => x"77",
          6080 => x"84",
          6081 => x"52",
          6082 => x"9d",
          6083 => x"d4",
          6084 => x"51",
          6085 => x"3f",
          6086 => x"55",
          6087 => x"81",
          6088 => x"34",
          6089 => x"16",
          6090 => x"16",
          6091 => x"16",
          6092 => x"05",
          6093 => x"c1",
          6094 => x"fe",
          6095 => x"fe",
          6096 => x"34",
          6097 => x"08",
          6098 => x"07",
          6099 => x"16",
          6100 => x"f0",
          6101 => x"34",
          6102 => x"c6",
          6103 => x"9c",
          6104 => x"52",
          6105 => x"51",
          6106 => x"3f",
          6107 => x"53",
          6108 => x"51",
          6109 => x"3f",
          6110 => x"fe",
          6111 => x"38",
          6112 => x"52",
          6113 => x"99",
          6114 => x"56",
          6115 => x"08",
          6116 => x"39",
          6117 => x"39",
          6118 => x"39",
          6119 => x"08",
          6120 => x"fe",
          6121 => x"3d",
          6122 => x"3d",
          6123 => x"5b",
          6124 => x"60",
          6125 => x"57",
          6126 => x"25",
          6127 => x"3d",
          6128 => x"55",
          6129 => x"15",
          6130 => x"c9",
          6131 => x"81",
          6132 => x"06",
          6133 => x"3d",
          6134 => x"8d",
          6135 => x"74",
          6136 => x"05",
          6137 => x"17",
          6138 => x"2e",
          6139 => x"c9",
          6140 => x"34",
          6141 => x"83",
          6142 => x"74",
          6143 => x"0c",
          6144 => x"04",
          6145 => x"7b",
          6146 => x"b3",
          6147 => x"57",
          6148 => x"09",
          6149 => x"38",
          6150 => x"51",
          6151 => x"17",
          6152 => x"76",
          6153 => x"88",
          6154 => x"17",
          6155 => x"59",
          6156 => x"81",
          6157 => x"76",
          6158 => x"8b",
          6159 => x"54",
          6160 => x"17",
          6161 => x"51",
          6162 => x"79",
          6163 => x"30",
          6164 => x"9f",
          6165 => x"53",
          6166 => x"75",
          6167 => x"81",
          6168 => x"0c",
          6169 => x"04",
          6170 => x"79",
          6171 => x"56",
          6172 => x"24",
          6173 => x"3d",
          6174 => x"74",
          6175 => x"52",
          6176 => x"cb",
          6177 => x"fe",
          6178 => x"38",
          6179 => x"78",
          6180 => x"06",
          6181 => x"16",
          6182 => x"39",
          6183 => x"81",
          6184 => x"89",
          6185 => x"fd",
          6186 => x"54",
          6187 => x"80",
          6188 => x"ff",
          6189 => x"76",
          6190 => x"3d",
          6191 => x"3d",
          6192 => x"e3",
          6193 => x"53",
          6194 => x"53",
          6195 => x"3f",
          6196 => x"51",
          6197 => x"72",
          6198 => x"3f",
          6199 => x"04",
          6200 => x"7a",
          6201 => x"56",
          6202 => x"80",
          6203 => x"38",
          6204 => x"15",
          6205 => x"16",
          6206 => x"d4",
          6207 => x"54",
          6208 => x"09",
          6209 => x"38",
          6210 => x"f1",
          6211 => x"76",
          6212 => x"fb",
          6213 => x"08",
          6214 => x"da",
          6215 => x"fe",
          6216 => x"fe",
          6217 => x"75",
          6218 => x"52",
          6219 => x"ff",
          6220 => x"f0",
          6221 => x"84",
          6222 => x"73",
          6223 => x"b2",
          6224 => x"70",
          6225 => x"58",
          6226 => x"27",
          6227 => x"54",
          6228 => x"f0",
          6229 => x"0d",
          6230 => x"0d",
          6231 => x"93",
          6232 => x"38",
          6233 => x"81",
          6234 => x"52",
          6235 => x"81",
          6236 => x"81",
          6237 => x"ee",
          6238 => x"f9",
          6239 => x"d8",
          6240 => x"39",
          6241 => x"51",
          6242 => x"81",
          6243 => x"80",
          6244 => x"ef",
          6245 => x"dd",
          6246 => x"a0",
          6247 => x"39",
          6248 => x"51",
          6249 => x"81",
          6250 => x"80",
          6251 => x"ef",
          6252 => x"c1",
          6253 => x"f8",
          6254 => x"81",
          6255 => x"b5",
          6256 => x"a8",
          6257 => x"81",
          6258 => x"a9",
          6259 => x"e8",
          6260 => x"81",
          6261 => x"9d",
          6262 => x"9c",
          6263 => x"81",
          6264 => x"91",
          6265 => x"cc",
          6266 => x"81",
          6267 => x"85",
          6268 => x"f0",
          6269 => x"ae",
          6270 => x"0d",
          6271 => x"0d",
          6272 => x"56",
          6273 => x"26",
          6274 => x"52",
          6275 => x"29",
          6276 => x"87",
          6277 => x"51",
          6278 => x"3f",
          6279 => x"08",
          6280 => x"fe",
          6281 => x"81",
          6282 => x"54",
          6283 => x"52",
          6284 => x"51",
          6285 => x"3f",
          6286 => x"04",
          6287 => x"66",
          6288 => x"80",
          6289 => x"5b",
          6290 => x"78",
          6291 => x"07",
          6292 => x"57",
          6293 => x"56",
          6294 => x"26",
          6295 => x"56",
          6296 => x"70",
          6297 => x"51",
          6298 => x"74",
          6299 => x"81",
          6300 => x"8c",
          6301 => x"56",
          6302 => x"3f",
          6303 => x"08",
          6304 => x"f0",
          6305 => x"81",
          6306 => x"87",
          6307 => x"0c",
          6308 => x"08",
          6309 => x"d4",
          6310 => x"80",
          6311 => x"75",
          6312 => x"3f",
          6313 => x"08",
          6314 => x"f0",
          6315 => x"7a",
          6316 => x"2e",
          6317 => x"19",
          6318 => x"59",
          6319 => x"3d",
          6320 => x"cb",
          6321 => x"30",
          6322 => x"80",
          6323 => x"70",
          6324 => x"06",
          6325 => x"56",
          6326 => x"90",
          6327 => x"a4",
          6328 => x"98",
          6329 => x"78",
          6330 => x"3f",
          6331 => x"81",
          6332 => x"96",
          6333 => x"f9",
          6334 => x"02",
          6335 => x"05",
          6336 => x"ff",
          6337 => x"7a",
          6338 => x"fe",
          6339 => x"fe",
          6340 => x"38",
          6341 => x"88",
          6342 => x"2e",
          6343 => x"39",
          6344 => x"54",
          6345 => x"53",
          6346 => x"51",
          6347 => x"fe",
          6348 => x"83",
          6349 => x"76",
          6350 => x"0c",
          6351 => x"04",
          6352 => x"7f",
          6353 => x"8c",
          6354 => x"05",
          6355 => x"15",
          6356 => x"5c",
          6357 => x"5e",
          6358 => x"f2",
          6359 => x"f5",
          6360 => x"f2",
          6361 => x"ef",
          6362 => x"55",
          6363 => x"80",
          6364 => x"90",
          6365 => x"7b",
          6366 => x"38",
          6367 => x"74",
          6368 => x"7a",
          6369 => x"72",
          6370 => x"f2",
          6371 => x"f4",
          6372 => x"39",
          6373 => x"51",
          6374 => x"3f",
          6375 => x"80",
          6376 => x"18",
          6377 => x"27",
          6378 => x"08",
          6379 => x"ac",
          6380 => x"d6",
          6381 => x"81",
          6382 => x"fe",
          6383 => x"84",
          6384 => x"39",
          6385 => x"72",
          6386 => x"38",
          6387 => x"81",
          6388 => x"fe",
          6389 => x"89",
          6390 => x"d4",
          6391 => x"c6",
          6392 => x"55",
          6393 => x"ed",
          6394 => x"80",
          6395 => x"d8",
          6396 => x"b2",
          6397 => x"74",
          6398 => x"38",
          6399 => x"33",
          6400 => x"56",
          6401 => x"83",
          6402 => x"80",
          6403 => x"27",
          6404 => x"53",
          6405 => x"70",
          6406 => x"51",
          6407 => x"2e",
          6408 => x"80",
          6409 => x"38",
          6410 => x"39",
          6411 => x"ed",
          6412 => x"15",
          6413 => x"81",
          6414 => x"fe",
          6415 => x"78",
          6416 => x"5c",
          6417 => x"96",
          6418 => x"f0",
          6419 => x"70",
          6420 => x"57",
          6421 => x"09",
          6422 => x"38",
          6423 => x"3f",
          6424 => x"08",
          6425 => x"98",
          6426 => x"32",
          6427 => x"9b",
          6428 => x"70",
          6429 => x"75",
          6430 => x"58",
          6431 => x"51",
          6432 => x"24",
          6433 => x"9b",
          6434 => x"06",
          6435 => x"53",
          6436 => x"1e",
          6437 => x"26",
          6438 => x"ff",
          6439 => x"fe",
          6440 => x"3d",
          6441 => x"3d",
          6442 => x"05",
          6443 => x"e0",
          6444 => x"e8",
          6445 => x"f2",
          6446 => x"fa",
          6447 => x"fe",
          6448 => x"81",
          6449 => x"81",
          6450 => x"81",
          6451 => x"52",
          6452 => x"51",
          6453 => x"3f",
          6454 => x"85",
          6455 => x"a2",
          6456 => x"0d",
          6457 => x"0d",
          6458 => x"80",
          6459 => x"e7",
          6460 => x"51",
          6461 => x"3f",
          6462 => x"51",
          6463 => x"3f",
          6464 => x"d8",
          6465 => x"81",
          6466 => x"06",
          6467 => x"80",
          6468 => x"81",
          6469 => x"da",
          6470 => x"c0",
          6471 => x"d2",
          6472 => x"fe",
          6473 => x"72",
          6474 => x"81",
          6475 => x"71",
          6476 => x"38",
          6477 => x"d8",
          6478 => x"f3",
          6479 => x"da",
          6480 => x"51",
          6481 => x"3f",
          6482 => x"70",
          6483 => x"52",
          6484 => x"95",
          6485 => x"fe",
          6486 => x"81",
          6487 => x"fe",
          6488 => x"80",
          6489 => x"8a",
          6490 => x"2a",
          6491 => x"51",
          6492 => x"2e",
          6493 => x"51",
          6494 => x"3f",
          6495 => x"51",
          6496 => x"3f",
          6497 => x"d7",
          6498 => x"85",
          6499 => x"06",
          6500 => x"80",
          6501 => x"81",
          6502 => x"d6",
          6503 => x"8c",
          6504 => x"ce",
          6505 => x"fe",
          6506 => x"72",
          6507 => x"81",
          6508 => x"71",
          6509 => x"38",
          6510 => x"d7",
          6511 => x"f4",
          6512 => x"d9",
          6513 => x"51",
          6514 => x"3f",
          6515 => x"70",
          6516 => x"52",
          6517 => x"95",
          6518 => x"fe",
          6519 => x"81",
          6520 => x"fe",
          6521 => x"80",
          6522 => x"86",
          6523 => x"2a",
          6524 => x"51",
          6525 => x"2e",
          6526 => x"51",
          6527 => x"3f",
          6528 => x"51",
          6529 => x"3f",
          6530 => x"d6",
          6531 => x"e5",
          6532 => x"3d",
          6533 => x"3d",
          6534 => x"84",
          6535 => x"33",
          6536 => x"56",
          6537 => x"51",
          6538 => x"3f",
          6539 => x"33",
          6540 => x"38",
          6541 => x"f5",
          6542 => x"96",
          6543 => x"b8",
          6544 => x"fe",
          6545 => x"70",
          6546 => x"08",
          6547 => x"82",
          6548 => x"51",
          6549 => x"fb",
          6550 => x"fb",
          6551 => x"73",
          6552 => x"81",
          6553 => x"82",
          6554 => x"74",
          6555 => x"f2",
          6556 => x"fe",
          6557 => x"2e",
          6558 => x"fe",
          6559 => x"fe",
          6560 => x"8e",
          6561 => x"88",
          6562 => x"3f",
          6563 => x"fb",
          6564 => x"fb",
          6565 => x"73",
          6566 => x"81",
          6567 => x"74",
          6568 => x"fe",
          6569 => x"80",
          6570 => x"f0",
          6571 => x"0d",
          6572 => x"0d",
          6573 => x"82",
          6574 => x"5f",
          6575 => x"7c",
          6576 => x"db",
          6577 => x"f0",
          6578 => x"06",
          6579 => x"2e",
          6580 => x"a2",
          6581 => x"98",
          6582 => x"70",
          6583 => x"ee",
          6584 => x"53",
          6585 => x"80",
          6586 => x"b5",
          6587 => x"fe",
          6588 => x"2e",
          6589 => x"f5",
          6590 => x"fe",
          6591 => x"5f",
          6592 => x"d4",
          6593 => x"9e",
          6594 => x"70",
          6595 => x"f8",
          6596 => x"fe",
          6597 => x"3d",
          6598 => x"51",
          6599 => x"81",
          6600 => x"90",
          6601 => x"2c",
          6602 => x"80",
          6603 => x"f1",
          6604 => x"c1",
          6605 => x"38",
          6606 => x"83",
          6607 => x"ab",
          6608 => x"78",
          6609 => x"b3",
          6610 => x"24",
          6611 => x"80",
          6612 => x"38",
          6613 => x"78",
          6614 => x"86",
          6615 => x"2e",
          6616 => x"8f",
          6617 => x"bd",
          6618 => x"38",
          6619 => x"90",
          6620 => x"2e",
          6621 => x"78",
          6622 => x"91",
          6623 => x"39",
          6624 => x"85",
          6625 => x"80",
          6626 => x"d2",
          6627 => x"39",
          6628 => x"2e",
          6629 => x"78",
          6630 => x"b0",
          6631 => x"d0",
          6632 => x"38",
          6633 => x"24",
          6634 => x"80",
          6635 => x"99",
          6636 => x"c3",
          6637 => x"38",
          6638 => x"78",
          6639 => x"8c",
          6640 => x"80",
          6641 => x"f3",
          6642 => x"39",
          6643 => x"2e",
          6644 => x"78",
          6645 => x"92",
          6646 => x"f8",
          6647 => x"38",
          6648 => x"2e",
          6649 => x"8e",
          6650 => x"81",
          6651 => x"f7",
          6652 => x"85",
          6653 => x"38",
          6654 => x"b4",
          6655 => x"11",
          6656 => x"05",
          6657 => x"f7",
          6658 => x"f0",
          6659 => x"81",
          6660 => x"8f",
          6661 => x"3d",
          6662 => x"53",
          6663 => x"51",
          6664 => x"3f",
          6665 => x"08",
          6666 => x"38",
          6667 => x"83",
          6668 => x"02",
          6669 => x"33",
          6670 => x"cf",
          6671 => x"ff",
          6672 => x"81",
          6673 => x"81",
          6674 => x"78",
          6675 => x"f5",
          6676 => x"e5",
          6677 => x"5e",
          6678 => x"81",
          6679 => x"87",
          6680 => x"3d",
          6681 => x"53",
          6682 => x"51",
          6683 => x"3f",
          6684 => x"08",
          6685 => x"89",
          6686 => x"80",
          6687 => x"cf",
          6688 => x"ff",
          6689 => x"81",
          6690 => x"52",
          6691 => x"51",
          6692 => x"b4",
          6693 => x"11",
          6694 => x"05",
          6695 => x"df",
          6696 => x"f0",
          6697 => x"87",
          6698 => x"26",
          6699 => x"b4",
          6700 => x"11",
          6701 => x"05",
          6702 => x"c3",
          6703 => x"f0",
          6704 => x"81",
          6705 => x"43",
          6706 => x"f6",
          6707 => x"51",
          6708 => x"3f",
          6709 => x"05",
          6710 => x"52",
          6711 => x"29",
          6712 => x"05",
          6713 => x"fb",
          6714 => x"f0",
          6715 => x"38",
          6716 => x"51",
          6717 => x"3f",
          6718 => x"85",
          6719 => x"ff",
          6720 => x"fe",
          6721 => x"81",
          6722 => x"b5",
          6723 => x"05",
          6724 => x"cd",
          6725 => x"53",
          6726 => x"08",
          6727 => x"f2",
          6728 => x"d5",
          6729 => x"ff",
          6730 => x"fe",
          6731 => x"81",
          6732 => x"b5",
          6733 => x"05",
          6734 => x"cd",
          6735 => x"fe",
          6736 => x"3d",
          6737 => x"52",
          6738 => x"b9",
          6739 => x"f0",
          6740 => x"ff",
          6741 => x"59",
          6742 => x"3f",
          6743 => x"58",
          6744 => x"57",
          6745 => x"55",
          6746 => x"08",
          6747 => x"54",
          6748 => x"52",
          6749 => x"ff",
          6750 => x"f0",
          6751 => x"fb",
          6752 => x"fe",
          6753 => x"ef",
          6754 => x"f5",
          6755 => x"ff",
          6756 => x"ff",
          6757 => x"fe",
          6758 => x"81",
          6759 => x"80",
          6760 => x"38",
          6761 => x"fc",
          6762 => x"84",
          6763 => x"ea",
          6764 => x"fe",
          6765 => x"2e",
          6766 => x"b4",
          6767 => x"11",
          6768 => x"05",
          6769 => x"b7",
          6770 => x"f0",
          6771 => x"81",
          6772 => x"42",
          6773 => x"51",
          6774 => x"3f",
          6775 => x"5a",
          6776 => x"81",
          6777 => x"59",
          6778 => x"84",
          6779 => x"7a",
          6780 => x"38",
          6781 => x"b4",
          6782 => x"11",
          6783 => x"05",
          6784 => x"fb",
          6785 => x"f0",
          6786 => x"f9",
          6787 => x"3d",
          6788 => x"53",
          6789 => x"51",
          6790 => x"3f",
          6791 => x"08",
          6792 => x"dd",
          6793 => x"fe",
          6794 => x"ff",
          6795 => x"fe",
          6796 => x"81",
          6797 => x"80",
          6798 => x"38",
          6799 => x"51",
          6800 => x"3f",
          6801 => x"63",
          6802 => x"38",
          6803 => x"70",
          6804 => x"33",
          6805 => x"81",
          6806 => x"39",
          6807 => x"80",
          6808 => x"84",
          6809 => x"e9",
          6810 => x"fe",
          6811 => x"2e",
          6812 => x"b4",
          6813 => x"11",
          6814 => x"05",
          6815 => x"ff",
          6816 => x"f0",
          6817 => x"f8",
          6818 => x"3d",
          6819 => x"53",
          6820 => x"51",
          6821 => x"3f",
          6822 => x"08",
          6823 => x"e1",
          6824 => x"b8",
          6825 => x"fe",
          6826 => x"79",
          6827 => x"38",
          6828 => x"7b",
          6829 => x"5b",
          6830 => x"92",
          6831 => x"7a",
          6832 => x"53",
          6833 => x"f6",
          6834 => x"e6",
          6835 => x"1a",
          6836 => x"43",
          6837 => x"81",
          6838 => x"82",
          6839 => x"3d",
          6840 => x"53",
          6841 => x"51",
          6842 => x"3f",
          6843 => x"08",
          6844 => x"81",
          6845 => x"59",
          6846 => x"89",
          6847 => x"ec",
          6848 => x"cd",
          6849 => x"b5",
          6850 => x"80",
          6851 => x"81",
          6852 => x"44",
          6853 => x"fa",
          6854 => x"78",
          6855 => x"38",
          6856 => x"08",
          6857 => x"81",
          6858 => x"59",
          6859 => x"88",
          6860 => x"84",
          6861 => x"39",
          6862 => x"33",
          6863 => x"2e",
          6864 => x"fa",
          6865 => x"89",
          6866 => x"9c",
          6867 => x"05",
          6868 => x"fe",
          6869 => x"ff",
          6870 => x"fe",
          6871 => x"81",
          6872 => x"80",
          6873 => x"fa",
          6874 => x"78",
          6875 => x"38",
          6876 => x"08",
          6877 => x"39",
          6878 => x"33",
          6879 => x"2e",
          6880 => x"f9",
          6881 => x"bb",
          6882 => x"b6",
          6883 => x"80",
          6884 => x"81",
          6885 => x"43",
          6886 => x"fa",
          6887 => x"78",
          6888 => x"38",
          6889 => x"08",
          6890 => x"81",
          6891 => x"59",
          6892 => x"88",
          6893 => x"90",
          6894 => x"39",
          6895 => x"08",
          6896 => x"b4",
          6897 => x"11",
          6898 => x"05",
          6899 => x"af",
          6900 => x"f0",
          6901 => x"a7",
          6902 => x"5c",
          6903 => x"2e",
          6904 => x"5c",
          6905 => x"70",
          6906 => x"07",
          6907 => x"7f",
          6908 => x"5a",
          6909 => x"2e",
          6910 => x"a0",
          6911 => x"88",
          6912 => x"e4",
          6913 => x"9e",
          6914 => x"63",
          6915 => x"62",
          6916 => x"ee",
          6917 => x"f6",
          6918 => x"de",
          6919 => x"e1",
          6920 => x"ff",
          6921 => x"ff",
          6922 => x"fe",
          6923 => x"81",
          6924 => x"80",
          6925 => x"38",
          6926 => x"fc",
          6927 => x"84",
          6928 => x"e5",
          6929 => x"fe",
          6930 => x"2e",
          6931 => x"59",
          6932 => x"05",
          6933 => x"63",
          6934 => x"b4",
          6935 => x"11",
          6936 => x"05",
          6937 => x"97",
          6938 => x"f0",
          6939 => x"f5",
          6940 => x"70",
          6941 => x"81",
          6942 => x"fe",
          6943 => x"80",
          6944 => x"51",
          6945 => x"3f",
          6946 => x"33",
          6947 => x"2e",
          6948 => x"9f",
          6949 => x"38",
          6950 => x"fc",
          6951 => x"84",
          6952 => x"e4",
          6953 => x"fe",
          6954 => x"2e",
          6955 => x"59",
          6956 => x"05",
          6957 => x"63",
          6958 => x"ff",
          6959 => x"f7",
          6960 => x"dc",
          6961 => x"aa",
          6962 => x"fe",
          6963 => x"ff",
          6964 => x"fe",
          6965 => x"81",
          6966 => x"80",
          6967 => x"38",
          6968 => x"f0",
          6969 => x"84",
          6970 => x"e6",
          6971 => x"fe",
          6972 => x"2e",
          6973 => x"59",
          6974 => x"22",
          6975 => x"05",
          6976 => x"41",
          6977 => x"f0",
          6978 => x"84",
          6979 => x"e5",
          6980 => x"fe",
          6981 => x"38",
          6982 => x"60",
          6983 => x"52",
          6984 => x"51",
          6985 => x"3f",
          6986 => x"79",
          6987 => x"b4",
          6988 => x"79",
          6989 => x"ae",
          6990 => x"38",
          6991 => x"87",
          6992 => x"05",
          6993 => x"b4",
          6994 => x"11",
          6995 => x"05",
          6996 => x"9d",
          6997 => x"f0",
          6998 => x"92",
          6999 => x"02",
          7000 => x"79",
          7001 => x"5b",
          7002 => x"ff",
          7003 => x"f7",
          7004 => x"db",
          7005 => x"a3",
          7006 => x"fe",
          7007 => x"ff",
          7008 => x"fe",
          7009 => x"81",
          7010 => x"80",
          7011 => x"38",
          7012 => x"f0",
          7013 => x"84",
          7014 => x"e4",
          7015 => x"fe",
          7016 => x"2e",
          7017 => x"60",
          7018 => x"60",
          7019 => x"b4",
          7020 => x"11",
          7021 => x"05",
          7022 => x"b5",
          7023 => x"f0",
          7024 => x"f2",
          7025 => x"70",
          7026 => x"81",
          7027 => x"fe",
          7028 => x"80",
          7029 => x"51",
          7030 => x"3f",
          7031 => x"33",
          7032 => x"2e",
          7033 => x"9f",
          7034 => x"38",
          7035 => x"f0",
          7036 => x"84",
          7037 => x"e3",
          7038 => x"fe",
          7039 => x"2e",
          7040 => x"60",
          7041 => x"60",
          7042 => x"ff",
          7043 => x"f7",
          7044 => x"da",
          7045 => x"ae",
          7046 => x"ac",
          7047 => x"86",
          7048 => x"fe",
          7049 => x"f1",
          7050 => x"f7",
          7051 => x"d9",
          7052 => x"51",
          7053 => x"3f",
          7054 => x"81",
          7055 => x"fe",
          7056 => x"84",
          7057 => x"87",
          7058 => x"0c",
          7059 => x"0b",
          7060 => x"94",
          7061 => x"39",
          7062 => x"51",
          7063 => x"3f",
          7064 => x"0b",
          7065 => x"84",
          7066 => x"83",
          7067 => x"94",
          7068 => x"8d",
          7069 => x"ff",
          7070 => x"ff",
          7071 => x"fe",
          7072 => x"81",
          7073 => x"80",
          7074 => x"38",
          7075 => x"f8",
          7076 => x"de",
          7077 => x"59",
          7078 => x"3d",
          7079 => x"53",
          7080 => x"51",
          7081 => x"3f",
          7082 => x"08",
          7083 => x"d1",
          7084 => x"81",
          7085 => x"fe",
          7086 => x"63",
          7087 => x"81",
          7088 => x"80",
          7089 => x"38",
          7090 => x"08",
          7091 => x"bc",
          7092 => x"b6",
          7093 => x"39",
          7094 => x"51",
          7095 => x"3f",
          7096 => x"3f",
          7097 => x"81",
          7098 => x"fe",
          7099 => x"80",
          7100 => x"39",
          7101 => x"3f",
          7102 => x"79",
          7103 => x"59",
          7104 => x"ef",
          7105 => x"7d",
          7106 => x"80",
          7107 => x"38",
          7108 => x"84",
          7109 => x"c1",
          7110 => x"fe",
          7111 => x"81",
          7112 => x"2e",
          7113 => x"82",
          7114 => x"7b",
          7115 => x"38",
          7116 => x"7b",
          7117 => x"38",
          7118 => x"81",
          7119 => x"7a",
          7120 => x"8c",
          7121 => x"81",
          7122 => x"b4",
          7123 => x"05",
          7124 => x"cc",
          7125 => x"81",
          7126 => x"b4",
          7127 => x"05",
          7128 => x"bc",
          7129 => x"7a",
          7130 => x"8c",
          7131 => x"81",
          7132 => x"b4",
          7133 => x"05",
          7134 => x"a4",
          7135 => x"7a",
          7136 => x"81",
          7137 => x"b4",
          7138 => x"05",
          7139 => x"90",
          7140 => x"ec",
          7141 => x"b8",
          7142 => x"64",
          7143 => x"83",
          7144 => x"83",
          7145 => x"b4",
          7146 => x"05",
          7147 => x"3f",
          7148 => x"08",
          7149 => x"08",
          7150 => x"70",
          7151 => x"25",
          7152 => x"5f",
          7153 => x"83",
          7154 => x"81",
          7155 => x"06",
          7156 => x"2e",
          7157 => x"1c",
          7158 => x"06",
          7159 => x"fe",
          7160 => x"81",
          7161 => x"32",
          7162 => x"8a",
          7163 => x"2e",
          7164 => x"ee",
          7165 => x"f9",
          7166 => x"dc",
          7167 => x"81",
          7168 => x"0d",
          7169 => x"ff",
          7170 => x"c0",
          7171 => x"08",
          7172 => x"84",
          7173 => x"51",
          7174 => x"3f",
          7175 => x"08",
          7176 => x"08",
          7177 => x"84",
          7178 => x"51",
          7179 => x"3f",
          7180 => x"f0",
          7181 => x"0c",
          7182 => x"9c",
          7183 => x"55",
          7184 => x"52",
          7185 => x"b2",
          7186 => x"fe",
          7187 => x"2b",
          7188 => x"53",
          7189 => x"52",
          7190 => x"b2",
          7191 => x"81",
          7192 => x"07",
          7193 => x"80",
          7194 => x"c0",
          7195 => x"8c",
          7196 => x"87",
          7197 => x"0c",
          7198 => x"81",
          7199 => x"a6",
          7200 => x"ff",
          7201 => x"c6",
          7202 => x"d0",
          7203 => x"f9",
          7204 => x"d5",
          7205 => x"f9",
          7206 => x"d5",
          7207 => x"c9",
          7208 => x"cf",
          7209 => x"51",
          7210 => x"ec",
          7211 => x"04",
          7212 => x"ff",
          7213 => x"ff",
          7214 => x"00",
          7215 => x"ff",
          7216 => x"18",
          7217 => x"18",
          7218 => x"18",
          7219 => x"18",
          7220 => x"18",
          7221 => x"25",
          7222 => x"26",
          7223 => x"27",
          7224 => x"27",
          7225 => x"27",
          7226 => x"28",
          7227 => x"24",
          7228 => x"24",
          7229 => x"28",
          7230 => x"29",
          7231 => x"29",
          7232 => x"29",
          7233 => x"61",
          7234 => x"61",
          7235 => x"61",
          7236 => x"61",
          7237 => x"61",
          7238 => x"61",
          7239 => x"61",
          7240 => x"61",
          7241 => x"61",
          7242 => x"61",
          7243 => x"61",
          7244 => x"61",
          7245 => x"61",
          7246 => x"61",
          7247 => x"61",
          7248 => x"61",
          7249 => x"61",
          7250 => x"61",
          7251 => x"61",
          7252 => x"61",
          7253 => x"2f",
          7254 => x"25",
          7255 => x"64",
          7256 => x"3a",
          7257 => x"25",
          7258 => x"0a",
          7259 => x"43",
          7260 => x"6e",
          7261 => x"75",
          7262 => x"69",
          7263 => x"00",
          7264 => x"66",
          7265 => x"20",
          7266 => x"20",
          7267 => x"66",
          7268 => x"00",
          7269 => x"44",
          7270 => x"63",
          7271 => x"69",
          7272 => x"65",
          7273 => x"74",
          7274 => x"0a",
          7275 => x"20",
          7276 => x"20",
          7277 => x"41",
          7278 => x"28",
          7279 => x"58",
          7280 => x"38",
          7281 => x"0a",
          7282 => x"20",
          7283 => x"52",
          7284 => x"20",
          7285 => x"28",
          7286 => x"58",
          7287 => x"38",
          7288 => x"0a",
          7289 => x"20",
          7290 => x"53",
          7291 => x"52",
          7292 => x"28",
          7293 => x"58",
          7294 => x"38",
          7295 => x"0a",
          7296 => x"20",
          7297 => x"41",
          7298 => x"20",
          7299 => x"28",
          7300 => x"58",
          7301 => x"38",
          7302 => x"0a",
          7303 => x"20",
          7304 => x"4d",
          7305 => x"20",
          7306 => x"28",
          7307 => x"58",
          7308 => x"38",
          7309 => x"0a",
          7310 => x"20",
          7311 => x"20",
          7312 => x"44",
          7313 => x"28",
          7314 => x"69",
          7315 => x"20",
          7316 => x"32",
          7317 => x"0a",
          7318 => x"20",
          7319 => x"4d",
          7320 => x"20",
          7321 => x"28",
          7322 => x"65",
          7323 => x"20",
          7324 => x"32",
          7325 => x"0a",
          7326 => x"20",
          7327 => x"54",
          7328 => x"54",
          7329 => x"28",
          7330 => x"6e",
          7331 => x"73",
          7332 => x"32",
          7333 => x"0a",
          7334 => x"20",
          7335 => x"53",
          7336 => x"4e",
          7337 => x"55",
          7338 => x"00",
          7339 => x"20",
          7340 => x"20",
          7341 => x"0a",
          7342 => x"20",
          7343 => x"43",
          7344 => x"00",
          7345 => x"20",
          7346 => x"32",
          7347 => x"00",
          7348 => x"20",
          7349 => x"49",
          7350 => x"00",
          7351 => x"64",
          7352 => x"73",
          7353 => x"0a",
          7354 => x"20",
          7355 => x"55",
          7356 => x"73",
          7357 => x"56",
          7358 => x"6f",
          7359 => x"64",
          7360 => x"73",
          7361 => x"20",
          7362 => x"58",
          7363 => x"00",
          7364 => x"20",
          7365 => x"55",
          7366 => x"6d",
          7367 => x"20",
          7368 => x"72",
          7369 => x"64",
          7370 => x"73",
          7371 => x"20",
          7372 => x"58",
          7373 => x"00",
          7374 => x"20",
          7375 => x"61",
          7376 => x"53",
          7377 => x"74",
          7378 => x"64",
          7379 => x"73",
          7380 => x"20",
          7381 => x"20",
          7382 => x"58",
          7383 => x"00",
          7384 => x"73",
          7385 => x"00",
          7386 => x"20",
          7387 => x"55",
          7388 => x"20",
          7389 => x"20",
          7390 => x"20",
          7391 => x"20",
          7392 => x"20",
          7393 => x"20",
          7394 => x"58",
          7395 => x"00",
          7396 => x"20",
          7397 => x"73",
          7398 => x"20",
          7399 => x"63",
          7400 => x"72",
          7401 => x"20",
          7402 => x"20",
          7403 => x"20",
          7404 => x"25",
          7405 => x"4d",
          7406 => x"00",
          7407 => x"20",
          7408 => x"52",
          7409 => x"43",
          7410 => x"6b",
          7411 => x"65",
          7412 => x"20",
          7413 => x"20",
          7414 => x"20",
          7415 => x"25",
          7416 => x"4d",
          7417 => x"00",
          7418 => x"20",
          7419 => x"73",
          7420 => x"6e",
          7421 => x"44",
          7422 => x"20",
          7423 => x"63",
          7424 => x"72",
          7425 => x"20",
          7426 => x"25",
          7427 => x"4d",
          7428 => x"00",
          7429 => x"61",
          7430 => x"00",
          7431 => x"64",
          7432 => x"00",
          7433 => x"65",
          7434 => x"00",
          7435 => x"4f",
          7436 => x"4f",
          7437 => x"00",
          7438 => x"6b",
          7439 => x"6e",
          7440 => x"73",
          7441 => x"79",
          7442 => x"74",
          7443 => x"73",
          7444 => x"79",
          7445 => x"73",
          7446 => x"00",
          7447 => x"00",
          7448 => x"34",
          7449 => x"25",
          7450 => x"00",
          7451 => x"69",
          7452 => x"20",
          7453 => x"72",
          7454 => x"74",
          7455 => x"65",
          7456 => x"73",
          7457 => x"79",
          7458 => x"6c",
          7459 => x"6f",
          7460 => x"46",
          7461 => x"00",
          7462 => x"6e",
          7463 => x"20",
          7464 => x"6e",
          7465 => x"65",
          7466 => x"20",
          7467 => x"74",
          7468 => x"20",
          7469 => x"65",
          7470 => x"69",
          7471 => x"6c",
          7472 => x"2e",
          7473 => x"00",
          7474 => x"75",
          7475 => x"00",
          7476 => x"00",
          7477 => x"75",
          7478 => x"00",
          7479 => x"00",
          7480 => x"75",
          7481 => x"00",
          7482 => x"00",
          7483 => x"75",
          7484 => x"00",
          7485 => x"00",
          7486 => x"75",
          7487 => x"00",
          7488 => x"00",
          7489 => x"75",
          7490 => x"00",
          7491 => x"00",
          7492 => x"75",
          7493 => x"00",
          7494 => x"00",
          7495 => x"75",
          7496 => x"00",
          7497 => x"00",
          7498 => x"75",
          7499 => x"00",
          7500 => x"00",
          7501 => x"75",
          7502 => x"00",
          7503 => x"00",
          7504 => x"75",
          7505 => x"00",
          7506 => x"00",
          7507 => x"44",
          7508 => x"43",
          7509 => x"42",
          7510 => x"41",
          7511 => x"36",
          7512 => x"35",
          7513 => x"34",
          7514 => x"33",
          7515 => x"31",
          7516 => x"00",
          7517 => x"00",
          7518 => x"00",
          7519 => x"2b",
          7520 => x"3c",
          7521 => x"5b",
          7522 => x"00",
          7523 => x"54",
          7524 => x"54",
          7525 => x"00",
          7526 => x"90",
          7527 => x"4f",
          7528 => x"30",
          7529 => x"20",
          7530 => x"45",
          7531 => x"20",
          7532 => x"33",
          7533 => x"20",
          7534 => x"20",
          7535 => x"45",
          7536 => x"20",
          7537 => x"20",
          7538 => x"20",
          7539 => x"75",
          7540 => x"00",
          7541 => x"00",
          7542 => x"00",
          7543 => x"45",
          7544 => x"8f",
          7545 => x"45",
          7546 => x"8e",
          7547 => x"92",
          7548 => x"55",
          7549 => x"9a",
          7550 => x"9e",
          7551 => x"4f",
          7552 => x"a6",
          7553 => x"aa",
          7554 => x"ae",
          7555 => x"b2",
          7556 => x"b6",
          7557 => x"ba",
          7558 => x"be",
          7559 => x"c2",
          7560 => x"c6",
          7561 => x"ca",
          7562 => x"ce",
          7563 => x"d2",
          7564 => x"d6",
          7565 => x"da",
          7566 => x"de",
          7567 => x"e2",
          7568 => x"e6",
          7569 => x"ea",
          7570 => x"ee",
          7571 => x"f2",
          7572 => x"f6",
          7573 => x"fa",
          7574 => x"fe",
          7575 => x"2c",
          7576 => x"5d",
          7577 => x"2a",
          7578 => x"3f",
          7579 => x"00",
          7580 => x"00",
          7581 => x"00",
          7582 => x"02",
          7583 => x"00",
          7584 => x"00",
          7585 => x"00",
          7586 => x"00",
          7587 => x"00",
          7588 => x"6e",
          7589 => x"00",
          7590 => x"6f",
          7591 => x"00",
          7592 => x"6e",
          7593 => x"00",
          7594 => x"6f",
          7595 => x"00",
          7596 => x"78",
          7597 => x"00",
          7598 => x"6c",
          7599 => x"00",
          7600 => x"6f",
          7601 => x"00",
          7602 => x"69",
          7603 => x"00",
          7604 => x"75",
          7605 => x"00",
          7606 => x"62",
          7607 => x"68",
          7608 => x"77",
          7609 => x"64",
          7610 => x"65",
          7611 => x"64",
          7612 => x"65",
          7613 => x"6c",
          7614 => x"00",
          7615 => x"70",
          7616 => x"73",
          7617 => x"74",
          7618 => x"73",
          7619 => x"00",
          7620 => x"66",
          7621 => x"00",
          7622 => x"73",
          7623 => x"00",
          7624 => x"61",
          7625 => x"00",
          7626 => x"61",
          7627 => x"00",
          7628 => x"6c",
          7629 => x"00",
          7630 => x"73",
          7631 => x"72",
          7632 => x"0a",
          7633 => x"74",
          7634 => x"61",
          7635 => x"72",
          7636 => x"2e",
          7637 => x"00",
          7638 => x"73",
          7639 => x"6f",
          7640 => x"65",
          7641 => x"2e",
          7642 => x"00",
          7643 => x"20",
          7644 => x"65",
          7645 => x"75",
          7646 => x"0a",
          7647 => x"20",
          7648 => x"68",
          7649 => x"75",
          7650 => x"0a",
          7651 => x"76",
          7652 => x"64",
          7653 => x"6c",
          7654 => x"6d",
          7655 => x"00",
          7656 => x"63",
          7657 => x"20",
          7658 => x"69",
          7659 => x"0a",
          7660 => x"6c",
          7661 => x"6c",
          7662 => x"64",
          7663 => x"78",
          7664 => x"73",
          7665 => x"00",
          7666 => x"6c",
          7667 => x"61",
          7668 => x"65",
          7669 => x"76",
          7670 => x"64",
          7671 => x"00",
          7672 => x"20",
          7673 => x"77",
          7674 => x"65",
          7675 => x"6f",
          7676 => x"74",
          7677 => x"0a",
          7678 => x"69",
          7679 => x"6e",
          7680 => x"65",
          7681 => x"73",
          7682 => x"76",
          7683 => x"64",
          7684 => x"00",
          7685 => x"73",
          7686 => x"6f",
          7687 => x"6e",
          7688 => x"65",
          7689 => x"00",
          7690 => x"20",
          7691 => x"70",
          7692 => x"62",
          7693 => x"66",
          7694 => x"73",
          7695 => x"65",
          7696 => x"6f",
          7697 => x"20",
          7698 => x"64",
          7699 => x"2e",
          7700 => x"00",
          7701 => x"72",
          7702 => x"20",
          7703 => x"72",
          7704 => x"2e",
          7705 => x"00",
          7706 => x"6d",
          7707 => x"74",
          7708 => x"70",
          7709 => x"74",
          7710 => x"20",
          7711 => x"63",
          7712 => x"65",
          7713 => x"00",
          7714 => x"6c",
          7715 => x"73",
          7716 => x"63",
          7717 => x"2e",
          7718 => x"00",
          7719 => x"73",
          7720 => x"69",
          7721 => x"6e",
          7722 => x"65",
          7723 => x"79",
          7724 => x"00",
          7725 => x"6f",
          7726 => x"6e",
          7727 => x"70",
          7728 => x"66",
          7729 => x"73",
          7730 => x"00",
          7731 => x"72",
          7732 => x"74",
          7733 => x"20",
          7734 => x"6f",
          7735 => x"63",
          7736 => x"00",
          7737 => x"63",
          7738 => x"73",
          7739 => x"00",
          7740 => x"6b",
          7741 => x"6e",
          7742 => x"72",
          7743 => x"0a",
          7744 => x"6c",
          7745 => x"79",
          7746 => x"20",
          7747 => x"61",
          7748 => x"6c",
          7749 => x"79",
          7750 => x"2f",
          7751 => x"2e",
          7752 => x"00",
          7753 => x"61",
          7754 => x"00",
          7755 => x"38",
          7756 => x"00",
          7757 => x"20",
          7758 => x"34",
          7759 => x"00",
          7760 => x"20",
          7761 => x"20",
          7762 => x"00",
          7763 => x"32",
          7764 => x"00",
          7765 => x"00",
          7766 => x"00",
          7767 => x"0a",
          7768 => x"55",
          7769 => x"00",
          7770 => x"2a",
          7771 => x"20",
          7772 => x"00",
          7773 => x"2f",
          7774 => x"32",
          7775 => x"00",
          7776 => x"2e",
          7777 => x"00",
          7778 => x"50",
          7779 => x"72",
          7780 => x"25",
          7781 => x"29",
          7782 => x"20",
          7783 => x"2a",
          7784 => x"00",
          7785 => x"55",
          7786 => x"49",
          7787 => x"72",
          7788 => x"74",
          7789 => x"6e",
          7790 => x"72",
          7791 => x"00",
          7792 => x"6d",
          7793 => x"69",
          7794 => x"72",
          7795 => x"74",
          7796 => x"00",
          7797 => x"32",
          7798 => x"74",
          7799 => x"75",
          7800 => x"00",
          7801 => x"43",
          7802 => x"52",
          7803 => x"6e",
          7804 => x"72",
          7805 => x"0a",
          7806 => x"43",
          7807 => x"57",
          7808 => x"6e",
          7809 => x"72",
          7810 => x"0a",
          7811 => x"52",
          7812 => x"52",
          7813 => x"6e",
          7814 => x"72",
          7815 => x"0a",
          7816 => x"52",
          7817 => x"54",
          7818 => x"6e",
          7819 => x"72",
          7820 => x"0a",
          7821 => x"52",
          7822 => x"52",
          7823 => x"6e",
          7824 => x"72",
          7825 => x"0a",
          7826 => x"52",
          7827 => x"54",
          7828 => x"6e",
          7829 => x"72",
          7830 => x"0a",
          7831 => x"74",
          7832 => x"67",
          7833 => x"20",
          7834 => x"65",
          7835 => x"2e",
          7836 => x"00",
          7837 => x"61",
          7838 => x"6e",
          7839 => x"69",
          7840 => x"2e",
          7841 => x"00",
          7842 => x"74",
          7843 => x"65",
          7844 => x"61",
          7845 => x"00",
          7846 => x"00",
          7847 => x"69",
          7848 => x"20",
          7849 => x"69",
          7850 => x"69",
          7851 => x"73",
          7852 => x"64",
          7853 => x"72",
          7854 => x"2c",
          7855 => x"65",
          7856 => x"20",
          7857 => x"74",
          7858 => x"6e",
          7859 => x"6c",
          7860 => x"00",
          7861 => x"00",
          7862 => x"64",
          7863 => x"73",
          7864 => x"64",
          7865 => x"00",
          7866 => x"69",
          7867 => x"6c",
          7868 => x"64",
          7869 => x"00",
          7870 => x"69",
          7871 => x"20",
          7872 => x"69",
          7873 => x"69",
          7874 => x"73",
          7875 => x"00",
          7876 => x"3d",
          7877 => x"00",
          7878 => x"3a",
          7879 => x"65",
          7880 => x"6e",
          7881 => x"2e",
          7882 => x"00",
          7883 => x"70",
          7884 => x"67",
          7885 => x"00",
          7886 => x"6d",
          7887 => x"69",
          7888 => x"2e",
          7889 => x"00",
          7890 => x"38",
          7891 => x"25",
          7892 => x"29",
          7893 => x"30",
          7894 => x"28",
          7895 => x"78",
          7896 => x"00",
          7897 => x"6d",
          7898 => x"65",
          7899 => x"79",
          7900 => x"00",
          7901 => x"6f",
          7902 => x"65",
          7903 => x"0a",
          7904 => x"38",
          7905 => x"30",
          7906 => x"00",
          7907 => x"3f",
          7908 => x"00",
          7909 => x"38",
          7910 => x"30",
          7911 => x"00",
          7912 => x"38",
          7913 => x"30",
          7914 => x"00",
          7915 => x"73",
          7916 => x"69",
          7917 => x"69",
          7918 => x"72",
          7919 => x"74",
          7920 => x"00",
          7921 => x"61",
          7922 => x"6e",
          7923 => x"6e",
          7924 => x"72",
          7925 => x"73",
          7926 => x"00",
          7927 => x"73",
          7928 => x"65",
          7929 => x"61",
          7930 => x"66",
          7931 => x"0a",
          7932 => x"61",
          7933 => x"6e",
          7934 => x"61",
          7935 => x"66",
          7936 => x"0a",
          7937 => x"65",
          7938 => x"69",
          7939 => x"63",
          7940 => x"20",
          7941 => x"30",
          7942 => x"2e",
          7943 => x"00",
          7944 => x"6c",
          7945 => x"67",
          7946 => x"64",
          7947 => x"20",
          7948 => x"78",
          7949 => x"2e",
          7950 => x"00",
          7951 => x"6c",
          7952 => x"65",
          7953 => x"6e",
          7954 => x"63",
          7955 => x"20",
          7956 => x"29",
          7957 => x"00",
          7958 => x"73",
          7959 => x"74",
          7960 => x"20",
          7961 => x"6c",
          7962 => x"74",
          7963 => x"2e",
          7964 => x"00",
          7965 => x"6c",
          7966 => x"65",
          7967 => x"74",
          7968 => x"2e",
          7969 => x"00",
          7970 => x"55",
          7971 => x"6e",
          7972 => x"3a",
          7973 => x"5c",
          7974 => x"25",
          7975 => x"00",
          7976 => x"3a",
          7977 => x"5c",
          7978 => x"00",
          7979 => x"3a",
          7980 => x"00",
          7981 => x"64",
          7982 => x"6d",
          7983 => x"64",
          7984 => x"00",
          7985 => x"6e",
          7986 => x"67",
          7987 => x"0a",
          7988 => x"61",
          7989 => x"6e",
          7990 => x"6e",
          7991 => x"72",
          7992 => x"73",
          7993 => x"0a",
          7994 => x"00",
          7995 => x"00",
          7996 => x"7f",
          7997 => x"00",
          7998 => x"7f",
          7999 => x"00",
          8000 => x"7f",
          8001 => x"00",
          8002 => x"00",
          8003 => x"00",
          8004 => x"ff",
          8005 => x"00",
          8006 => x"00",
          8007 => x"78",
          8008 => x"00",
          8009 => x"e1",
          8010 => x"e1",
          8011 => x"e1",
          8012 => x"00",
          8013 => x"01",
          8014 => x"01",
          8015 => x"10",
          8016 => x"00",
          8017 => x"00",
          8018 => x"00",
          8019 => x"00",
          8020 => x"7d",
          8021 => x"7d",
          8022 => x"7d",
          8023 => x"7d",
          8024 => x"74",
          8025 => x"00",
          8026 => x"00",
          8027 => x"00",
          8028 => x"00",
          8029 => x"00",
          8030 => x"00",
          8031 => x"00",
          8032 => x"00",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"74",
          8049 => x"00",
          8050 => x"74",
          8051 => x"00",
          8052 => x"74",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"76",
          8057 => x"01",
          8058 => x"00",
          8059 => x"00",
          8060 => x"76",
          8061 => x"01",
          8062 => x"00",
          8063 => x"00",
          8064 => x"76",
          8065 => x"03",
          8066 => x"00",
          8067 => x"00",
          8068 => x"76",
          8069 => x"03",
          8070 => x"00",
          8071 => x"00",
          8072 => x"76",
          8073 => x"03",
          8074 => x"00",
          8075 => x"00",
          8076 => x"76",
          8077 => x"04",
          8078 => x"00",
          8079 => x"00",
          8080 => x"76",
          8081 => x"04",
          8082 => x"00",
          8083 => x"00",
          8084 => x"76",
          8085 => x"04",
          8086 => x"00",
          8087 => x"00",
          8088 => x"76",
          8089 => x"04",
          8090 => x"00",
          8091 => x"00",
          8092 => x"76",
          8093 => x"04",
          8094 => x"00",
          8095 => x"00",
          8096 => x"76",
          8097 => x"04",
          8098 => x"00",
          8099 => x"00",
          8100 => x"76",
          8101 => x"04",
          8102 => x"00",
          8103 => x"00",
          8104 => x"76",
          8105 => x"05",
          8106 => x"00",
          8107 => x"00",
          8108 => x"76",
          8109 => x"05",
          8110 => x"00",
          8111 => x"00",
          8112 => x"76",
          8113 => x"05",
          8114 => x"00",
          8115 => x"00",
          8116 => x"76",
          8117 => x"05",
          8118 => x"00",
          8119 => x"00",
          8120 => x"76",
          8121 => x"07",
          8122 => x"00",
          8123 => x"00",
          8124 => x"76",
          8125 => x"07",
          8126 => x"00",
          8127 => x"00",
          8128 => x"77",
          8129 => x"08",
          8130 => x"00",
          8131 => x"00",
          8132 => x"77",
          8133 => x"08",
          8134 => x"00",
          8135 => x"00",
          8136 => x"77",
          8137 => x"08",
          8138 => x"00",
          8139 => x"00",
          8140 => x"77",
          8141 => x"08",
          8142 => x"00",
          8143 => x"00",
          8144 => x"77",
          8145 => x"09",
          8146 => x"00",
          8147 => x"00",
          8148 => x"77",
          8149 => x"09",
          8150 => x"00",
          8151 => x"00",
          8152 => x"77",
          8153 => x"09",
          8154 => x"00",
          8155 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"d8",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8c",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"81",
           386 => x"a3",
           387 => x"fe",
           388 => x"80",
           389 => x"fe",
           390 => x"c8",
           391 => x"fc",
           392 => x"90",
           393 => x"fc",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"81",
           399 => x"83",
           400 => x"81",
           401 => x"bc",
           402 => x"fe",
           403 => x"80",
           404 => x"fe",
           405 => x"e1",
           406 => x"fc",
           407 => x"90",
           408 => x"fc",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"81",
           414 => x"83",
           415 => x"81",
           416 => x"bf",
           417 => x"fe",
           418 => x"80",
           419 => x"fe",
           420 => x"89",
           421 => x"fc",
           422 => x"90",
           423 => x"fc",
           424 => x"2d",
           425 => x"08",
           426 => x"04",
           427 => x"0c",
           428 => x"81",
           429 => x"83",
           430 => x"81",
           431 => x"bc",
           432 => x"fe",
           433 => x"80",
           434 => x"fe",
           435 => x"8c",
           436 => x"fc",
           437 => x"90",
           438 => x"fc",
           439 => x"2d",
           440 => x"08",
           441 => x"04",
           442 => x"0c",
           443 => x"81",
           444 => x"83",
           445 => x"81",
           446 => x"a0",
           447 => x"fe",
           448 => x"80",
           449 => x"fe",
           450 => x"e1",
           451 => x"fc",
           452 => x"90",
           453 => x"fc",
           454 => x"c3",
           455 => x"fc",
           456 => x"90",
           457 => x"fc",
           458 => x"b4",
           459 => x"fc",
           460 => x"90",
           461 => x"fc",
           462 => x"a8",
           463 => x"fc",
           464 => x"90",
           465 => x"fc",
           466 => x"a5",
           467 => x"fc",
           468 => x"90",
           469 => x"fc",
           470 => x"c3",
           471 => x"fc",
           472 => x"90",
           473 => x"fc",
           474 => x"a3",
           475 => x"fc",
           476 => x"90",
           477 => x"fc",
           478 => x"96",
           479 => x"fc",
           480 => x"90",
           481 => x"fc",
           482 => x"e2",
           483 => x"fc",
           484 => x"90",
           485 => x"fc",
           486 => x"81",
           487 => x"fc",
           488 => x"90",
           489 => x"fc",
           490 => x"a0",
           491 => x"fc",
           492 => x"90",
           493 => x"fc",
           494 => x"8a",
           495 => x"fc",
           496 => x"90",
           497 => x"fc",
           498 => x"f0",
           499 => x"fc",
           500 => x"90",
           501 => x"fc",
           502 => x"de",
           503 => x"fc",
           504 => x"90",
           505 => x"fc",
           506 => x"a4",
           507 => x"fc",
           508 => x"90",
           509 => x"fc",
           510 => x"de",
           511 => x"fc",
           512 => x"90",
           513 => x"fc",
           514 => x"df",
           515 => x"fc",
           516 => x"90",
           517 => x"fc",
           518 => x"94",
           519 => x"fc",
           520 => x"90",
           521 => x"fc",
           522 => x"ed",
           523 => x"fc",
           524 => x"90",
           525 => x"fc",
           526 => x"98",
           527 => x"fc",
           528 => x"90",
           529 => x"fc",
           530 => x"fb",
           531 => x"fc",
           532 => x"90",
           533 => x"fc",
           534 => x"d0",
           535 => x"fc",
           536 => x"90",
           537 => x"fc",
           538 => x"da",
           539 => x"fc",
           540 => x"90",
           541 => x"fc",
           542 => x"9c",
           543 => x"fc",
           544 => x"90",
           545 => x"fc",
           546 => x"e2",
           547 => x"fc",
           548 => x"90",
           549 => x"fc",
           550 => x"88",
           551 => x"fc",
           552 => x"90",
           553 => x"fc",
           554 => x"bd",
           555 => x"fc",
           556 => x"90",
           557 => x"fc",
           558 => x"a9",
           559 => x"fc",
           560 => x"90",
           561 => x"fc",
           562 => x"9d",
           563 => x"fc",
           564 => x"90",
           565 => x"fc",
           566 => x"87",
           567 => x"fc",
           568 => x"90",
           569 => x"fc",
           570 => x"eb",
           571 => x"fc",
           572 => x"90",
           573 => x"fc",
           574 => x"2d",
           575 => x"08",
           576 => x"04",
           577 => x"0c",
           578 => x"81",
           579 => x"83",
           580 => x"81",
           581 => x"a2",
           582 => x"fe",
           583 => x"80",
           584 => x"fe",
           585 => x"c2",
           586 => x"fe",
           587 => x"80",
           588 => x"04",
           589 => x"10",
           590 => x"10",
           591 => x"10",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"04",
           598 => x"81",
           599 => x"83",
           600 => x"05",
           601 => x"10",
           602 => x"72",
           603 => x"51",
           604 => x"72",
           605 => x"06",
           606 => x"72",
           607 => x"10",
           608 => x"10",
           609 => x"ed",
           610 => x"53",
           611 => x"fe",
           612 => x"96",
           613 => x"38",
           614 => x"84",
           615 => x"0b",
           616 => x"8f",
           617 => x"51",
           618 => x"04",
           619 => x"fc",
           620 => x"fe",
           621 => x"3d",
           622 => x"81",
           623 => x"8c",
           624 => x"81",
           625 => x"88",
           626 => x"83",
           627 => x"fe",
           628 => x"81",
           629 => x"54",
           630 => x"81",
           631 => x"04",
           632 => x"08",
           633 => x"fc",
           634 => x"0d",
           635 => x"fe",
           636 => x"05",
           637 => x"fe",
           638 => x"05",
           639 => x"a1",
           640 => x"f0",
           641 => x"fe",
           642 => x"85",
           643 => x"fe",
           644 => x"81",
           645 => x"02",
           646 => x"0c",
           647 => x"80",
           648 => x"fc",
           649 => x"0c",
           650 => x"08",
           651 => x"80",
           652 => x"81",
           653 => x"88",
           654 => x"81",
           655 => x"88",
           656 => x"0b",
           657 => x"08",
           658 => x"81",
           659 => x"fc",
           660 => x"38",
           661 => x"fe",
           662 => x"05",
           663 => x"fc",
           664 => x"08",
           665 => x"08",
           666 => x"81",
           667 => x"8c",
           668 => x"25",
           669 => x"fe",
           670 => x"05",
           671 => x"fe",
           672 => x"05",
           673 => x"81",
           674 => x"f0",
           675 => x"fe",
           676 => x"05",
           677 => x"81",
           678 => x"fc",
           679 => x"0c",
           680 => x"08",
           681 => x"81",
           682 => x"fc",
           683 => x"53",
           684 => x"08",
           685 => x"52",
           686 => x"08",
           687 => x"51",
           688 => x"81",
           689 => x"70",
           690 => x"08",
           691 => x"54",
           692 => x"08",
           693 => x"80",
           694 => x"81",
           695 => x"f8",
           696 => x"81",
           697 => x"f8",
           698 => x"fe",
           699 => x"05",
           700 => x"fe",
           701 => x"89",
           702 => x"fe",
           703 => x"81",
           704 => x"02",
           705 => x"0c",
           706 => x"80",
           707 => x"fc",
           708 => x"0c",
           709 => x"08",
           710 => x"80",
           711 => x"81",
           712 => x"88",
           713 => x"81",
           714 => x"88",
           715 => x"0b",
           716 => x"08",
           717 => x"81",
           718 => x"8c",
           719 => x"25",
           720 => x"fe",
           721 => x"05",
           722 => x"fe",
           723 => x"05",
           724 => x"81",
           725 => x"8c",
           726 => x"81",
           727 => x"88",
           728 => x"bd",
           729 => x"f0",
           730 => x"fe",
           731 => x"05",
           732 => x"fe",
           733 => x"05",
           734 => x"90",
           735 => x"fc",
           736 => x"08",
           737 => x"fc",
           738 => x"0c",
           739 => x"08",
           740 => x"70",
           741 => x"0c",
           742 => x"0d",
           743 => x"0c",
           744 => x"fc",
           745 => x"fe",
           746 => x"3d",
           747 => x"81",
           748 => x"fc",
           749 => x"0b",
           750 => x"08",
           751 => x"81",
           752 => x"8c",
           753 => x"fe",
           754 => x"05",
           755 => x"38",
           756 => x"08",
           757 => x"80",
           758 => x"80",
           759 => x"fc",
           760 => x"08",
           761 => x"81",
           762 => x"8c",
           763 => x"81",
           764 => x"8c",
           765 => x"fe",
           766 => x"05",
           767 => x"fe",
           768 => x"05",
           769 => x"39",
           770 => x"08",
           771 => x"80",
           772 => x"38",
           773 => x"08",
           774 => x"81",
           775 => x"88",
           776 => x"ad",
           777 => x"fc",
           778 => x"08",
           779 => x"08",
           780 => x"31",
           781 => x"08",
           782 => x"81",
           783 => x"f8",
           784 => x"fe",
           785 => x"05",
           786 => x"fe",
           787 => x"05",
           788 => x"fc",
           789 => x"08",
           790 => x"fe",
           791 => x"05",
           792 => x"fc",
           793 => x"08",
           794 => x"fe",
           795 => x"05",
           796 => x"39",
           797 => x"08",
           798 => x"80",
           799 => x"81",
           800 => x"88",
           801 => x"81",
           802 => x"f4",
           803 => x"91",
           804 => x"fc",
           805 => x"08",
           806 => x"fc",
           807 => x"0c",
           808 => x"fc",
           809 => x"08",
           810 => x"0c",
           811 => x"81",
           812 => x"04",
           813 => x"76",
           814 => x"55",
           815 => x"8f",
           816 => x"38",
           817 => x"83",
           818 => x"80",
           819 => x"ff",
           820 => x"ff",
           821 => x"72",
           822 => x"54",
           823 => x"81",
           824 => x"ff",
           825 => x"ff",
           826 => x"06",
           827 => x"81",
           828 => x"86",
           829 => x"74",
           830 => x"84",
           831 => x"71",
           832 => x"53",
           833 => x"84",
           834 => x"71",
           835 => x"53",
           836 => x"84",
           837 => x"71",
           838 => x"53",
           839 => x"84",
           840 => x"71",
           841 => x"53",
           842 => x"52",
           843 => x"c9",
           844 => x"27",
           845 => x"70",
           846 => x"08",
           847 => x"05",
           848 => x"12",
           849 => x"26",
           850 => x"54",
           851 => x"fc",
           852 => x"79",
           853 => x"05",
           854 => x"57",
           855 => x"83",
           856 => x"38",
           857 => x"51",
           858 => x"a4",
           859 => x"52",
           860 => x"93",
           861 => x"70",
           862 => x"34",
           863 => x"71",
           864 => x"81",
           865 => x"74",
           866 => x"0c",
           867 => x"04",
           868 => x"2b",
           869 => x"71",
           870 => x"51",
           871 => x"72",
           872 => x"72",
           873 => x"05",
           874 => x"71",
           875 => x"53",
           876 => x"70",
           877 => x"0c",
           878 => x"84",
           879 => x"f0",
           880 => x"8f",
           881 => x"83",
           882 => x"38",
           883 => x"84",
           884 => x"fc",
           885 => x"83",
           886 => x"70",
           887 => x"39",
           888 => x"76",
           889 => x"73",
           890 => x"54",
           891 => x"70",
           892 => x"71",
           893 => x"09",
           894 => x"fd",
           895 => x"70",
           896 => x"81",
           897 => x"51",
           898 => x"70",
           899 => x"14",
           900 => x"84",
           901 => x"70",
           902 => x"70",
           903 => x"ff",
           904 => x"f8",
           905 => x"80",
           906 => x"53",
           907 => x"80",
           908 => x"73",
           909 => x"81",
           910 => x"51",
           911 => x"81",
           912 => x"70",
           913 => x"81",
           914 => x"86",
           915 => x"fd",
           916 => x"70",
           917 => x"53",
           918 => x"b8",
           919 => x"08",
           920 => x"fb",
           921 => x"06",
           922 => x"82",
           923 => x"51",
           924 => x"70",
           925 => x"13",
           926 => x"09",
           927 => x"ff",
           928 => x"f8",
           929 => x"80",
           930 => x"52",
           931 => x"2e",
           932 => x"52",
           933 => x"70",
           934 => x"38",
           935 => x"33",
           936 => x"f8",
           937 => x"31",
           938 => x"0c",
           939 => x"04",
           940 => x"78",
           941 => x"54",
           942 => x"72",
           943 => x"d9",
           944 => x"07",
           945 => x"70",
           946 => x"d6",
           947 => x"53",
           948 => x"b1",
           949 => x"74",
           950 => x"74",
           951 => x"81",
           952 => x"72",
           953 => x"89",
           954 => x"ff",
           955 => x"80",
           956 => x"38",
           957 => x"15",
           958 => x"55",
           959 => x"2e",
           960 => x"d1",
           961 => x"74",
           962 => x"70",
           963 => x"75",
           964 => x"71",
           965 => x"52",
           966 => x"fe",
           967 => x"3d",
           968 => x"74",
           969 => x"73",
           970 => x"71",
           971 => x"2e",
           972 => x"76",
           973 => x"95",
           974 => x"53",
           975 => x"b1",
           976 => x"70",
           977 => x"fd",
           978 => x"70",
           979 => x"81",
           980 => x"51",
           981 => x"38",
           982 => x"17",
           983 => x"73",
           984 => x"74",
           985 => x"2e",
           986 => x"76",
           987 => x"dd",
           988 => x"81",
           989 => x"88",
           990 => x"fe",
           991 => x"52",
           992 => x"88",
           993 => x"86",
           994 => x"f0",
           995 => x"06",
           996 => x"14",
           997 => x"80",
           998 => x"71",
           999 => x"0c",
          1000 => x"04",
          1001 => x"77",
          1002 => x"53",
          1003 => x"80",
          1004 => x"38",
          1005 => x"70",
          1006 => x"81",
          1007 => x"81",
          1008 => x"39",
          1009 => x"39",
          1010 => x"80",
          1011 => x"81",
          1012 => x"55",
          1013 => x"2e",
          1014 => x"55",
          1015 => x"84",
          1016 => x"38",
          1017 => x"06",
          1018 => x"2e",
          1019 => x"88",
          1020 => x"70",
          1021 => x"34",
          1022 => x"71",
          1023 => x"fe",
          1024 => x"3d",
          1025 => x"3d",
          1026 => x"72",
          1027 => x"91",
          1028 => x"fc",
          1029 => x"51",
          1030 => x"81",
          1031 => x"85",
          1032 => x"83",
          1033 => x"72",
          1034 => x"0c",
          1035 => x"04",
          1036 => x"76",
          1037 => x"ff",
          1038 => x"81",
          1039 => x"26",
          1040 => x"83",
          1041 => x"05",
          1042 => x"70",
          1043 => x"8a",
          1044 => x"33",
          1045 => x"70",
          1046 => x"fe",
          1047 => x"33",
          1048 => x"70",
          1049 => x"f2",
          1050 => x"33",
          1051 => x"70",
          1052 => x"e6",
          1053 => x"22",
          1054 => x"74",
          1055 => x"80",
          1056 => x"13",
          1057 => x"52",
          1058 => x"26",
          1059 => x"81",
          1060 => x"98",
          1061 => x"22",
          1062 => x"bc",
          1063 => x"33",
          1064 => x"b8",
          1065 => x"33",
          1066 => x"b4",
          1067 => x"33",
          1068 => x"b0",
          1069 => x"33",
          1070 => x"ac",
          1071 => x"33",
          1072 => x"a8",
          1073 => x"c0",
          1074 => x"73",
          1075 => x"a0",
          1076 => x"87",
          1077 => x"0c",
          1078 => x"81",
          1079 => x"86",
          1080 => x"f3",
          1081 => x"5b",
          1082 => x"9c",
          1083 => x"0c",
          1084 => x"bc",
          1085 => x"7b",
          1086 => x"98",
          1087 => x"79",
          1088 => x"87",
          1089 => x"08",
          1090 => x"1c",
          1091 => x"98",
          1092 => x"79",
          1093 => x"87",
          1094 => x"08",
          1095 => x"1c",
          1096 => x"98",
          1097 => x"79",
          1098 => x"87",
          1099 => x"08",
          1100 => x"1c",
          1101 => x"98",
          1102 => x"79",
          1103 => x"80",
          1104 => x"83",
          1105 => x"59",
          1106 => x"ff",
          1107 => x"1b",
          1108 => x"1b",
          1109 => x"1b",
          1110 => x"1b",
          1111 => x"1b",
          1112 => x"83",
          1113 => x"52",
          1114 => x"51",
          1115 => x"8f",
          1116 => x"ff",
          1117 => x"8f",
          1118 => x"30",
          1119 => x"51",
          1120 => x"0b",
          1121 => x"e8",
          1122 => x"0d",
          1123 => x"0d",
          1124 => x"81",
          1125 => x"70",
          1126 => x"57",
          1127 => x"c0",
          1128 => x"74",
          1129 => x"38",
          1130 => x"94",
          1131 => x"70",
          1132 => x"81",
          1133 => x"52",
          1134 => x"8c",
          1135 => x"2a",
          1136 => x"51",
          1137 => x"38",
          1138 => x"70",
          1139 => x"51",
          1140 => x"8d",
          1141 => x"2a",
          1142 => x"51",
          1143 => x"be",
          1144 => x"ff",
          1145 => x"c0",
          1146 => x"70",
          1147 => x"38",
          1148 => x"90",
          1149 => x"0c",
          1150 => x"f0",
          1151 => x"0d",
          1152 => x"0d",
          1153 => x"33",
          1154 => x"f9",
          1155 => x"81",
          1156 => x"55",
          1157 => x"94",
          1158 => x"80",
          1159 => x"87",
          1160 => x"51",
          1161 => x"96",
          1162 => x"06",
          1163 => x"70",
          1164 => x"38",
          1165 => x"70",
          1166 => x"51",
          1167 => x"72",
          1168 => x"81",
          1169 => x"70",
          1170 => x"38",
          1171 => x"70",
          1172 => x"51",
          1173 => x"38",
          1174 => x"06",
          1175 => x"94",
          1176 => x"80",
          1177 => x"87",
          1178 => x"52",
          1179 => x"87",
          1180 => x"f9",
          1181 => x"54",
          1182 => x"70",
          1183 => x"53",
          1184 => x"77",
          1185 => x"38",
          1186 => x"06",
          1187 => x"0b",
          1188 => x"33",
          1189 => x"06",
          1190 => x"58",
          1191 => x"84",
          1192 => x"2e",
          1193 => x"c0",
          1194 => x"70",
          1195 => x"2a",
          1196 => x"53",
          1197 => x"80",
          1198 => x"71",
          1199 => x"81",
          1200 => x"70",
          1201 => x"81",
          1202 => x"06",
          1203 => x"80",
          1204 => x"71",
          1205 => x"81",
          1206 => x"70",
          1207 => x"74",
          1208 => x"51",
          1209 => x"80",
          1210 => x"2e",
          1211 => x"c0",
          1212 => x"77",
          1213 => x"17",
          1214 => x"81",
          1215 => x"53",
          1216 => x"84",
          1217 => x"fe",
          1218 => x"3d",
          1219 => x"3d",
          1220 => x"81",
          1221 => x"70",
          1222 => x"54",
          1223 => x"94",
          1224 => x"80",
          1225 => x"87",
          1226 => x"51",
          1227 => x"82",
          1228 => x"06",
          1229 => x"70",
          1230 => x"38",
          1231 => x"06",
          1232 => x"94",
          1233 => x"80",
          1234 => x"87",
          1235 => x"52",
          1236 => x"81",
          1237 => x"fe",
          1238 => x"84",
          1239 => x"fe",
          1240 => x"0b",
          1241 => x"33",
          1242 => x"06",
          1243 => x"c0",
          1244 => x"70",
          1245 => x"38",
          1246 => x"94",
          1247 => x"70",
          1248 => x"81",
          1249 => x"51",
          1250 => x"80",
          1251 => x"72",
          1252 => x"51",
          1253 => x"80",
          1254 => x"2e",
          1255 => x"c0",
          1256 => x"71",
          1257 => x"2b",
          1258 => x"51",
          1259 => x"81",
          1260 => x"84",
          1261 => x"ff",
          1262 => x"c0",
          1263 => x"70",
          1264 => x"06",
          1265 => x"80",
          1266 => x"38",
          1267 => x"a4",
          1268 => x"ec",
          1269 => x"9e",
          1270 => x"f9",
          1271 => x"c0",
          1272 => x"81",
          1273 => x"87",
          1274 => x"08",
          1275 => x"0c",
          1276 => x"9c",
          1277 => x"fc",
          1278 => x"9e",
          1279 => x"fa",
          1280 => x"c0",
          1281 => x"81",
          1282 => x"87",
          1283 => x"08",
          1284 => x"0c",
          1285 => x"b4",
          1286 => x"8c",
          1287 => x"9e",
          1288 => x"fa",
          1289 => x"c0",
          1290 => x"81",
          1291 => x"87",
          1292 => x"08",
          1293 => x"0c",
          1294 => x"c4",
          1295 => x"9c",
          1296 => x"9e",
          1297 => x"70",
          1298 => x"23",
          1299 => x"84",
          1300 => x"a4",
          1301 => x"9e",
          1302 => x"fa",
          1303 => x"c0",
          1304 => x"81",
          1305 => x"81",
          1306 => x"b0",
          1307 => x"87",
          1308 => x"08",
          1309 => x"0a",
          1310 => x"52",
          1311 => x"83",
          1312 => x"71",
          1313 => x"34",
          1314 => x"c0",
          1315 => x"70",
          1316 => x"06",
          1317 => x"70",
          1318 => x"38",
          1319 => x"81",
          1320 => x"80",
          1321 => x"9e",
          1322 => x"90",
          1323 => x"51",
          1324 => x"80",
          1325 => x"81",
          1326 => x"fa",
          1327 => x"0b",
          1328 => x"90",
          1329 => x"80",
          1330 => x"52",
          1331 => x"2e",
          1332 => x"52",
          1333 => x"b4",
          1334 => x"87",
          1335 => x"08",
          1336 => x"80",
          1337 => x"52",
          1338 => x"83",
          1339 => x"71",
          1340 => x"34",
          1341 => x"c0",
          1342 => x"70",
          1343 => x"06",
          1344 => x"70",
          1345 => x"38",
          1346 => x"81",
          1347 => x"80",
          1348 => x"9e",
          1349 => x"84",
          1350 => x"51",
          1351 => x"80",
          1352 => x"81",
          1353 => x"fa",
          1354 => x"0b",
          1355 => x"90",
          1356 => x"80",
          1357 => x"52",
          1358 => x"2e",
          1359 => x"52",
          1360 => x"b8",
          1361 => x"87",
          1362 => x"08",
          1363 => x"80",
          1364 => x"52",
          1365 => x"83",
          1366 => x"71",
          1367 => x"34",
          1368 => x"c0",
          1369 => x"70",
          1370 => x"06",
          1371 => x"70",
          1372 => x"38",
          1373 => x"81",
          1374 => x"80",
          1375 => x"9e",
          1376 => x"a0",
          1377 => x"52",
          1378 => x"2e",
          1379 => x"52",
          1380 => x"bb",
          1381 => x"9e",
          1382 => x"98",
          1383 => x"8a",
          1384 => x"51",
          1385 => x"bc",
          1386 => x"87",
          1387 => x"08",
          1388 => x"06",
          1389 => x"70",
          1390 => x"38",
          1391 => x"81",
          1392 => x"87",
          1393 => x"08",
          1394 => x"06",
          1395 => x"51",
          1396 => x"81",
          1397 => x"80",
          1398 => x"9e",
          1399 => x"88",
          1400 => x"52",
          1401 => x"83",
          1402 => x"71",
          1403 => x"34",
          1404 => x"90",
          1405 => x"06",
          1406 => x"81",
          1407 => x"83",
          1408 => x"fb",
          1409 => x"e2",
          1410 => x"9b",
          1411 => x"b0",
          1412 => x"80",
          1413 => x"81",
          1414 => x"8a",
          1415 => x"e3",
          1416 => x"83",
          1417 => x"b2",
          1418 => x"80",
          1419 => x"81",
          1420 => x"81",
          1421 => x"11",
          1422 => x"e3",
          1423 => x"cb",
          1424 => x"b7",
          1425 => x"80",
          1426 => x"81",
          1427 => x"81",
          1428 => x"11",
          1429 => x"e3",
          1430 => x"af",
          1431 => x"b4",
          1432 => x"80",
          1433 => x"81",
          1434 => x"81",
          1435 => x"11",
          1436 => x"e3",
          1437 => x"93",
          1438 => x"b5",
          1439 => x"80",
          1440 => x"81",
          1441 => x"81",
          1442 => x"11",
          1443 => x"e4",
          1444 => x"f7",
          1445 => x"b6",
          1446 => x"80",
          1447 => x"81",
          1448 => x"81",
          1449 => x"11",
          1450 => x"e4",
          1451 => x"db",
          1452 => x"bb",
          1453 => x"80",
          1454 => x"81",
          1455 => x"52",
          1456 => x"51",
          1457 => x"81",
          1458 => x"54",
          1459 => x"8d",
          1460 => x"c0",
          1461 => x"e4",
          1462 => x"af",
          1463 => x"bd",
          1464 => x"80",
          1465 => x"81",
          1466 => x"52",
          1467 => x"51",
          1468 => x"81",
          1469 => x"54",
          1470 => x"88",
          1471 => x"98",
          1472 => x"3f",
          1473 => x"33",
          1474 => x"2e",
          1475 => x"e5",
          1476 => x"93",
          1477 => x"b8",
          1478 => x"80",
          1479 => x"81",
          1480 => x"88",
          1481 => x"fa",
          1482 => x"73",
          1483 => x"38",
          1484 => x"51",
          1485 => x"81",
          1486 => x"54",
          1487 => x"88",
          1488 => x"d0",
          1489 => x"3f",
          1490 => x"51",
          1491 => x"81",
          1492 => x"52",
          1493 => x"51",
          1494 => x"81",
          1495 => x"52",
          1496 => x"51",
          1497 => x"81",
          1498 => x"52",
          1499 => x"51",
          1500 => x"81",
          1501 => x"87",
          1502 => x"fa",
          1503 => x"81",
          1504 => x"8d",
          1505 => x"fa",
          1506 => x"bd",
          1507 => x"75",
          1508 => x"3f",
          1509 => x"08",
          1510 => x"29",
          1511 => x"54",
          1512 => x"f0",
          1513 => x"e7",
          1514 => x"df",
          1515 => x"b7",
          1516 => x"80",
          1517 => x"81",
          1518 => x"56",
          1519 => x"52",
          1520 => x"e9",
          1521 => x"f0",
          1522 => x"c0",
          1523 => x"31",
          1524 => x"fe",
          1525 => x"81",
          1526 => x"8c",
          1527 => x"fa",
          1528 => x"73",
          1529 => x"38",
          1530 => x"08",
          1531 => x"c0",
          1532 => x"e3",
          1533 => x"fe",
          1534 => x"84",
          1535 => x"71",
          1536 => x"81",
          1537 => x"52",
          1538 => x"51",
          1539 => x"81",
          1540 => x"86",
          1541 => x"3d",
          1542 => x"3d",
          1543 => x"05",
          1544 => x"52",
          1545 => x"aa",
          1546 => x"29",
          1547 => x"05",
          1548 => x"04",
          1549 => x"51",
          1550 => x"e8",
          1551 => x"39",
          1552 => x"51",
          1553 => x"e8",
          1554 => x"39",
          1555 => x"51",
          1556 => x"e8",
          1557 => x"cf",
          1558 => x"0d",
          1559 => x"80",
          1560 => x"3d",
          1561 => x"96",
          1562 => x"52",
          1563 => x"0c",
          1564 => x"70",
          1565 => x"0c",
          1566 => x"3d",
          1567 => x"3d",
          1568 => x"96",
          1569 => x"81",
          1570 => x"52",
          1571 => x"73",
          1572 => x"fa",
          1573 => x"70",
          1574 => x"0c",
          1575 => x"83",
          1576 => x"80",
          1577 => x"96",
          1578 => x"81",
          1579 => x"87",
          1580 => x"0c",
          1581 => x"0d",
          1582 => x"08",
          1583 => x"96",
          1584 => x"ff",
          1585 => x"ff",
          1586 => x"11",
          1587 => x"53",
          1588 => x"f8",
          1589 => x"70",
          1590 => x"0c",
          1591 => x"81",
          1592 => x"84",
          1593 => x"f9",
          1594 => x"7b",
          1595 => x"a0",
          1596 => x"08",
          1597 => x"90",
          1598 => x"58",
          1599 => x"53",
          1600 => x"ba",
          1601 => x"88",
          1602 => x"51",
          1603 => x"76",
          1604 => x"12",
          1605 => x"0c",
          1606 => x"0c",
          1607 => x"0c",
          1608 => x"0c",
          1609 => x"0c",
          1610 => x"0c",
          1611 => x"0c",
          1612 => x"0c",
          1613 => x"0c",
          1614 => x"0c",
          1615 => x"73",
          1616 => x"16",
          1617 => x"15",
          1618 => x"fe",
          1619 => x"3d",
          1620 => x"3d",
          1621 => x"11",
          1622 => x"08",
          1623 => x"71",
          1624 => x"09",
          1625 => x"38",
          1626 => x"70",
          1627 => x"70",
          1628 => x"81",
          1629 => x"84",
          1630 => x"84",
          1631 => x"88",
          1632 => x"8c",
          1633 => x"53",
          1634 => x"73",
          1635 => x"d8",
          1636 => x"0c",
          1637 => x"0b",
          1638 => x"72",
          1639 => x"0c",
          1640 => x"73",
          1641 => x"51",
          1642 => x"2e",
          1643 => x"b3",
          1644 => x"08",
          1645 => x"52",
          1646 => x"09",
          1647 => x"38",
          1648 => x"12",
          1649 => x"94",
          1650 => x"15",
          1651 => x"13",
          1652 => x"12",
          1653 => x"08",
          1654 => x"70",
          1655 => x"52",
          1656 => x"72",
          1657 => x"0c",
          1658 => x"04",
          1659 => x"79",
          1660 => x"76",
          1661 => x"b5",
          1662 => x"f0",
          1663 => x"d8",
          1664 => x"75",
          1665 => x"8f",
          1666 => x"08",
          1667 => x"c7",
          1668 => x"08",
          1669 => x"83",
          1670 => x"fc",
          1671 => x"70",
          1672 => x"91",
          1673 => x"f0",
          1674 => x"f0",
          1675 => x"81",
          1676 => x"07",
          1677 => x"fe",
          1678 => x"70",
          1679 => x"07",
          1680 => x"07",
          1681 => x"51",
          1682 => x"54",
          1683 => x"09",
          1684 => x"d9",
          1685 => x"76",
          1686 => x"80",
          1687 => x"0b",
          1688 => x"08",
          1689 => x"fe",
          1690 => x"05",
          1691 => x"d4",
          1692 => x"08",
          1693 => x"38",
          1694 => x"87",
          1695 => x"08",
          1696 => x"88",
          1697 => x"17",
          1698 => x"17",
          1699 => x"14",
          1700 => x"08",
          1701 => x"0c",
          1702 => x"fd",
          1703 => x"52",
          1704 => x"08",
          1705 => x"3f",
          1706 => x"08",
          1707 => x"fe",
          1708 => x"3d",
          1709 => x"3d",
          1710 => x"71",
          1711 => x"38",
          1712 => x"fd",
          1713 => x"3d",
          1714 => x"3d",
          1715 => x"05",
          1716 => x"8a",
          1717 => x"06",
          1718 => x"51",
          1719 => x"ff",
          1720 => x"71",
          1721 => x"38",
          1722 => x"81",
          1723 => x"81",
          1724 => x"8c",
          1725 => x"81",
          1726 => x"52",
          1727 => x"85",
          1728 => x"71",
          1729 => x"0d",
          1730 => x"0d",
          1731 => x"33",
          1732 => x"08",
          1733 => x"84",
          1734 => x"ff",
          1735 => x"81",
          1736 => x"84",
          1737 => x"fd",
          1738 => x"54",
          1739 => x"81",
          1740 => x"53",
          1741 => x"8e",
          1742 => x"ff",
          1743 => x"14",
          1744 => x"3f",
          1745 => x"3d",
          1746 => x"3d",
          1747 => x"ff",
          1748 => x"81",
          1749 => x"56",
          1750 => x"70",
          1751 => x"53",
          1752 => x"2e",
          1753 => x"81",
          1754 => x"81",
          1755 => x"da",
          1756 => x"74",
          1757 => x"0c",
          1758 => x"04",
          1759 => x"66",
          1760 => x"78",
          1761 => x"5a",
          1762 => x"80",
          1763 => x"38",
          1764 => x"09",
          1765 => x"de",
          1766 => x"7a",
          1767 => x"5c",
          1768 => x"5b",
          1769 => x"09",
          1770 => x"38",
          1771 => x"39",
          1772 => x"09",
          1773 => x"38",
          1774 => x"70",
          1775 => x"33",
          1776 => x"2e",
          1777 => x"92",
          1778 => x"19",
          1779 => x"70",
          1780 => x"33",
          1781 => x"53",
          1782 => x"16",
          1783 => x"26",
          1784 => x"88",
          1785 => x"05",
          1786 => x"05",
          1787 => x"05",
          1788 => x"5b",
          1789 => x"80",
          1790 => x"30",
          1791 => x"80",
          1792 => x"cc",
          1793 => x"70",
          1794 => x"25",
          1795 => x"54",
          1796 => x"53",
          1797 => x"8c",
          1798 => x"07",
          1799 => x"05",
          1800 => x"5a",
          1801 => x"83",
          1802 => x"54",
          1803 => x"27",
          1804 => x"16",
          1805 => x"06",
          1806 => x"80",
          1807 => x"aa",
          1808 => x"cf",
          1809 => x"73",
          1810 => x"81",
          1811 => x"80",
          1812 => x"38",
          1813 => x"2e",
          1814 => x"81",
          1815 => x"80",
          1816 => x"8a",
          1817 => x"39",
          1818 => x"2e",
          1819 => x"73",
          1820 => x"8a",
          1821 => x"d3",
          1822 => x"80",
          1823 => x"80",
          1824 => x"ee",
          1825 => x"39",
          1826 => x"71",
          1827 => x"53",
          1828 => x"54",
          1829 => x"2e",
          1830 => x"15",
          1831 => x"33",
          1832 => x"72",
          1833 => x"81",
          1834 => x"39",
          1835 => x"56",
          1836 => x"27",
          1837 => x"51",
          1838 => x"75",
          1839 => x"72",
          1840 => x"38",
          1841 => x"df",
          1842 => x"16",
          1843 => x"7b",
          1844 => x"38",
          1845 => x"f2",
          1846 => x"77",
          1847 => x"12",
          1848 => x"53",
          1849 => x"5c",
          1850 => x"5c",
          1851 => x"5c",
          1852 => x"5c",
          1853 => x"51",
          1854 => x"fd",
          1855 => x"82",
          1856 => x"06",
          1857 => x"80",
          1858 => x"77",
          1859 => x"53",
          1860 => x"18",
          1861 => x"72",
          1862 => x"c4",
          1863 => x"70",
          1864 => x"25",
          1865 => x"55",
          1866 => x"8d",
          1867 => x"2e",
          1868 => x"30",
          1869 => x"5b",
          1870 => x"8f",
          1871 => x"7b",
          1872 => x"d9",
          1873 => x"fe",
          1874 => x"ff",
          1875 => x"75",
          1876 => x"d9",
          1877 => x"f0",
          1878 => x"74",
          1879 => x"a7",
          1880 => x"80",
          1881 => x"38",
          1882 => x"72",
          1883 => x"54",
          1884 => x"72",
          1885 => x"05",
          1886 => x"17",
          1887 => x"77",
          1888 => x"51",
          1889 => x"9f",
          1890 => x"72",
          1891 => x"79",
          1892 => x"81",
          1893 => x"72",
          1894 => x"38",
          1895 => x"05",
          1896 => x"ad",
          1897 => x"17",
          1898 => x"81",
          1899 => x"b0",
          1900 => x"38",
          1901 => x"81",
          1902 => x"06",
          1903 => x"9f",
          1904 => x"55",
          1905 => x"97",
          1906 => x"f9",
          1907 => x"81",
          1908 => x"8b",
          1909 => x"16",
          1910 => x"73",
          1911 => x"96",
          1912 => x"e0",
          1913 => x"17",
          1914 => x"33",
          1915 => x"f9",
          1916 => x"f2",
          1917 => x"16",
          1918 => x"7b",
          1919 => x"38",
          1920 => x"c6",
          1921 => x"96",
          1922 => x"fd",
          1923 => x"3d",
          1924 => x"05",
          1925 => x"52",
          1926 => x"e0",
          1927 => x"0d",
          1928 => x"0d",
          1929 => x"8c",
          1930 => x"88",
          1931 => x"51",
          1932 => x"81",
          1933 => x"53",
          1934 => x"80",
          1935 => x"8c",
          1936 => x"0d",
          1937 => x"0d",
          1938 => x"08",
          1939 => x"84",
          1940 => x"88",
          1941 => x"52",
          1942 => x"3f",
          1943 => x"84",
          1944 => x"0d",
          1945 => x"0d",
          1946 => x"ff",
          1947 => x"56",
          1948 => x"80",
          1949 => x"2e",
          1950 => x"81",
          1951 => x"52",
          1952 => x"fe",
          1953 => x"ff",
          1954 => x"80",
          1955 => x"38",
          1956 => x"b9",
          1957 => x"32",
          1958 => x"80",
          1959 => x"52",
          1960 => x"8b",
          1961 => x"2e",
          1962 => x"14",
          1963 => x"9f",
          1964 => x"38",
          1965 => x"73",
          1966 => x"38",
          1967 => x"72",
          1968 => x"14",
          1969 => x"f8",
          1970 => x"af",
          1971 => x"52",
          1972 => x"8a",
          1973 => x"3f",
          1974 => x"81",
          1975 => x"87",
          1976 => x"fe",
          1977 => x"ff",
          1978 => x"81",
          1979 => x"77",
          1980 => x"53",
          1981 => x"72",
          1982 => x"0c",
          1983 => x"04",
          1984 => x"7a",
          1985 => x"80",
          1986 => x"58",
          1987 => x"33",
          1988 => x"a0",
          1989 => x"06",
          1990 => x"13",
          1991 => x"39",
          1992 => x"09",
          1993 => x"38",
          1994 => x"11",
          1995 => x"08",
          1996 => x"54",
          1997 => x"2e",
          1998 => x"80",
          1999 => x"08",
          2000 => x"0c",
          2001 => x"33",
          2002 => x"80",
          2003 => x"38",
          2004 => x"80",
          2005 => x"38",
          2006 => x"57",
          2007 => x"0c",
          2008 => x"33",
          2009 => x"39",
          2010 => x"74",
          2011 => x"38",
          2012 => x"80",
          2013 => x"89",
          2014 => x"38",
          2015 => x"d0",
          2016 => x"55",
          2017 => x"80",
          2018 => x"39",
          2019 => x"d9",
          2020 => x"80",
          2021 => x"27",
          2022 => x"80",
          2023 => x"89",
          2024 => x"70",
          2025 => x"55",
          2026 => x"70",
          2027 => x"55",
          2028 => x"27",
          2029 => x"14",
          2030 => x"06",
          2031 => x"74",
          2032 => x"73",
          2033 => x"38",
          2034 => x"14",
          2035 => x"05",
          2036 => x"08",
          2037 => x"54",
          2038 => x"39",
          2039 => x"84",
          2040 => x"55",
          2041 => x"81",
          2042 => x"fe",
          2043 => x"3d",
          2044 => x"3d",
          2045 => x"5a",
          2046 => x"7a",
          2047 => x"08",
          2048 => x"53",
          2049 => x"09",
          2050 => x"38",
          2051 => x"0c",
          2052 => x"ad",
          2053 => x"06",
          2054 => x"76",
          2055 => x"0c",
          2056 => x"33",
          2057 => x"73",
          2058 => x"81",
          2059 => x"38",
          2060 => x"05",
          2061 => x"08",
          2062 => x"53",
          2063 => x"2e",
          2064 => x"57",
          2065 => x"2e",
          2066 => x"39",
          2067 => x"13",
          2068 => x"08",
          2069 => x"53",
          2070 => x"55",
          2071 => x"80",
          2072 => x"14",
          2073 => x"88",
          2074 => x"27",
          2075 => x"eb",
          2076 => x"53",
          2077 => x"89",
          2078 => x"38",
          2079 => x"55",
          2080 => x"8a",
          2081 => x"a0",
          2082 => x"c2",
          2083 => x"74",
          2084 => x"e0",
          2085 => x"ff",
          2086 => x"d0",
          2087 => x"ff",
          2088 => x"90",
          2089 => x"38",
          2090 => x"81",
          2091 => x"53",
          2092 => x"ca",
          2093 => x"27",
          2094 => x"77",
          2095 => x"08",
          2096 => x"0c",
          2097 => x"33",
          2098 => x"ff",
          2099 => x"80",
          2100 => x"74",
          2101 => x"79",
          2102 => x"74",
          2103 => x"0c",
          2104 => x"04",
          2105 => x"76",
          2106 => x"98",
          2107 => x"2b",
          2108 => x"72",
          2109 => x"82",
          2110 => x"51",
          2111 => x"80",
          2112 => x"cc",
          2113 => x"53",
          2114 => x"9c",
          2115 => x"c8",
          2116 => x"02",
          2117 => x"05",
          2118 => x"52",
          2119 => x"72",
          2120 => x"06",
          2121 => x"53",
          2122 => x"f0",
          2123 => x"0d",
          2124 => x"0d",
          2125 => x"05",
          2126 => x"71",
          2127 => x"53",
          2128 => x"9f",
          2129 => x"f3",
          2130 => x"51",
          2131 => x"88",
          2132 => x"3f",
          2133 => x"05",
          2134 => x"34",
          2135 => x"06",
          2136 => x"76",
          2137 => x"3f",
          2138 => x"86",
          2139 => x"f6",
          2140 => x"02",
          2141 => x"05",
          2142 => x"05",
          2143 => x"81",
          2144 => x"70",
          2145 => x"fa",
          2146 => x"08",
          2147 => x"5a",
          2148 => x"80",
          2149 => x"74",
          2150 => x"3f",
          2151 => x"33",
          2152 => x"81",
          2153 => x"81",
          2154 => x"58",
          2155 => x"bc",
          2156 => x"f0",
          2157 => x"81",
          2158 => x"70",
          2159 => x"fa",
          2160 => x"08",
          2161 => x"74",
          2162 => x"38",
          2163 => x"52",
          2164 => x"e0",
          2165 => x"bc",
          2166 => x"55",
          2167 => x"bc",
          2168 => x"ff",
          2169 => x"75",
          2170 => x"80",
          2171 => x"bc",
          2172 => x"2e",
          2173 => x"fb",
          2174 => x"75",
          2175 => x"38",
          2176 => x"33",
          2177 => x"38",
          2178 => x"05",
          2179 => x"78",
          2180 => x"80",
          2181 => x"81",
          2182 => x"52",
          2183 => x"fd",
          2184 => x"fb",
          2185 => x"80",
          2186 => x"8c",
          2187 => x"dc",
          2188 => x"57",
          2189 => x"fb",
          2190 => x"80",
          2191 => x"81",
          2192 => x"80",
          2193 => x"fb",
          2194 => x"80",
          2195 => x"3d",
          2196 => x"80",
          2197 => x"81",
          2198 => x"80",
          2199 => x"75",
          2200 => x"3f",
          2201 => x"08",
          2202 => x"81",
          2203 => x"25",
          2204 => x"fe",
          2205 => x"05",
          2206 => x"55",
          2207 => x"75",
          2208 => x"81",
          2209 => x"e0",
          2210 => x"ff",
          2211 => x"2e",
          2212 => x"ff",
          2213 => x"3d",
          2214 => x"3d",
          2215 => x"08",
          2216 => x"5a",
          2217 => x"58",
          2218 => x"81",
          2219 => x"51",
          2220 => x"3f",
          2221 => x"08",
          2222 => x"ff",
          2223 => x"b8",
          2224 => x"80",
          2225 => x"3d",
          2226 => x"80",
          2227 => x"81",
          2228 => x"80",
          2229 => x"75",
          2230 => x"3f",
          2231 => x"08",
          2232 => x"55",
          2233 => x"fe",
          2234 => x"8e",
          2235 => x"f0",
          2236 => x"70",
          2237 => x"80",
          2238 => x"09",
          2239 => x"72",
          2240 => x"51",
          2241 => x"77",
          2242 => x"73",
          2243 => x"81",
          2244 => x"8c",
          2245 => x"51",
          2246 => x"3f",
          2247 => x"08",
          2248 => x"38",
          2249 => x"51",
          2250 => x"78",
          2251 => x"81",
          2252 => x"75",
          2253 => x"d5",
          2254 => x"51",
          2255 => x"ab",
          2256 => x"81",
          2257 => x"74",
          2258 => x"77",
          2259 => x"0c",
          2260 => x"04",
          2261 => x"7c",
          2262 => x"71",
          2263 => x"59",
          2264 => x"a0",
          2265 => x"06",
          2266 => x"33",
          2267 => x"77",
          2268 => x"38",
          2269 => x"5b",
          2270 => x"56",
          2271 => x"a0",
          2272 => x"06",
          2273 => x"75",
          2274 => x"80",
          2275 => x"29",
          2276 => x"05",
          2277 => x"55",
          2278 => x"81",
          2279 => x"53",
          2280 => x"08",
          2281 => x"3f",
          2282 => x"08",
          2283 => x"84",
          2284 => x"74",
          2285 => x"38",
          2286 => x"88",
          2287 => x"fc",
          2288 => x"39",
          2289 => x"8c",
          2290 => x"53",
          2291 => x"f6",
          2292 => x"fe",
          2293 => x"2e",
          2294 => x"53",
          2295 => x"51",
          2296 => x"81",
          2297 => x"81",
          2298 => x"74",
          2299 => x"54",
          2300 => x"14",
          2301 => x"06",
          2302 => x"74",
          2303 => x"38",
          2304 => x"81",
          2305 => x"8c",
          2306 => x"d3",
          2307 => x"3d",
          2308 => x"05",
          2309 => x"33",
          2310 => x"0b",
          2311 => x"81",
          2312 => x"5b",
          2313 => x"08",
          2314 => x"81",
          2315 => x"54",
          2316 => x"38",
          2317 => x"b4",
          2318 => x"f0",
          2319 => x"b8",
          2320 => x"f0",
          2321 => x"80",
          2322 => x"53",
          2323 => x"08",
          2324 => x"f0",
          2325 => x"ed",
          2326 => x"f0",
          2327 => x"8b",
          2328 => x"98",
          2329 => x"3f",
          2330 => x"81",
          2331 => x"53",
          2332 => x"90",
          2333 => x"54",
          2334 => x"3f",
          2335 => x"08",
          2336 => x"f0",
          2337 => x"09",
          2338 => x"c1",
          2339 => x"f0",
          2340 => x"bb",
          2341 => x"f0",
          2342 => x"0b",
          2343 => x"08",
          2344 => x"81",
          2345 => x"ff",
          2346 => x"55",
          2347 => x"34",
          2348 => x"81",
          2349 => x"75",
          2350 => x"3f",
          2351 => x"09",
          2352 => x"a7",
          2353 => x"81",
          2354 => x"b4",
          2355 => x"5d",
          2356 => x"81",
          2357 => x"98",
          2358 => x"2c",
          2359 => x"ff",
          2360 => x"78",
          2361 => x"81",
          2362 => x"70",
          2363 => x"98",
          2364 => x"90",
          2365 => x"2b",
          2366 => x"71",
          2367 => x"70",
          2368 => x"e9",
          2369 => x"08",
          2370 => x"51",
          2371 => x"59",
          2372 => x"5d",
          2373 => x"73",
          2374 => x"e9",
          2375 => x"27",
          2376 => x"81",
          2377 => x"81",
          2378 => x"70",
          2379 => x"55",
          2380 => x"80",
          2381 => x"53",
          2382 => x"51",
          2383 => x"81",
          2384 => x"81",
          2385 => x"73",
          2386 => x"38",
          2387 => x"90",
          2388 => x"b1",
          2389 => x"80",
          2390 => x"80",
          2391 => x"98",
          2392 => x"ff",
          2393 => x"55",
          2394 => x"97",
          2395 => x"74",
          2396 => x"f6",
          2397 => x"fe",
          2398 => x"ff",
          2399 => x"cc",
          2400 => x"80",
          2401 => x"2e",
          2402 => x"81",
          2403 => x"81",
          2404 => x"74",
          2405 => x"98",
          2406 => x"90",
          2407 => x"2b",
          2408 => x"70",
          2409 => x"82",
          2410 => x"cc",
          2411 => x"51",
          2412 => x"58",
          2413 => x"77",
          2414 => x"06",
          2415 => x"81",
          2416 => x"08",
          2417 => x"0b",
          2418 => x"34",
          2419 => x"ff",
          2420 => x"39",
          2421 => x"94",
          2422 => x"ff",
          2423 => x"af",
          2424 => x"7d",
          2425 => x"73",
          2426 => x"e1",
          2427 => x"29",
          2428 => x"05",
          2429 => x"04",
          2430 => x"33",
          2431 => x"2e",
          2432 => x"81",
          2433 => x"55",
          2434 => x"ab",
          2435 => x"2b",
          2436 => x"51",
          2437 => x"24",
          2438 => x"1a",
          2439 => x"81",
          2440 => x"81",
          2441 => x"81",
          2442 => x"70",
          2443 => x"ff",
          2444 => x"51",
          2445 => x"81",
          2446 => x"81",
          2447 => x"74",
          2448 => x"34",
          2449 => x"ae",
          2450 => x"34",
          2451 => x"33",
          2452 => x"27",
          2453 => x"14",
          2454 => x"ff",
          2455 => x"ff",
          2456 => x"81",
          2457 => x"81",
          2458 => x"70",
          2459 => x"ff",
          2460 => x"51",
          2461 => x"77",
          2462 => x"74",
          2463 => x"52",
          2464 => x"3f",
          2465 => x"0a",
          2466 => x"0a",
          2467 => x"2c",
          2468 => x"33",
          2469 => x"73",
          2470 => x"38",
          2471 => x"33",
          2472 => x"70",
          2473 => x"ff",
          2474 => x"51",
          2475 => x"77",
          2476 => x"38",
          2477 => x"92",
          2478 => x"80",
          2479 => x"80",
          2480 => x"98",
          2481 => x"98",
          2482 => x"55",
          2483 => x"e4",
          2484 => x"39",
          2485 => x"33",
          2486 => x"06",
          2487 => x"80",
          2488 => x"38",
          2489 => x"33",
          2490 => x"73",
          2491 => x"34",
          2492 => x"73",
          2493 => x"34",
          2494 => x"ce",
          2495 => x"9c",
          2496 => x"2b",
          2497 => x"81",
          2498 => x"57",
          2499 => x"74",
          2500 => x"38",
          2501 => x"81",
          2502 => x"34",
          2503 => x"e7",
          2504 => x"81",
          2505 => x"81",
          2506 => x"70",
          2507 => x"ff",
          2508 => x"51",
          2509 => x"24",
          2510 => x"51",
          2511 => x"81",
          2512 => x"70",
          2513 => x"98",
          2514 => x"98",
          2515 => x"56",
          2516 => x"24",
          2517 => x"88",
          2518 => x"3f",
          2519 => x"0a",
          2520 => x"0a",
          2521 => x"2c",
          2522 => x"33",
          2523 => x"75",
          2524 => x"38",
          2525 => x"81",
          2526 => x"7a",
          2527 => x"74",
          2528 => x"e6",
          2529 => x"ff",
          2530 => x"51",
          2531 => x"81",
          2532 => x"81",
          2533 => x"73",
          2534 => x"ff",
          2535 => x"73",
          2536 => x"c9",
          2537 => x"73",
          2538 => x"f3",
          2539 => x"bd",
          2540 => x"34",
          2541 => x"81",
          2542 => x"54",
          2543 => x"fa",
          2544 => x"51",
          2545 => x"81",
          2546 => x"ff",
          2547 => x"81",
          2548 => x"73",
          2549 => x"54",
          2550 => x"ff",
          2551 => x"ff",
          2552 => x"55",
          2553 => x"f9",
          2554 => x"14",
          2555 => x"ff",
          2556 => x"98",
          2557 => x"2c",
          2558 => x"06",
          2559 => x"74",
          2560 => x"38",
          2561 => x"81",
          2562 => x"34",
          2563 => x"e5",
          2564 => x"81",
          2565 => x"81",
          2566 => x"70",
          2567 => x"ff",
          2568 => x"51",
          2569 => x"24",
          2570 => x"51",
          2571 => x"81",
          2572 => x"70",
          2573 => x"98",
          2574 => x"98",
          2575 => x"56",
          2576 => x"24",
          2577 => x"88",
          2578 => x"3f",
          2579 => x"0a",
          2580 => x"0a",
          2581 => x"2c",
          2582 => x"33",
          2583 => x"75",
          2584 => x"38",
          2585 => x"81",
          2586 => x"70",
          2587 => x"81",
          2588 => x"59",
          2589 => x"77",
          2590 => x"38",
          2591 => x"73",
          2592 => x"34",
          2593 => x"33",
          2594 => x"be",
          2595 => x"9c",
          2596 => x"ff",
          2597 => x"98",
          2598 => x"54",
          2599 => x"dc",
          2600 => x"39",
          2601 => x"81",
          2602 => x"55",
          2603 => x"a4",
          2604 => x"cb",
          2605 => x"fe",
          2606 => x"ff",
          2607 => x"fe",
          2608 => x"ff",
          2609 => x"53",
          2610 => x"51",
          2611 => x"93",
          2612 => x"39",
          2613 => x"81",
          2614 => x"fc",
          2615 => x"54",
          2616 => x"a5",
          2617 => x"ca",
          2618 => x"fe",
          2619 => x"ff",
          2620 => x"fe",
          2621 => x"ff",
          2622 => x"53",
          2623 => x"51",
          2624 => x"ff",
          2625 => x"de",
          2626 => x"55",
          2627 => x"f7",
          2628 => x"51",
          2629 => x"80",
          2630 => x"93",
          2631 => x"06",
          2632 => x"fa",
          2633 => x"74",
          2634 => x"38",
          2635 => x"9f",
          2636 => x"39",
          2637 => x"81",
          2638 => x"84",
          2639 => x"54",
          2640 => x"a9",
          2641 => x"ca",
          2642 => x"fe",
          2643 => x"ff",
          2644 => x"fe",
          2645 => x"ff",
          2646 => x"53",
          2647 => x"51",
          2648 => x"81",
          2649 => x"81",
          2650 => x"a8",
          2651 => x"55",
          2652 => x"f6",
          2653 => x"51",
          2654 => x"81",
          2655 => x"81",
          2656 => x"81",
          2657 => x"81",
          2658 => x"05",
          2659 => x"79",
          2660 => x"3f",
          2661 => x"53",
          2662 => x"33",
          2663 => x"ef",
          2664 => x"a9",
          2665 => x"9c",
          2666 => x"ff",
          2667 => x"98",
          2668 => x"54",
          2669 => x"f6",
          2670 => x"14",
          2671 => x"ff",
          2672 => x"1a",
          2673 => x"54",
          2674 => x"f6",
          2675 => x"ff",
          2676 => x"73",
          2677 => x"f5",
          2678 => x"e1",
          2679 => x"ff",
          2680 => x"05",
          2681 => x"ff",
          2682 => x"e1",
          2683 => x"81",
          2684 => x"80",
          2685 => x"98",
          2686 => x"fe",
          2687 => x"3d",
          2688 => x"3d",
          2689 => x"05",
          2690 => x"52",
          2691 => x"87",
          2692 => x"d8",
          2693 => x"71",
          2694 => x"0c",
          2695 => x"04",
          2696 => x"02",
          2697 => x"02",
          2698 => x"05",
          2699 => x"83",
          2700 => x"26",
          2701 => x"72",
          2702 => x"c0",
          2703 => x"53",
          2704 => x"74",
          2705 => x"38",
          2706 => x"73",
          2707 => x"c0",
          2708 => x"51",
          2709 => x"85",
          2710 => x"98",
          2711 => x"52",
          2712 => x"82",
          2713 => x"70",
          2714 => x"38",
          2715 => x"8c",
          2716 => x"ec",
          2717 => x"fc",
          2718 => x"52",
          2719 => x"87",
          2720 => x"08",
          2721 => x"2e",
          2722 => x"81",
          2723 => x"34",
          2724 => x"13",
          2725 => x"81",
          2726 => x"86",
          2727 => x"f3",
          2728 => x"62",
          2729 => x"05",
          2730 => x"57",
          2731 => x"83",
          2732 => x"fe",
          2733 => x"fe",
          2734 => x"06",
          2735 => x"71",
          2736 => x"71",
          2737 => x"2b",
          2738 => x"80",
          2739 => x"92",
          2740 => x"c0",
          2741 => x"41",
          2742 => x"5a",
          2743 => x"87",
          2744 => x"0c",
          2745 => x"84",
          2746 => x"08",
          2747 => x"70",
          2748 => x"53",
          2749 => x"2e",
          2750 => x"08",
          2751 => x"70",
          2752 => x"34",
          2753 => x"80",
          2754 => x"53",
          2755 => x"2e",
          2756 => x"53",
          2757 => x"26",
          2758 => x"80",
          2759 => x"87",
          2760 => x"08",
          2761 => x"38",
          2762 => x"8c",
          2763 => x"80",
          2764 => x"78",
          2765 => x"99",
          2766 => x"0c",
          2767 => x"8c",
          2768 => x"08",
          2769 => x"51",
          2770 => x"38",
          2771 => x"8d",
          2772 => x"17",
          2773 => x"81",
          2774 => x"53",
          2775 => x"2e",
          2776 => x"fc",
          2777 => x"52",
          2778 => x"7d",
          2779 => x"ed",
          2780 => x"80",
          2781 => x"71",
          2782 => x"38",
          2783 => x"53",
          2784 => x"f0",
          2785 => x"0d",
          2786 => x"0d",
          2787 => x"02",
          2788 => x"05",
          2789 => x"58",
          2790 => x"80",
          2791 => x"fc",
          2792 => x"fe",
          2793 => x"06",
          2794 => x"71",
          2795 => x"81",
          2796 => x"38",
          2797 => x"2b",
          2798 => x"80",
          2799 => x"92",
          2800 => x"c0",
          2801 => x"40",
          2802 => x"5a",
          2803 => x"c0",
          2804 => x"76",
          2805 => x"76",
          2806 => x"75",
          2807 => x"2a",
          2808 => x"51",
          2809 => x"80",
          2810 => x"7a",
          2811 => x"5c",
          2812 => x"81",
          2813 => x"81",
          2814 => x"06",
          2815 => x"80",
          2816 => x"87",
          2817 => x"08",
          2818 => x"38",
          2819 => x"8c",
          2820 => x"80",
          2821 => x"77",
          2822 => x"99",
          2823 => x"0c",
          2824 => x"8c",
          2825 => x"08",
          2826 => x"51",
          2827 => x"38",
          2828 => x"8d",
          2829 => x"70",
          2830 => x"84",
          2831 => x"5b",
          2832 => x"2e",
          2833 => x"fc",
          2834 => x"52",
          2835 => x"7d",
          2836 => x"f8",
          2837 => x"80",
          2838 => x"71",
          2839 => x"38",
          2840 => x"53",
          2841 => x"f0",
          2842 => x"0d",
          2843 => x"0d",
          2844 => x"05",
          2845 => x"02",
          2846 => x"05",
          2847 => x"54",
          2848 => x"fe",
          2849 => x"f0",
          2850 => x"53",
          2851 => x"80",
          2852 => x"0b",
          2853 => x"8c",
          2854 => x"71",
          2855 => x"dc",
          2856 => x"24",
          2857 => x"84",
          2858 => x"92",
          2859 => x"54",
          2860 => x"8d",
          2861 => x"39",
          2862 => x"80",
          2863 => x"cb",
          2864 => x"70",
          2865 => x"81",
          2866 => x"52",
          2867 => x"8a",
          2868 => x"98",
          2869 => x"71",
          2870 => x"c0",
          2871 => x"52",
          2872 => x"81",
          2873 => x"c0",
          2874 => x"53",
          2875 => x"82",
          2876 => x"71",
          2877 => x"39",
          2878 => x"39",
          2879 => x"77",
          2880 => x"81",
          2881 => x"72",
          2882 => x"84",
          2883 => x"73",
          2884 => x"0c",
          2885 => x"04",
          2886 => x"74",
          2887 => x"71",
          2888 => x"2b",
          2889 => x"f0",
          2890 => x"84",
          2891 => x"fd",
          2892 => x"83",
          2893 => x"12",
          2894 => x"2b",
          2895 => x"07",
          2896 => x"70",
          2897 => x"2b",
          2898 => x"07",
          2899 => x"0c",
          2900 => x"56",
          2901 => x"3d",
          2902 => x"3d",
          2903 => x"84",
          2904 => x"22",
          2905 => x"72",
          2906 => x"54",
          2907 => x"2a",
          2908 => x"34",
          2909 => x"04",
          2910 => x"73",
          2911 => x"70",
          2912 => x"05",
          2913 => x"88",
          2914 => x"72",
          2915 => x"54",
          2916 => x"2a",
          2917 => x"70",
          2918 => x"34",
          2919 => x"51",
          2920 => x"83",
          2921 => x"fe",
          2922 => x"75",
          2923 => x"51",
          2924 => x"92",
          2925 => x"81",
          2926 => x"73",
          2927 => x"55",
          2928 => x"51",
          2929 => x"3d",
          2930 => x"3d",
          2931 => x"76",
          2932 => x"72",
          2933 => x"05",
          2934 => x"11",
          2935 => x"38",
          2936 => x"04",
          2937 => x"78",
          2938 => x"56",
          2939 => x"81",
          2940 => x"74",
          2941 => x"56",
          2942 => x"31",
          2943 => x"52",
          2944 => x"80",
          2945 => x"71",
          2946 => x"38",
          2947 => x"f0",
          2948 => x"0d",
          2949 => x"0d",
          2950 => x"51",
          2951 => x"73",
          2952 => x"81",
          2953 => x"33",
          2954 => x"38",
          2955 => x"fe",
          2956 => x"3d",
          2957 => x"0b",
          2958 => x"0c",
          2959 => x"81",
          2960 => x"04",
          2961 => x"7b",
          2962 => x"83",
          2963 => x"5a",
          2964 => x"80",
          2965 => x"54",
          2966 => x"53",
          2967 => x"53",
          2968 => x"52",
          2969 => x"3f",
          2970 => x"08",
          2971 => x"81",
          2972 => x"81",
          2973 => x"83",
          2974 => x"16",
          2975 => x"18",
          2976 => x"18",
          2977 => x"58",
          2978 => x"9f",
          2979 => x"33",
          2980 => x"2e",
          2981 => x"93",
          2982 => x"76",
          2983 => x"52",
          2984 => x"51",
          2985 => x"83",
          2986 => x"79",
          2987 => x"0c",
          2988 => x"04",
          2989 => x"78",
          2990 => x"80",
          2991 => x"17",
          2992 => x"38",
          2993 => x"fc",
          2994 => x"f0",
          2995 => x"fe",
          2996 => x"38",
          2997 => x"53",
          2998 => x"81",
          2999 => x"f7",
          3000 => x"fe",
          3001 => x"2e",
          3002 => x"55",
          3003 => x"b0",
          3004 => x"81",
          3005 => x"88",
          3006 => x"f8",
          3007 => x"70",
          3008 => x"c0",
          3009 => x"f0",
          3010 => x"fe",
          3011 => x"91",
          3012 => x"55",
          3013 => x"09",
          3014 => x"f0",
          3015 => x"33",
          3016 => x"2e",
          3017 => x"80",
          3018 => x"80",
          3019 => x"f0",
          3020 => x"17",
          3021 => x"fd",
          3022 => x"d4",
          3023 => x"b2",
          3024 => x"96",
          3025 => x"85",
          3026 => x"75",
          3027 => x"3f",
          3028 => x"e4",
          3029 => x"98",
          3030 => x"9c",
          3031 => x"08",
          3032 => x"17",
          3033 => x"3f",
          3034 => x"52",
          3035 => x"51",
          3036 => x"a0",
          3037 => x"05",
          3038 => x"0c",
          3039 => x"75",
          3040 => x"33",
          3041 => x"3f",
          3042 => x"34",
          3043 => x"52",
          3044 => x"51",
          3045 => x"81",
          3046 => x"80",
          3047 => x"81",
          3048 => x"fe",
          3049 => x"3d",
          3050 => x"3d",
          3051 => x"1a",
          3052 => x"fe",
          3053 => x"54",
          3054 => x"73",
          3055 => x"8a",
          3056 => x"71",
          3057 => x"08",
          3058 => x"75",
          3059 => x"0c",
          3060 => x"04",
          3061 => x"7a",
          3062 => x"56",
          3063 => x"77",
          3064 => x"38",
          3065 => x"08",
          3066 => x"38",
          3067 => x"54",
          3068 => x"2e",
          3069 => x"72",
          3070 => x"38",
          3071 => x"8d",
          3072 => x"39",
          3073 => x"81",
          3074 => x"b6",
          3075 => x"2a",
          3076 => x"2a",
          3077 => x"05",
          3078 => x"55",
          3079 => x"81",
          3080 => x"81",
          3081 => x"83",
          3082 => x"b4",
          3083 => x"17",
          3084 => x"a4",
          3085 => x"55",
          3086 => x"57",
          3087 => x"3f",
          3088 => x"08",
          3089 => x"74",
          3090 => x"14",
          3091 => x"70",
          3092 => x"07",
          3093 => x"71",
          3094 => x"52",
          3095 => x"72",
          3096 => x"75",
          3097 => x"58",
          3098 => x"76",
          3099 => x"15",
          3100 => x"73",
          3101 => x"3f",
          3102 => x"08",
          3103 => x"76",
          3104 => x"06",
          3105 => x"05",
          3106 => x"3f",
          3107 => x"08",
          3108 => x"06",
          3109 => x"76",
          3110 => x"15",
          3111 => x"73",
          3112 => x"3f",
          3113 => x"08",
          3114 => x"82",
          3115 => x"06",
          3116 => x"05",
          3117 => x"3f",
          3118 => x"08",
          3119 => x"58",
          3120 => x"58",
          3121 => x"f0",
          3122 => x"0d",
          3123 => x"0d",
          3124 => x"5a",
          3125 => x"59",
          3126 => x"82",
          3127 => x"98",
          3128 => x"82",
          3129 => x"33",
          3130 => x"2e",
          3131 => x"72",
          3132 => x"38",
          3133 => x"8d",
          3134 => x"39",
          3135 => x"81",
          3136 => x"f7",
          3137 => x"2a",
          3138 => x"2a",
          3139 => x"05",
          3140 => x"55",
          3141 => x"81",
          3142 => x"59",
          3143 => x"08",
          3144 => x"74",
          3145 => x"16",
          3146 => x"16",
          3147 => x"59",
          3148 => x"53",
          3149 => x"8f",
          3150 => x"2b",
          3151 => x"74",
          3152 => x"71",
          3153 => x"72",
          3154 => x"0b",
          3155 => x"74",
          3156 => x"17",
          3157 => x"75",
          3158 => x"3f",
          3159 => x"08",
          3160 => x"f0",
          3161 => x"38",
          3162 => x"06",
          3163 => x"78",
          3164 => x"54",
          3165 => x"77",
          3166 => x"33",
          3167 => x"71",
          3168 => x"51",
          3169 => x"34",
          3170 => x"76",
          3171 => x"17",
          3172 => x"75",
          3173 => x"3f",
          3174 => x"08",
          3175 => x"f0",
          3176 => x"38",
          3177 => x"ff",
          3178 => x"10",
          3179 => x"76",
          3180 => x"51",
          3181 => x"be",
          3182 => x"2a",
          3183 => x"05",
          3184 => x"f9",
          3185 => x"fe",
          3186 => x"81",
          3187 => x"ab",
          3188 => x"0a",
          3189 => x"2b",
          3190 => x"70",
          3191 => x"70",
          3192 => x"54",
          3193 => x"81",
          3194 => x"8f",
          3195 => x"07",
          3196 => x"f7",
          3197 => x"0b",
          3198 => x"78",
          3199 => x"0c",
          3200 => x"04",
          3201 => x"7a",
          3202 => x"08",
          3203 => x"59",
          3204 => x"a4",
          3205 => x"17",
          3206 => x"38",
          3207 => x"aa",
          3208 => x"73",
          3209 => x"fd",
          3210 => x"fe",
          3211 => x"81",
          3212 => x"80",
          3213 => x"39",
          3214 => x"eb",
          3215 => x"80",
          3216 => x"fe",
          3217 => x"80",
          3218 => x"52",
          3219 => x"84",
          3220 => x"f0",
          3221 => x"fe",
          3222 => x"2e",
          3223 => x"81",
          3224 => x"81",
          3225 => x"81",
          3226 => x"ff",
          3227 => x"80",
          3228 => x"75",
          3229 => x"3f",
          3230 => x"08",
          3231 => x"16",
          3232 => x"90",
          3233 => x"55",
          3234 => x"27",
          3235 => x"15",
          3236 => x"84",
          3237 => x"07",
          3238 => x"17",
          3239 => x"76",
          3240 => x"a6",
          3241 => x"73",
          3242 => x"0c",
          3243 => x"04",
          3244 => x"7c",
          3245 => x"59",
          3246 => x"95",
          3247 => x"08",
          3248 => x"2e",
          3249 => x"17",
          3250 => x"b2",
          3251 => x"ae",
          3252 => x"7a",
          3253 => x"3f",
          3254 => x"81",
          3255 => x"27",
          3256 => x"81",
          3257 => x"55",
          3258 => x"08",
          3259 => x"d2",
          3260 => x"08",
          3261 => x"08",
          3262 => x"38",
          3263 => x"17",
          3264 => x"54",
          3265 => x"82",
          3266 => x"7a",
          3267 => x"06",
          3268 => x"81",
          3269 => x"17",
          3270 => x"83",
          3271 => x"75",
          3272 => x"f9",
          3273 => x"59",
          3274 => x"08",
          3275 => x"81",
          3276 => x"81",
          3277 => x"59",
          3278 => x"08",
          3279 => x"70",
          3280 => x"25",
          3281 => x"81",
          3282 => x"54",
          3283 => x"55",
          3284 => x"38",
          3285 => x"08",
          3286 => x"38",
          3287 => x"54",
          3288 => x"90",
          3289 => x"18",
          3290 => x"38",
          3291 => x"39",
          3292 => x"38",
          3293 => x"16",
          3294 => x"08",
          3295 => x"38",
          3296 => x"78",
          3297 => x"38",
          3298 => x"51",
          3299 => x"81",
          3300 => x"80",
          3301 => x"80",
          3302 => x"f0",
          3303 => x"09",
          3304 => x"38",
          3305 => x"08",
          3306 => x"f0",
          3307 => x"30",
          3308 => x"80",
          3309 => x"07",
          3310 => x"55",
          3311 => x"38",
          3312 => x"09",
          3313 => x"ae",
          3314 => x"80",
          3315 => x"53",
          3316 => x"51",
          3317 => x"81",
          3318 => x"81",
          3319 => x"30",
          3320 => x"f0",
          3321 => x"25",
          3322 => x"79",
          3323 => x"38",
          3324 => x"8f",
          3325 => x"79",
          3326 => x"f9",
          3327 => x"fe",
          3328 => x"74",
          3329 => x"8c",
          3330 => x"17",
          3331 => x"90",
          3332 => x"54",
          3333 => x"86",
          3334 => x"90",
          3335 => x"17",
          3336 => x"54",
          3337 => x"34",
          3338 => x"56",
          3339 => x"90",
          3340 => x"80",
          3341 => x"81",
          3342 => x"55",
          3343 => x"56",
          3344 => x"81",
          3345 => x"8c",
          3346 => x"f8",
          3347 => x"70",
          3348 => x"f0",
          3349 => x"f0",
          3350 => x"56",
          3351 => x"08",
          3352 => x"7b",
          3353 => x"f6",
          3354 => x"fe",
          3355 => x"fe",
          3356 => x"17",
          3357 => x"80",
          3358 => x"b4",
          3359 => x"57",
          3360 => x"77",
          3361 => x"81",
          3362 => x"15",
          3363 => x"78",
          3364 => x"81",
          3365 => x"53",
          3366 => x"15",
          3367 => x"e9",
          3368 => x"f0",
          3369 => x"df",
          3370 => x"22",
          3371 => x"30",
          3372 => x"70",
          3373 => x"51",
          3374 => x"81",
          3375 => x"8a",
          3376 => x"f8",
          3377 => x"7c",
          3378 => x"56",
          3379 => x"80",
          3380 => x"f1",
          3381 => x"06",
          3382 => x"e9",
          3383 => x"18",
          3384 => x"08",
          3385 => x"38",
          3386 => x"82",
          3387 => x"38",
          3388 => x"54",
          3389 => x"74",
          3390 => x"82",
          3391 => x"22",
          3392 => x"79",
          3393 => x"38",
          3394 => x"98",
          3395 => x"cd",
          3396 => x"22",
          3397 => x"54",
          3398 => x"26",
          3399 => x"52",
          3400 => x"b0",
          3401 => x"f0",
          3402 => x"fe",
          3403 => x"2e",
          3404 => x"0b",
          3405 => x"08",
          3406 => x"98",
          3407 => x"fe",
          3408 => x"85",
          3409 => x"bd",
          3410 => x"31",
          3411 => x"73",
          3412 => x"f4",
          3413 => x"fe",
          3414 => x"18",
          3415 => x"18",
          3416 => x"08",
          3417 => x"72",
          3418 => x"38",
          3419 => x"58",
          3420 => x"89",
          3421 => x"18",
          3422 => x"ff",
          3423 => x"05",
          3424 => x"80",
          3425 => x"fe",
          3426 => x"3d",
          3427 => x"3d",
          3428 => x"08",
          3429 => x"a0",
          3430 => x"54",
          3431 => x"77",
          3432 => x"80",
          3433 => x"0c",
          3434 => x"53",
          3435 => x"80",
          3436 => x"38",
          3437 => x"06",
          3438 => x"b5",
          3439 => x"98",
          3440 => x"14",
          3441 => x"92",
          3442 => x"2a",
          3443 => x"56",
          3444 => x"26",
          3445 => x"80",
          3446 => x"16",
          3447 => x"77",
          3448 => x"53",
          3449 => x"38",
          3450 => x"51",
          3451 => x"81",
          3452 => x"53",
          3453 => x"0b",
          3454 => x"08",
          3455 => x"38",
          3456 => x"fe",
          3457 => x"2e",
          3458 => x"98",
          3459 => x"fe",
          3460 => x"80",
          3461 => x"8a",
          3462 => x"15",
          3463 => x"80",
          3464 => x"14",
          3465 => x"51",
          3466 => x"81",
          3467 => x"53",
          3468 => x"fe",
          3469 => x"2e",
          3470 => x"82",
          3471 => x"f0",
          3472 => x"ba",
          3473 => x"81",
          3474 => x"ff",
          3475 => x"81",
          3476 => x"52",
          3477 => x"f3",
          3478 => x"f0",
          3479 => x"72",
          3480 => x"72",
          3481 => x"f2",
          3482 => x"fe",
          3483 => x"15",
          3484 => x"15",
          3485 => x"b4",
          3486 => x"0c",
          3487 => x"81",
          3488 => x"8a",
          3489 => x"f7",
          3490 => x"7d",
          3491 => x"5b",
          3492 => x"76",
          3493 => x"3f",
          3494 => x"08",
          3495 => x"f0",
          3496 => x"38",
          3497 => x"08",
          3498 => x"08",
          3499 => x"f0",
          3500 => x"fe",
          3501 => x"81",
          3502 => x"80",
          3503 => x"fe",
          3504 => x"18",
          3505 => x"51",
          3506 => x"81",
          3507 => x"81",
          3508 => x"81",
          3509 => x"f0",
          3510 => x"83",
          3511 => x"77",
          3512 => x"72",
          3513 => x"38",
          3514 => x"75",
          3515 => x"81",
          3516 => x"a5",
          3517 => x"f0",
          3518 => x"52",
          3519 => x"8e",
          3520 => x"f0",
          3521 => x"fe",
          3522 => x"2e",
          3523 => x"73",
          3524 => x"81",
          3525 => x"87",
          3526 => x"fe",
          3527 => x"3d",
          3528 => x"3d",
          3529 => x"11",
          3530 => x"ec",
          3531 => x"f0",
          3532 => x"ff",
          3533 => x"33",
          3534 => x"71",
          3535 => x"81",
          3536 => x"94",
          3537 => x"d0",
          3538 => x"f0",
          3539 => x"73",
          3540 => x"81",
          3541 => x"85",
          3542 => x"fc",
          3543 => x"79",
          3544 => x"ff",
          3545 => x"12",
          3546 => x"eb",
          3547 => x"70",
          3548 => x"72",
          3549 => x"81",
          3550 => x"73",
          3551 => x"94",
          3552 => x"d6",
          3553 => x"0d",
          3554 => x"0d",
          3555 => x"55",
          3556 => x"5a",
          3557 => x"08",
          3558 => x"8a",
          3559 => x"08",
          3560 => x"ee",
          3561 => x"fe",
          3562 => x"81",
          3563 => x"80",
          3564 => x"15",
          3565 => x"55",
          3566 => x"38",
          3567 => x"e6",
          3568 => x"33",
          3569 => x"70",
          3570 => x"58",
          3571 => x"86",
          3572 => x"fe",
          3573 => x"73",
          3574 => x"83",
          3575 => x"73",
          3576 => x"38",
          3577 => x"06",
          3578 => x"80",
          3579 => x"75",
          3580 => x"38",
          3581 => x"08",
          3582 => x"54",
          3583 => x"2e",
          3584 => x"83",
          3585 => x"73",
          3586 => x"38",
          3587 => x"51",
          3588 => x"81",
          3589 => x"58",
          3590 => x"08",
          3591 => x"15",
          3592 => x"38",
          3593 => x"0b",
          3594 => x"77",
          3595 => x"0c",
          3596 => x"04",
          3597 => x"77",
          3598 => x"54",
          3599 => x"51",
          3600 => x"81",
          3601 => x"55",
          3602 => x"08",
          3603 => x"14",
          3604 => x"51",
          3605 => x"81",
          3606 => x"55",
          3607 => x"08",
          3608 => x"53",
          3609 => x"08",
          3610 => x"08",
          3611 => x"3f",
          3612 => x"14",
          3613 => x"08",
          3614 => x"3f",
          3615 => x"17",
          3616 => x"fe",
          3617 => x"3d",
          3618 => x"3d",
          3619 => x"08",
          3620 => x"54",
          3621 => x"53",
          3622 => x"81",
          3623 => x"8d",
          3624 => x"08",
          3625 => x"34",
          3626 => x"15",
          3627 => x"0d",
          3628 => x"0d",
          3629 => x"57",
          3630 => x"17",
          3631 => x"08",
          3632 => x"82",
          3633 => x"89",
          3634 => x"55",
          3635 => x"14",
          3636 => x"16",
          3637 => x"71",
          3638 => x"38",
          3639 => x"09",
          3640 => x"38",
          3641 => x"73",
          3642 => x"81",
          3643 => x"ae",
          3644 => x"05",
          3645 => x"15",
          3646 => x"70",
          3647 => x"34",
          3648 => x"8a",
          3649 => x"38",
          3650 => x"05",
          3651 => x"81",
          3652 => x"17",
          3653 => x"12",
          3654 => x"34",
          3655 => x"9c",
          3656 => x"e8",
          3657 => x"fe",
          3658 => x"0c",
          3659 => x"e7",
          3660 => x"fe",
          3661 => x"17",
          3662 => x"51",
          3663 => x"81",
          3664 => x"84",
          3665 => x"3d",
          3666 => x"3d",
          3667 => x"08",
          3668 => x"61",
          3669 => x"55",
          3670 => x"2e",
          3671 => x"55",
          3672 => x"2e",
          3673 => x"80",
          3674 => x"94",
          3675 => x"1c",
          3676 => x"81",
          3677 => x"61",
          3678 => x"56",
          3679 => x"2e",
          3680 => x"83",
          3681 => x"73",
          3682 => x"70",
          3683 => x"25",
          3684 => x"51",
          3685 => x"38",
          3686 => x"0c",
          3687 => x"51",
          3688 => x"26",
          3689 => x"80",
          3690 => x"34",
          3691 => x"51",
          3692 => x"81",
          3693 => x"55",
          3694 => x"91",
          3695 => x"1d",
          3696 => x"8b",
          3697 => x"79",
          3698 => x"3f",
          3699 => x"57",
          3700 => x"55",
          3701 => x"2e",
          3702 => x"80",
          3703 => x"18",
          3704 => x"1a",
          3705 => x"70",
          3706 => x"2a",
          3707 => x"07",
          3708 => x"5a",
          3709 => x"8c",
          3710 => x"54",
          3711 => x"81",
          3712 => x"39",
          3713 => x"70",
          3714 => x"2a",
          3715 => x"75",
          3716 => x"8c",
          3717 => x"2e",
          3718 => x"a0",
          3719 => x"38",
          3720 => x"0c",
          3721 => x"76",
          3722 => x"38",
          3723 => x"b8",
          3724 => x"70",
          3725 => x"5a",
          3726 => x"76",
          3727 => x"38",
          3728 => x"70",
          3729 => x"dc",
          3730 => x"72",
          3731 => x"80",
          3732 => x"51",
          3733 => x"73",
          3734 => x"38",
          3735 => x"18",
          3736 => x"1a",
          3737 => x"55",
          3738 => x"2e",
          3739 => x"83",
          3740 => x"73",
          3741 => x"70",
          3742 => x"25",
          3743 => x"51",
          3744 => x"38",
          3745 => x"75",
          3746 => x"81",
          3747 => x"81",
          3748 => x"27",
          3749 => x"73",
          3750 => x"38",
          3751 => x"70",
          3752 => x"32",
          3753 => x"80",
          3754 => x"2a",
          3755 => x"56",
          3756 => x"81",
          3757 => x"57",
          3758 => x"f5",
          3759 => x"2b",
          3760 => x"25",
          3761 => x"80",
          3762 => x"eb",
          3763 => x"57",
          3764 => x"e6",
          3765 => x"fe",
          3766 => x"2e",
          3767 => x"18",
          3768 => x"1a",
          3769 => x"56",
          3770 => x"3f",
          3771 => x"08",
          3772 => x"e8",
          3773 => x"54",
          3774 => x"80",
          3775 => x"17",
          3776 => x"34",
          3777 => x"11",
          3778 => x"74",
          3779 => x"75",
          3780 => x"fc",
          3781 => x"3f",
          3782 => x"08",
          3783 => x"9f",
          3784 => x"99",
          3785 => x"e0",
          3786 => x"ff",
          3787 => x"79",
          3788 => x"74",
          3789 => x"57",
          3790 => x"77",
          3791 => x"76",
          3792 => x"38",
          3793 => x"73",
          3794 => x"09",
          3795 => x"38",
          3796 => x"84",
          3797 => x"27",
          3798 => x"39",
          3799 => x"f2",
          3800 => x"80",
          3801 => x"54",
          3802 => x"34",
          3803 => x"58",
          3804 => x"f2",
          3805 => x"fe",
          3806 => x"81",
          3807 => x"80",
          3808 => x"1b",
          3809 => x"51",
          3810 => x"81",
          3811 => x"56",
          3812 => x"08",
          3813 => x"9c",
          3814 => x"33",
          3815 => x"80",
          3816 => x"38",
          3817 => x"bf",
          3818 => x"86",
          3819 => x"15",
          3820 => x"2a",
          3821 => x"51",
          3822 => x"92",
          3823 => x"79",
          3824 => x"e4",
          3825 => x"fe",
          3826 => x"2e",
          3827 => x"52",
          3828 => x"ba",
          3829 => x"39",
          3830 => x"33",
          3831 => x"80",
          3832 => x"74",
          3833 => x"81",
          3834 => x"38",
          3835 => x"70",
          3836 => x"82",
          3837 => x"54",
          3838 => x"96",
          3839 => x"06",
          3840 => x"2e",
          3841 => x"ff",
          3842 => x"1c",
          3843 => x"80",
          3844 => x"81",
          3845 => x"ba",
          3846 => x"b6",
          3847 => x"2a",
          3848 => x"51",
          3849 => x"38",
          3850 => x"70",
          3851 => x"81",
          3852 => x"55",
          3853 => x"e1",
          3854 => x"08",
          3855 => x"1d",
          3856 => x"7c",
          3857 => x"3f",
          3858 => x"08",
          3859 => x"fa",
          3860 => x"81",
          3861 => x"8f",
          3862 => x"f6",
          3863 => x"5b",
          3864 => x"70",
          3865 => x"59",
          3866 => x"73",
          3867 => x"c6",
          3868 => x"81",
          3869 => x"70",
          3870 => x"52",
          3871 => x"8d",
          3872 => x"38",
          3873 => x"09",
          3874 => x"a5",
          3875 => x"d0",
          3876 => x"ff",
          3877 => x"53",
          3878 => x"91",
          3879 => x"73",
          3880 => x"d0",
          3881 => x"71",
          3882 => x"f7",
          3883 => x"81",
          3884 => x"55",
          3885 => x"55",
          3886 => x"81",
          3887 => x"74",
          3888 => x"56",
          3889 => x"12",
          3890 => x"70",
          3891 => x"38",
          3892 => x"81",
          3893 => x"51",
          3894 => x"51",
          3895 => x"89",
          3896 => x"70",
          3897 => x"53",
          3898 => x"70",
          3899 => x"51",
          3900 => x"09",
          3901 => x"38",
          3902 => x"38",
          3903 => x"77",
          3904 => x"70",
          3905 => x"2a",
          3906 => x"07",
          3907 => x"51",
          3908 => x"8f",
          3909 => x"84",
          3910 => x"83",
          3911 => x"94",
          3912 => x"74",
          3913 => x"38",
          3914 => x"0c",
          3915 => x"86",
          3916 => x"b4",
          3917 => x"81",
          3918 => x"8c",
          3919 => x"fa",
          3920 => x"56",
          3921 => x"17",
          3922 => x"b0",
          3923 => x"52",
          3924 => x"e0",
          3925 => x"81",
          3926 => x"81",
          3927 => x"b2",
          3928 => x"b4",
          3929 => x"f0",
          3930 => x"ff",
          3931 => x"55",
          3932 => x"d5",
          3933 => x"06",
          3934 => x"80",
          3935 => x"33",
          3936 => x"81",
          3937 => x"81",
          3938 => x"81",
          3939 => x"eb",
          3940 => x"70",
          3941 => x"07",
          3942 => x"73",
          3943 => x"81",
          3944 => x"81",
          3945 => x"83",
          3946 => x"8c",
          3947 => x"16",
          3948 => x"3f",
          3949 => x"08",
          3950 => x"f0",
          3951 => x"9d",
          3952 => x"81",
          3953 => x"81",
          3954 => x"e0",
          3955 => x"fe",
          3956 => x"81",
          3957 => x"80",
          3958 => x"82",
          3959 => x"fe",
          3960 => x"3d",
          3961 => x"3d",
          3962 => x"84",
          3963 => x"05",
          3964 => x"80",
          3965 => x"51",
          3966 => x"81",
          3967 => x"58",
          3968 => x"0b",
          3969 => x"08",
          3970 => x"38",
          3971 => x"08",
          3972 => x"ff",
          3973 => x"08",
          3974 => x"56",
          3975 => x"86",
          3976 => x"75",
          3977 => x"fe",
          3978 => x"54",
          3979 => x"2e",
          3980 => x"14",
          3981 => x"ca",
          3982 => x"f0",
          3983 => x"06",
          3984 => x"54",
          3985 => x"38",
          3986 => x"86",
          3987 => x"82",
          3988 => x"06",
          3989 => x"56",
          3990 => x"38",
          3991 => x"80",
          3992 => x"81",
          3993 => x"52",
          3994 => x"51",
          3995 => x"81",
          3996 => x"81",
          3997 => x"81",
          3998 => x"83",
          3999 => x"87",
          4000 => x"2e",
          4001 => x"82",
          4002 => x"06",
          4003 => x"56",
          4004 => x"38",
          4005 => x"74",
          4006 => x"a3",
          4007 => x"f0",
          4008 => x"06",
          4009 => x"2e",
          4010 => x"80",
          4011 => x"3d",
          4012 => x"83",
          4013 => x"15",
          4014 => x"53",
          4015 => x"8d",
          4016 => x"15",
          4017 => x"3f",
          4018 => x"08",
          4019 => x"70",
          4020 => x"0c",
          4021 => x"16",
          4022 => x"80",
          4023 => x"80",
          4024 => x"54",
          4025 => x"84",
          4026 => x"5b",
          4027 => x"80",
          4028 => x"7a",
          4029 => x"fc",
          4030 => x"fe",
          4031 => x"ff",
          4032 => x"77",
          4033 => x"81",
          4034 => x"76",
          4035 => x"81",
          4036 => x"2e",
          4037 => x"8d",
          4038 => x"26",
          4039 => x"bf",
          4040 => x"f4",
          4041 => x"f0",
          4042 => x"ff",
          4043 => x"84",
          4044 => x"81",
          4045 => x"38",
          4046 => x"51",
          4047 => x"81",
          4048 => x"83",
          4049 => x"58",
          4050 => x"80",
          4051 => x"db",
          4052 => x"fe",
          4053 => x"77",
          4054 => x"80",
          4055 => x"82",
          4056 => x"c4",
          4057 => x"11",
          4058 => x"06",
          4059 => x"8d",
          4060 => x"26",
          4061 => x"74",
          4062 => x"78",
          4063 => x"c1",
          4064 => x"59",
          4065 => x"15",
          4066 => x"2e",
          4067 => x"13",
          4068 => x"72",
          4069 => x"38",
          4070 => x"eb",
          4071 => x"14",
          4072 => x"3f",
          4073 => x"08",
          4074 => x"f0",
          4075 => x"23",
          4076 => x"57",
          4077 => x"83",
          4078 => x"c7",
          4079 => x"d8",
          4080 => x"f0",
          4081 => x"ff",
          4082 => x"8d",
          4083 => x"14",
          4084 => x"3f",
          4085 => x"08",
          4086 => x"14",
          4087 => x"3f",
          4088 => x"08",
          4089 => x"06",
          4090 => x"72",
          4091 => x"97",
          4092 => x"22",
          4093 => x"84",
          4094 => x"5a",
          4095 => x"83",
          4096 => x"14",
          4097 => x"79",
          4098 => x"93",
          4099 => x"fe",
          4100 => x"81",
          4101 => x"80",
          4102 => x"38",
          4103 => x"08",
          4104 => x"ff",
          4105 => x"38",
          4106 => x"83",
          4107 => x"83",
          4108 => x"74",
          4109 => x"85",
          4110 => x"89",
          4111 => x"76",
          4112 => x"c3",
          4113 => x"70",
          4114 => x"7b",
          4115 => x"73",
          4116 => x"17",
          4117 => x"ac",
          4118 => x"55",
          4119 => x"09",
          4120 => x"38",
          4121 => x"51",
          4122 => x"81",
          4123 => x"83",
          4124 => x"53",
          4125 => x"82",
          4126 => x"82",
          4127 => x"e0",
          4128 => x"ab",
          4129 => x"f0",
          4130 => x"0c",
          4131 => x"53",
          4132 => x"56",
          4133 => x"81",
          4134 => x"13",
          4135 => x"74",
          4136 => x"82",
          4137 => x"74",
          4138 => x"81",
          4139 => x"06",
          4140 => x"83",
          4141 => x"2a",
          4142 => x"72",
          4143 => x"26",
          4144 => x"ff",
          4145 => x"0c",
          4146 => x"15",
          4147 => x"0b",
          4148 => x"76",
          4149 => x"81",
          4150 => x"38",
          4151 => x"51",
          4152 => x"81",
          4153 => x"83",
          4154 => x"53",
          4155 => x"09",
          4156 => x"f9",
          4157 => x"52",
          4158 => x"b8",
          4159 => x"f0",
          4160 => x"38",
          4161 => x"08",
          4162 => x"84",
          4163 => x"d8",
          4164 => x"fe",
          4165 => x"ff",
          4166 => x"72",
          4167 => x"2e",
          4168 => x"80",
          4169 => x"14",
          4170 => x"3f",
          4171 => x"08",
          4172 => x"a4",
          4173 => x"81",
          4174 => x"84",
          4175 => x"d7",
          4176 => x"fe",
          4177 => x"8a",
          4178 => x"2e",
          4179 => x"9d",
          4180 => x"14",
          4181 => x"3f",
          4182 => x"08",
          4183 => x"84",
          4184 => x"d7",
          4185 => x"fe",
          4186 => x"15",
          4187 => x"34",
          4188 => x"22",
          4189 => x"72",
          4190 => x"23",
          4191 => x"23",
          4192 => x"15",
          4193 => x"75",
          4194 => x"0c",
          4195 => x"04",
          4196 => x"77",
          4197 => x"73",
          4198 => x"38",
          4199 => x"72",
          4200 => x"38",
          4201 => x"71",
          4202 => x"38",
          4203 => x"84",
          4204 => x"52",
          4205 => x"09",
          4206 => x"38",
          4207 => x"51",
          4208 => x"81",
          4209 => x"81",
          4210 => x"88",
          4211 => x"08",
          4212 => x"39",
          4213 => x"73",
          4214 => x"74",
          4215 => x"0c",
          4216 => x"04",
          4217 => x"02",
          4218 => x"7a",
          4219 => x"fc",
          4220 => x"f4",
          4221 => x"54",
          4222 => x"fe",
          4223 => x"bc",
          4224 => x"f0",
          4225 => x"81",
          4226 => x"70",
          4227 => x"73",
          4228 => x"38",
          4229 => x"78",
          4230 => x"2e",
          4231 => x"74",
          4232 => x"0c",
          4233 => x"80",
          4234 => x"80",
          4235 => x"70",
          4236 => x"51",
          4237 => x"81",
          4238 => x"54",
          4239 => x"f0",
          4240 => x"0d",
          4241 => x"0d",
          4242 => x"05",
          4243 => x"33",
          4244 => x"54",
          4245 => x"84",
          4246 => x"bf",
          4247 => x"98",
          4248 => x"53",
          4249 => x"05",
          4250 => x"fa",
          4251 => x"f0",
          4252 => x"fe",
          4253 => x"a4",
          4254 => x"68",
          4255 => x"70",
          4256 => x"c6",
          4257 => x"f0",
          4258 => x"fe",
          4259 => x"38",
          4260 => x"05",
          4261 => x"2b",
          4262 => x"80",
          4263 => x"86",
          4264 => x"06",
          4265 => x"2e",
          4266 => x"74",
          4267 => x"38",
          4268 => x"09",
          4269 => x"38",
          4270 => x"f8",
          4271 => x"f0",
          4272 => x"39",
          4273 => x"33",
          4274 => x"73",
          4275 => x"77",
          4276 => x"81",
          4277 => x"73",
          4278 => x"38",
          4279 => x"bc",
          4280 => x"07",
          4281 => x"b4",
          4282 => x"2a",
          4283 => x"51",
          4284 => x"2e",
          4285 => x"62",
          4286 => x"e8",
          4287 => x"fe",
          4288 => x"82",
          4289 => x"52",
          4290 => x"51",
          4291 => x"62",
          4292 => x"8b",
          4293 => x"53",
          4294 => x"51",
          4295 => x"80",
          4296 => x"05",
          4297 => x"3f",
          4298 => x"0b",
          4299 => x"75",
          4300 => x"f1",
          4301 => x"11",
          4302 => x"80",
          4303 => x"97",
          4304 => x"51",
          4305 => x"81",
          4306 => x"55",
          4307 => x"08",
          4308 => x"b7",
          4309 => x"c4",
          4310 => x"05",
          4311 => x"2a",
          4312 => x"51",
          4313 => x"80",
          4314 => x"84",
          4315 => x"39",
          4316 => x"70",
          4317 => x"54",
          4318 => x"a9",
          4319 => x"06",
          4320 => x"2e",
          4321 => x"55",
          4322 => x"73",
          4323 => x"d6",
          4324 => x"fe",
          4325 => x"ff",
          4326 => x"0c",
          4327 => x"fe",
          4328 => x"f8",
          4329 => x"2a",
          4330 => x"51",
          4331 => x"2e",
          4332 => x"80",
          4333 => x"7a",
          4334 => x"a0",
          4335 => x"a4",
          4336 => x"53",
          4337 => x"e6",
          4338 => x"fe",
          4339 => x"fe",
          4340 => x"1b",
          4341 => x"05",
          4342 => x"d3",
          4343 => x"f0",
          4344 => x"f0",
          4345 => x"0c",
          4346 => x"56",
          4347 => x"84",
          4348 => x"90",
          4349 => x"0b",
          4350 => x"80",
          4351 => x"0c",
          4352 => x"1a",
          4353 => x"2a",
          4354 => x"51",
          4355 => x"2e",
          4356 => x"81",
          4357 => x"80",
          4358 => x"38",
          4359 => x"08",
          4360 => x"8a",
          4361 => x"89",
          4362 => x"59",
          4363 => x"76",
          4364 => x"d7",
          4365 => x"fe",
          4366 => x"81",
          4367 => x"81",
          4368 => x"82",
          4369 => x"f0",
          4370 => x"09",
          4371 => x"38",
          4372 => x"78",
          4373 => x"30",
          4374 => x"80",
          4375 => x"77",
          4376 => x"38",
          4377 => x"06",
          4378 => x"c3",
          4379 => x"1a",
          4380 => x"38",
          4381 => x"06",
          4382 => x"2e",
          4383 => x"52",
          4384 => x"a6",
          4385 => x"f0",
          4386 => x"82",
          4387 => x"75",
          4388 => x"fe",
          4389 => x"9c",
          4390 => x"39",
          4391 => x"74",
          4392 => x"fe",
          4393 => x"3d",
          4394 => x"3d",
          4395 => x"65",
          4396 => x"5d",
          4397 => x"0c",
          4398 => x"05",
          4399 => x"f9",
          4400 => x"fe",
          4401 => x"81",
          4402 => x"8a",
          4403 => x"33",
          4404 => x"2e",
          4405 => x"56",
          4406 => x"90",
          4407 => x"06",
          4408 => x"74",
          4409 => x"b6",
          4410 => x"82",
          4411 => x"34",
          4412 => x"aa",
          4413 => x"91",
          4414 => x"56",
          4415 => x"8c",
          4416 => x"1a",
          4417 => x"74",
          4418 => x"38",
          4419 => x"80",
          4420 => x"38",
          4421 => x"70",
          4422 => x"56",
          4423 => x"b2",
          4424 => x"11",
          4425 => x"77",
          4426 => x"5b",
          4427 => x"38",
          4428 => x"88",
          4429 => x"8f",
          4430 => x"08",
          4431 => x"d5",
          4432 => x"fe",
          4433 => x"81",
          4434 => x"9f",
          4435 => x"2e",
          4436 => x"74",
          4437 => x"98",
          4438 => x"7e",
          4439 => x"3f",
          4440 => x"08",
          4441 => x"83",
          4442 => x"f0",
          4443 => x"89",
          4444 => x"77",
          4445 => x"d6",
          4446 => x"7f",
          4447 => x"58",
          4448 => x"75",
          4449 => x"75",
          4450 => x"77",
          4451 => x"7c",
          4452 => x"33",
          4453 => x"3f",
          4454 => x"08",
          4455 => x"7e",
          4456 => x"56",
          4457 => x"2e",
          4458 => x"16",
          4459 => x"55",
          4460 => x"94",
          4461 => x"53",
          4462 => x"b0",
          4463 => x"31",
          4464 => x"05",
          4465 => x"3f",
          4466 => x"56",
          4467 => x"9c",
          4468 => x"19",
          4469 => x"06",
          4470 => x"31",
          4471 => x"76",
          4472 => x"7b",
          4473 => x"08",
          4474 => x"d1",
          4475 => x"fe",
          4476 => x"81",
          4477 => x"94",
          4478 => x"ff",
          4479 => x"05",
          4480 => x"cf",
          4481 => x"76",
          4482 => x"17",
          4483 => x"1e",
          4484 => x"18",
          4485 => x"5e",
          4486 => x"39",
          4487 => x"81",
          4488 => x"90",
          4489 => x"f2",
          4490 => x"63",
          4491 => x"40",
          4492 => x"7e",
          4493 => x"fc",
          4494 => x"51",
          4495 => x"81",
          4496 => x"55",
          4497 => x"08",
          4498 => x"18",
          4499 => x"80",
          4500 => x"74",
          4501 => x"39",
          4502 => x"70",
          4503 => x"81",
          4504 => x"56",
          4505 => x"80",
          4506 => x"38",
          4507 => x"0b",
          4508 => x"82",
          4509 => x"39",
          4510 => x"19",
          4511 => x"83",
          4512 => x"18",
          4513 => x"56",
          4514 => x"27",
          4515 => x"09",
          4516 => x"2e",
          4517 => x"94",
          4518 => x"83",
          4519 => x"56",
          4520 => x"38",
          4521 => x"22",
          4522 => x"89",
          4523 => x"55",
          4524 => x"75",
          4525 => x"18",
          4526 => x"9c",
          4527 => x"85",
          4528 => x"08",
          4529 => x"d7",
          4530 => x"fe",
          4531 => x"81",
          4532 => x"80",
          4533 => x"38",
          4534 => x"ff",
          4535 => x"ff",
          4536 => x"38",
          4537 => x"0c",
          4538 => x"85",
          4539 => x"19",
          4540 => x"b0",
          4541 => x"19",
          4542 => x"81",
          4543 => x"74",
          4544 => x"3f",
          4545 => x"08",
          4546 => x"98",
          4547 => x"7e",
          4548 => x"3f",
          4549 => x"08",
          4550 => x"d2",
          4551 => x"f0",
          4552 => x"89",
          4553 => x"78",
          4554 => x"d5",
          4555 => x"7f",
          4556 => x"58",
          4557 => x"75",
          4558 => x"75",
          4559 => x"78",
          4560 => x"7c",
          4561 => x"33",
          4562 => x"3f",
          4563 => x"08",
          4564 => x"7e",
          4565 => x"78",
          4566 => x"74",
          4567 => x"38",
          4568 => x"b0",
          4569 => x"31",
          4570 => x"05",
          4571 => x"51",
          4572 => x"7e",
          4573 => x"83",
          4574 => x"89",
          4575 => x"db",
          4576 => x"08",
          4577 => x"26",
          4578 => x"51",
          4579 => x"81",
          4580 => x"fd",
          4581 => x"77",
          4582 => x"55",
          4583 => x"0c",
          4584 => x"83",
          4585 => x"80",
          4586 => x"55",
          4587 => x"83",
          4588 => x"9c",
          4589 => x"7e",
          4590 => x"3f",
          4591 => x"08",
          4592 => x"75",
          4593 => x"94",
          4594 => x"ff",
          4595 => x"05",
          4596 => x"3f",
          4597 => x"0b",
          4598 => x"7b",
          4599 => x"08",
          4600 => x"76",
          4601 => x"08",
          4602 => x"1c",
          4603 => x"08",
          4604 => x"5c",
          4605 => x"83",
          4606 => x"74",
          4607 => x"fd",
          4608 => x"18",
          4609 => x"07",
          4610 => x"19",
          4611 => x"75",
          4612 => x"0c",
          4613 => x"04",
          4614 => x"7a",
          4615 => x"05",
          4616 => x"56",
          4617 => x"81",
          4618 => x"57",
          4619 => x"08",
          4620 => x"90",
          4621 => x"86",
          4622 => x"06",
          4623 => x"73",
          4624 => x"e9",
          4625 => x"08",
          4626 => x"cc",
          4627 => x"fe",
          4628 => x"81",
          4629 => x"80",
          4630 => x"16",
          4631 => x"33",
          4632 => x"55",
          4633 => x"34",
          4634 => x"53",
          4635 => x"08",
          4636 => x"3f",
          4637 => x"52",
          4638 => x"c9",
          4639 => x"88",
          4640 => x"96",
          4641 => x"f0",
          4642 => x"92",
          4643 => x"ca",
          4644 => x"81",
          4645 => x"34",
          4646 => x"df",
          4647 => x"f0",
          4648 => x"33",
          4649 => x"55",
          4650 => x"17",
          4651 => x"fe",
          4652 => x"3d",
          4653 => x"3d",
          4654 => x"52",
          4655 => x"3f",
          4656 => x"08",
          4657 => x"f0",
          4658 => x"86",
          4659 => x"52",
          4660 => x"bc",
          4661 => x"f0",
          4662 => x"fe",
          4663 => x"38",
          4664 => x"08",
          4665 => x"81",
          4666 => x"86",
          4667 => x"ff",
          4668 => x"3d",
          4669 => x"3f",
          4670 => x"0b",
          4671 => x"08",
          4672 => x"81",
          4673 => x"81",
          4674 => x"80",
          4675 => x"fe",
          4676 => x"3d",
          4677 => x"3d",
          4678 => x"93",
          4679 => x"52",
          4680 => x"e9",
          4681 => x"fe",
          4682 => x"81",
          4683 => x"80",
          4684 => x"58",
          4685 => x"3d",
          4686 => x"e0",
          4687 => x"fe",
          4688 => x"81",
          4689 => x"bc",
          4690 => x"c7",
          4691 => x"98",
          4692 => x"73",
          4693 => x"38",
          4694 => x"12",
          4695 => x"39",
          4696 => x"33",
          4697 => x"70",
          4698 => x"55",
          4699 => x"2e",
          4700 => x"7f",
          4701 => x"54",
          4702 => x"81",
          4703 => x"94",
          4704 => x"39",
          4705 => x"08",
          4706 => x"81",
          4707 => x"85",
          4708 => x"fe",
          4709 => x"3d",
          4710 => x"3d",
          4711 => x"5b",
          4712 => x"34",
          4713 => x"3d",
          4714 => x"52",
          4715 => x"e8",
          4716 => x"fe",
          4717 => x"81",
          4718 => x"82",
          4719 => x"43",
          4720 => x"11",
          4721 => x"58",
          4722 => x"80",
          4723 => x"38",
          4724 => x"3d",
          4725 => x"d5",
          4726 => x"fe",
          4727 => x"81",
          4728 => x"82",
          4729 => x"52",
          4730 => x"c8",
          4731 => x"f0",
          4732 => x"fe",
          4733 => x"c1",
          4734 => x"7b",
          4735 => x"3f",
          4736 => x"08",
          4737 => x"74",
          4738 => x"3f",
          4739 => x"08",
          4740 => x"f0",
          4741 => x"38",
          4742 => x"51",
          4743 => x"81",
          4744 => x"57",
          4745 => x"08",
          4746 => x"52",
          4747 => x"f2",
          4748 => x"fe",
          4749 => x"a6",
          4750 => x"74",
          4751 => x"3f",
          4752 => x"08",
          4753 => x"f0",
          4754 => x"cc",
          4755 => x"2e",
          4756 => x"86",
          4757 => x"81",
          4758 => x"81",
          4759 => x"3d",
          4760 => x"52",
          4761 => x"c9",
          4762 => x"3d",
          4763 => x"11",
          4764 => x"5a",
          4765 => x"2e",
          4766 => x"b9",
          4767 => x"16",
          4768 => x"33",
          4769 => x"73",
          4770 => x"16",
          4771 => x"26",
          4772 => x"75",
          4773 => x"38",
          4774 => x"05",
          4775 => x"6f",
          4776 => x"ff",
          4777 => x"55",
          4778 => x"74",
          4779 => x"38",
          4780 => x"11",
          4781 => x"74",
          4782 => x"39",
          4783 => x"09",
          4784 => x"38",
          4785 => x"11",
          4786 => x"74",
          4787 => x"81",
          4788 => x"70",
          4789 => x"eb",
          4790 => x"08",
          4791 => x"5c",
          4792 => x"73",
          4793 => x"38",
          4794 => x"1a",
          4795 => x"55",
          4796 => x"38",
          4797 => x"73",
          4798 => x"38",
          4799 => x"76",
          4800 => x"74",
          4801 => x"33",
          4802 => x"05",
          4803 => x"15",
          4804 => x"ba",
          4805 => x"05",
          4806 => x"ff",
          4807 => x"06",
          4808 => x"57",
          4809 => x"18",
          4810 => x"54",
          4811 => x"70",
          4812 => x"34",
          4813 => x"ee",
          4814 => x"34",
          4815 => x"f0",
          4816 => x"0d",
          4817 => x"0d",
          4818 => x"3d",
          4819 => x"71",
          4820 => x"ec",
          4821 => x"fe",
          4822 => x"81",
          4823 => x"82",
          4824 => x"15",
          4825 => x"82",
          4826 => x"15",
          4827 => x"76",
          4828 => x"90",
          4829 => x"81",
          4830 => x"06",
          4831 => x"72",
          4832 => x"56",
          4833 => x"54",
          4834 => x"17",
          4835 => x"78",
          4836 => x"38",
          4837 => x"22",
          4838 => x"59",
          4839 => x"78",
          4840 => x"76",
          4841 => x"51",
          4842 => x"3f",
          4843 => x"08",
          4844 => x"54",
          4845 => x"53",
          4846 => x"3f",
          4847 => x"08",
          4848 => x"38",
          4849 => x"75",
          4850 => x"18",
          4851 => x"31",
          4852 => x"57",
          4853 => x"b1",
          4854 => x"08",
          4855 => x"38",
          4856 => x"51",
          4857 => x"81",
          4858 => x"54",
          4859 => x"08",
          4860 => x"9a",
          4861 => x"f0",
          4862 => x"81",
          4863 => x"fe",
          4864 => x"16",
          4865 => x"16",
          4866 => x"2e",
          4867 => x"76",
          4868 => x"dc",
          4869 => x"31",
          4870 => x"18",
          4871 => x"90",
          4872 => x"81",
          4873 => x"06",
          4874 => x"56",
          4875 => x"9a",
          4876 => x"74",
          4877 => x"3f",
          4878 => x"08",
          4879 => x"f0",
          4880 => x"81",
          4881 => x"56",
          4882 => x"52",
          4883 => x"84",
          4884 => x"f0",
          4885 => x"ff",
          4886 => x"81",
          4887 => x"38",
          4888 => x"98",
          4889 => x"a6",
          4890 => x"16",
          4891 => x"39",
          4892 => x"16",
          4893 => x"75",
          4894 => x"53",
          4895 => x"aa",
          4896 => x"79",
          4897 => x"3f",
          4898 => x"08",
          4899 => x"0b",
          4900 => x"82",
          4901 => x"39",
          4902 => x"16",
          4903 => x"bb",
          4904 => x"2a",
          4905 => x"08",
          4906 => x"15",
          4907 => x"15",
          4908 => x"90",
          4909 => x"16",
          4910 => x"33",
          4911 => x"53",
          4912 => x"34",
          4913 => x"06",
          4914 => x"2e",
          4915 => x"9c",
          4916 => x"85",
          4917 => x"16",
          4918 => x"72",
          4919 => x"0c",
          4920 => x"04",
          4921 => x"79",
          4922 => x"75",
          4923 => x"8a",
          4924 => x"89",
          4925 => x"52",
          4926 => x"05",
          4927 => x"3f",
          4928 => x"08",
          4929 => x"f0",
          4930 => x"38",
          4931 => x"7a",
          4932 => x"d8",
          4933 => x"fe",
          4934 => x"81",
          4935 => x"80",
          4936 => x"16",
          4937 => x"2b",
          4938 => x"74",
          4939 => x"86",
          4940 => x"84",
          4941 => x"06",
          4942 => x"73",
          4943 => x"38",
          4944 => x"52",
          4945 => x"da",
          4946 => x"f0",
          4947 => x"0c",
          4948 => x"14",
          4949 => x"23",
          4950 => x"51",
          4951 => x"81",
          4952 => x"55",
          4953 => x"09",
          4954 => x"38",
          4955 => x"39",
          4956 => x"84",
          4957 => x"0c",
          4958 => x"81",
          4959 => x"89",
          4960 => x"fc",
          4961 => x"87",
          4962 => x"53",
          4963 => x"e7",
          4964 => x"fe",
          4965 => x"38",
          4966 => x"08",
          4967 => x"3d",
          4968 => x"3d",
          4969 => x"89",
          4970 => x"54",
          4971 => x"54",
          4972 => x"81",
          4973 => x"53",
          4974 => x"08",
          4975 => x"74",
          4976 => x"fe",
          4977 => x"73",
          4978 => x"3f",
          4979 => x"08",
          4980 => x"39",
          4981 => x"08",
          4982 => x"d3",
          4983 => x"fe",
          4984 => x"81",
          4985 => x"84",
          4986 => x"06",
          4987 => x"53",
          4988 => x"fe",
          4989 => x"38",
          4990 => x"51",
          4991 => x"72",
          4992 => x"cf",
          4993 => x"fe",
          4994 => x"32",
          4995 => x"72",
          4996 => x"70",
          4997 => x"08",
          4998 => x"54",
          4999 => x"fe",
          5000 => x"3d",
          5001 => x"3d",
          5002 => x"80",
          5003 => x"70",
          5004 => x"52",
          5005 => x"3f",
          5006 => x"08",
          5007 => x"f0",
          5008 => x"64",
          5009 => x"d6",
          5010 => x"fe",
          5011 => x"81",
          5012 => x"a0",
          5013 => x"cb",
          5014 => x"98",
          5015 => x"73",
          5016 => x"38",
          5017 => x"39",
          5018 => x"88",
          5019 => x"75",
          5020 => x"3f",
          5021 => x"f0",
          5022 => x"0d",
          5023 => x"0d",
          5024 => x"5c",
          5025 => x"3d",
          5026 => x"93",
          5027 => x"d6",
          5028 => x"f0",
          5029 => x"fe",
          5030 => x"80",
          5031 => x"0c",
          5032 => x"11",
          5033 => x"90",
          5034 => x"56",
          5035 => x"74",
          5036 => x"75",
          5037 => x"e4",
          5038 => x"81",
          5039 => x"5b",
          5040 => x"81",
          5041 => x"75",
          5042 => x"73",
          5043 => x"81",
          5044 => x"82",
          5045 => x"76",
          5046 => x"f0",
          5047 => x"f4",
          5048 => x"f0",
          5049 => x"d1",
          5050 => x"f0",
          5051 => x"ce",
          5052 => x"f0",
          5053 => x"81",
          5054 => x"07",
          5055 => x"05",
          5056 => x"53",
          5057 => x"98",
          5058 => x"26",
          5059 => x"f9",
          5060 => x"08",
          5061 => x"08",
          5062 => x"98",
          5063 => x"81",
          5064 => x"58",
          5065 => x"3f",
          5066 => x"08",
          5067 => x"f0",
          5068 => x"38",
          5069 => x"77",
          5070 => x"5d",
          5071 => x"74",
          5072 => x"81",
          5073 => x"b4",
          5074 => x"bb",
          5075 => x"fe",
          5076 => x"ff",
          5077 => x"30",
          5078 => x"1b",
          5079 => x"5b",
          5080 => x"39",
          5081 => x"ff",
          5082 => x"81",
          5083 => x"f0",
          5084 => x"30",
          5085 => x"1b",
          5086 => x"5b",
          5087 => x"83",
          5088 => x"58",
          5089 => x"92",
          5090 => x"0c",
          5091 => x"12",
          5092 => x"33",
          5093 => x"54",
          5094 => x"34",
          5095 => x"f0",
          5096 => x"0d",
          5097 => x"0d",
          5098 => x"fc",
          5099 => x"52",
          5100 => x"3f",
          5101 => x"08",
          5102 => x"f0",
          5103 => x"38",
          5104 => x"56",
          5105 => x"38",
          5106 => x"70",
          5107 => x"81",
          5108 => x"55",
          5109 => x"80",
          5110 => x"38",
          5111 => x"54",
          5112 => x"08",
          5113 => x"38",
          5114 => x"81",
          5115 => x"53",
          5116 => x"52",
          5117 => x"8c",
          5118 => x"f0",
          5119 => x"19",
          5120 => x"c9",
          5121 => x"08",
          5122 => x"ff",
          5123 => x"81",
          5124 => x"ff",
          5125 => x"06",
          5126 => x"56",
          5127 => x"08",
          5128 => x"81",
          5129 => x"82",
          5130 => x"75",
          5131 => x"54",
          5132 => x"08",
          5133 => x"27",
          5134 => x"17",
          5135 => x"fe",
          5136 => x"76",
          5137 => x"3f",
          5138 => x"08",
          5139 => x"08",
          5140 => x"90",
          5141 => x"c0",
          5142 => x"90",
          5143 => x"80",
          5144 => x"75",
          5145 => x"75",
          5146 => x"fe",
          5147 => x"3d",
          5148 => x"3d",
          5149 => x"a0",
          5150 => x"05",
          5151 => x"51",
          5152 => x"81",
          5153 => x"55",
          5154 => x"08",
          5155 => x"78",
          5156 => x"08",
          5157 => x"70",
          5158 => x"ae",
          5159 => x"f0",
          5160 => x"fe",
          5161 => x"db",
          5162 => x"fb",
          5163 => x"85",
          5164 => x"06",
          5165 => x"86",
          5166 => x"c7",
          5167 => x"2b",
          5168 => x"24",
          5169 => x"02",
          5170 => x"33",
          5171 => x"58",
          5172 => x"76",
          5173 => x"6b",
          5174 => x"cc",
          5175 => x"fe",
          5176 => x"84",
          5177 => x"06",
          5178 => x"73",
          5179 => x"d4",
          5180 => x"81",
          5181 => x"94",
          5182 => x"81",
          5183 => x"5a",
          5184 => x"08",
          5185 => x"8a",
          5186 => x"54",
          5187 => x"81",
          5188 => x"55",
          5189 => x"08",
          5190 => x"81",
          5191 => x"52",
          5192 => x"e5",
          5193 => x"f0",
          5194 => x"fe",
          5195 => x"38",
          5196 => x"cf",
          5197 => x"f0",
          5198 => x"88",
          5199 => x"f0",
          5200 => x"38",
          5201 => x"c2",
          5202 => x"f0",
          5203 => x"f0",
          5204 => x"81",
          5205 => x"07",
          5206 => x"55",
          5207 => x"2e",
          5208 => x"80",
          5209 => x"80",
          5210 => x"77",
          5211 => x"3f",
          5212 => x"08",
          5213 => x"38",
          5214 => x"ba",
          5215 => x"fe",
          5216 => x"74",
          5217 => x"0c",
          5218 => x"04",
          5219 => x"82",
          5220 => x"c0",
          5221 => x"3d",
          5222 => x"3f",
          5223 => x"08",
          5224 => x"f0",
          5225 => x"38",
          5226 => x"52",
          5227 => x"52",
          5228 => x"3f",
          5229 => x"08",
          5230 => x"f0",
          5231 => x"88",
          5232 => x"39",
          5233 => x"08",
          5234 => x"81",
          5235 => x"38",
          5236 => x"05",
          5237 => x"2a",
          5238 => x"55",
          5239 => x"81",
          5240 => x"5a",
          5241 => x"3d",
          5242 => x"c1",
          5243 => x"fe",
          5244 => x"55",
          5245 => x"f0",
          5246 => x"87",
          5247 => x"f0",
          5248 => x"09",
          5249 => x"38",
          5250 => x"fe",
          5251 => x"2e",
          5252 => x"86",
          5253 => x"81",
          5254 => x"81",
          5255 => x"fe",
          5256 => x"78",
          5257 => x"3f",
          5258 => x"08",
          5259 => x"f0",
          5260 => x"38",
          5261 => x"52",
          5262 => x"ff",
          5263 => x"78",
          5264 => x"b4",
          5265 => x"54",
          5266 => x"15",
          5267 => x"b2",
          5268 => x"ca",
          5269 => x"b6",
          5270 => x"53",
          5271 => x"53",
          5272 => x"3f",
          5273 => x"b4",
          5274 => x"d4",
          5275 => x"b6",
          5276 => x"54",
          5277 => x"d5",
          5278 => x"53",
          5279 => x"11",
          5280 => x"d7",
          5281 => x"81",
          5282 => x"34",
          5283 => x"a4",
          5284 => x"f0",
          5285 => x"fe",
          5286 => x"38",
          5287 => x"0a",
          5288 => x"05",
          5289 => x"d0",
          5290 => x"64",
          5291 => x"c9",
          5292 => x"54",
          5293 => x"15",
          5294 => x"81",
          5295 => x"34",
          5296 => x"b8",
          5297 => x"fe",
          5298 => x"8b",
          5299 => x"75",
          5300 => x"ff",
          5301 => x"73",
          5302 => x"0c",
          5303 => x"04",
          5304 => x"a9",
          5305 => x"51",
          5306 => x"82",
          5307 => x"ff",
          5308 => x"a9",
          5309 => x"ee",
          5310 => x"f0",
          5311 => x"fe",
          5312 => x"d3",
          5313 => x"a9",
          5314 => x"9d",
          5315 => x"58",
          5316 => x"81",
          5317 => x"55",
          5318 => x"08",
          5319 => x"02",
          5320 => x"33",
          5321 => x"54",
          5322 => x"82",
          5323 => x"53",
          5324 => x"52",
          5325 => x"88",
          5326 => x"b4",
          5327 => x"53",
          5328 => x"3d",
          5329 => x"ff",
          5330 => x"aa",
          5331 => x"73",
          5332 => x"3f",
          5333 => x"08",
          5334 => x"f0",
          5335 => x"63",
          5336 => x"81",
          5337 => x"65",
          5338 => x"2e",
          5339 => x"55",
          5340 => x"81",
          5341 => x"84",
          5342 => x"06",
          5343 => x"73",
          5344 => x"3f",
          5345 => x"08",
          5346 => x"f0",
          5347 => x"38",
          5348 => x"53",
          5349 => x"95",
          5350 => x"16",
          5351 => x"87",
          5352 => x"05",
          5353 => x"34",
          5354 => x"70",
          5355 => x"81",
          5356 => x"55",
          5357 => x"74",
          5358 => x"73",
          5359 => x"78",
          5360 => x"83",
          5361 => x"16",
          5362 => x"2a",
          5363 => x"51",
          5364 => x"80",
          5365 => x"38",
          5366 => x"80",
          5367 => x"52",
          5368 => x"be",
          5369 => x"f0",
          5370 => x"51",
          5371 => x"3f",
          5372 => x"fe",
          5373 => x"2e",
          5374 => x"81",
          5375 => x"52",
          5376 => x"b5",
          5377 => x"fe",
          5378 => x"80",
          5379 => x"58",
          5380 => x"f0",
          5381 => x"38",
          5382 => x"54",
          5383 => x"09",
          5384 => x"38",
          5385 => x"52",
          5386 => x"af",
          5387 => x"81",
          5388 => x"34",
          5389 => x"fe",
          5390 => x"38",
          5391 => x"ca",
          5392 => x"f0",
          5393 => x"fe",
          5394 => x"38",
          5395 => x"b5",
          5396 => x"fe",
          5397 => x"74",
          5398 => x"0c",
          5399 => x"04",
          5400 => x"02",
          5401 => x"33",
          5402 => x"80",
          5403 => x"57",
          5404 => x"95",
          5405 => x"52",
          5406 => x"d2",
          5407 => x"fe",
          5408 => x"81",
          5409 => x"80",
          5410 => x"5a",
          5411 => x"3d",
          5412 => x"c9",
          5413 => x"fe",
          5414 => x"81",
          5415 => x"b8",
          5416 => x"cf",
          5417 => x"a0",
          5418 => x"55",
          5419 => x"75",
          5420 => x"71",
          5421 => x"33",
          5422 => x"74",
          5423 => x"57",
          5424 => x"8b",
          5425 => x"54",
          5426 => x"15",
          5427 => x"ff",
          5428 => x"81",
          5429 => x"55",
          5430 => x"f0",
          5431 => x"0d",
          5432 => x"0d",
          5433 => x"53",
          5434 => x"05",
          5435 => x"51",
          5436 => x"81",
          5437 => x"55",
          5438 => x"08",
          5439 => x"76",
          5440 => x"93",
          5441 => x"51",
          5442 => x"81",
          5443 => x"55",
          5444 => x"08",
          5445 => x"80",
          5446 => x"81",
          5447 => x"86",
          5448 => x"38",
          5449 => x"86",
          5450 => x"90",
          5451 => x"54",
          5452 => x"ff",
          5453 => x"76",
          5454 => x"83",
          5455 => x"51",
          5456 => x"3f",
          5457 => x"08",
          5458 => x"fe",
          5459 => x"3d",
          5460 => x"3d",
          5461 => x"5c",
          5462 => x"98",
          5463 => x"52",
          5464 => x"d1",
          5465 => x"fe",
          5466 => x"fe",
          5467 => x"70",
          5468 => x"08",
          5469 => x"51",
          5470 => x"80",
          5471 => x"38",
          5472 => x"06",
          5473 => x"80",
          5474 => x"38",
          5475 => x"5f",
          5476 => x"3d",
          5477 => x"ff",
          5478 => x"81",
          5479 => x"57",
          5480 => x"08",
          5481 => x"74",
          5482 => x"c3",
          5483 => x"fe",
          5484 => x"81",
          5485 => x"bf",
          5486 => x"f0",
          5487 => x"f0",
          5488 => x"59",
          5489 => x"81",
          5490 => x"56",
          5491 => x"33",
          5492 => x"16",
          5493 => x"27",
          5494 => x"56",
          5495 => x"80",
          5496 => x"80",
          5497 => x"ff",
          5498 => x"70",
          5499 => x"56",
          5500 => x"e8",
          5501 => x"76",
          5502 => x"81",
          5503 => x"80",
          5504 => x"57",
          5505 => x"78",
          5506 => x"51",
          5507 => x"2e",
          5508 => x"73",
          5509 => x"38",
          5510 => x"08",
          5511 => x"b1",
          5512 => x"fe",
          5513 => x"81",
          5514 => x"a7",
          5515 => x"33",
          5516 => x"c3",
          5517 => x"2e",
          5518 => x"e4",
          5519 => x"2e",
          5520 => x"56",
          5521 => x"05",
          5522 => x"e3",
          5523 => x"f0",
          5524 => x"76",
          5525 => x"0c",
          5526 => x"04",
          5527 => x"82",
          5528 => x"ff",
          5529 => x"9d",
          5530 => x"fa",
          5531 => x"f0",
          5532 => x"f0",
          5533 => x"81",
          5534 => x"83",
          5535 => x"53",
          5536 => x"3d",
          5537 => x"ff",
          5538 => x"73",
          5539 => x"70",
          5540 => x"52",
          5541 => x"9f",
          5542 => x"bc",
          5543 => x"74",
          5544 => x"6d",
          5545 => x"70",
          5546 => x"af",
          5547 => x"fe",
          5548 => x"2e",
          5549 => x"70",
          5550 => x"57",
          5551 => x"fd",
          5552 => x"f0",
          5553 => x"8d",
          5554 => x"2b",
          5555 => x"81",
          5556 => x"86",
          5557 => x"f0",
          5558 => x"9f",
          5559 => x"ff",
          5560 => x"54",
          5561 => x"8a",
          5562 => x"70",
          5563 => x"06",
          5564 => x"ff",
          5565 => x"38",
          5566 => x"15",
          5567 => x"80",
          5568 => x"74",
          5569 => x"dc",
          5570 => x"89",
          5571 => x"f0",
          5572 => x"81",
          5573 => x"88",
          5574 => x"26",
          5575 => x"39",
          5576 => x"86",
          5577 => x"81",
          5578 => x"ff",
          5579 => x"38",
          5580 => x"54",
          5581 => x"81",
          5582 => x"81",
          5583 => x"78",
          5584 => x"5a",
          5585 => x"6d",
          5586 => x"81",
          5587 => x"57",
          5588 => x"9f",
          5589 => x"38",
          5590 => x"54",
          5591 => x"81",
          5592 => x"b1",
          5593 => x"2e",
          5594 => x"a7",
          5595 => x"15",
          5596 => x"54",
          5597 => x"09",
          5598 => x"38",
          5599 => x"76",
          5600 => x"41",
          5601 => x"52",
          5602 => x"52",
          5603 => x"b3",
          5604 => x"f0",
          5605 => x"fe",
          5606 => x"f7",
          5607 => x"74",
          5608 => x"e5",
          5609 => x"f0",
          5610 => x"fe",
          5611 => x"38",
          5612 => x"38",
          5613 => x"74",
          5614 => x"39",
          5615 => x"08",
          5616 => x"81",
          5617 => x"38",
          5618 => x"74",
          5619 => x"38",
          5620 => x"51",
          5621 => x"3f",
          5622 => x"08",
          5623 => x"f0",
          5624 => x"a0",
          5625 => x"f0",
          5626 => x"51",
          5627 => x"3f",
          5628 => x"0b",
          5629 => x"8b",
          5630 => x"67",
          5631 => x"a7",
          5632 => x"81",
          5633 => x"34",
          5634 => x"ad",
          5635 => x"fe",
          5636 => x"73",
          5637 => x"fe",
          5638 => x"3d",
          5639 => x"3d",
          5640 => x"02",
          5641 => x"cb",
          5642 => x"3d",
          5643 => x"72",
          5644 => x"5a",
          5645 => x"81",
          5646 => x"58",
          5647 => x"08",
          5648 => x"91",
          5649 => x"77",
          5650 => x"7c",
          5651 => x"38",
          5652 => x"59",
          5653 => x"90",
          5654 => x"81",
          5655 => x"06",
          5656 => x"73",
          5657 => x"54",
          5658 => x"82",
          5659 => x"39",
          5660 => x"8b",
          5661 => x"11",
          5662 => x"2b",
          5663 => x"54",
          5664 => x"fe",
          5665 => x"ff",
          5666 => x"70",
          5667 => x"07",
          5668 => x"fe",
          5669 => x"8c",
          5670 => x"40",
          5671 => x"55",
          5672 => x"88",
          5673 => x"08",
          5674 => x"38",
          5675 => x"77",
          5676 => x"56",
          5677 => x"51",
          5678 => x"3f",
          5679 => x"55",
          5680 => x"08",
          5681 => x"38",
          5682 => x"fe",
          5683 => x"2e",
          5684 => x"81",
          5685 => x"ff",
          5686 => x"38",
          5687 => x"08",
          5688 => x"16",
          5689 => x"2e",
          5690 => x"87",
          5691 => x"74",
          5692 => x"74",
          5693 => x"81",
          5694 => x"38",
          5695 => x"ff",
          5696 => x"2e",
          5697 => x"7b",
          5698 => x"80",
          5699 => x"81",
          5700 => x"81",
          5701 => x"06",
          5702 => x"56",
          5703 => x"52",
          5704 => x"af",
          5705 => x"fe",
          5706 => x"81",
          5707 => x"80",
          5708 => x"81",
          5709 => x"56",
          5710 => x"d3",
          5711 => x"ff",
          5712 => x"7c",
          5713 => x"55",
          5714 => x"b3",
          5715 => x"1b",
          5716 => x"1b",
          5717 => x"33",
          5718 => x"54",
          5719 => x"34",
          5720 => x"fe",
          5721 => x"08",
          5722 => x"74",
          5723 => x"75",
          5724 => x"16",
          5725 => x"33",
          5726 => x"73",
          5727 => x"77",
          5728 => x"fe",
          5729 => x"3d",
          5730 => x"3d",
          5731 => x"02",
          5732 => x"eb",
          5733 => x"3d",
          5734 => x"59",
          5735 => x"8b",
          5736 => x"81",
          5737 => x"24",
          5738 => x"81",
          5739 => x"84",
          5740 => x"a0",
          5741 => x"51",
          5742 => x"2e",
          5743 => x"75",
          5744 => x"f0",
          5745 => x"06",
          5746 => x"7e",
          5747 => x"d0",
          5748 => x"f0",
          5749 => x"06",
          5750 => x"56",
          5751 => x"74",
          5752 => x"76",
          5753 => x"81",
          5754 => x"8a",
          5755 => x"b2",
          5756 => x"fc",
          5757 => x"52",
          5758 => x"a4",
          5759 => x"fe",
          5760 => x"38",
          5761 => x"80",
          5762 => x"74",
          5763 => x"26",
          5764 => x"15",
          5765 => x"74",
          5766 => x"38",
          5767 => x"80",
          5768 => x"84",
          5769 => x"92",
          5770 => x"80",
          5771 => x"38",
          5772 => x"06",
          5773 => x"2e",
          5774 => x"56",
          5775 => x"78",
          5776 => x"89",
          5777 => x"2b",
          5778 => x"43",
          5779 => x"38",
          5780 => x"30",
          5781 => x"77",
          5782 => x"91",
          5783 => x"c2",
          5784 => x"f8",
          5785 => x"52",
          5786 => x"a4",
          5787 => x"56",
          5788 => x"08",
          5789 => x"77",
          5790 => x"77",
          5791 => x"f0",
          5792 => x"45",
          5793 => x"bf",
          5794 => x"8e",
          5795 => x"26",
          5796 => x"74",
          5797 => x"48",
          5798 => x"75",
          5799 => x"38",
          5800 => x"81",
          5801 => x"fa",
          5802 => x"2a",
          5803 => x"56",
          5804 => x"2e",
          5805 => x"87",
          5806 => x"82",
          5807 => x"38",
          5808 => x"55",
          5809 => x"83",
          5810 => x"81",
          5811 => x"56",
          5812 => x"80",
          5813 => x"38",
          5814 => x"83",
          5815 => x"06",
          5816 => x"78",
          5817 => x"91",
          5818 => x"0b",
          5819 => x"22",
          5820 => x"80",
          5821 => x"74",
          5822 => x"38",
          5823 => x"56",
          5824 => x"17",
          5825 => x"57",
          5826 => x"2e",
          5827 => x"75",
          5828 => x"79",
          5829 => x"fe",
          5830 => x"81",
          5831 => x"84",
          5832 => x"05",
          5833 => x"5e",
          5834 => x"80",
          5835 => x"f0",
          5836 => x"8a",
          5837 => x"fd",
          5838 => x"75",
          5839 => x"38",
          5840 => x"78",
          5841 => x"8c",
          5842 => x"0b",
          5843 => x"22",
          5844 => x"80",
          5845 => x"74",
          5846 => x"38",
          5847 => x"56",
          5848 => x"17",
          5849 => x"57",
          5850 => x"2e",
          5851 => x"75",
          5852 => x"79",
          5853 => x"fe",
          5854 => x"81",
          5855 => x"10",
          5856 => x"81",
          5857 => x"9f",
          5858 => x"38",
          5859 => x"fe",
          5860 => x"81",
          5861 => x"05",
          5862 => x"2a",
          5863 => x"56",
          5864 => x"17",
          5865 => x"81",
          5866 => x"60",
          5867 => x"65",
          5868 => x"12",
          5869 => x"30",
          5870 => x"74",
          5871 => x"59",
          5872 => x"7d",
          5873 => x"81",
          5874 => x"76",
          5875 => x"41",
          5876 => x"76",
          5877 => x"90",
          5878 => x"62",
          5879 => x"51",
          5880 => x"26",
          5881 => x"75",
          5882 => x"31",
          5883 => x"65",
          5884 => x"fe",
          5885 => x"81",
          5886 => x"58",
          5887 => x"09",
          5888 => x"38",
          5889 => x"08",
          5890 => x"26",
          5891 => x"78",
          5892 => x"79",
          5893 => x"78",
          5894 => x"86",
          5895 => x"82",
          5896 => x"06",
          5897 => x"83",
          5898 => x"81",
          5899 => x"27",
          5900 => x"8f",
          5901 => x"55",
          5902 => x"26",
          5903 => x"59",
          5904 => x"62",
          5905 => x"74",
          5906 => x"38",
          5907 => x"88",
          5908 => x"f0",
          5909 => x"26",
          5910 => x"86",
          5911 => x"1a",
          5912 => x"79",
          5913 => x"38",
          5914 => x"80",
          5915 => x"2e",
          5916 => x"83",
          5917 => x"9f",
          5918 => x"8b",
          5919 => x"06",
          5920 => x"74",
          5921 => x"84",
          5922 => x"52",
          5923 => x"a2",
          5924 => x"53",
          5925 => x"52",
          5926 => x"a2",
          5927 => x"80",
          5928 => x"51",
          5929 => x"3f",
          5930 => x"34",
          5931 => x"ff",
          5932 => x"1b",
          5933 => x"a2",
          5934 => x"90",
          5935 => x"83",
          5936 => x"70",
          5937 => x"80",
          5938 => x"55",
          5939 => x"ff",
          5940 => x"66",
          5941 => x"ff",
          5942 => x"38",
          5943 => x"ff",
          5944 => x"1b",
          5945 => x"f2",
          5946 => x"74",
          5947 => x"51",
          5948 => x"3f",
          5949 => x"1c",
          5950 => x"98",
          5951 => x"a0",
          5952 => x"ff",
          5953 => x"51",
          5954 => x"3f",
          5955 => x"1b",
          5956 => x"e4",
          5957 => x"2e",
          5958 => x"80",
          5959 => x"88",
          5960 => x"80",
          5961 => x"ff",
          5962 => x"7c",
          5963 => x"51",
          5964 => x"3f",
          5965 => x"1b",
          5966 => x"bc",
          5967 => x"b0",
          5968 => x"a0",
          5969 => x"52",
          5970 => x"ff",
          5971 => x"ff",
          5972 => x"c0",
          5973 => x"0b",
          5974 => x"34",
          5975 => x"eb",
          5976 => x"c7",
          5977 => x"39",
          5978 => x"0a",
          5979 => x"51",
          5980 => x"3f",
          5981 => x"ff",
          5982 => x"1b",
          5983 => x"da",
          5984 => x"0b",
          5985 => x"a9",
          5986 => x"34",
          5987 => x"eb",
          5988 => x"1b",
          5989 => x"8f",
          5990 => x"d5",
          5991 => x"1b",
          5992 => x"ff",
          5993 => x"81",
          5994 => x"7a",
          5995 => x"ff",
          5996 => x"81",
          5997 => x"f0",
          5998 => x"38",
          5999 => x"09",
          6000 => x"ee",
          6001 => x"60",
          6002 => x"7a",
          6003 => x"ff",
          6004 => x"84",
          6005 => x"52",
          6006 => x"9f",
          6007 => x"8b",
          6008 => x"52",
          6009 => x"9f",
          6010 => x"8a",
          6011 => x"52",
          6012 => x"51",
          6013 => x"3f",
          6014 => x"83",
          6015 => x"ff",
          6016 => x"82",
          6017 => x"1b",
          6018 => x"ec",
          6019 => x"d5",
          6020 => x"ff",
          6021 => x"75",
          6022 => x"05",
          6023 => x"7e",
          6024 => x"e5",
          6025 => x"60",
          6026 => x"52",
          6027 => x"9a",
          6028 => x"53",
          6029 => x"51",
          6030 => x"3f",
          6031 => x"58",
          6032 => x"09",
          6033 => x"38",
          6034 => x"51",
          6035 => x"3f",
          6036 => x"1b",
          6037 => x"a0",
          6038 => x"52",
          6039 => x"91",
          6040 => x"ff",
          6041 => x"81",
          6042 => x"f8",
          6043 => x"7a",
          6044 => x"84",
          6045 => x"61",
          6046 => x"26",
          6047 => x"57",
          6048 => x"53",
          6049 => x"51",
          6050 => x"3f",
          6051 => x"08",
          6052 => x"84",
          6053 => x"fe",
          6054 => x"7a",
          6055 => x"aa",
          6056 => x"75",
          6057 => x"56",
          6058 => x"81",
          6059 => x"80",
          6060 => x"38",
          6061 => x"83",
          6062 => x"63",
          6063 => x"74",
          6064 => x"38",
          6065 => x"54",
          6066 => x"52",
          6067 => x"99",
          6068 => x"fe",
          6069 => x"c1",
          6070 => x"75",
          6071 => x"56",
          6072 => x"8c",
          6073 => x"2e",
          6074 => x"56",
          6075 => x"ff",
          6076 => x"84",
          6077 => x"2e",
          6078 => x"56",
          6079 => x"58",
          6080 => x"38",
          6081 => x"77",
          6082 => x"ff",
          6083 => x"82",
          6084 => x"78",
          6085 => x"c2",
          6086 => x"1b",
          6087 => x"34",
          6088 => x"16",
          6089 => x"82",
          6090 => x"83",
          6091 => x"84",
          6092 => x"67",
          6093 => x"fd",
          6094 => x"51",
          6095 => x"3f",
          6096 => x"16",
          6097 => x"f0",
          6098 => x"bf",
          6099 => x"86",
          6100 => x"fe",
          6101 => x"16",
          6102 => x"83",
          6103 => x"ff",
          6104 => x"66",
          6105 => x"1b",
          6106 => x"8c",
          6107 => x"77",
          6108 => x"7e",
          6109 => x"91",
          6110 => x"81",
          6111 => x"a2",
          6112 => x"80",
          6113 => x"ff",
          6114 => x"81",
          6115 => x"f0",
          6116 => x"89",
          6117 => x"8a",
          6118 => x"86",
          6119 => x"f0",
          6120 => x"81",
          6121 => x"99",
          6122 => x"f5",
          6123 => x"60",
          6124 => x"79",
          6125 => x"5a",
          6126 => x"78",
          6127 => x"8d",
          6128 => x"55",
          6129 => x"fc",
          6130 => x"51",
          6131 => x"7a",
          6132 => x"81",
          6133 => x"8c",
          6134 => x"74",
          6135 => x"38",
          6136 => x"81",
          6137 => x"81",
          6138 => x"8a",
          6139 => x"06",
          6140 => x"76",
          6141 => x"76",
          6142 => x"55",
          6143 => x"f0",
          6144 => x"0d",
          6145 => x"0d",
          6146 => x"05",
          6147 => x"59",
          6148 => x"2e",
          6149 => x"87",
          6150 => x"76",
          6151 => x"84",
          6152 => x"80",
          6153 => x"38",
          6154 => x"77",
          6155 => x"56",
          6156 => x"34",
          6157 => x"bb",
          6158 => x"38",
          6159 => x"05",
          6160 => x"8c",
          6161 => x"08",
          6162 => x"3f",
          6163 => x"70",
          6164 => x"07",
          6165 => x"30",
          6166 => x"56",
          6167 => x"0c",
          6168 => x"18",
          6169 => x"0d",
          6170 => x"0d",
          6171 => x"08",
          6172 => x"75",
          6173 => x"89",
          6174 => x"54",
          6175 => x"16",
          6176 => x"51",
          6177 => x"81",
          6178 => x"91",
          6179 => x"08",
          6180 => x"81",
          6181 => x"88",
          6182 => x"83",
          6183 => x"74",
          6184 => x"0c",
          6185 => x"04",
          6186 => x"75",
          6187 => x"53",
          6188 => x"51",
          6189 => x"3f",
          6190 => x"85",
          6191 => x"ea",
          6192 => x"80",
          6193 => x"6a",
          6194 => x"70",
          6195 => x"d8",
          6196 => x"72",
          6197 => x"3f",
          6198 => x"8d",
          6199 => x"0d",
          6200 => x"0d",
          6201 => x"70",
          6202 => x"74",
          6203 => x"e1",
          6204 => x"77",
          6205 => x"85",
          6206 => x"80",
          6207 => x"33",
          6208 => x"2e",
          6209 => x"86",
          6210 => x"55",
          6211 => x"57",
          6212 => x"81",
          6213 => x"70",
          6214 => x"fe",
          6215 => x"81",
          6216 => x"81",
          6217 => x"54",
          6218 => x"08",
          6219 => x"da",
          6220 => x"fe",
          6221 => x"38",
          6222 => x"54",
          6223 => x"ff",
          6224 => x"17",
          6225 => x"06",
          6226 => x"77",
          6227 => x"ff",
          6228 => x"fe",
          6229 => x"3d",
          6230 => x"3d",
          6231 => x"71",
          6232 => x"8e",
          6233 => x"29",
          6234 => x"05",
          6235 => x"04",
          6236 => x"51",
          6237 => x"81",
          6238 => x"80",
          6239 => x"ee",
          6240 => x"f2",
          6241 => x"ec",
          6242 => x"39",
          6243 => x"51",
          6244 => x"81",
          6245 => x"80",
          6246 => x"ef",
          6247 => x"d6",
          6248 => x"b0",
          6249 => x"39",
          6250 => x"51",
          6251 => x"81",
          6252 => x"80",
          6253 => x"ef",
          6254 => x"39",
          6255 => x"51",
          6256 => x"f0",
          6257 => x"39",
          6258 => x"51",
          6259 => x"f0",
          6260 => x"39",
          6261 => x"51",
          6262 => x"f1",
          6263 => x"39",
          6264 => x"51",
          6265 => x"f1",
          6266 => x"39",
          6267 => x"51",
          6268 => x"f1",
          6269 => x"f2",
          6270 => x"3d",
          6271 => x"3d",
          6272 => x"56",
          6273 => x"e7",
          6274 => x"74",
          6275 => x"e8",
          6276 => x"39",
          6277 => x"74",
          6278 => x"91",
          6279 => x"f0",
          6280 => x"51",
          6281 => x"3f",
          6282 => x"08",
          6283 => x"75",
          6284 => x"80",
          6285 => x"d3",
          6286 => x"0d",
          6287 => x"0d",
          6288 => x"05",
          6289 => x"33",
          6290 => x"68",
          6291 => x"7a",
          6292 => x"51",
          6293 => x"78",
          6294 => x"ff",
          6295 => x"81",
          6296 => x"07",
          6297 => x"06",
          6298 => x"56",
          6299 => x"38",
          6300 => x"52",
          6301 => x"52",
          6302 => x"c9",
          6303 => x"f0",
          6304 => x"fe",
          6305 => x"38",
          6306 => x"08",
          6307 => x"88",
          6308 => x"f0",
          6309 => x"3d",
          6310 => x"84",
          6311 => x"52",
          6312 => x"86",
          6313 => x"f0",
          6314 => x"fe",
          6315 => x"38",
          6316 => x"80",
          6317 => x"74",
          6318 => x"59",
          6319 => x"96",
          6320 => x"51",
          6321 => x"76",
          6322 => x"07",
          6323 => x"30",
          6324 => x"72",
          6325 => x"51",
          6326 => x"2e",
          6327 => x"f2",
          6328 => x"c0",
          6329 => x"52",
          6330 => x"92",
          6331 => x"75",
          6332 => x"0c",
          6333 => x"04",
          6334 => x"7b",
          6335 => x"b3",
          6336 => x"58",
          6337 => x"53",
          6338 => x"51",
          6339 => x"81",
          6340 => x"a4",
          6341 => x"2e",
          6342 => x"81",
          6343 => x"98",
          6344 => x"7f",
          6345 => x"f0",
          6346 => x"7d",
          6347 => x"81",
          6348 => x"57",
          6349 => x"04",
          6350 => x"f0",
          6351 => x"0d",
          6352 => x"0d",
          6353 => x"02",
          6354 => x"cf",
          6355 => x"73",
          6356 => x"5f",
          6357 => x"5e",
          6358 => x"81",
          6359 => x"fe",
          6360 => x"81",
          6361 => x"fe",
          6362 => x"80",
          6363 => x"27",
          6364 => x"7b",
          6365 => x"38",
          6366 => x"a7",
          6367 => x"39",
          6368 => x"72",
          6369 => x"38",
          6370 => x"81",
          6371 => x"fe",
          6372 => x"89",
          6373 => x"c4",
          6374 => x"8b",
          6375 => x"55",
          6376 => x"74",
          6377 => x"7a",
          6378 => x"72",
          6379 => x"f2",
          6380 => x"f4",
          6381 => x"39",
          6382 => x"51",
          6383 => x"3f",
          6384 => x"a1",
          6385 => x"53",
          6386 => x"8e",
          6387 => x"52",
          6388 => x"51",
          6389 => x"3f",
          6390 => x"f2",
          6391 => x"ee",
          6392 => x"15",
          6393 => x"fe",
          6394 => x"ff",
          6395 => x"f2",
          6396 => x"ee",
          6397 => x"55",
          6398 => x"bc",
          6399 => x"70",
          6400 => x"80",
          6401 => x"27",
          6402 => x"56",
          6403 => x"74",
          6404 => x"81",
          6405 => x"06",
          6406 => x"06",
          6407 => x"80",
          6408 => x"73",
          6409 => x"85",
          6410 => x"83",
          6411 => x"fe",
          6412 => x"81",
          6413 => x"39",
          6414 => x"51",
          6415 => x"3f",
          6416 => x"1c",
          6417 => x"de",
          6418 => x"fe",
          6419 => x"2b",
          6420 => x"51",
          6421 => x"2e",
          6422 => x"ab",
          6423 => x"ff",
          6424 => x"f0",
          6425 => x"70",
          6426 => x"a0",
          6427 => x"72",
          6428 => x"30",
          6429 => x"73",
          6430 => x"51",
          6431 => x"57",
          6432 => x"73",
          6433 => x"76",
          6434 => x"81",
          6435 => x"80",
          6436 => x"7c",
          6437 => x"78",
          6438 => x"38",
          6439 => x"81",
          6440 => x"8f",
          6441 => x"fc",
          6442 => x"9b",
          6443 => x"f2",
          6444 => x"f2",
          6445 => x"fe",
          6446 => x"81",
          6447 => x"51",
          6448 => x"3f",
          6449 => x"54",
          6450 => x"53",
          6451 => x"33",
          6452 => x"88",
          6453 => x"b3",
          6454 => x"2e",
          6455 => x"e2",
          6456 => x"3d",
          6457 => x"3d",
          6458 => x"96",
          6459 => x"fe",
          6460 => x"81",
          6461 => x"fb",
          6462 => x"a4",
          6463 => x"f3",
          6464 => x"fe",
          6465 => x"72",
          6466 => x"81",
          6467 => x"71",
          6468 => x"38",
          6469 => x"d8",
          6470 => x"f3",
          6471 => x"da",
          6472 => x"51",
          6473 => x"3f",
          6474 => x"70",
          6475 => x"52",
          6476 => x"95",
          6477 => x"fe",
          6478 => x"81",
          6479 => x"fe",
          6480 => x"80",
          6481 => x"ab",
          6482 => x"2a",
          6483 => x"51",
          6484 => x"2e",
          6485 => x"51",
          6486 => x"3f",
          6487 => x"51",
          6488 => x"3f",
          6489 => x"d8",
          6490 => x"84",
          6491 => x"06",
          6492 => x"80",
          6493 => x"81",
          6494 => x"f7",
          6495 => x"f8",
          6496 => x"ef",
          6497 => x"fe",
          6498 => x"72",
          6499 => x"81",
          6500 => x"71",
          6501 => x"38",
          6502 => x"d7",
          6503 => x"f4",
          6504 => x"d9",
          6505 => x"51",
          6506 => x"3f",
          6507 => x"70",
          6508 => x"52",
          6509 => x"95",
          6510 => x"fe",
          6511 => x"81",
          6512 => x"fe",
          6513 => x"80",
          6514 => x"a7",
          6515 => x"2a",
          6516 => x"51",
          6517 => x"2e",
          6518 => x"51",
          6519 => x"3f",
          6520 => x"51",
          6521 => x"3f",
          6522 => x"d7",
          6523 => x"88",
          6524 => x"06",
          6525 => x"80",
          6526 => x"81",
          6527 => x"f3",
          6528 => x"c8",
          6529 => x"eb",
          6530 => x"fe",
          6531 => x"fe",
          6532 => x"84",
          6533 => x"fb",
          6534 => x"02",
          6535 => x"05",
          6536 => x"56",
          6537 => x"75",
          6538 => x"a3",
          6539 => x"dc",
          6540 => x"a7",
          6541 => x"81",
          6542 => x"82",
          6543 => x"ff",
          6544 => x"81",
          6545 => x"30",
          6546 => x"f0",
          6547 => x"25",
          6548 => x"51",
          6549 => x"81",
          6550 => x"81",
          6551 => x"54",
          6552 => x"09",
          6553 => x"38",
          6554 => x"53",
          6555 => x"51",
          6556 => x"81",
          6557 => x"80",
          6558 => x"81",
          6559 => x"51",
          6560 => x"3f",
          6561 => x"96",
          6562 => x"aa",
          6563 => x"81",
          6564 => x"81",
          6565 => x"54",
          6566 => x"09",
          6567 => x"38",
          6568 => x"51",
          6569 => x"3f",
          6570 => x"fe",
          6571 => x"3d",
          6572 => x"3d",
          6573 => x"71",
          6574 => x"0c",
          6575 => x"52",
          6576 => x"86",
          6577 => x"fe",
          6578 => x"ff",
          6579 => x"7d",
          6580 => x"06",
          6581 => x"f5",
          6582 => x"3d",
          6583 => x"fe",
          6584 => x"7c",
          6585 => x"82",
          6586 => x"ff",
          6587 => x"81",
          6588 => x"7d",
          6589 => x"81",
          6590 => x"91",
          6591 => x"70",
          6592 => x"f5",
          6593 => x"e8",
          6594 => x"3d",
          6595 => x"80",
          6596 => x"51",
          6597 => x"b4",
          6598 => x"05",
          6599 => x"3f",
          6600 => x"08",
          6601 => x"90",
          6602 => x"78",
          6603 => x"89",
          6604 => x"80",
          6605 => x"d9",
          6606 => x"2e",
          6607 => x"78",
          6608 => x"38",
          6609 => x"81",
          6610 => x"82",
          6611 => x"78",
          6612 => x"ae",
          6613 => x"39",
          6614 => x"82",
          6615 => x"94",
          6616 => x"38",
          6617 => x"78",
          6618 => x"8c",
          6619 => x"24",
          6620 => x"b0",
          6621 => x"38",
          6622 => x"84",
          6623 => x"fc",
          6624 => x"2e",
          6625 => x"78",
          6626 => x"86",
          6627 => x"ec",
          6628 => x"d5",
          6629 => x"38",
          6630 => x"24",
          6631 => x"80",
          6632 => x"f6",
          6633 => x"d0",
          6634 => x"78",
          6635 => x"8a",
          6636 => x"80",
          6637 => x"c2",
          6638 => x"39",
          6639 => x"2e",
          6640 => x"78",
          6641 => x"8c",
          6642 => x"b0",
          6643 => x"82",
          6644 => x"38",
          6645 => x"24",
          6646 => x"80",
          6647 => x"96",
          6648 => x"f9",
          6649 => x"38",
          6650 => x"78",
          6651 => x"8d",
          6652 => x"81",
          6653 => x"fd",
          6654 => x"39",
          6655 => x"80",
          6656 => x"84",
          6657 => x"ed",
          6658 => x"fe",
          6659 => x"38",
          6660 => x"51",
          6661 => x"b4",
          6662 => x"11",
          6663 => x"05",
          6664 => x"dc",
          6665 => x"f0",
          6666 => x"88",
          6667 => x"25",
          6668 => x"43",
          6669 => x"05",
          6670 => x"80",
          6671 => x"51",
          6672 => x"3f",
          6673 => x"08",
          6674 => x"59",
          6675 => x"81",
          6676 => x"fe",
          6677 => x"81",
          6678 => x"39",
          6679 => x"51",
          6680 => x"b4",
          6681 => x"11",
          6682 => x"05",
          6683 => x"90",
          6684 => x"f0",
          6685 => x"fd",
          6686 => x"53",
          6687 => x"80",
          6688 => x"51",
          6689 => x"3f",
          6690 => x"08",
          6691 => x"90",
          6692 => x"39",
          6693 => x"80",
          6694 => x"84",
          6695 => x"ec",
          6696 => x"fe",
          6697 => x"2e",
          6698 => x"89",
          6699 => x"38",
          6700 => x"fc",
          6701 => x"84",
          6702 => x"ec",
          6703 => x"fe",
          6704 => x"38",
          6705 => x"08",
          6706 => x"81",
          6707 => x"79",
          6708 => x"cd",
          6709 => x"cb",
          6710 => x"79",
          6711 => x"b4",
          6712 => x"b4",
          6713 => x"b1",
          6714 => x"fe",
          6715 => x"93",
          6716 => x"e8",
          6717 => x"af",
          6718 => x"fc",
          6719 => x"3d",
          6720 => x"51",
          6721 => x"3f",
          6722 => x"08",
          6723 => x"84",
          6724 => x"fe",
          6725 => x"81",
          6726 => x"f0",
          6727 => x"51",
          6728 => x"80",
          6729 => x"3d",
          6730 => x"51",
          6731 => x"3f",
          6732 => x"08",
          6733 => x"84",
          6734 => x"fe",
          6735 => x"81",
          6736 => x"b5",
          6737 => x"05",
          6738 => x"cd",
          6739 => x"fe",
          6740 => x"3d",
          6741 => x"52",
          6742 => x"aa",
          6743 => x"ec",
          6744 => x"b8",
          6745 => x"80",
          6746 => x"f0",
          6747 => x"06",
          6748 => x"79",
          6749 => x"f2",
          6750 => x"fe",
          6751 => x"2e",
          6752 => x"81",
          6753 => x"51",
          6754 => x"fa",
          6755 => x"3d",
          6756 => x"53",
          6757 => x"51",
          6758 => x"3f",
          6759 => x"08",
          6760 => x"de",
          6761 => x"fe",
          6762 => x"ff",
          6763 => x"fe",
          6764 => x"81",
          6765 => x"80",
          6766 => x"38",
          6767 => x"f8",
          6768 => x"84",
          6769 => x"ea",
          6770 => x"fe",
          6771 => x"38",
          6772 => x"08",
          6773 => x"9c",
          6774 => x"cb",
          6775 => x"5c",
          6776 => x"27",
          6777 => x"61",
          6778 => x"70",
          6779 => x"0c",
          6780 => x"f5",
          6781 => x"39",
          6782 => x"80",
          6783 => x"84",
          6784 => x"e9",
          6785 => x"fe",
          6786 => x"2e",
          6787 => x"b4",
          6788 => x"11",
          6789 => x"05",
          6790 => x"e4",
          6791 => x"f0",
          6792 => x"f9",
          6793 => x"3d",
          6794 => x"53",
          6795 => x"51",
          6796 => x"3f",
          6797 => x"08",
          6798 => x"c6",
          6799 => x"ac",
          6800 => x"e3",
          6801 => x"79",
          6802 => x"8c",
          6803 => x"79",
          6804 => x"5b",
          6805 => x"61",
          6806 => x"eb",
          6807 => x"ff",
          6808 => x"ff",
          6809 => x"fe",
          6810 => x"81",
          6811 => x"80",
          6812 => x"38",
          6813 => x"fc",
          6814 => x"84",
          6815 => x"e8",
          6816 => x"fe",
          6817 => x"2e",
          6818 => x"b4",
          6819 => x"11",
          6820 => x"05",
          6821 => x"e8",
          6822 => x"f0",
          6823 => x"f8",
          6824 => x"f6",
          6825 => x"e0",
          6826 => x"5a",
          6827 => x"a8",
          6828 => x"33",
          6829 => x"5a",
          6830 => x"2e",
          6831 => x"55",
          6832 => x"33",
          6833 => x"81",
          6834 => x"fe",
          6835 => x"81",
          6836 => x"05",
          6837 => x"39",
          6838 => x"51",
          6839 => x"b4",
          6840 => x"11",
          6841 => x"05",
          6842 => x"94",
          6843 => x"f0",
          6844 => x"38",
          6845 => x"33",
          6846 => x"2e",
          6847 => x"f9",
          6848 => x"80",
          6849 => x"fa",
          6850 => x"78",
          6851 => x"38",
          6852 => x"08",
          6853 => x"81",
          6854 => x"59",
          6855 => x"88",
          6856 => x"fc",
          6857 => x"39",
          6858 => x"33",
          6859 => x"2e",
          6860 => x"fa",
          6861 => x"9a",
          6862 => x"b2",
          6863 => x"80",
          6864 => x"81",
          6865 => x"44",
          6866 => x"fa",
          6867 => x"80",
          6868 => x"3d",
          6869 => x"53",
          6870 => x"51",
          6871 => x"3f",
          6872 => x"08",
          6873 => x"81",
          6874 => x"59",
          6875 => x"89",
          6876 => x"f0",
          6877 => x"cc",
          6878 => x"b5",
          6879 => x"80",
          6880 => x"81",
          6881 => x"43",
          6882 => x"fa",
          6883 => x"78",
          6884 => x"38",
          6885 => x"08",
          6886 => x"81",
          6887 => x"59",
          6888 => x"88",
          6889 => x"88",
          6890 => x"39",
          6891 => x"33",
          6892 => x"2e",
          6893 => x"fa",
          6894 => x"88",
          6895 => x"9c",
          6896 => x"43",
          6897 => x"f8",
          6898 => x"84",
          6899 => x"e6",
          6900 => x"fe",
          6901 => x"2e",
          6902 => x"62",
          6903 => x"88",
          6904 => x"81",
          6905 => x"32",
          6906 => x"72",
          6907 => x"70",
          6908 => x"51",
          6909 => x"80",
          6910 => x"7a",
          6911 => x"38",
          6912 => x"f6",
          6913 => x"de",
          6914 => x"55",
          6915 => x"53",
          6916 => x"51",
          6917 => x"81",
          6918 => x"fe",
          6919 => x"f5",
          6920 => x"3d",
          6921 => x"53",
          6922 => x"51",
          6923 => x"3f",
          6924 => x"08",
          6925 => x"ca",
          6926 => x"fe",
          6927 => x"ff",
          6928 => x"fe",
          6929 => x"81",
          6930 => x"80",
          6931 => x"63",
          6932 => x"cb",
          6933 => x"34",
          6934 => x"44",
          6935 => x"fc",
          6936 => x"84",
          6937 => x"e5",
          6938 => x"fe",
          6939 => x"38",
          6940 => x"63",
          6941 => x"52",
          6942 => x"51",
          6943 => x"3f",
          6944 => x"79",
          6945 => x"dd",
          6946 => x"79",
          6947 => x"ae",
          6948 => x"38",
          6949 => x"a0",
          6950 => x"fe",
          6951 => x"ff",
          6952 => x"fe",
          6953 => x"81",
          6954 => x"80",
          6955 => x"63",
          6956 => x"cb",
          6957 => x"34",
          6958 => x"44",
          6959 => x"81",
          6960 => x"fe",
          6961 => x"ff",
          6962 => x"3d",
          6963 => x"53",
          6964 => x"51",
          6965 => x"3f",
          6966 => x"08",
          6967 => x"a2",
          6968 => x"fe",
          6969 => x"ff",
          6970 => x"fe",
          6971 => x"81",
          6972 => x"80",
          6973 => x"60",
          6974 => x"05",
          6975 => x"82",
          6976 => x"78",
          6977 => x"fe",
          6978 => x"ff",
          6979 => x"fe",
          6980 => x"81",
          6981 => x"df",
          6982 => x"39",
          6983 => x"54",
          6984 => x"94",
          6985 => x"e3",
          6986 => x"52",
          6987 => x"e2",
          6988 => x"45",
          6989 => x"78",
          6990 => x"c6",
          6991 => x"26",
          6992 => x"82",
          6993 => x"39",
          6994 => x"f0",
          6995 => x"84",
          6996 => x"e5",
          6997 => x"fe",
          6998 => x"2e",
          6999 => x"59",
          7000 => x"22",
          7001 => x"05",
          7002 => x"41",
          7003 => x"81",
          7004 => x"fe",
          7005 => x"ff",
          7006 => x"3d",
          7007 => x"53",
          7008 => x"51",
          7009 => x"3f",
          7010 => x"08",
          7011 => x"f2",
          7012 => x"fe",
          7013 => x"ff",
          7014 => x"fe",
          7015 => x"81",
          7016 => x"80",
          7017 => x"60",
          7018 => x"59",
          7019 => x"41",
          7020 => x"f0",
          7021 => x"84",
          7022 => x"e4",
          7023 => x"fe",
          7024 => x"38",
          7025 => x"60",
          7026 => x"52",
          7027 => x"51",
          7028 => x"3f",
          7029 => x"79",
          7030 => x"89",
          7031 => x"79",
          7032 => x"ae",
          7033 => x"38",
          7034 => x"9c",
          7035 => x"fe",
          7036 => x"ff",
          7037 => x"fe",
          7038 => x"81",
          7039 => x"80",
          7040 => x"60",
          7041 => x"59",
          7042 => x"41",
          7043 => x"81",
          7044 => x"fe",
          7045 => x"ff",
          7046 => x"f7",
          7047 => x"da",
          7048 => x"51",
          7049 => x"3f",
          7050 => x"81",
          7051 => x"fe",
          7052 => x"a2",
          7053 => x"aa",
          7054 => x"39",
          7055 => x"51",
          7056 => x"3f",
          7057 => x"0b",
          7058 => x"84",
          7059 => x"81",
          7060 => x"94",
          7061 => x"aa",
          7062 => x"f0",
          7063 => x"c7",
          7064 => x"83",
          7065 => x"94",
          7066 => x"80",
          7067 => x"c0",
          7068 => x"f1",
          7069 => x"3d",
          7070 => x"53",
          7071 => x"51",
          7072 => x"3f",
          7073 => x"08",
          7074 => x"f6",
          7075 => x"81",
          7076 => x"fe",
          7077 => x"63",
          7078 => x"b4",
          7079 => x"11",
          7080 => x"05",
          7081 => x"d8",
          7082 => x"f0",
          7083 => x"f0",
          7084 => x"52",
          7085 => x"51",
          7086 => x"3f",
          7087 => x"2d",
          7088 => x"08",
          7089 => x"ba",
          7090 => x"f0",
          7091 => x"f8",
          7092 => x"de",
          7093 => x"aa",
          7094 => x"d8",
          7095 => x"c7",
          7096 => x"aa",
          7097 => x"39",
          7098 => x"51",
          7099 => x"3f",
          7100 => x"a5",
          7101 => x"8b",
          7102 => x"39",
          7103 => x"33",
          7104 => x"2e",
          7105 => x"7d",
          7106 => x"78",
          7107 => x"d3",
          7108 => x"ff",
          7109 => x"fe",
          7110 => x"81",
          7111 => x"5b",
          7112 => x"82",
          7113 => x"7b",
          7114 => x"38",
          7115 => x"8c",
          7116 => x"39",
          7117 => x"b0",
          7118 => x"39",
          7119 => x"56",
          7120 => x"f9",
          7121 => x"53",
          7122 => x"52",
          7123 => x"b0",
          7124 => x"dd",
          7125 => x"39",
          7126 => x"52",
          7127 => x"b0",
          7128 => x"dd",
          7129 => x"39",
          7130 => x"f9",
          7131 => x"53",
          7132 => x"52",
          7133 => x"b0",
          7134 => x"dd",
          7135 => x"39",
          7136 => x"53",
          7137 => x"52",
          7138 => x"b0",
          7139 => x"dd",
          7140 => x"f9",
          7141 => x"ff",
          7142 => x"56",
          7143 => x"54",
          7144 => x"53",
          7145 => x"52",
          7146 => x"b0",
          7147 => x"c8",
          7148 => x"f0",
          7149 => x"f0",
          7150 => x"30",
          7151 => x"80",
          7152 => x"5b",
          7153 => x"7b",
          7154 => x"38",
          7155 => x"7a",
          7156 => x"80",
          7157 => x"81",
          7158 => x"ff",
          7159 => x"7b",
          7160 => x"7d",
          7161 => x"81",
          7162 => x"78",
          7163 => x"ff",
          7164 => x"06",
          7165 => x"81",
          7166 => x"fe",
          7167 => x"ee",
          7168 => x"3d",
          7169 => x"81",
          7170 => x"87",
          7171 => x"70",
          7172 => x"87",
          7173 => x"72",
          7174 => x"91",
          7175 => x"f0",
          7176 => x"75",
          7177 => x"87",
          7178 => x"73",
          7179 => x"fd",
          7180 => x"fe",
          7181 => x"75",
          7182 => x"94",
          7183 => x"54",
          7184 => x"80",
          7185 => x"fe",
          7186 => x"81",
          7187 => x"90",
          7188 => x"55",
          7189 => x"80",
          7190 => x"fe",
          7191 => x"72",
          7192 => x"08",
          7193 => x"8c",
          7194 => x"87",
          7195 => x"0c",
          7196 => x"0b",
          7197 => x"94",
          7198 => x"0b",
          7199 => x"0c",
          7200 => x"81",
          7201 => x"fe",
          7202 => x"fe",
          7203 => x"81",
          7204 => x"fe",
          7205 => x"81",
          7206 => x"fe",
          7207 => x"81",
          7208 => x"fe",
          7209 => x"81",
          7210 => x"3f",
          7211 => x"80",
          7212 => x"ff",
          7213 => x"00",
          7214 => x"ff",
          7215 => x"ff",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"64",
          7254 => x"2f",
          7255 => x"25",
          7256 => x"64",
          7257 => x"2e",
          7258 => x"64",
          7259 => x"6f",
          7260 => x"6f",
          7261 => x"67",
          7262 => x"74",
          7263 => x"00",
          7264 => x"28",
          7265 => x"6d",
          7266 => x"43",
          7267 => x"6e",
          7268 => x"29",
          7269 => x"0a",
          7270 => x"69",
          7271 => x"20",
          7272 => x"6c",
          7273 => x"6e",
          7274 => x"3a",
          7275 => x"20",
          7276 => x"42",
          7277 => x"52",
          7278 => x"20",
          7279 => x"38",
          7280 => x"30",
          7281 => x"2e",
          7282 => x"20",
          7283 => x"44",
          7284 => x"20",
          7285 => x"20",
          7286 => x"38",
          7287 => x"30",
          7288 => x"2e",
          7289 => x"20",
          7290 => x"4e",
          7291 => x"42",
          7292 => x"20",
          7293 => x"38",
          7294 => x"30",
          7295 => x"2e",
          7296 => x"20",
          7297 => x"52",
          7298 => x"20",
          7299 => x"20",
          7300 => x"38",
          7301 => x"30",
          7302 => x"2e",
          7303 => x"20",
          7304 => x"41",
          7305 => x"20",
          7306 => x"20",
          7307 => x"38",
          7308 => x"30",
          7309 => x"2e",
          7310 => x"20",
          7311 => x"44",
          7312 => x"52",
          7313 => x"20",
          7314 => x"76",
          7315 => x"73",
          7316 => x"30",
          7317 => x"2e",
          7318 => x"20",
          7319 => x"49",
          7320 => x"31",
          7321 => x"20",
          7322 => x"6d",
          7323 => x"20",
          7324 => x"30",
          7325 => x"2e",
          7326 => x"20",
          7327 => x"4e",
          7328 => x"43",
          7329 => x"20",
          7330 => x"61",
          7331 => x"6c",
          7332 => x"30",
          7333 => x"2e",
          7334 => x"20",
          7335 => x"49",
          7336 => x"4f",
          7337 => x"42",
          7338 => x"00",
          7339 => x"20",
          7340 => x"42",
          7341 => x"43",
          7342 => x"20",
          7343 => x"4f",
          7344 => x"0a",
          7345 => x"20",
          7346 => x"53",
          7347 => x"00",
          7348 => x"20",
          7349 => x"50",
          7350 => x"00",
          7351 => x"64",
          7352 => x"73",
          7353 => x"3a",
          7354 => x"20",
          7355 => x"50",
          7356 => x"65",
          7357 => x"20",
          7358 => x"74",
          7359 => x"41",
          7360 => x"65",
          7361 => x"3d",
          7362 => x"38",
          7363 => x"00",
          7364 => x"20",
          7365 => x"50",
          7366 => x"65",
          7367 => x"79",
          7368 => x"61",
          7369 => x"41",
          7370 => x"65",
          7371 => x"3d",
          7372 => x"38",
          7373 => x"00",
          7374 => x"20",
          7375 => x"74",
          7376 => x"20",
          7377 => x"72",
          7378 => x"64",
          7379 => x"73",
          7380 => x"20",
          7381 => x"3d",
          7382 => x"38",
          7383 => x"00",
          7384 => x"69",
          7385 => x"0a",
          7386 => x"20",
          7387 => x"50",
          7388 => x"64",
          7389 => x"20",
          7390 => x"20",
          7391 => x"20",
          7392 => x"20",
          7393 => x"3d",
          7394 => x"34",
          7395 => x"00",
          7396 => x"20",
          7397 => x"79",
          7398 => x"6d",
          7399 => x"6f",
          7400 => x"46",
          7401 => x"20",
          7402 => x"20",
          7403 => x"3d",
          7404 => x"2e",
          7405 => x"64",
          7406 => x"0a",
          7407 => x"20",
          7408 => x"44",
          7409 => x"20",
          7410 => x"63",
          7411 => x"72",
          7412 => x"20",
          7413 => x"20",
          7414 => x"3d",
          7415 => x"2e",
          7416 => x"64",
          7417 => x"0a",
          7418 => x"20",
          7419 => x"69",
          7420 => x"6f",
          7421 => x"53",
          7422 => x"4d",
          7423 => x"6f",
          7424 => x"46",
          7425 => x"3d",
          7426 => x"2e",
          7427 => x"64",
          7428 => x"0a",
          7429 => x"6d",
          7430 => x"00",
          7431 => x"65",
          7432 => x"6d",
          7433 => x"6c",
          7434 => x"00",
          7435 => x"56",
          7436 => x"56",
          7437 => x"6e",
          7438 => x"6e",
          7439 => x"77",
          7440 => x"69",
          7441 => x"72",
          7442 => x"78",
          7443 => x"69",
          7444 => x"72",
          7445 => x"69",
          7446 => x"00",
          7447 => x"00",
          7448 => x"30",
          7449 => x"20",
          7450 => x"00",
          7451 => x"61",
          7452 => x"64",
          7453 => x"20",
          7454 => x"65",
          7455 => x"68",
          7456 => x"69",
          7457 => x"72",
          7458 => x"69",
          7459 => x"74",
          7460 => x"4f",
          7461 => x"00",
          7462 => x"61",
          7463 => x"74",
          7464 => x"65",
          7465 => x"72",
          7466 => x"65",
          7467 => x"73",
          7468 => x"79",
          7469 => x"6c",
          7470 => x"64",
          7471 => x"62",
          7472 => x"67",
          7473 => x"00",
          7474 => x"00",
          7475 => x"00",
          7476 => x"00",
          7477 => x"00",
          7478 => x"00",
          7479 => x"00",
          7480 => x"00",
          7481 => x"00",
          7482 => x"00",
          7483 => x"00",
          7484 => x"00",
          7485 => x"00",
          7486 => x"00",
          7487 => x"00",
          7488 => x"00",
          7489 => x"00",
          7490 => x"00",
          7491 => x"00",
          7492 => x"00",
          7493 => x"00",
          7494 => x"00",
          7495 => x"00",
          7496 => x"00",
          7497 => x"00",
          7498 => x"00",
          7499 => x"00",
          7500 => x"00",
          7501 => x"00",
          7502 => x"00",
          7503 => x"00",
          7504 => x"00",
          7505 => x"00",
          7506 => x"00",
          7507 => x"5b",
          7508 => x"5b",
          7509 => x"5b",
          7510 => x"5b",
          7511 => x"5b",
          7512 => x"5b",
          7513 => x"5b",
          7514 => x"5b",
          7515 => x"5b",
          7516 => x"00",
          7517 => x"00",
          7518 => x"44",
          7519 => x"2a",
          7520 => x"3b",
          7521 => x"3f",
          7522 => x"7f",
          7523 => x"41",
          7524 => x"41",
          7525 => x"00",
          7526 => x"fe",
          7527 => x"44",
          7528 => x"2e",
          7529 => x"4f",
          7530 => x"4d",
          7531 => x"20",
          7532 => x"54",
          7533 => x"20",
          7534 => x"4f",
          7535 => x"4d",
          7536 => x"20",
          7537 => x"54",
          7538 => x"20",
          7539 => x"00",
          7540 => x"00",
          7541 => x"00",
          7542 => x"00",
          7543 => x"9a",
          7544 => x"41",
          7545 => x"45",
          7546 => x"49",
          7547 => x"92",
          7548 => x"4f",
          7549 => x"99",
          7550 => x"9d",
          7551 => x"49",
          7552 => x"a5",
          7553 => x"a9",
          7554 => x"ad",
          7555 => x"b1",
          7556 => x"b5",
          7557 => x"b9",
          7558 => x"bd",
          7559 => x"c1",
          7560 => x"c5",
          7561 => x"c9",
          7562 => x"cd",
          7563 => x"d1",
          7564 => x"d5",
          7565 => x"d9",
          7566 => x"dd",
          7567 => x"e1",
          7568 => x"e5",
          7569 => x"e9",
          7570 => x"ed",
          7571 => x"f1",
          7572 => x"f5",
          7573 => x"f9",
          7574 => x"fd",
          7575 => x"2e",
          7576 => x"5b",
          7577 => x"22",
          7578 => x"3e",
          7579 => x"00",
          7580 => x"01",
          7581 => x"10",
          7582 => x"00",
          7583 => x"00",
          7584 => x"01",
          7585 => x"04",
          7586 => x"10",
          7587 => x"00",
          7588 => x"69",
          7589 => x"00",
          7590 => x"69",
          7591 => x"6c",
          7592 => x"69",
          7593 => x"00",
          7594 => x"6c",
          7595 => x"00",
          7596 => x"65",
          7597 => x"00",
          7598 => x"63",
          7599 => x"72",
          7600 => x"63",
          7601 => x"00",
          7602 => x"64",
          7603 => x"00",
          7604 => x"64",
          7605 => x"00",
          7606 => x"65",
          7607 => x"65",
          7608 => x"65",
          7609 => x"69",
          7610 => x"69",
          7611 => x"66",
          7612 => x"66",
          7613 => x"61",
          7614 => x"00",
          7615 => x"6d",
          7616 => x"65",
          7617 => x"72",
          7618 => x"65",
          7619 => x"00",
          7620 => x"6e",
          7621 => x"00",
          7622 => x"65",
          7623 => x"00",
          7624 => x"62",
          7625 => x"63",
          7626 => x"62",
          7627 => x"63",
          7628 => x"69",
          7629 => x"00",
          7630 => x"69",
          7631 => x"45",
          7632 => x"72",
          7633 => x"6e",
          7634 => x"6e",
          7635 => x"65",
          7636 => x"72",
          7637 => x"00",
          7638 => x"69",
          7639 => x"6e",
          7640 => x"72",
          7641 => x"79",
          7642 => x"00",
          7643 => x"6f",
          7644 => x"6c",
          7645 => x"6f",
          7646 => x"2e",
          7647 => x"6f",
          7648 => x"74",
          7649 => x"6f",
          7650 => x"2e",
          7651 => x"6e",
          7652 => x"69",
          7653 => x"69",
          7654 => x"61",
          7655 => x"0a",
          7656 => x"63",
          7657 => x"73",
          7658 => x"6e",
          7659 => x"2e",
          7660 => x"69",
          7661 => x"61",
          7662 => x"61",
          7663 => x"65",
          7664 => x"74",
          7665 => x"00",
          7666 => x"69",
          7667 => x"68",
          7668 => x"6c",
          7669 => x"6e",
          7670 => x"69",
          7671 => x"00",
          7672 => x"44",
          7673 => x"20",
          7674 => x"74",
          7675 => x"72",
          7676 => x"63",
          7677 => x"2e",
          7678 => x"72",
          7679 => x"20",
          7680 => x"62",
          7681 => x"69",
          7682 => x"6e",
          7683 => x"69",
          7684 => x"00",
          7685 => x"69",
          7686 => x"6e",
          7687 => x"65",
          7688 => x"6c",
          7689 => x"0a",
          7690 => x"6f",
          7691 => x"6d",
          7692 => x"69",
          7693 => x"20",
          7694 => x"65",
          7695 => x"74",
          7696 => x"66",
          7697 => x"64",
          7698 => x"20",
          7699 => x"6b",
          7700 => x"00",
          7701 => x"6f",
          7702 => x"74",
          7703 => x"6f",
          7704 => x"64",
          7705 => x"00",
          7706 => x"69",
          7707 => x"75",
          7708 => x"6f",
          7709 => x"61",
          7710 => x"6e",
          7711 => x"6e",
          7712 => x"6c",
          7713 => x"0a",
          7714 => x"69",
          7715 => x"69",
          7716 => x"6f",
          7717 => x"64",
          7718 => x"00",
          7719 => x"6e",
          7720 => x"66",
          7721 => x"65",
          7722 => x"6d",
          7723 => x"72",
          7724 => x"00",
          7725 => x"6f",
          7726 => x"61",
          7727 => x"6f",
          7728 => x"20",
          7729 => x"65",
          7730 => x"00",
          7731 => x"61",
          7732 => x"65",
          7733 => x"73",
          7734 => x"63",
          7735 => x"65",
          7736 => x"0a",
          7737 => x"75",
          7738 => x"73",
          7739 => x"00",
          7740 => x"6e",
          7741 => x"77",
          7742 => x"72",
          7743 => x"2e",
          7744 => x"25",
          7745 => x"62",
          7746 => x"73",
          7747 => x"20",
          7748 => x"25",
          7749 => x"62",
          7750 => x"73",
          7751 => x"63",
          7752 => x"00",
          7753 => x"65",
          7754 => x"00",
          7755 => x"30",
          7756 => x"00",
          7757 => x"20",
          7758 => x"30",
          7759 => x"00",
          7760 => x"20",
          7761 => x"20",
          7762 => x"00",
          7763 => x"30",
          7764 => x"00",
          7765 => x"20",
          7766 => x"7c",
          7767 => x"0d",
          7768 => x"50",
          7769 => x"00",
          7770 => x"2a",
          7771 => x"73",
          7772 => x"00",
          7773 => x"31",
          7774 => x"2f",
          7775 => x"30",
          7776 => x"31",
          7777 => x"00",
          7778 => x"5a",
          7779 => x"20",
          7780 => x"20",
          7781 => x"78",
          7782 => x"73",
          7783 => x"20",
          7784 => x"0a",
          7785 => x"50",
          7786 => x"20",
          7787 => x"65",
          7788 => x"70",
          7789 => x"61",
          7790 => x"65",
          7791 => x"00",
          7792 => x"69",
          7793 => x"20",
          7794 => x"65",
          7795 => x"70",
          7796 => x"00",
          7797 => x"53",
          7798 => x"6e",
          7799 => x"72",
          7800 => x"0a",
          7801 => x"4f",
          7802 => x"20",
          7803 => x"69",
          7804 => x"72",
          7805 => x"74",
          7806 => x"4f",
          7807 => x"20",
          7808 => x"69",
          7809 => x"72",
          7810 => x"74",
          7811 => x"41",
          7812 => x"20",
          7813 => x"69",
          7814 => x"72",
          7815 => x"74",
          7816 => x"41",
          7817 => x"20",
          7818 => x"69",
          7819 => x"72",
          7820 => x"74",
          7821 => x"41",
          7822 => x"20",
          7823 => x"69",
          7824 => x"72",
          7825 => x"74",
          7826 => x"41",
          7827 => x"20",
          7828 => x"69",
          7829 => x"72",
          7830 => x"74",
          7831 => x"65",
          7832 => x"6e",
          7833 => x"70",
          7834 => x"6d",
          7835 => x"2e",
          7836 => x"00",
          7837 => x"6e",
          7838 => x"69",
          7839 => x"74",
          7840 => x"72",
          7841 => x"0a",
          7842 => x"75",
          7843 => x"78",
          7844 => x"62",
          7845 => x"00",
          7846 => x"3a",
          7847 => x"61",
          7848 => x"64",
          7849 => x"20",
          7850 => x"74",
          7851 => x"69",
          7852 => x"73",
          7853 => x"61",
          7854 => x"30",
          7855 => x"6c",
          7856 => x"65",
          7857 => x"69",
          7858 => x"61",
          7859 => x"6c",
          7860 => x"0a",
          7861 => x"20",
          7862 => x"61",
          7863 => x"69",
          7864 => x"69",
          7865 => x"00",
          7866 => x"6e",
          7867 => x"61",
          7868 => x"65",
          7869 => x"00",
          7870 => x"61",
          7871 => x"64",
          7872 => x"20",
          7873 => x"74",
          7874 => x"69",
          7875 => x"0a",
          7876 => x"63",
          7877 => x"0a",
          7878 => x"75",
          7879 => x"6c",
          7880 => x"69",
          7881 => x"2e",
          7882 => x"00",
          7883 => x"6f",
          7884 => x"6e",
          7885 => x"2e",
          7886 => x"6f",
          7887 => x"72",
          7888 => x"2e",
          7889 => x"00",
          7890 => x"30",
          7891 => x"28",
          7892 => x"78",
          7893 => x"25",
          7894 => x"78",
          7895 => x"38",
          7896 => x"00",
          7897 => x"75",
          7898 => x"4d",
          7899 => x"72",
          7900 => x"00",
          7901 => x"43",
          7902 => x"6c",
          7903 => x"2e",
          7904 => x"30",
          7905 => x"25",
          7906 => x"2d",
          7907 => x"3f",
          7908 => x"00",
          7909 => x"30",
          7910 => x"25",
          7911 => x"2d",
          7912 => x"30",
          7913 => x"25",
          7914 => x"2d",
          7915 => x"69",
          7916 => x"6c",
          7917 => x"20",
          7918 => x"65",
          7919 => x"70",
          7920 => x"00",
          7921 => x"6e",
          7922 => x"69",
          7923 => x"69",
          7924 => x"72",
          7925 => x"74",
          7926 => x"00",
          7927 => x"69",
          7928 => x"6c",
          7929 => x"75",
          7930 => x"20",
          7931 => x"6f",
          7932 => x"6e",
          7933 => x"69",
          7934 => x"75",
          7935 => x"20",
          7936 => x"6f",
          7937 => x"78",
          7938 => x"74",
          7939 => x"20",
          7940 => x"65",
          7941 => x"25",
          7942 => x"20",
          7943 => x"0a",
          7944 => x"61",
          7945 => x"6e",
          7946 => x"6f",
          7947 => x"40",
          7948 => x"38",
          7949 => x"2e",
          7950 => x"00",
          7951 => x"61",
          7952 => x"72",
          7953 => x"72",
          7954 => x"20",
          7955 => x"65",
          7956 => x"64",
          7957 => x"00",
          7958 => x"65",
          7959 => x"72",
          7960 => x"67",
          7961 => x"70",
          7962 => x"61",
          7963 => x"6e",
          7964 => x"0a",
          7965 => x"6f",
          7966 => x"72",
          7967 => x"6f",
          7968 => x"67",
          7969 => x"0a",
          7970 => x"50",
          7971 => x"69",
          7972 => x"64",
          7973 => x"73",
          7974 => x"2e",
          7975 => x"00",
          7976 => x"64",
          7977 => x"73",
          7978 => x"00",
          7979 => x"64",
          7980 => x"73",
          7981 => x"61",
          7982 => x"6f",
          7983 => x"6e",
          7984 => x"00",
          7985 => x"75",
          7986 => x"6e",
          7987 => x"2e",
          7988 => x"6e",
          7989 => x"69",
          7990 => x"69",
          7991 => x"72",
          7992 => x"74",
          7993 => x"2e",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"01",
          8000 => x"00",
          8001 => x"01",
          8002 => x"81",
          8003 => x"00",
          8004 => x"7f",
          8005 => x"00",
          8006 => x"00",
          8007 => x"00",
          8008 => x"00",
          8009 => x"f5",
          8010 => x"f5",
          8011 => x"f5",
          8012 => x"00",
          8013 => x"01",
          8014 => x"01",
          8015 => x"01",
          8016 => x"00",
          8017 => x"00",
          8018 => x"00",
          8019 => x"00",
          8020 => x"00",
          8021 => x"00",
          8022 => x"00",
          8023 => x"00",
          8024 => x"00",
          8025 => x"00",
          8026 => x"00",
          8027 => x"00",
          8028 => x"00",
          8029 => x"00",
          8030 => x"00",
          8031 => x"00",
          8032 => x"00",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"02",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"04",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"14",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"2b",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"30",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"3c",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"3d",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"3f",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"40",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"41",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"42",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"43",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"50",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"51",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"54",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"55",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"79",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"78",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"82",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"83",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"85",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"87",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"8c",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"8d",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"8e",
          8154 => x"00",
          8155 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"8c",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"f0",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"b0",
           163 => x"10",
           164 => x"06",
           165 => x"92",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"91",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"fd",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"94",
           269 => x"0b",
           270 => x"0b",
           271 => x"b2",
           272 => x"0b",
           273 => x"0b",
           274 => x"d0",
           275 => x"0b",
           276 => x"0b",
           277 => x"ee",
           278 => x"0b",
           279 => x"0b",
           280 => x"8c",
           281 => x"0b",
           282 => x"0b",
           283 => x"aa",
           284 => x"0b",
           285 => x"0b",
           286 => x"c8",
           287 => x"0b",
           288 => x"0b",
           289 => x"e6",
           290 => x"0b",
           291 => x"0b",
           292 => x"84",
           293 => x"0b",
           294 => x"0b",
           295 => x"a3",
           296 => x"0b",
           297 => x"0b",
           298 => x"c3",
           299 => x"0b",
           300 => x"0b",
           301 => x"e3",
           302 => x"0b",
           303 => x"0b",
           304 => x"83",
           305 => x"0b",
           306 => x"0b",
           307 => x"a3",
           308 => x"0b",
           309 => x"0b",
           310 => x"c3",
           311 => x"0b",
           312 => x"0b",
           313 => x"e3",
           314 => x"0b",
           315 => x"0b",
           316 => x"83",
           317 => x"0b",
           318 => x"0b",
           319 => x"a3",
           320 => x"0b",
           321 => x"0b",
           322 => x"c3",
           323 => x"0b",
           324 => x"0b",
           325 => x"e3",
           326 => x"0b",
           327 => x"0b",
           328 => x"83",
           329 => x"0b",
           330 => x"0b",
           331 => x"a3",
           332 => x"0b",
           333 => x"0b",
           334 => x"c3",
           335 => x"0b",
           336 => x"0b",
           337 => x"e3",
           338 => x"0b",
           339 => x"0b",
           340 => x"82",
           341 => x"0b",
           342 => x"0b",
           343 => x"a0",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"81",
           388 => x"83",
           389 => x"81",
           390 => x"b5",
           391 => x"fe",
           392 => x"80",
           393 => x"fe",
           394 => x"87",
           395 => x"fc",
           396 => x"90",
           397 => x"fc",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"81",
           403 => x"83",
           404 => x"81",
           405 => x"bd",
           406 => x"fe",
           407 => x"80",
           408 => x"fe",
           409 => x"c8",
           410 => x"fc",
           411 => x"90",
           412 => x"fc",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"81",
           418 => x"83",
           419 => x"81",
           420 => x"bc",
           421 => x"fe",
           422 => x"80",
           423 => x"fe",
           424 => x"fa",
           425 => x"fc",
           426 => x"90",
           427 => x"fc",
           428 => x"2d",
           429 => x"08",
           430 => x"04",
           431 => x"0c",
           432 => x"81",
           433 => x"83",
           434 => x"81",
           435 => x"a6",
           436 => x"fe",
           437 => x"80",
           438 => x"fe",
           439 => x"dd",
           440 => x"fc",
           441 => x"90",
           442 => x"fc",
           443 => x"2d",
           444 => x"08",
           445 => x"04",
           446 => x"0c",
           447 => x"81",
           448 => x"83",
           449 => x"81",
           450 => x"a1",
           451 => x"fe",
           452 => x"80",
           453 => x"fe",
           454 => x"84",
           455 => x"fe",
           456 => x"80",
           457 => x"fe",
           458 => x"91",
           459 => x"fe",
           460 => x"80",
           461 => x"fe",
           462 => x"89",
           463 => x"fe",
           464 => x"80",
           465 => x"fe",
           466 => x"8c",
           467 => x"fe",
           468 => x"80",
           469 => x"fe",
           470 => x"96",
           471 => x"fe",
           472 => x"80",
           473 => x"fe",
           474 => x"9f",
           475 => x"fe",
           476 => x"80",
           477 => x"fe",
           478 => x"90",
           479 => x"fe",
           480 => x"80",
           481 => x"fe",
           482 => x"99",
           483 => x"fe",
           484 => x"80",
           485 => x"fe",
           486 => x"9b",
           487 => x"fe",
           488 => x"80",
           489 => x"fe",
           490 => x"9b",
           491 => x"fe",
           492 => x"80",
           493 => x"fe",
           494 => x"a3",
           495 => x"fe",
           496 => x"80",
           497 => x"fe",
           498 => x"a0",
           499 => x"fe",
           500 => x"80",
           501 => x"fe",
           502 => x"a5",
           503 => x"fe",
           504 => x"80",
           505 => x"fe",
           506 => x"9c",
           507 => x"fe",
           508 => x"80",
           509 => x"fe",
           510 => x"a8",
           511 => x"fe",
           512 => x"80",
           513 => x"fe",
           514 => x"a9",
           515 => x"fe",
           516 => x"80",
           517 => x"fe",
           518 => x"92",
           519 => x"fe",
           520 => x"80",
           521 => x"fe",
           522 => x"91",
           523 => x"fe",
           524 => x"80",
           525 => x"fe",
           526 => x"93",
           527 => x"fe",
           528 => x"80",
           529 => x"fe",
           530 => x"9c",
           531 => x"fe",
           532 => x"80",
           533 => x"fe",
           534 => x"aa",
           535 => x"fe",
           536 => x"80",
           537 => x"fe",
           538 => x"ac",
           539 => x"fe",
           540 => x"80",
           541 => x"fe",
           542 => x"b0",
           543 => x"fe",
           544 => x"80",
           545 => x"fe",
           546 => x"83",
           547 => x"fe",
           548 => x"80",
           549 => x"fe",
           550 => x"b3",
           551 => x"fe",
           552 => x"80",
           553 => x"fe",
           554 => x"c1",
           555 => x"fe",
           556 => x"80",
           557 => x"fe",
           558 => x"bf",
           559 => x"fe",
           560 => x"80",
           561 => x"fe",
           562 => x"d5",
           563 => x"fe",
           564 => x"80",
           565 => x"fe",
           566 => x"d7",
           567 => x"fe",
           568 => x"80",
           569 => x"fe",
           570 => x"d8",
           571 => x"fe",
           572 => x"80",
           573 => x"fe",
           574 => x"a2",
           575 => x"fc",
           576 => x"90",
           577 => x"fc",
           578 => x"2d",
           579 => x"08",
           580 => x"04",
           581 => x"0c",
           582 => x"81",
           583 => x"83",
           584 => x"81",
           585 => x"81",
           586 => x"81",
           587 => x"83",
           588 => x"3c",
           589 => x"10",
           590 => x"10",
           591 => x"10",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"51",
           598 => x"73",
           599 => x"73",
           600 => x"81",
           601 => x"10",
           602 => x"07",
           603 => x"0c",
           604 => x"72",
           605 => x"81",
           606 => x"09",
           607 => x"71",
           608 => x"0a",
           609 => x"72",
           610 => x"51",
           611 => x"81",
           612 => x"82",
           613 => x"8e",
           614 => x"70",
           615 => x"0c",
           616 => x"93",
           617 => x"81",
           618 => x"80",
           619 => x"fe",
           620 => x"81",
           621 => x"fd",
           622 => x"53",
           623 => x"08",
           624 => x"52",
           625 => x"08",
           626 => x"51",
           627 => x"81",
           628 => x"70",
           629 => x"0c",
           630 => x"0d",
           631 => x"0c",
           632 => x"fc",
           633 => x"fe",
           634 => x"3d",
           635 => x"81",
           636 => x"8c",
           637 => x"81",
           638 => x"88",
           639 => x"83",
           640 => x"fe",
           641 => x"81",
           642 => x"54",
           643 => x"81",
           644 => x"04",
           645 => x"08",
           646 => x"fc",
           647 => x"0d",
           648 => x"fe",
           649 => x"05",
           650 => x"fc",
           651 => x"08",
           652 => x"38",
           653 => x"08",
           654 => x"30",
           655 => x"08",
           656 => x"80",
           657 => x"fc",
           658 => x"0c",
           659 => x"08",
           660 => x"8a",
           661 => x"81",
           662 => x"f4",
           663 => x"fe",
           664 => x"05",
           665 => x"fc",
           666 => x"0c",
           667 => x"08",
           668 => x"80",
           669 => x"81",
           670 => x"8c",
           671 => x"81",
           672 => x"8c",
           673 => x"0b",
           674 => x"08",
           675 => x"81",
           676 => x"fc",
           677 => x"38",
           678 => x"fe",
           679 => x"05",
           680 => x"fc",
           681 => x"08",
           682 => x"08",
           683 => x"80",
           684 => x"fc",
           685 => x"08",
           686 => x"fc",
           687 => x"08",
           688 => x"3f",
           689 => x"08",
           690 => x"fc",
           691 => x"0c",
           692 => x"fc",
           693 => x"08",
           694 => x"38",
           695 => x"08",
           696 => x"30",
           697 => x"08",
           698 => x"81",
           699 => x"f8",
           700 => x"81",
           701 => x"54",
           702 => x"81",
           703 => x"04",
           704 => x"08",
           705 => x"fc",
           706 => x"0d",
           707 => x"fe",
           708 => x"05",
           709 => x"fc",
           710 => x"08",
           711 => x"38",
           712 => x"08",
           713 => x"30",
           714 => x"08",
           715 => x"81",
           716 => x"fc",
           717 => x"0c",
           718 => x"08",
           719 => x"80",
           720 => x"81",
           721 => x"8c",
           722 => x"81",
           723 => x"8c",
           724 => x"53",
           725 => x"08",
           726 => x"52",
           727 => x"08",
           728 => x"51",
           729 => x"fe",
           730 => x"81",
           731 => x"f8",
           732 => x"81",
           733 => x"fc",
           734 => x"2e",
           735 => x"fe",
           736 => x"05",
           737 => x"fe",
           738 => x"05",
           739 => x"fc",
           740 => x"08",
           741 => x"f0",
           742 => x"3d",
           743 => x"fc",
           744 => x"fe",
           745 => x"81",
           746 => x"fd",
           747 => x"0b",
           748 => x"08",
           749 => x"80",
           750 => x"fc",
           751 => x"0c",
           752 => x"08",
           753 => x"81",
           754 => x"88",
           755 => x"b9",
           756 => x"fc",
           757 => x"08",
           758 => x"38",
           759 => x"fe",
           760 => x"05",
           761 => x"38",
           762 => x"08",
           763 => x"10",
           764 => x"08",
           765 => x"81",
           766 => x"fc",
           767 => x"81",
           768 => x"fc",
           769 => x"b8",
           770 => x"fc",
           771 => x"08",
           772 => x"e1",
           773 => x"fc",
           774 => x"08",
           775 => x"08",
           776 => x"26",
           777 => x"fe",
           778 => x"05",
           779 => x"fc",
           780 => x"08",
           781 => x"fc",
           782 => x"0c",
           783 => x"08",
           784 => x"81",
           785 => x"fc",
           786 => x"81",
           787 => x"f8",
           788 => x"fe",
           789 => x"05",
           790 => x"81",
           791 => x"fc",
           792 => x"fe",
           793 => x"05",
           794 => x"81",
           795 => x"8c",
           796 => x"95",
           797 => x"fc",
           798 => x"08",
           799 => x"38",
           800 => x"08",
           801 => x"70",
           802 => x"08",
           803 => x"51",
           804 => x"fe",
           805 => x"05",
           806 => x"fe",
           807 => x"05",
           808 => x"fe",
           809 => x"05",
           810 => x"f0",
           811 => x"0d",
           812 => x"0c",
           813 => x"0d",
           814 => x"7b",
           815 => x"55",
           816 => x"8c",
           817 => x"07",
           818 => x"70",
           819 => x"38",
           820 => x"71",
           821 => x"38",
           822 => x"05",
           823 => x"70",
           824 => x"34",
           825 => x"71",
           826 => x"81",
           827 => x"74",
           828 => x"0c",
           829 => x"04",
           830 => x"70",
           831 => x"08",
           832 => x"05",
           833 => x"70",
           834 => x"08",
           835 => x"05",
           836 => x"70",
           837 => x"08",
           838 => x"05",
           839 => x"70",
           840 => x"08",
           841 => x"05",
           842 => x"12",
           843 => x"26",
           844 => x"72",
           845 => x"72",
           846 => x"54",
           847 => x"84",
           848 => x"fc",
           849 => x"83",
           850 => x"70",
           851 => x"39",
           852 => x"76",
           853 => x"8c",
           854 => x"33",
           855 => x"55",
           856 => x"8a",
           857 => x"06",
           858 => x"2e",
           859 => x"12",
           860 => x"2e",
           861 => x"73",
           862 => x"55",
           863 => x"52",
           864 => x"09",
           865 => x"38",
           866 => x"f0",
           867 => x"0d",
           868 => x"88",
           869 => x"70",
           870 => x"07",
           871 => x"8f",
           872 => x"38",
           873 => x"84",
           874 => x"72",
           875 => x"05",
           876 => x"71",
           877 => x"53",
           878 => x"70",
           879 => x"0c",
           880 => x"71",
           881 => x"38",
           882 => x"90",
           883 => x"70",
           884 => x"0c",
           885 => x"71",
           886 => x"38",
           887 => x"8e",
           888 => x"0d",
           889 => x"70",
           890 => x"06",
           891 => x"55",
           892 => x"38",
           893 => x"70",
           894 => x"fb",
           895 => x"06",
           896 => x"82",
           897 => x"51",
           898 => x"54",
           899 => x"84",
           900 => x"70",
           901 => x"0c",
           902 => x"09",
           903 => x"fd",
           904 => x"70",
           905 => x"81",
           906 => x"51",
           907 => x"70",
           908 => x"38",
           909 => x"70",
           910 => x"33",
           911 => x"70",
           912 => x"34",
           913 => x"74",
           914 => x"0c",
           915 => x"04",
           916 => x"75",
           917 => x"06",
           918 => x"70",
           919 => x"70",
           920 => x"f7",
           921 => x"12",
           922 => x"84",
           923 => x"06",
           924 => x"53",
           925 => x"84",
           926 => x"70",
           927 => x"fd",
           928 => x"70",
           929 => x"81",
           930 => x"51",
           931 => x"80",
           932 => x"72",
           933 => x"51",
           934 => x"8a",
           935 => x"70",
           936 => x"70",
           937 => x"74",
           938 => x"f0",
           939 => x"0d",
           940 => x"0d",
           941 => x"70",
           942 => x"52",
           943 => x"80",
           944 => x"74",
           945 => x"51",
           946 => x"80",
           947 => x"13",
           948 => x"2e",
           949 => x"33",
           950 => x"51",
           951 => x"09",
           952 => x"38",
           953 => x"81",
           954 => x"81",
           955 => x"70",
           956 => x"fe",
           957 => x"81",
           958 => x"55",
           959 => x"ff",
           960 => x"06",
           961 => x"33",
           962 => x"51",
           963 => x"06",
           964 => x"06",
           965 => x"51",
           966 => x"81",
           967 => x"88",
           968 => x"71",
           969 => x"83",
           970 => x"38",
           971 => x"08",
           972 => x"74",
           973 => x"ff",
           974 => x"13",
           975 => x"2e",
           976 => x"08",
           977 => x"fb",
           978 => x"06",
           979 => x"82",
           980 => x"51",
           981 => x"9a",
           982 => x"84",
           983 => x"83",
           984 => x"38",
           985 => x"08",
           986 => x"74",
           987 => x"fe",
           988 => x"0b",
           989 => x"0c",
           990 => x"04",
           991 => x"80",
           992 => x"71",
           993 => x"87",
           994 => x"fe",
           995 => x"ff",
           996 => x"ff",
           997 => x"72",
           998 => x"38",
           999 => x"f0",
          1000 => x"0d",
          1001 => x"0d",
          1002 => x"70",
          1003 => x"71",
          1004 => x"ca",
          1005 => x"51",
          1006 => x"09",
          1007 => x"38",
          1008 => x"f1",
          1009 => x"84",
          1010 => x"53",
          1011 => x"70",
          1012 => x"53",
          1013 => x"a0",
          1014 => x"81",
          1015 => x"2e",
          1016 => x"e5",
          1017 => x"ff",
          1018 => x"a0",
          1019 => x"06",
          1020 => x"73",
          1021 => x"55",
          1022 => x"0c",
          1023 => x"81",
          1024 => x"87",
          1025 => x"fc",
          1026 => x"53",
          1027 => x"2e",
          1028 => x"3d",
          1029 => x"72",
          1030 => x"3f",
          1031 => x"08",
          1032 => x"53",
          1033 => x"53",
          1034 => x"f0",
          1035 => x"0d",
          1036 => x"0d",
          1037 => x"33",
          1038 => x"53",
          1039 => x"8b",
          1040 => x"38",
          1041 => x"ff",
          1042 => x"52",
          1043 => x"81",
          1044 => x"13",
          1045 => x"52",
          1046 => x"80",
          1047 => x"13",
          1048 => x"52",
          1049 => x"80",
          1050 => x"13",
          1051 => x"52",
          1052 => x"80",
          1053 => x"13",
          1054 => x"52",
          1055 => x"26",
          1056 => x"8a",
          1057 => x"87",
          1058 => x"e7",
          1059 => x"38",
          1060 => x"c0",
          1061 => x"72",
          1062 => x"98",
          1063 => x"13",
          1064 => x"98",
          1065 => x"13",
          1066 => x"98",
          1067 => x"13",
          1068 => x"98",
          1069 => x"13",
          1070 => x"98",
          1071 => x"13",
          1072 => x"98",
          1073 => x"87",
          1074 => x"0c",
          1075 => x"98",
          1076 => x"0b",
          1077 => x"9c",
          1078 => x"71",
          1079 => x"0c",
          1080 => x"04",
          1081 => x"7f",
          1082 => x"98",
          1083 => x"7d",
          1084 => x"98",
          1085 => x"7d",
          1086 => x"c0",
          1087 => x"5a",
          1088 => x"34",
          1089 => x"b4",
          1090 => x"83",
          1091 => x"c0",
          1092 => x"5a",
          1093 => x"34",
          1094 => x"ac",
          1095 => x"85",
          1096 => x"c0",
          1097 => x"5a",
          1098 => x"34",
          1099 => x"a4",
          1100 => x"88",
          1101 => x"c0",
          1102 => x"5a",
          1103 => x"23",
          1104 => x"79",
          1105 => x"06",
          1106 => x"ff",
          1107 => x"86",
          1108 => x"85",
          1109 => x"84",
          1110 => x"83",
          1111 => x"82",
          1112 => x"7d",
          1113 => x"06",
          1114 => x"d4",
          1115 => x"3f",
          1116 => x"04",
          1117 => x"02",
          1118 => x"70",
          1119 => x"2a",
          1120 => x"70",
          1121 => x"f9",
          1122 => x"3d",
          1123 => x"3d",
          1124 => x"0b",
          1125 => x"33",
          1126 => x"06",
          1127 => x"87",
          1128 => x"51",
          1129 => x"86",
          1130 => x"94",
          1131 => x"08",
          1132 => x"70",
          1133 => x"54",
          1134 => x"2e",
          1135 => x"91",
          1136 => x"06",
          1137 => x"d7",
          1138 => x"32",
          1139 => x"51",
          1140 => x"2e",
          1141 => x"93",
          1142 => x"06",
          1143 => x"ff",
          1144 => x"81",
          1145 => x"87",
          1146 => x"52",
          1147 => x"86",
          1148 => x"94",
          1149 => x"72",
          1150 => x"fe",
          1151 => x"3d",
          1152 => x"3d",
          1153 => x"05",
          1154 => x"81",
          1155 => x"70",
          1156 => x"57",
          1157 => x"c0",
          1158 => x"74",
          1159 => x"38",
          1160 => x"94",
          1161 => x"70",
          1162 => x"81",
          1163 => x"52",
          1164 => x"8c",
          1165 => x"2a",
          1166 => x"51",
          1167 => x"38",
          1168 => x"70",
          1169 => x"51",
          1170 => x"8d",
          1171 => x"2a",
          1172 => x"51",
          1173 => x"be",
          1174 => x"ff",
          1175 => x"c0",
          1176 => x"70",
          1177 => x"38",
          1178 => x"90",
          1179 => x"0c",
          1180 => x"04",
          1181 => x"79",
          1182 => x"33",
          1183 => x"06",
          1184 => x"70",
          1185 => x"fe",
          1186 => x"ff",
          1187 => x"0b",
          1188 => x"e8",
          1189 => x"ff",
          1190 => x"55",
          1191 => x"94",
          1192 => x"80",
          1193 => x"87",
          1194 => x"51",
          1195 => x"96",
          1196 => x"06",
          1197 => x"70",
          1198 => x"38",
          1199 => x"70",
          1200 => x"51",
          1201 => x"72",
          1202 => x"81",
          1203 => x"70",
          1204 => x"38",
          1205 => x"70",
          1206 => x"51",
          1207 => x"38",
          1208 => x"06",
          1209 => x"94",
          1210 => x"80",
          1211 => x"87",
          1212 => x"52",
          1213 => x"81",
          1214 => x"70",
          1215 => x"53",
          1216 => x"ff",
          1217 => x"81",
          1218 => x"89",
          1219 => x"fe",
          1220 => x"0b",
          1221 => x"33",
          1222 => x"06",
          1223 => x"c0",
          1224 => x"72",
          1225 => x"38",
          1226 => x"94",
          1227 => x"70",
          1228 => x"81",
          1229 => x"51",
          1230 => x"e2",
          1231 => x"ff",
          1232 => x"c0",
          1233 => x"70",
          1234 => x"38",
          1235 => x"90",
          1236 => x"70",
          1237 => x"81",
          1238 => x"51",
          1239 => x"04",
          1240 => x"0b",
          1241 => x"e8",
          1242 => x"ff",
          1243 => x"87",
          1244 => x"52",
          1245 => x"86",
          1246 => x"94",
          1247 => x"08",
          1248 => x"70",
          1249 => x"51",
          1250 => x"70",
          1251 => x"38",
          1252 => x"06",
          1253 => x"94",
          1254 => x"80",
          1255 => x"87",
          1256 => x"52",
          1257 => x"98",
          1258 => x"2c",
          1259 => x"71",
          1260 => x"0c",
          1261 => x"04",
          1262 => x"87",
          1263 => x"08",
          1264 => x"8a",
          1265 => x"70",
          1266 => x"b4",
          1267 => x"9e",
          1268 => x"f9",
          1269 => x"c0",
          1270 => x"81",
          1271 => x"87",
          1272 => x"08",
          1273 => x"0c",
          1274 => x"98",
          1275 => x"f8",
          1276 => x"9e",
          1277 => x"f9",
          1278 => x"c0",
          1279 => x"81",
          1280 => x"87",
          1281 => x"08",
          1282 => x"0c",
          1283 => x"b0",
          1284 => x"88",
          1285 => x"9e",
          1286 => x"fa",
          1287 => x"c0",
          1288 => x"81",
          1289 => x"87",
          1290 => x"08",
          1291 => x"0c",
          1292 => x"c0",
          1293 => x"98",
          1294 => x"9e",
          1295 => x"fa",
          1296 => x"c0",
          1297 => x"51",
          1298 => x"a0",
          1299 => x"9e",
          1300 => x"fa",
          1301 => x"c0",
          1302 => x"81",
          1303 => x"87",
          1304 => x"08",
          1305 => x"0c",
          1306 => x"fa",
          1307 => x"0b",
          1308 => x"90",
          1309 => x"80",
          1310 => x"52",
          1311 => x"2e",
          1312 => x"52",
          1313 => x"b1",
          1314 => x"87",
          1315 => x"08",
          1316 => x"0a",
          1317 => x"52",
          1318 => x"83",
          1319 => x"71",
          1320 => x"34",
          1321 => x"c0",
          1322 => x"70",
          1323 => x"06",
          1324 => x"70",
          1325 => x"38",
          1326 => x"81",
          1327 => x"80",
          1328 => x"9e",
          1329 => x"88",
          1330 => x"51",
          1331 => x"80",
          1332 => x"81",
          1333 => x"fa",
          1334 => x"0b",
          1335 => x"90",
          1336 => x"80",
          1337 => x"52",
          1338 => x"2e",
          1339 => x"52",
          1340 => x"b5",
          1341 => x"87",
          1342 => x"08",
          1343 => x"80",
          1344 => x"52",
          1345 => x"83",
          1346 => x"71",
          1347 => x"34",
          1348 => x"c0",
          1349 => x"70",
          1350 => x"06",
          1351 => x"70",
          1352 => x"38",
          1353 => x"81",
          1354 => x"80",
          1355 => x"9e",
          1356 => x"82",
          1357 => x"51",
          1358 => x"80",
          1359 => x"81",
          1360 => x"fa",
          1361 => x"0b",
          1362 => x"90",
          1363 => x"80",
          1364 => x"52",
          1365 => x"2e",
          1366 => x"52",
          1367 => x"b9",
          1368 => x"87",
          1369 => x"08",
          1370 => x"80",
          1371 => x"52",
          1372 => x"83",
          1373 => x"71",
          1374 => x"34",
          1375 => x"c0",
          1376 => x"70",
          1377 => x"51",
          1378 => x"80",
          1379 => x"81",
          1380 => x"fa",
          1381 => x"c0",
          1382 => x"70",
          1383 => x"70",
          1384 => x"51",
          1385 => x"fa",
          1386 => x"0b",
          1387 => x"90",
          1388 => x"80",
          1389 => x"52",
          1390 => x"83",
          1391 => x"71",
          1392 => x"34",
          1393 => x"90",
          1394 => x"f0",
          1395 => x"2a",
          1396 => x"70",
          1397 => x"34",
          1398 => x"c0",
          1399 => x"70",
          1400 => x"52",
          1401 => x"2e",
          1402 => x"52",
          1403 => x"bf",
          1404 => x"9e",
          1405 => x"87",
          1406 => x"70",
          1407 => x"34",
          1408 => x"04",
          1409 => x"81",
          1410 => x"8a",
          1411 => x"fa",
          1412 => x"73",
          1413 => x"38",
          1414 => x"51",
          1415 => x"81",
          1416 => x"8a",
          1417 => x"fa",
          1418 => x"73",
          1419 => x"38",
          1420 => x"08",
          1421 => x"08",
          1422 => x"81",
          1423 => x"8f",
          1424 => x"fa",
          1425 => x"73",
          1426 => x"38",
          1427 => x"08",
          1428 => x"08",
          1429 => x"81",
          1430 => x"8f",
          1431 => x"fa",
          1432 => x"73",
          1433 => x"38",
          1434 => x"08",
          1435 => x"08",
          1436 => x"81",
          1437 => x"8f",
          1438 => x"fa",
          1439 => x"73",
          1440 => x"38",
          1441 => x"08",
          1442 => x"08",
          1443 => x"81",
          1444 => x"8e",
          1445 => x"fa",
          1446 => x"73",
          1447 => x"38",
          1448 => x"08",
          1449 => x"08",
          1450 => x"81",
          1451 => x"8e",
          1452 => x"fa",
          1453 => x"73",
          1454 => x"38",
          1455 => x"33",
          1456 => x"b8",
          1457 => x"3f",
          1458 => x"33",
          1459 => x"2e",
          1460 => x"fa",
          1461 => x"81",
          1462 => x"8e",
          1463 => x"fa",
          1464 => x"73",
          1465 => x"38",
          1466 => x"33",
          1467 => x"f8",
          1468 => x"3f",
          1469 => x"33",
          1470 => x"2e",
          1471 => x"e5",
          1472 => x"a4",
          1473 => x"b3",
          1474 => x"80",
          1475 => x"81",
          1476 => x"88",
          1477 => x"fa",
          1478 => x"73",
          1479 => x"38",
          1480 => x"51",
          1481 => x"81",
          1482 => x"54",
          1483 => x"88",
          1484 => x"c4",
          1485 => x"3f",
          1486 => x"33",
          1487 => x"2e",
          1488 => x"e5",
          1489 => x"e0",
          1490 => x"dc",
          1491 => x"3f",
          1492 => x"08",
          1493 => x"e8",
          1494 => x"3f",
          1495 => x"08",
          1496 => x"90",
          1497 => x"3f",
          1498 => x"08",
          1499 => x"b8",
          1500 => x"3f",
          1501 => x"51",
          1502 => x"81",
          1503 => x"52",
          1504 => x"51",
          1505 => x"81",
          1506 => x"56",
          1507 => x"52",
          1508 => x"9a",
          1509 => x"f0",
          1510 => x"c0",
          1511 => x"31",
          1512 => x"fe",
          1513 => x"81",
          1514 => x"8c",
          1515 => x"fa",
          1516 => x"73",
          1517 => x"38",
          1518 => x"08",
          1519 => x"c0",
          1520 => x"e3",
          1521 => x"fe",
          1522 => x"84",
          1523 => x"71",
          1524 => x"81",
          1525 => x"52",
          1526 => x"51",
          1527 => x"81",
          1528 => x"54",
          1529 => x"a8",
          1530 => x"ac",
          1531 => x"84",
          1532 => x"51",
          1533 => x"81",
          1534 => x"bd",
          1535 => x"76",
          1536 => x"54",
          1537 => x"08",
          1538 => x"e8",
          1539 => x"3f",
          1540 => x"51",
          1541 => x"87",
          1542 => x"fe",
          1543 => x"92",
          1544 => x"05",
          1545 => x"26",
          1546 => x"84",
          1547 => x"c0",
          1548 => x"08",
          1549 => x"94",
          1550 => x"81",
          1551 => x"97",
          1552 => x"a4",
          1553 => x"81",
          1554 => x"8b",
          1555 => x"b0",
          1556 => x"81",
          1557 => x"85",
          1558 => x"3d",
          1559 => x"88",
          1560 => x"ff",
          1561 => x"c0",
          1562 => x"08",
          1563 => x"72",
          1564 => x"07",
          1565 => x"c4",
          1566 => x"83",
          1567 => x"ff",
          1568 => x"c0",
          1569 => x"08",
          1570 => x"0c",
          1571 => x"0c",
          1572 => x"81",
          1573 => x"06",
          1574 => x"c4",
          1575 => x"51",
          1576 => x"04",
          1577 => x"c0",
          1578 => x"04",
          1579 => x"08",
          1580 => x"84",
          1581 => x"3d",
          1582 => x"80",
          1583 => x"82",
          1584 => x"81",
          1585 => x"81",
          1586 => x"75",
          1587 => x"ff",
          1588 => x"b7",
          1589 => x"38",
          1590 => x"80",
          1591 => x"72",
          1592 => x"0c",
          1593 => x"04",
          1594 => x"79",
          1595 => x"08",
          1596 => x"14",
          1597 => x"08",
          1598 => x"5a",
          1599 => x"57",
          1600 => x"26",
          1601 => x"13",
          1602 => x"53",
          1603 => x"0c",
          1604 => x"84",
          1605 => x"73",
          1606 => x"14",
          1607 => x"12",
          1608 => x"12",
          1609 => x"13",
          1610 => x"14",
          1611 => x"12",
          1612 => x"12",
          1613 => x"15",
          1614 => x"16",
          1615 => x"80",
          1616 => x"90",
          1617 => x"94",
          1618 => x"81",
          1619 => x"89",
          1620 => x"fc",
          1621 => x"8c",
          1622 => x"12",
          1623 => x"53",
          1624 => x"2e",
          1625 => x"a3",
          1626 => x"08",
          1627 => x"55",
          1628 => x"09",
          1629 => x"38",
          1630 => x"15",
          1631 => x"73",
          1632 => x"71",
          1633 => x"71",
          1634 => x"81",
          1635 => x"fa",
          1636 => x"14",
          1637 => x"c8",
          1638 => x"0c",
          1639 => x"d8",
          1640 => x"08",
          1641 => x"0c",
          1642 => x"81",
          1643 => x"06",
          1644 => x"13",
          1645 => x"52",
          1646 => x"2e",
          1647 => x"a4",
          1648 => x"08",
          1649 => x"0c",
          1650 => x"90",
          1651 => x"90",
          1652 => x"94",
          1653 => x"14",
          1654 => x"08",
          1655 => x"0c",
          1656 => x"0c",
          1657 => x"f0",
          1658 => x"0d",
          1659 => x"0d",
          1660 => x"57",
          1661 => x"81",
          1662 => x"17",
          1663 => x"fa",
          1664 => x"57",
          1665 => x"2e",
          1666 => x"16",
          1667 => x"80",
          1668 => x"16",
          1669 => x"39",
          1670 => x"17",
          1671 => x"06",
          1672 => x"fd",
          1673 => x"fe",
          1674 => x"fe",
          1675 => x"70",
          1676 => x"08",
          1677 => x"81",
          1678 => x"09",
          1679 => x"72",
          1680 => x"73",
          1681 => x"58",
          1682 => x"80",
          1683 => x"2e",
          1684 => x"80",
          1685 => x"39",
          1686 => x"51",
          1687 => x"81",
          1688 => x"f0",
          1689 => x"81",
          1690 => x"84",
          1691 => x"fa",
          1692 => x"72",
          1693 => x"8c",
          1694 => x"26",
          1695 => x"13",
          1696 => x"39",
          1697 => x"88",
          1698 => x"8c",
          1699 => x"88",
          1700 => x"16",
          1701 => x"12",
          1702 => x"51",
          1703 => x"76",
          1704 => x"f0",
          1705 => x"c0",
          1706 => x"f0",
          1707 => x"81",
          1708 => x"89",
          1709 => x"ff",
          1710 => x"52",
          1711 => x"87",
          1712 => x"51",
          1713 => x"83",
          1714 => x"fe",
          1715 => x"93",
          1716 => x"72",
          1717 => x"81",
          1718 => x"8d",
          1719 => x"81",
          1720 => x"52",
          1721 => x"90",
          1722 => x"34",
          1723 => x"08",
          1724 => x"ff",
          1725 => x"39",
          1726 => x"08",
          1727 => x"2e",
          1728 => x"51",
          1729 => x"3d",
          1730 => x"3d",
          1731 => x"05",
          1732 => x"84",
          1733 => x"ff",
          1734 => x"51",
          1735 => x"72",
          1736 => x"0c",
          1737 => x"04",
          1738 => x"75",
          1739 => x"70",
          1740 => x"53",
          1741 => x"2e",
          1742 => x"81",
          1743 => x"81",
          1744 => x"87",
          1745 => x"85",
          1746 => x"fc",
          1747 => x"81",
          1748 => x"78",
          1749 => x"0c",
          1750 => x"33",
          1751 => x"06",
          1752 => x"80",
          1753 => x"72",
          1754 => x"51",
          1755 => x"fe",
          1756 => x"39",
          1757 => x"84",
          1758 => x"0d",
          1759 => x"0d",
          1760 => x"59",
          1761 => x"05",
          1762 => x"75",
          1763 => x"f8",
          1764 => x"2e",
          1765 => x"82",
          1766 => x"70",
          1767 => x"05",
          1768 => x"5b",
          1769 => x"2e",
          1770 => x"85",
          1771 => x"8b",
          1772 => x"2e",
          1773 => x"8a",
          1774 => x"78",
          1775 => x"5a",
          1776 => x"aa",
          1777 => x"06",
          1778 => x"84",
          1779 => x"7b",
          1780 => x"5d",
          1781 => x"59",
          1782 => x"d0",
          1783 => x"89",
          1784 => x"7a",
          1785 => x"10",
          1786 => x"d0",
          1787 => x"81",
          1788 => x"57",
          1789 => x"75",
          1790 => x"70",
          1791 => x"07",
          1792 => x"80",
          1793 => x"30",
          1794 => x"80",
          1795 => x"53",
          1796 => x"55",
          1797 => x"2e",
          1798 => x"84",
          1799 => x"81",
          1800 => x"57",
          1801 => x"2e",
          1802 => x"75",
          1803 => x"76",
          1804 => x"e0",
          1805 => x"ff",
          1806 => x"73",
          1807 => x"81",
          1808 => x"80",
          1809 => x"38",
          1810 => x"2e",
          1811 => x"73",
          1812 => x"8b",
          1813 => x"c2",
          1814 => x"38",
          1815 => x"73",
          1816 => x"81",
          1817 => x"8f",
          1818 => x"d5",
          1819 => x"38",
          1820 => x"24",
          1821 => x"80",
          1822 => x"38",
          1823 => x"73",
          1824 => x"80",
          1825 => x"ef",
          1826 => x"19",
          1827 => x"59",
          1828 => x"33",
          1829 => x"75",
          1830 => x"81",
          1831 => x"70",
          1832 => x"55",
          1833 => x"79",
          1834 => x"90",
          1835 => x"16",
          1836 => x"7b",
          1837 => x"a0",
          1838 => x"3f",
          1839 => x"53",
          1840 => x"e9",
          1841 => x"fc",
          1842 => x"81",
          1843 => x"72",
          1844 => x"b0",
          1845 => x"fb",
          1846 => x"39",
          1847 => x"83",
          1848 => x"59",
          1849 => x"82",
          1850 => x"88",
          1851 => x"8a",
          1852 => x"90",
          1853 => x"75",
          1854 => x"3f",
          1855 => x"79",
          1856 => x"81",
          1857 => x"72",
          1858 => x"38",
          1859 => x"59",
          1860 => x"84",
          1861 => x"58",
          1862 => x"80",
          1863 => x"30",
          1864 => x"80",
          1865 => x"55",
          1866 => x"25",
          1867 => x"80",
          1868 => x"74",
          1869 => x"07",
          1870 => x"0b",
          1871 => x"57",
          1872 => x"51",
          1873 => x"81",
          1874 => x"81",
          1875 => x"53",
          1876 => x"d8",
          1877 => x"fe",
          1878 => x"89",
          1879 => x"38",
          1880 => x"75",
          1881 => x"84",
          1882 => x"53",
          1883 => x"06",
          1884 => x"53",
          1885 => x"81",
          1886 => x"81",
          1887 => x"70",
          1888 => x"2a",
          1889 => x"76",
          1890 => x"38",
          1891 => x"38",
          1892 => x"70",
          1893 => x"53",
          1894 => x"8e",
          1895 => x"77",
          1896 => x"53",
          1897 => x"81",
          1898 => x"7a",
          1899 => x"55",
          1900 => x"83",
          1901 => x"79",
          1902 => x"81",
          1903 => x"72",
          1904 => x"17",
          1905 => x"27",
          1906 => x"51",
          1907 => x"75",
          1908 => x"72",
          1909 => x"81",
          1910 => x"7a",
          1911 => x"38",
          1912 => x"05",
          1913 => x"ff",
          1914 => x"70",
          1915 => x"57",
          1916 => x"76",
          1917 => x"81",
          1918 => x"72",
          1919 => x"84",
          1920 => x"f9",
          1921 => x"39",
          1922 => x"04",
          1923 => x"86",
          1924 => x"84",
          1925 => x"55",
          1926 => x"fa",
          1927 => x"3d",
          1928 => x"3d",
          1929 => x"ff",
          1930 => x"3d",
          1931 => x"75",
          1932 => x"3f",
          1933 => x"08",
          1934 => x"34",
          1935 => x"ff",
          1936 => x"3d",
          1937 => x"3d",
          1938 => x"84",
          1939 => x"ff",
          1940 => x"3d",
          1941 => x"77",
          1942 => x"a1",
          1943 => x"ff",
          1944 => x"3d",
          1945 => x"3d",
          1946 => x"81",
          1947 => x"70",
          1948 => x"55",
          1949 => x"80",
          1950 => x"38",
          1951 => x"08",
          1952 => x"81",
          1953 => x"81",
          1954 => x"72",
          1955 => x"cb",
          1956 => x"2e",
          1957 => x"88",
          1958 => x"70",
          1959 => x"51",
          1960 => x"2e",
          1961 => x"80",
          1962 => x"ff",
          1963 => x"39",
          1964 => x"c8",
          1965 => x"52",
          1966 => x"c0",
          1967 => x"52",
          1968 => x"81",
          1969 => x"51",
          1970 => x"ff",
          1971 => x"15",
          1972 => x"34",
          1973 => x"f3",
          1974 => x"72",
          1975 => x"0c",
          1976 => x"04",
          1977 => x"81",
          1978 => x"75",
          1979 => x"0c",
          1980 => x"52",
          1981 => x"3f",
          1982 => x"88",
          1983 => x"0d",
          1984 => x"0d",
          1985 => x"56",
          1986 => x"0c",
          1987 => x"70",
          1988 => x"73",
          1989 => x"81",
          1990 => x"81",
          1991 => x"ed",
          1992 => x"2e",
          1993 => x"8e",
          1994 => x"08",
          1995 => x"76",
          1996 => x"56",
          1997 => x"b0",
          1998 => x"06",
          1999 => x"75",
          2000 => x"76",
          2001 => x"70",
          2002 => x"73",
          2003 => x"8b",
          2004 => x"73",
          2005 => x"85",
          2006 => x"82",
          2007 => x"76",
          2008 => x"70",
          2009 => x"ac",
          2010 => x"a0",
          2011 => x"fa",
          2012 => x"53",
          2013 => x"57",
          2014 => x"98",
          2015 => x"39",
          2016 => x"80",
          2017 => x"26",
          2018 => x"86",
          2019 => x"80",
          2020 => x"57",
          2021 => x"74",
          2022 => x"38",
          2023 => x"27",
          2024 => x"14",
          2025 => x"06",
          2026 => x"14",
          2027 => x"06",
          2028 => x"74",
          2029 => x"f9",
          2030 => x"ff",
          2031 => x"89",
          2032 => x"38",
          2033 => x"c5",
          2034 => x"29",
          2035 => x"81",
          2036 => x"76",
          2037 => x"56",
          2038 => x"ba",
          2039 => x"2e",
          2040 => x"30",
          2041 => x"0c",
          2042 => x"81",
          2043 => x"8a",
          2044 => x"f8",
          2045 => x"7c",
          2046 => x"70",
          2047 => x"75",
          2048 => x"55",
          2049 => x"2e",
          2050 => x"87",
          2051 => x"76",
          2052 => x"73",
          2053 => x"81",
          2054 => x"81",
          2055 => x"77",
          2056 => x"70",
          2057 => x"58",
          2058 => x"09",
          2059 => x"c2",
          2060 => x"81",
          2061 => x"75",
          2062 => x"55",
          2063 => x"e2",
          2064 => x"90",
          2065 => x"f8",
          2066 => x"8f",
          2067 => x"81",
          2068 => x"75",
          2069 => x"55",
          2070 => x"81",
          2071 => x"27",
          2072 => x"d0",
          2073 => x"55",
          2074 => x"73",
          2075 => x"80",
          2076 => x"14",
          2077 => x"72",
          2078 => x"e0",
          2079 => x"80",
          2080 => x"39",
          2081 => x"55",
          2082 => x"80",
          2083 => x"e0",
          2084 => x"38",
          2085 => x"81",
          2086 => x"53",
          2087 => x"81",
          2088 => x"53",
          2089 => x"8e",
          2090 => x"70",
          2091 => x"55",
          2092 => x"27",
          2093 => x"77",
          2094 => x"74",
          2095 => x"76",
          2096 => x"77",
          2097 => x"70",
          2098 => x"55",
          2099 => x"77",
          2100 => x"38",
          2101 => x"74",
          2102 => x"55",
          2103 => x"f0",
          2104 => x"0d",
          2105 => x"0d",
          2106 => x"70",
          2107 => x"98",
          2108 => x"2c",
          2109 => x"70",
          2110 => x"53",
          2111 => x"51",
          2112 => x"e9",
          2113 => x"55",
          2114 => x"25",
          2115 => x"e9",
          2116 => x"12",
          2117 => x"97",
          2118 => x"33",
          2119 => x"70",
          2120 => x"81",
          2121 => x"81",
          2122 => x"fe",
          2123 => x"3d",
          2124 => x"3d",
          2125 => x"84",
          2126 => x"33",
          2127 => x"55",
          2128 => x"2e",
          2129 => x"51",
          2130 => x"a0",
          2131 => x"3f",
          2132 => x"f7",
          2133 => x"ff",
          2134 => x"73",
          2135 => x"ff",
          2136 => x"39",
          2137 => x"c0",
          2138 => x"34",
          2139 => x"04",
          2140 => x"7c",
          2141 => x"b7",
          2142 => x"88",
          2143 => x"33",
          2144 => x"33",
          2145 => x"81",
          2146 => x"70",
          2147 => x"59",
          2148 => x"74",
          2149 => x"38",
          2150 => x"9b",
          2151 => x"bc",
          2152 => x"29",
          2153 => x"05",
          2154 => x"54",
          2155 => x"f0",
          2156 => x"fe",
          2157 => x"0c",
          2158 => x"33",
          2159 => x"81",
          2160 => x"70",
          2161 => x"5a",
          2162 => x"a6",
          2163 => x"78",
          2164 => x"d5",
          2165 => x"fb",
          2166 => x"05",
          2167 => x"fb",
          2168 => x"81",
          2169 => x"93",
          2170 => x"38",
          2171 => x"fb",
          2172 => x"80",
          2173 => x"81",
          2174 => x"56",
          2175 => x"ac",
          2176 => x"b4",
          2177 => x"a4",
          2178 => x"fc",
          2179 => x"53",
          2180 => x"51",
          2181 => x"3f",
          2182 => x"08",
          2183 => x"80",
          2184 => x"81",
          2185 => x"51",
          2186 => x"3f",
          2187 => x"04",
          2188 => x"81",
          2189 => x"81",
          2190 => x"51",
          2191 => x"3f",
          2192 => x"08",
          2193 => x"81",
          2194 => x"53",
          2195 => x"88",
          2196 => x"56",
          2197 => x"3f",
          2198 => x"08",
          2199 => x"38",
          2200 => x"ec",
          2201 => x"f0",
          2202 => x"0b",
          2203 => x"08",
          2204 => x"81",
          2205 => x"ff",
          2206 => x"55",
          2207 => x"34",
          2208 => x"52",
          2209 => x"e8",
          2210 => x"f6",
          2211 => x"ff",
          2212 => x"06",
          2213 => x"a6",
          2214 => x"d9",
          2215 => x"3d",
          2216 => x"08",
          2217 => x"70",
          2218 => x"52",
          2219 => x"08",
          2220 => x"92",
          2221 => x"f0",
          2222 => x"38",
          2223 => x"fb",
          2224 => x"55",
          2225 => x"8b",
          2226 => x"56",
          2227 => x"3f",
          2228 => x"08",
          2229 => x"38",
          2230 => x"f4",
          2231 => x"f0",
          2232 => x"58",
          2233 => x"81",
          2234 => x"25",
          2235 => x"fe",
          2236 => x"05",
          2237 => x"55",
          2238 => x"74",
          2239 => x"70",
          2240 => x"2a",
          2241 => x"78",
          2242 => x"38",
          2243 => x"38",
          2244 => x"08",
          2245 => x"53",
          2246 => x"aa",
          2247 => x"f0",
          2248 => x"88",
          2249 => x"ec",
          2250 => x"3f",
          2251 => x"09",
          2252 => x"38",
          2253 => x"51",
          2254 => x"79",
          2255 => x"3f",
          2256 => x"54",
          2257 => x"08",
          2258 => x"58",
          2259 => x"f0",
          2260 => x"0d",
          2261 => x"0d",
          2262 => x"5c",
          2263 => x"57",
          2264 => x"73",
          2265 => x"81",
          2266 => x"78",
          2267 => x"56",
          2268 => x"98",
          2269 => x"70",
          2270 => x"33",
          2271 => x"73",
          2272 => x"81",
          2273 => x"75",
          2274 => x"38",
          2275 => x"88",
          2276 => x"c0",
          2277 => x"52",
          2278 => x"3f",
          2279 => x"08",
          2280 => x"74",
          2281 => x"89",
          2282 => x"f0",
          2283 => x"38",
          2284 => x"55",
          2285 => x"88",
          2286 => x"2e",
          2287 => x"39",
          2288 => x"ab",
          2289 => x"5a",
          2290 => x"11",
          2291 => x"51",
          2292 => x"81",
          2293 => x"80",
          2294 => x"7a",
          2295 => x"77",
          2296 => x"3f",
          2297 => x"08",
          2298 => x"55",
          2299 => x"74",
          2300 => x"81",
          2301 => x"ff",
          2302 => x"82",
          2303 => x"8e",
          2304 => x"73",
          2305 => x"0c",
          2306 => x"04",
          2307 => x"b0",
          2308 => x"84",
          2309 => x"05",
          2310 => x"80",
          2311 => x"34",
          2312 => x"33",
          2313 => x"b8",
          2314 => x"38",
          2315 => x"33",
          2316 => x"9a",
          2317 => x"eb",
          2318 => x"fe",
          2319 => x"fb",
          2320 => x"fe",
          2321 => x"2e",
          2322 => x"93",
          2323 => x"e0",
          2324 => x"fe",
          2325 => x"bb",
          2326 => x"fe",
          2327 => x"2e",
          2328 => x"e9",
          2329 => x"a4",
          2330 => x"39",
          2331 => x"08",
          2332 => x"52",
          2333 => x"52",
          2334 => x"b0",
          2335 => x"f0",
          2336 => x"fe",
          2337 => x"2e",
          2338 => x"80",
          2339 => x"fe",
          2340 => x"d3",
          2341 => x"fe",
          2342 => x"80",
          2343 => x"f0",
          2344 => x"38",
          2345 => x"08",
          2346 => x"17",
          2347 => x"74",
          2348 => x"74",
          2349 => x"52",
          2350 => x"b4",
          2351 => x"2e",
          2352 => x"ff",
          2353 => x"39",
          2354 => x"fb",
          2355 => x"3d",
          2356 => x"3f",
          2357 => x"08",
          2358 => x"98",
          2359 => x"78",
          2360 => x"38",
          2361 => x"06",
          2362 => x"33",
          2363 => x"70",
          2364 => x"ff",
          2365 => x"98",
          2366 => x"2c",
          2367 => x"05",
          2368 => x"81",
          2369 => x"70",
          2370 => x"33",
          2371 => x"51",
          2372 => x"59",
          2373 => x"56",
          2374 => x"80",
          2375 => x"74",
          2376 => x"74",
          2377 => x"29",
          2378 => x"05",
          2379 => x"51",
          2380 => x"24",
          2381 => x"76",
          2382 => x"77",
          2383 => x"3f",
          2384 => x"08",
          2385 => x"54",
          2386 => x"d7",
          2387 => x"ff",
          2388 => x"56",
          2389 => x"81",
          2390 => x"81",
          2391 => x"70",
          2392 => x"81",
          2393 => x"51",
          2394 => x"26",
          2395 => x"53",
          2396 => x"51",
          2397 => x"81",
          2398 => x"81",
          2399 => x"73",
          2400 => x"39",
          2401 => x"80",
          2402 => x"38",
          2403 => x"74",
          2404 => x"34",
          2405 => x"70",
          2406 => x"ff",
          2407 => x"98",
          2408 => x"2c",
          2409 => x"70",
          2410 => x"e9",
          2411 => x"5e",
          2412 => x"57",
          2413 => x"74",
          2414 => x"81",
          2415 => x"38",
          2416 => x"14",
          2417 => x"80",
          2418 => x"94",
          2419 => x"81",
          2420 => x"92",
          2421 => x"ff",
          2422 => x"81",
          2423 => x"78",
          2424 => x"75",
          2425 => x"54",
          2426 => x"fd",
          2427 => x"84",
          2428 => x"d4",
          2429 => x"08",
          2430 => x"9c",
          2431 => x"7e",
          2432 => x"38",
          2433 => x"33",
          2434 => x"27",
          2435 => x"98",
          2436 => x"2c",
          2437 => x"75",
          2438 => x"74",
          2439 => x"33",
          2440 => x"74",
          2441 => x"29",
          2442 => x"05",
          2443 => x"81",
          2444 => x"56",
          2445 => x"39",
          2446 => x"33",
          2447 => x"54",
          2448 => x"9c",
          2449 => x"54",
          2450 => x"74",
          2451 => x"98",
          2452 => x"7e",
          2453 => x"81",
          2454 => x"81",
          2455 => x"81",
          2456 => x"70",
          2457 => x"29",
          2458 => x"05",
          2459 => x"81",
          2460 => x"5a",
          2461 => x"74",
          2462 => x"38",
          2463 => x"33",
          2464 => x"c7",
          2465 => x"80",
          2466 => x"80",
          2467 => x"98",
          2468 => x"98",
          2469 => x"55",
          2470 => x"e0",
          2471 => x"9c",
          2472 => x"2b",
          2473 => x"81",
          2474 => x"5a",
          2475 => x"74",
          2476 => x"9a",
          2477 => x"e8",
          2478 => x"81",
          2479 => x"81",
          2480 => x"70",
          2481 => x"ff",
          2482 => x"51",
          2483 => x"24",
          2484 => x"fa",
          2485 => x"9c",
          2486 => x"ff",
          2487 => x"73",
          2488 => x"ea",
          2489 => x"98",
          2490 => x"54",
          2491 => x"98",
          2492 => x"54",
          2493 => x"9c",
          2494 => x"e7",
          2495 => x"ff",
          2496 => x"98",
          2497 => x"2c",
          2498 => x"33",
          2499 => x"57",
          2500 => x"a7",
          2501 => x"54",
          2502 => x"74",
          2503 => x"51",
          2504 => x"74",
          2505 => x"29",
          2506 => x"05",
          2507 => x"81",
          2508 => x"58",
          2509 => x"75",
          2510 => x"a0",
          2511 => x"3f",
          2512 => x"33",
          2513 => x"70",
          2514 => x"ff",
          2515 => x"51",
          2516 => x"74",
          2517 => x"38",
          2518 => x"ef",
          2519 => x"80",
          2520 => x"80",
          2521 => x"98",
          2522 => x"98",
          2523 => x"55",
          2524 => x"e4",
          2525 => x"39",
          2526 => x"33",
          2527 => x"80",
          2528 => x"51",
          2529 => x"81",
          2530 => x"79",
          2531 => x"3f",
          2532 => x"08",
          2533 => x"54",
          2534 => x"81",
          2535 => x"54",
          2536 => x"84",
          2537 => x"53",
          2538 => x"51",
          2539 => x"84",
          2540 => x"7a",
          2541 => x"39",
          2542 => x"33",
          2543 => x"2e",
          2544 => x"88",
          2545 => x"3f",
          2546 => x"33",
          2547 => x"73",
          2548 => x"34",
          2549 => x"06",
          2550 => x"81",
          2551 => x"81",
          2552 => x"55",
          2553 => x"2e",
          2554 => x"ff",
          2555 => x"81",
          2556 => x"74",
          2557 => x"98",
          2558 => x"ff",
          2559 => x"55",
          2560 => x"a7",
          2561 => x"54",
          2562 => x"74",
          2563 => x"51",
          2564 => x"74",
          2565 => x"29",
          2566 => x"05",
          2567 => x"81",
          2568 => x"58",
          2569 => x"75",
          2570 => x"a0",
          2571 => x"3f",
          2572 => x"33",
          2573 => x"70",
          2574 => x"ff",
          2575 => x"51",
          2576 => x"74",
          2577 => x"38",
          2578 => x"ff",
          2579 => x"80",
          2580 => x"80",
          2581 => x"98",
          2582 => x"98",
          2583 => x"55",
          2584 => x"e4",
          2585 => x"39",
          2586 => x"33",
          2587 => x"06",
          2588 => x"33",
          2589 => x"74",
          2590 => x"d2",
          2591 => x"54",
          2592 => x"9c",
          2593 => x"70",
          2594 => x"e4",
          2595 => x"ff",
          2596 => x"81",
          2597 => x"ff",
          2598 => x"56",
          2599 => x"26",
          2600 => x"aa",
          2601 => x"38",
          2602 => x"08",
          2603 => x"2e",
          2604 => x"51",
          2605 => x"81",
          2606 => x"81",
          2607 => x"81",
          2608 => x"81",
          2609 => x"05",
          2610 => x"79",
          2611 => x"3f",
          2612 => x"c1",
          2613 => x"29",
          2614 => x"05",
          2615 => x"56",
          2616 => x"2e",
          2617 => x"51",
          2618 => x"81",
          2619 => x"81",
          2620 => x"81",
          2621 => x"81",
          2622 => x"05",
          2623 => x"79",
          2624 => x"3f",
          2625 => x"80",
          2626 => x"08",
          2627 => x"2e",
          2628 => x"74",
          2629 => x"3f",
          2630 => x"7a",
          2631 => x"81",
          2632 => x"81",
          2633 => x"55",
          2634 => x"89",
          2635 => x"ca",
          2636 => x"c8",
          2637 => x"29",
          2638 => x"05",
          2639 => x"56",
          2640 => x"2e",
          2641 => x"51",
          2642 => x"81",
          2643 => x"81",
          2644 => x"81",
          2645 => x"81",
          2646 => x"05",
          2647 => x"79",
          2648 => x"3f",
          2649 => x"73",
          2650 => x"5b",
          2651 => x"08",
          2652 => x"2e",
          2653 => x"74",
          2654 => x"3f",
          2655 => x"08",
          2656 => x"34",
          2657 => x"08",
          2658 => x"81",
          2659 => x"52",
          2660 => x"a1",
          2661 => x"9c",
          2662 => x"98",
          2663 => x"51",
          2664 => x"f6",
          2665 => x"ff",
          2666 => x"81",
          2667 => x"ff",
          2668 => x"56",
          2669 => x"27",
          2670 => x"81",
          2671 => x"81",
          2672 => x"74",
          2673 => x"52",
          2674 => x"3f",
          2675 => x"81",
          2676 => x"54",
          2677 => x"f5",
          2678 => x"51",
          2679 => x"81",
          2680 => x"ff",
          2681 => x"81",
          2682 => x"f5",
          2683 => x"0b",
          2684 => x"34",
          2685 => x"ff",
          2686 => x"81",
          2687 => x"af",
          2688 => x"ff",
          2689 => x"8f",
          2690 => x"81",
          2691 => x"26",
          2692 => x"fb",
          2693 => x"52",
          2694 => x"f0",
          2695 => x"0d",
          2696 => x"0d",
          2697 => x"33",
          2698 => x"9f",
          2699 => x"53",
          2700 => x"81",
          2701 => x"38",
          2702 => x"87",
          2703 => x"11",
          2704 => x"54",
          2705 => x"84",
          2706 => x"54",
          2707 => x"87",
          2708 => x"11",
          2709 => x"0c",
          2710 => x"c0",
          2711 => x"70",
          2712 => x"70",
          2713 => x"51",
          2714 => x"8a",
          2715 => x"98",
          2716 => x"70",
          2717 => x"08",
          2718 => x"06",
          2719 => x"38",
          2720 => x"8c",
          2721 => x"80",
          2722 => x"71",
          2723 => x"14",
          2724 => x"d8",
          2725 => x"70",
          2726 => x"0c",
          2727 => x"04",
          2728 => x"60",
          2729 => x"8c",
          2730 => x"33",
          2731 => x"5b",
          2732 => x"5a",
          2733 => x"81",
          2734 => x"81",
          2735 => x"52",
          2736 => x"38",
          2737 => x"84",
          2738 => x"92",
          2739 => x"c0",
          2740 => x"87",
          2741 => x"13",
          2742 => x"57",
          2743 => x"0b",
          2744 => x"8c",
          2745 => x"0c",
          2746 => x"75",
          2747 => x"2a",
          2748 => x"51",
          2749 => x"80",
          2750 => x"7b",
          2751 => x"7b",
          2752 => x"5d",
          2753 => x"59",
          2754 => x"06",
          2755 => x"73",
          2756 => x"81",
          2757 => x"ff",
          2758 => x"72",
          2759 => x"38",
          2760 => x"8c",
          2761 => x"c3",
          2762 => x"98",
          2763 => x"71",
          2764 => x"38",
          2765 => x"2e",
          2766 => x"76",
          2767 => x"92",
          2768 => x"72",
          2769 => x"06",
          2770 => x"f7",
          2771 => x"5a",
          2772 => x"80",
          2773 => x"70",
          2774 => x"5a",
          2775 => x"80",
          2776 => x"73",
          2777 => x"06",
          2778 => x"38",
          2779 => x"fe",
          2780 => x"fc",
          2781 => x"52",
          2782 => x"83",
          2783 => x"71",
          2784 => x"fe",
          2785 => x"3d",
          2786 => x"3d",
          2787 => x"64",
          2788 => x"bf",
          2789 => x"40",
          2790 => x"59",
          2791 => x"58",
          2792 => x"81",
          2793 => x"81",
          2794 => x"52",
          2795 => x"09",
          2796 => x"b1",
          2797 => x"84",
          2798 => x"92",
          2799 => x"c0",
          2800 => x"87",
          2801 => x"13",
          2802 => x"56",
          2803 => x"87",
          2804 => x"0c",
          2805 => x"82",
          2806 => x"58",
          2807 => x"84",
          2808 => x"06",
          2809 => x"71",
          2810 => x"38",
          2811 => x"05",
          2812 => x"0c",
          2813 => x"73",
          2814 => x"81",
          2815 => x"71",
          2816 => x"38",
          2817 => x"8c",
          2818 => x"d0",
          2819 => x"98",
          2820 => x"71",
          2821 => x"38",
          2822 => x"2e",
          2823 => x"76",
          2824 => x"92",
          2825 => x"72",
          2826 => x"06",
          2827 => x"f7",
          2828 => x"59",
          2829 => x"1a",
          2830 => x"06",
          2831 => x"59",
          2832 => x"80",
          2833 => x"73",
          2834 => x"06",
          2835 => x"38",
          2836 => x"fe",
          2837 => x"fc",
          2838 => x"52",
          2839 => x"83",
          2840 => x"71",
          2841 => x"fe",
          2842 => x"3d",
          2843 => x"3d",
          2844 => x"84",
          2845 => x"33",
          2846 => x"a7",
          2847 => x"54",
          2848 => x"fa",
          2849 => x"fe",
          2850 => x"06",
          2851 => x"72",
          2852 => x"85",
          2853 => x"98",
          2854 => x"56",
          2855 => x"80",
          2856 => x"76",
          2857 => x"74",
          2858 => x"c0",
          2859 => x"54",
          2860 => x"2e",
          2861 => x"d4",
          2862 => x"2e",
          2863 => x"80",
          2864 => x"08",
          2865 => x"70",
          2866 => x"51",
          2867 => x"2e",
          2868 => x"c0",
          2869 => x"52",
          2870 => x"87",
          2871 => x"08",
          2872 => x"38",
          2873 => x"87",
          2874 => x"14",
          2875 => x"70",
          2876 => x"52",
          2877 => x"96",
          2878 => x"92",
          2879 => x"0a",
          2880 => x"39",
          2881 => x"0c",
          2882 => x"39",
          2883 => x"54",
          2884 => x"f0",
          2885 => x"0d",
          2886 => x"0d",
          2887 => x"33",
          2888 => x"88",
          2889 => x"fe",
          2890 => x"51",
          2891 => x"04",
          2892 => x"75",
          2893 => x"82",
          2894 => x"90",
          2895 => x"2b",
          2896 => x"33",
          2897 => x"88",
          2898 => x"71",
          2899 => x"f0",
          2900 => x"54",
          2901 => x"85",
          2902 => x"ff",
          2903 => x"02",
          2904 => x"05",
          2905 => x"70",
          2906 => x"05",
          2907 => x"88",
          2908 => x"72",
          2909 => x"0d",
          2910 => x"0d",
          2911 => x"52",
          2912 => x"81",
          2913 => x"70",
          2914 => x"70",
          2915 => x"05",
          2916 => x"88",
          2917 => x"72",
          2918 => x"54",
          2919 => x"2a",
          2920 => x"34",
          2921 => x"04",
          2922 => x"76",
          2923 => x"54",
          2924 => x"2e",
          2925 => x"70",
          2926 => x"33",
          2927 => x"05",
          2928 => x"11",
          2929 => x"84",
          2930 => x"fe",
          2931 => x"77",
          2932 => x"53",
          2933 => x"81",
          2934 => x"ff",
          2935 => x"f4",
          2936 => x"0d",
          2937 => x"0d",
          2938 => x"56",
          2939 => x"70",
          2940 => x"33",
          2941 => x"05",
          2942 => x"71",
          2943 => x"56",
          2944 => x"72",
          2945 => x"38",
          2946 => x"e2",
          2947 => x"fe",
          2948 => x"3d",
          2949 => x"3d",
          2950 => x"54",
          2951 => x"71",
          2952 => x"38",
          2953 => x"70",
          2954 => x"f3",
          2955 => x"81",
          2956 => x"84",
          2957 => x"80",
          2958 => x"f0",
          2959 => x"0b",
          2960 => x"0c",
          2961 => x"0d",
          2962 => x"0b",
          2963 => x"56",
          2964 => x"2e",
          2965 => x"81",
          2966 => x"08",
          2967 => x"70",
          2968 => x"33",
          2969 => x"a2",
          2970 => x"f0",
          2971 => x"09",
          2972 => x"38",
          2973 => x"08",
          2974 => x"b0",
          2975 => x"a4",
          2976 => x"9c",
          2977 => x"56",
          2978 => x"27",
          2979 => x"16",
          2980 => x"82",
          2981 => x"06",
          2982 => x"54",
          2983 => x"78",
          2984 => x"33",
          2985 => x"3f",
          2986 => x"5a",
          2987 => x"f0",
          2988 => x"0d",
          2989 => x"0d",
          2990 => x"56",
          2991 => x"b0",
          2992 => x"af",
          2993 => x"fe",
          2994 => x"fe",
          2995 => x"81",
          2996 => x"9f",
          2997 => x"74",
          2998 => x"52",
          2999 => x"51",
          3000 => x"81",
          3001 => x"80",
          3002 => x"ff",
          3003 => x"74",
          3004 => x"76",
          3005 => x"0c",
          3006 => x"04",
          3007 => x"7a",
          3008 => x"fe",
          3009 => x"fe",
          3010 => x"81",
          3011 => x"81",
          3012 => x"33",
          3013 => x"2e",
          3014 => x"80",
          3015 => x"17",
          3016 => x"81",
          3017 => x"06",
          3018 => x"84",
          3019 => x"fe",
          3020 => x"b4",
          3021 => x"56",
          3022 => x"82",
          3023 => x"84",
          3024 => x"fc",
          3025 => x"8b",
          3026 => x"52",
          3027 => x"a9",
          3028 => x"85",
          3029 => x"84",
          3030 => x"fc",
          3031 => x"17",
          3032 => x"9c",
          3033 => x"91",
          3034 => x"08",
          3035 => x"17",
          3036 => x"3f",
          3037 => x"81",
          3038 => x"19",
          3039 => x"53",
          3040 => x"17",
          3041 => x"82",
          3042 => x"18",
          3043 => x"80",
          3044 => x"33",
          3045 => x"3f",
          3046 => x"08",
          3047 => x"38",
          3048 => x"81",
          3049 => x"8a",
          3050 => x"fb",
          3051 => x"fe",
          3052 => x"08",
          3053 => x"56",
          3054 => x"74",
          3055 => x"38",
          3056 => x"75",
          3057 => x"16",
          3058 => x"53",
          3059 => x"f0",
          3060 => x"0d",
          3061 => x"0d",
          3062 => x"08",
          3063 => x"81",
          3064 => x"df",
          3065 => x"15",
          3066 => x"d7",
          3067 => x"33",
          3068 => x"82",
          3069 => x"38",
          3070 => x"89",
          3071 => x"2e",
          3072 => x"bf",
          3073 => x"2e",
          3074 => x"81",
          3075 => x"81",
          3076 => x"89",
          3077 => x"08",
          3078 => x"52",
          3079 => x"3f",
          3080 => x"08",
          3081 => x"74",
          3082 => x"14",
          3083 => x"81",
          3084 => x"2a",
          3085 => x"05",
          3086 => x"57",
          3087 => x"f5",
          3088 => x"f0",
          3089 => x"38",
          3090 => x"06",
          3091 => x"33",
          3092 => x"78",
          3093 => x"06",
          3094 => x"5c",
          3095 => x"53",
          3096 => x"38",
          3097 => x"06",
          3098 => x"39",
          3099 => x"a4",
          3100 => x"52",
          3101 => x"bd",
          3102 => x"f0",
          3103 => x"38",
          3104 => x"fe",
          3105 => x"b4",
          3106 => x"8d",
          3107 => x"f0",
          3108 => x"ff",
          3109 => x"39",
          3110 => x"a4",
          3111 => x"52",
          3112 => x"91",
          3113 => x"f0",
          3114 => x"76",
          3115 => x"fc",
          3116 => x"b4",
          3117 => x"f8",
          3118 => x"f0",
          3119 => x"06",
          3120 => x"81",
          3121 => x"fe",
          3122 => x"3d",
          3123 => x"3d",
          3124 => x"7e",
          3125 => x"82",
          3126 => x"27",
          3127 => x"76",
          3128 => x"27",
          3129 => x"75",
          3130 => x"79",
          3131 => x"38",
          3132 => x"89",
          3133 => x"2e",
          3134 => x"80",
          3135 => x"2e",
          3136 => x"81",
          3137 => x"81",
          3138 => x"89",
          3139 => x"08",
          3140 => x"52",
          3141 => x"3f",
          3142 => x"08",
          3143 => x"f0",
          3144 => x"38",
          3145 => x"06",
          3146 => x"81",
          3147 => x"06",
          3148 => x"77",
          3149 => x"2e",
          3150 => x"84",
          3151 => x"06",
          3152 => x"06",
          3153 => x"53",
          3154 => x"81",
          3155 => x"34",
          3156 => x"a4",
          3157 => x"52",
          3158 => x"d9",
          3159 => x"f0",
          3160 => x"fe",
          3161 => x"94",
          3162 => x"ff",
          3163 => x"05",
          3164 => x"54",
          3165 => x"38",
          3166 => x"74",
          3167 => x"06",
          3168 => x"07",
          3169 => x"74",
          3170 => x"39",
          3171 => x"a4",
          3172 => x"52",
          3173 => x"9d",
          3174 => x"f0",
          3175 => x"fe",
          3176 => x"d8",
          3177 => x"ff",
          3178 => x"76",
          3179 => x"06",
          3180 => x"05",
          3181 => x"3f",
          3182 => x"87",
          3183 => x"08",
          3184 => x"51",
          3185 => x"81",
          3186 => x"59",
          3187 => x"08",
          3188 => x"f0",
          3189 => x"82",
          3190 => x"06",
          3191 => x"05",
          3192 => x"54",
          3193 => x"3f",
          3194 => x"08",
          3195 => x"74",
          3196 => x"51",
          3197 => x"81",
          3198 => x"34",
          3199 => x"f0",
          3200 => x"0d",
          3201 => x"0d",
          3202 => x"72",
          3203 => x"56",
          3204 => x"27",
          3205 => x"98",
          3206 => x"9d",
          3207 => x"2e",
          3208 => x"53",
          3209 => x"51",
          3210 => x"81",
          3211 => x"54",
          3212 => x"08",
          3213 => x"93",
          3214 => x"80",
          3215 => x"54",
          3216 => x"81",
          3217 => x"54",
          3218 => x"74",
          3219 => x"fb",
          3220 => x"fe",
          3221 => x"81",
          3222 => x"80",
          3223 => x"38",
          3224 => x"08",
          3225 => x"38",
          3226 => x"08",
          3227 => x"38",
          3228 => x"52",
          3229 => x"d6",
          3230 => x"f0",
          3231 => x"98",
          3232 => x"11",
          3233 => x"57",
          3234 => x"74",
          3235 => x"81",
          3236 => x"0c",
          3237 => x"81",
          3238 => x"84",
          3239 => x"55",
          3240 => x"ff",
          3241 => x"54",
          3242 => x"f0",
          3243 => x"0d",
          3244 => x"0d",
          3245 => x"08",
          3246 => x"79",
          3247 => x"17",
          3248 => x"80",
          3249 => x"98",
          3250 => x"26",
          3251 => x"58",
          3252 => x"52",
          3253 => x"fd",
          3254 => x"74",
          3255 => x"08",
          3256 => x"38",
          3257 => x"08",
          3258 => x"f0",
          3259 => x"82",
          3260 => x"17",
          3261 => x"f0",
          3262 => x"c7",
          3263 => x"90",
          3264 => x"56",
          3265 => x"2e",
          3266 => x"77",
          3267 => x"81",
          3268 => x"38",
          3269 => x"98",
          3270 => x"26",
          3271 => x"56",
          3272 => x"51",
          3273 => x"80",
          3274 => x"f0",
          3275 => x"09",
          3276 => x"38",
          3277 => x"08",
          3278 => x"f0",
          3279 => x"30",
          3280 => x"80",
          3281 => x"07",
          3282 => x"08",
          3283 => x"55",
          3284 => x"ef",
          3285 => x"f0",
          3286 => x"95",
          3287 => x"08",
          3288 => x"27",
          3289 => x"98",
          3290 => x"89",
          3291 => x"85",
          3292 => x"db",
          3293 => x"81",
          3294 => x"17",
          3295 => x"89",
          3296 => x"75",
          3297 => x"ac",
          3298 => x"7a",
          3299 => x"3f",
          3300 => x"08",
          3301 => x"38",
          3302 => x"fe",
          3303 => x"2e",
          3304 => x"86",
          3305 => x"f0",
          3306 => x"fe",
          3307 => x"70",
          3308 => x"07",
          3309 => x"7c",
          3310 => x"55",
          3311 => x"f8",
          3312 => x"2e",
          3313 => x"ff",
          3314 => x"55",
          3315 => x"ff",
          3316 => x"76",
          3317 => x"3f",
          3318 => x"08",
          3319 => x"08",
          3320 => x"fe",
          3321 => x"80",
          3322 => x"55",
          3323 => x"94",
          3324 => x"2e",
          3325 => x"53",
          3326 => x"51",
          3327 => x"81",
          3328 => x"55",
          3329 => x"75",
          3330 => x"98",
          3331 => x"05",
          3332 => x"56",
          3333 => x"26",
          3334 => x"15",
          3335 => x"84",
          3336 => x"07",
          3337 => x"18",
          3338 => x"ff",
          3339 => x"2e",
          3340 => x"39",
          3341 => x"39",
          3342 => x"08",
          3343 => x"81",
          3344 => x"74",
          3345 => x"0c",
          3346 => x"04",
          3347 => x"7a",
          3348 => x"f3",
          3349 => x"fe",
          3350 => x"81",
          3351 => x"f0",
          3352 => x"38",
          3353 => x"51",
          3354 => x"81",
          3355 => x"81",
          3356 => x"b0",
          3357 => x"84",
          3358 => x"52",
          3359 => x"52",
          3360 => x"3f",
          3361 => x"39",
          3362 => x"8a",
          3363 => x"75",
          3364 => x"38",
          3365 => x"19",
          3366 => x"81",
          3367 => x"ed",
          3368 => x"fe",
          3369 => x"2e",
          3370 => x"15",
          3371 => x"70",
          3372 => x"07",
          3373 => x"53",
          3374 => x"75",
          3375 => x"0c",
          3376 => x"04",
          3377 => x"7a",
          3378 => x"58",
          3379 => x"f0",
          3380 => x"80",
          3381 => x"9f",
          3382 => x"80",
          3383 => x"90",
          3384 => x"17",
          3385 => x"aa",
          3386 => x"53",
          3387 => x"88",
          3388 => x"08",
          3389 => x"38",
          3390 => x"53",
          3391 => x"17",
          3392 => x"72",
          3393 => x"fe",
          3394 => x"08",
          3395 => x"80",
          3396 => x"16",
          3397 => x"2b",
          3398 => x"75",
          3399 => x"73",
          3400 => x"f5",
          3401 => x"fe",
          3402 => x"81",
          3403 => x"ff",
          3404 => x"81",
          3405 => x"f0",
          3406 => x"38",
          3407 => x"81",
          3408 => x"26",
          3409 => x"58",
          3410 => x"73",
          3411 => x"39",
          3412 => x"51",
          3413 => x"81",
          3414 => x"98",
          3415 => x"94",
          3416 => x"17",
          3417 => x"58",
          3418 => x"9a",
          3419 => x"81",
          3420 => x"74",
          3421 => x"98",
          3422 => x"83",
          3423 => x"b4",
          3424 => x"0c",
          3425 => x"81",
          3426 => x"8a",
          3427 => x"f8",
          3428 => x"70",
          3429 => x"08",
          3430 => x"57",
          3431 => x"0a",
          3432 => x"38",
          3433 => x"15",
          3434 => x"08",
          3435 => x"72",
          3436 => x"cb",
          3437 => x"ff",
          3438 => x"81",
          3439 => x"13",
          3440 => x"94",
          3441 => x"74",
          3442 => x"85",
          3443 => x"22",
          3444 => x"73",
          3445 => x"38",
          3446 => x"8a",
          3447 => x"05",
          3448 => x"06",
          3449 => x"8a",
          3450 => x"73",
          3451 => x"3f",
          3452 => x"08",
          3453 => x"81",
          3454 => x"f0",
          3455 => x"ff",
          3456 => x"81",
          3457 => x"ff",
          3458 => x"38",
          3459 => x"81",
          3460 => x"26",
          3461 => x"7b",
          3462 => x"98",
          3463 => x"55",
          3464 => x"94",
          3465 => x"73",
          3466 => x"3f",
          3467 => x"08",
          3468 => x"81",
          3469 => x"80",
          3470 => x"38",
          3471 => x"fe",
          3472 => x"2e",
          3473 => x"55",
          3474 => x"08",
          3475 => x"38",
          3476 => x"08",
          3477 => x"fb",
          3478 => x"fe",
          3479 => x"38",
          3480 => x"0c",
          3481 => x"51",
          3482 => x"81",
          3483 => x"98",
          3484 => x"90",
          3485 => x"16",
          3486 => x"15",
          3487 => x"74",
          3488 => x"0c",
          3489 => x"04",
          3490 => x"7b",
          3491 => x"5b",
          3492 => x"52",
          3493 => x"ac",
          3494 => x"f0",
          3495 => x"fe",
          3496 => x"ec",
          3497 => x"f0",
          3498 => x"17",
          3499 => x"51",
          3500 => x"81",
          3501 => x"54",
          3502 => x"08",
          3503 => x"81",
          3504 => x"9c",
          3505 => x"33",
          3506 => x"72",
          3507 => x"09",
          3508 => x"38",
          3509 => x"fe",
          3510 => x"72",
          3511 => x"55",
          3512 => x"53",
          3513 => x"8e",
          3514 => x"56",
          3515 => x"09",
          3516 => x"38",
          3517 => x"fe",
          3518 => x"81",
          3519 => x"fd",
          3520 => x"fe",
          3521 => x"81",
          3522 => x"80",
          3523 => x"38",
          3524 => x"09",
          3525 => x"38",
          3526 => x"81",
          3527 => x"8b",
          3528 => x"fd",
          3529 => x"9a",
          3530 => x"eb",
          3531 => x"fe",
          3532 => x"ff",
          3533 => x"70",
          3534 => x"53",
          3535 => x"09",
          3536 => x"38",
          3537 => x"eb",
          3538 => x"fe",
          3539 => x"2b",
          3540 => x"72",
          3541 => x"0c",
          3542 => x"04",
          3543 => x"77",
          3544 => x"ff",
          3545 => x"9a",
          3546 => x"55",
          3547 => x"76",
          3548 => x"53",
          3549 => x"09",
          3550 => x"38",
          3551 => x"52",
          3552 => x"eb",
          3553 => x"3d",
          3554 => x"3d",
          3555 => x"5b",
          3556 => x"08",
          3557 => x"15",
          3558 => x"81",
          3559 => x"15",
          3560 => x"51",
          3561 => x"81",
          3562 => x"58",
          3563 => x"08",
          3564 => x"9c",
          3565 => x"33",
          3566 => x"86",
          3567 => x"80",
          3568 => x"13",
          3569 => x"06",
          3570 => x"06",
          3571 => x"72",
          3572 => x"81",
          3573 => x"53",
          3574 => x"2e",
          3575 => x"53",
          3576 => x"a9",
          3577 => x"74",
          3578 => x"72",
          3579 => x"38",
          3580 => x"99",
          3581 => x"f0",
          3582 => x"06",
          3583 => x"88",
          3584 => x"06",
          3585 => x"54",
          3586 => x"a0",
          3587 => x"74",
          3588 => x"3f",
          3589 => x"08",
          3590 => x"f0",
          3591 => x"98",
          3592 => x"fa",
          3593 => x"80",
          3594 => x"0c",
          3595 => x"f0",
          3596 => x"0d",
          3597 => x"0d",
          3598 => x"57",
          3599 => x"73",
          3600 => x"3f",
          3601 => x"08",
          3602 => x"f0",
          3603 => x"98",
          3604 => x"75",
          3605 => x"3f",
          3606 => x"08",
          3607 => x"f0",
          3608 => x"a0",
          3609 => x"f0",
          3610 => x"14",
          3611 => x"db",
          3612 => x"a0",
          3613 => x"14",
          3614 => x"ac",
          3615 => x"83",
          3616 => x"81",
          3617 => x"87",
          3618 => x"fd",
          3619 => x"70",
          3620 => x"08",
          3621 => x"55",
          3622 => x"3f",
          3623 => x"08",
          3624 => x"13",
          3625 => x"73",
          3626 => x"83",
          3627 => x"3d",
          3628 => x"3d",
          3629 => x"57",
          3630 => x"89",
          3631 => x"17",
          3632 => x"81",
          3633 => x"70",
          3634 => x"55",
          3635 => x"08",
          3636 => x"81",
          3637 => x"52",
          3638 => x"a8",
          3639 => x"2e",
          3640 => x"84",
          3641 => x"52",
          3642 => x"09",
          3643 => x"38",
          3644 => x"81",
          3645 => x"81",
          3646 => x"73",
          3647 => x"55",
          3648 => x"55",
          3649 => x"c5",
          3650 => x"88",
          3651 => x"0b",
          3652 => x"9c",
          3653 => x"8b",
          3654 => x"17",
          3655 => x"08",
          3656 => x"52",
          3657 => x"81",
          3658 => x"76",
          3659 => x"51",
          3660 => x"81",
          3661 => x"86",
          3662 => x"12",
          3663 => x"3f",
          3664 => x"08",
          3665 => x"88",
          3666 => x"f3",
          3667 => x"70",
          3668 => x"80",
          3669 => x"51",
          3670 => x"af",
          3671 => x"81",
          3672 => x"dc",
          3673 => x"74",
          3674 => x"38",
          3675 => x"88",
          3676 => x"39",
          3677 => x"80",
          3678 => x"56",
          3679 => x"af",
          3680 => x"06",
          3681 => x"56",
          3682 => x"32",
          3683 => x"80",
          3684 => x"51",
          3685 => x"dc",
          3686 => x"1c",
          3687 => x"33",
          3688 => x"9f",
          3689 => x"ff",
          3690 => x"1c",
          3691 => x"7a",
          3692 => x"3f",
          3693 => x"08",
          3694 => x"39",
          3695 => x"a0",
          3696 => x"5e",
          3697 => x"52",
          3698 => x"ff",
          3699 => x"59",
          3700 => x"33",
          3701 => x"ae",
          3702 => x"06",
          3703 => x"78",
          3704 => x"81",
          3705 => x"32",
          3706 => x"9f",
          3707 => x"26",
          3708 => x"53",
          3709 => x"73",
          3710 => x"17",
          3711 => x"34",
          3712 => x"db",
          3713 => x"32",
          3714 => x"9f",
          3715 => x"54",
          3716 => x"2e",
          3717 => x"80",
          3718 => x"75",
          3719 => x"bd",
          3720 => x"7e",
          3721 => x"a0",
          3722 => x"bd",
          3723 => x"82",
          3724 => x"18",
          3725 => x"1a",
          3726 => x"a0",
          3727 => x"fc",
          3728 => x"32",
          3729 => x"80",
          3730 => x"30",
          3731 => x"71",
          3732 => x"51",
          3733 => x"55",
          3734 => x"ac",
          3735 => x"81",
          3736 => x"78",
          3737 => x"51",
          3738 => x"af",
          3739 => x"06",
          3740 => x"55",
          3741 => x"32",
          3742 => x"80",
          3743 => x"51",
          3744 => x"db",
          3745 => x"39",
          3746 => x"09",
          3747 => x"38",
          3748 => x"7c",
          3749 => x"54",
          3750 => x"a2",
          3751 => x"32",
          3752 => x"ae",
          3753 => x"72",
          3754 => x"9f",
          3755 => x"51",
          3756 => x"74",
          3757 => x"88",
          3758 => x"fe",
          3759 => x"98",
          3760 => x"80",
          3761 => x"75",
          3762 => x"81",
          3763 => x"33",
          3764 => x"51",
          3765 => x"81",
          3766 => x"80",
          3767 => x"78",
          3768 => x"81",
          3769 => x"5a",
          3770 => x"d2",
          3771 => x"f0",
          3772 => x"80",
          3773 => x"1c",
          3774 => x"27",
          3775 => x"79",
          3776 => x"74",
          3777 => x"7a",
          3778 => x"74",
          3779 => x"39",
          3780 => x"ea",
          3781 => x"fe",
          3782 => x"f0",
          3783 => x"ff",
          3784 => x"73",
          3785 => x"38",
          3786 => x"81",
          3787 => x"54",
          3788 => x"75",
          3789 => x"17",
          3790 => x"39",
          3791 => x"0c",
          3792 => x"99",
          3793 => x"54",
          3794 => x"2e",
          3795 => x"84",
          3796 => x"34",
          3797 => x"76",
          3798 => x"8b",
          3799 => x"81",
          3800 => x"56",
          3801 => x"80",
          3802 => x"1b",
          3803 => x"08",
          3804 => x"51",
          3805 => x"81",
          3806 => x"56",
          3807 => x"08",
          3808 => x"98",
          3809 => x"76",
          3810 => x"3f",
          3811 => x"08",
          3812 => x"f0",
          3813 => x"38",
          3814 => x"70",
          3815 => x"73",
          3816 => x"be",
          3817 => x"33",
          3818 => x"73",
          3819 => x"8b",
          3820 => x"83",
          3821 => x"06",
          3822 => x"73",
          3823 => x"53",
          3824 => x"51",
          3825 => x"81",
          3826 => x"80",
          3827 => x"75",
          3828 => x"f3",
          3829 => x"9f",
          3830 => x"1c",
          3831 => x"74",
          3832 => x"38",
          3833 => x"09",
          3834 => x"e7",
          3835 => x"2a",
          3836 => x"77",
          3837 => x"51",
          3838 => x"2e",
          3839 => x"81",
          3840 => x"80",
          3841 => x"38",
          3842 => x"ab",
          3843 => x"55",
          3844 => x"75",
          3845 => x"73",
          3846 => x"55",
          3847 => x"82",
          3848 => x"06",
          3849 => x"ab",
          3850 => x"33",
          3851 => x"70",
          3852 => x"55",
          3853 => x"2e",
          3854 => x"1b",
          3855 => x"06",
          3856 => x"52",
          3857 => x"db",
          3858 => x"f0",
          3859 => x"0c",
          3860 => x"74",
          3861 => x"0c",
          3862 => x"04",
          3863 => x"7c",
          3864 => x"08",
          3865 => x"55",
          3866 => x"59",
          3867 => x"81",
          3868 => x"70",
          3869 => x"33",
          3870 => x"52",
          3871 => x"2e",
          3872 => x"ee",
          3873 => x"2e",
          3874 => x"81",
          3875 => x"33",
          3876 => x"81",
          3877 => x"52",
          3878 => x"26",
          3879 => x"14",
          3880 => x"06",
          3881 => x"52",
          3882 => x"80",
          3883 => x"0b",
          3884 => x"59",
          3885 => x"7a",
          3886 => x"70",
          3887 => x"33",
          3888 => x"05",
          3889 => x"9f",
          3890 => x"53",
          3891 => x"89",
          3892 => x"70",
          3893 => x"54",
          3894 => x"12",
          3895 => x"26",
          3896 => x"12",
          3897 => x"06",
          3898 => x"30",
          3899 => x"51",
          3900 => x"2e",
          3901 => x"85",
          3902 => x"be",
          3903 => x"74",
          3904 => x"30",
          3905 => x"9f",
          3906 => x"2a",
          3907 => x"54",
          3908 => x"2e",
          3909 => x"15",
          3910 => x"55",
          3911 => x"ff",
          3912 => x"39",
          3913 => x"86",
          3914 => x"7c",
          3915 => x"51",
          3916 => x"ff",
          3917 => x"70",
          3918 => x"0c",
          3919 => x"04",
          3920 => x"78",
          3921 => x"83",
          3922 => x"0b",
          3923 => x"79",
          3924 => x"e2",
          3925 => x"55",
          3926 => x"08",
          3927 => x"84",
          3928 => x"df",
          3929 => x"fe",
          3930 => x"ff",
          3931 => x"83",
          3932 => x"d4",
          3933 => x"81",
          3934 => x"38",
          3935 => x"17",
          3936 => x"74",
          3937 => x"09",
          3938 => x"38",
          3939 => x"81",
          3940 => x"30",
          3941 => x"79",
          3942 => x"54",
          3943 => x"74",
          3944 => x"09",
          3945 => x"38",
          3946 => x"eb",
          3947 => x"ea",
          3948 => x"b1",
          3949 => x"f0",
          3950 => x"fe",
          3951 => x"2e",
          3952 => x"53",
          3953 => x"52",
          3954 => x"51",
          3955 => x"81",
          3956 => x"55",
          3957 => x"08",
          3958 => x"38",
          3959 => x"81",
          3960 => x"88",
          3961 => x"f2",
          3962 => x"02",
          3963 => x"cb",
          3964 => x"55",
          3965 => x"60",
          3966 => x"3f",
          3967 => x"08",
          3968 => x"80",
          3969 => x"f0",
          3970 => x"fc",
          3971 => x"f0",
          3972 => x"81",
          3973 => x"70",
          3974 => x"8c",
          3975 => x"2e",
          3976 => x"73",
          3977 => x"81",
          3978 => x"33",
          3979 => x"80",
          3980 => x"81",
          3981 => x"d7",
          3982 => x"fe",
          3983 => x"ff",
          3984 => x"06",
          3985 => x"98",
          3986 => x"2e",
          3987 => x"74",
          3988 => x"81",
          3989 => x"8a",
          3990 => x"ac",
          3991 => x"39",
          3992 => x"77",
          3993 => x"81",
          3994 => x"33",
          3995 => x"3f",
          3996 => x"08",
          3997 => x"70",
          3998 => x"55",
          3999 => x"86",
          4000 => x"80",
          4001 => x"74",
          4002 => x"81",
          4003 => x"8a",
          4004 => x"f4",
          4005 => x"53",
          4006 => x"fd",
          4007 => x"fe",
          4008 => x"ff",
          4009 => x"82",
          4010 => x"06",
          4011 => x"8c",
          4012 => x"58",
          4013 => x"f6",
          4014 => x"58",
          4015 => x"2e",
          4016 => x"fa",
          4017 => x"e8",
          4018 => x"f0",
          4019 => x"78",
          4020 => x"5a",
          4021 => x"90",
          4022 => x"75",
          4023 => x"38",
          4024 => x"3d",
          4025 => x"70",
          4026 => x"08",
          4027 => x"7a",
          4028 => x"38",
          4029 => x"51",
          4030 => x"81",
          4031 => x"81",
          4032 => x"81",
          4033 => x"38",
          4034 => x"83",
          4035 => x"38",
          4036 => x"84",
          4037 => x"38",
          4038 => x"81",
          4039 => x"38",
          4040 => x"db",
          4041 => x"fe",
          4042 => x"ff",
          4043 => x"72",
          4044 => x"09",
          4045 => x"d0",
          4046 => x"14",
          4047 => x"3f",
          4048 => x"08",
          4049 => x"06",
          4050 => x"38",
          4051 => x"51",
          4052 => x"81",
          4053 => x"58",
          4054 => x"0c",
          4055 => x"33",
          4056 => x"80",
          4057 => x"ff",
          4058 => x"ff",
          4059 => x"55",
          4060 => x"81",
          4061 => x"38",
          4062 => x"06",
          4063 => x"80",
          4064 => x"52",
          4065 => x"8a",
          4066 => x"80",
          4067 => x"ff",
          4068 => x"53",
          4069 => x"86",
          4070 => x"83",
          4071 => x"c5",
          4072 => x"f5",
          4073 => x"f0",
          4074 => x"fe",
          4075 => x"15",
          4076 => x"06",
          4077 => x"76",
          4078 => x"80",
          4079 => x"da",
          4080 => x"fe",
          4081 => x"ff",
          4082 => x"74",
          4083 => x"d4",
          4084 => x"dc",
          4085 => x"f0",
          4086 => x"c2",
          4087 => x"b9",
          4088 => x"f0",
          4089 => x"ff",
          4090 => x"56",
          4091 => x"83",
          4092 => x"14",
          4093 => x"71",
          4094 => x"5a",
          4095 => x"26",
          4096 => x"8a",
          4097 => x"74",
          4098 => x"ff",
          4099 => x"81",
          4100 => x"55",
          4101 => x"08",
          4102 => x"ec",
          4103 => x"f0",
          4104 => x"ff",
          4105 => x"83",
          4106 => x"74",
          4107 => x"26",
          4108 => x"57",
          4109 => x"26",
          4110 => x"57",
          4111 => x"56",
          4112 => x"82",
          4113 => x"15",
          4114 => x"0c",
          4115 => x"0c",
          4116 => x"a4",
          4117 => x"1d",
          4118 => x"54",
          4119 => x"2e",
          4120 => x"af",
          4121 => x"14",
          4122 => x"3f",
          4123 => x"08",
          4124 => x"06",
          4125 => x"72",
          4126 => x"79",
          4127 => x"80",
          4128 => x"d9",
          4129 => x"fe",
          4130 => x"15",
          4131 => x"2b",
          4132 => x"8d",
          4133 => x"2e",
          4134 => x"77",
          4135 => x"0c",
          4136 => x"76",
          4137 => x"38",
          4138 => x"70",
          4139 => x"81",
          4140 => x"53",
          4141 => x"89",
          4142 => x"56",
          4143 => x"08",
          4144 => x"38",
          4145 => x"15",
          4146 => x"8c",
          4147 => x"80",
          4148 => x"34",
          4149 => x"09",
          4150 => x"92",
          4151 => x"14",
          4152 => x"3f",
          4153 => x"08",
          4154 => x"06",
          4155 => x"2e",
          4156 => x"80",
          4157 => x"1b",
          4158 => x"db",
          4159 => x"fe",
          4160 => x"ea",
          4161 => x"f0",
          4162 => x"34",
          4163 => x"51",
          4164 => x"81",
          4165 => x"83",
          4166 => x"53",
          4167 => x"d5",
          4168 => x"06",
          4169 => x"b4",
          4170 => x"84",
          4171 => x"f0",
          4172 => x"85",
          4173 => x"09",
          4174 => x"38",
          4175 => x"51",
          4176 => x"81",
          4177 => x"86",
          4178 => x"f2",
          4179 => x"06",
          4180 => x"9c",
          4181 => x"d8",
          4182 => x"f0",
          4183 => x"0c",
          4184 => x"51",
          4185 => x"81",
          4186 => x"8c",
          4187 => x"74",
          4188 => x"b0",
          4189 => x"53",
          4190 => x"b0",
          4191 => x"15",
          4192 => x"94",
          4193 => x"56",
          4194 => x"f0",
          4195 => x"0d",
          4196 => x"0d",
          4197 => x"55",
          4198 => x"b9",
          4199 => x"53",
          4200 => x"b1",
          4201 => x"52",
          4202 => x"a9",
          4203 => x"22",
          4204 => x"57",
          4205 => x"2e",
          4206 => x"99",
          4207 => x"33",
          4208 => x"3f",
          4209 => x"08",
          4210 => x"71",
          4211 => x"74",
          4212 => x"83",
          4213 => x"78",
          4214 => x"52",
          4215 => x"f0",
          4216 => x"0d",
          4217 => x"0d",
          4218 => x"33",
          4219 => x"3d",
          4220 => x"56",
          4221 => x"8b",
          4222 => x"81",
          4223 => x"24",
          4224 => x"fe",
          4225 => x"29",
          4226 => x"05",
          4227 => x"55",
          4228 => x"84",
          4229 => x"34",
          4230 => x"80",
          4231 => x"80",
          4232 => x"75",
          4233 => x"75",
          4234 => x"38",
          4235 => x"3d",
          4236 => x"05",
          4237 => x"3f",
          4238 => x"08",
          4239 => x"fe",
          4240 => x"3d",
          4241 => x"3d",
          4242 => x"84",
          4243 => x"05",
          4244 => x"89",
          4245 => x"2e",
          4246 => x"77",
          4247 => x"54",
          4248 => x"05",
          4249 => x"84",
          4250 => x"f6",
          4251 => x"fe",
          4252 => x"81",
          4253 => x"84",
          4254 => x"5c",
          4255 => x"3d",
          4256 => x"ed",
          4257 => x"fe",
          4258 => x"81",
          4259 => x"92",
          4260 => x"d7",
          4261 => x"98",
          4262 => x"73",
          4263 => x"38",
          4264 => x"9c",
          4265 => x"80",
          4266 => x"38",
          4267 => x"95",
          4268 => x"2e",
          4269 => x"aa",
          4270 => x"ea",
          4271 => x"fe",
          4272 => x"9e",
          4273 => x"05",
          4274 => x"54",
          4275 => x"38",
          4276 => x"70",
          4277 => x"54",
          4278 => x"8e",
          4279 => x"83",
          4280 => x"88",
          4281 => x"83",
          4282 => x"83",
          4283 => x"06",
          4284 => x"80",
          4285 => x"38",
          4286 => x"51",
          4287 => x"81",
          4288 => x"56",
          4289 => x"0a",
          4290 => x"05",
          4291 => x"3f",
          4292 => x"0b",
          4293 => x"80",
          4294 => x"7a",
          4295 => x"3f",
          4296 => x"9c",
          4297 => x"d1",
          4298 => x"81",
          4299 => x"34",
          4300 => x"80",
          4301 => x"b0",
          4302 => x"54",
          4303 => x"52",
          4304 => x"05",
          4305 => x"3f",
          4306 => x"08",
          4307 => x"f0",
          4308 => x"38",
          4309 => x"82",
          4310 => x"b2",
          4311 => x"84",
          4312 => x"06",
          4313 => x"73",
          4314 => x"38",
          4315 => x"ad",
          4316 => x"2a",
          4317 => x"51",
          4318 => x"2e",
          4319 => x"81",
          4320 => x"80",
          4321 => x"87",
          4322 => x"39",
          4323 => x"51",
          4324 => x"81",
          4325 => x"7b",
          4326 => x"12",
          4327 => x"81",
          4328 => x"81",
          4329 => x"83",
          4330 => x"06",
          4331 => x"80",
          4332 => x"77",
          4333 => x"58",
          4334 => x"08",
          4335 => x"63",
          4336 => x"63",
          4337 => x"57",
          4338 => x"81",
          4339 => x"81",
          4340 => x"88",
          4341 => x"9c",
          4342 => x"d2",
          4343 => x"fe",
          4344 => x"fe",
          4345 => x"1b",
          4346 => x"0c",
          4347 => x"22",
          4348 => x"77",
          4349 => x"80",
          4350 => x"34",
          4351 => x"1a",
          4352 => x"94",
          4353 => x"85",
          4354 => x"06",
          4355 => x"80",
          4356 => x"38",
          4357 => x"08",
          4358 => x"84",
          4359 => x"f0",
          4360 => x"0c",
          4361 => x"70",
          4362 => x"52",
          4363 => x"39",
          4364 => x"51",
          4365 => x"81",
          4366 => x"57",
          4367 => x"08",
          4368 => x"38",
          4369 => x"fe",
          4370 => x"2e",
          4371 => x"83",
          4372 => x"75",
          4373 => x"74",
          4374 => x"07",
          4375 => x"54",
          4376 => x"8a",
          4377 => x"75",
          4378 => x"73",
          4379 => x"98",
          4380 => x"a9",
          4381 => x"ff",
          4382 => x"80",
          4383 => x"76",
          4384 => x"d6",
          4385 => x"fe",
          4386 => x"38",
          4387 => x"39",
          4388 => x"81",
          4389 => x"05",
          4390 => x"84",
          4391 => x"0c",
          4392 => x"81",
          4393 => x"97",
          4394 => x"f2",
          4395 => x"63",
          4396 => x"40",
          4397 => x"7e",
          4398 => x"fc",
          4399 => x"51",
          4400 => x"81",
          4401 => x"55",
          4402 => x"08",
          4403 => x"19",
          4404 => x"80",
          4405 => x"74",
          4406 => x"39",
          4407 => x"81",
          4408 => x"56",
          4409 => x"82",
          4410 => x"39",
          4411 => x"1a",
          4412 => x"82",
          4413 => x"0b",
          4414 => x"81",
          4415 => x"39",
          4416 => x"94",
          4417 => x"55",
          4418 => x"83",
          4419 => x"7b",
          4420 => x"89",
          4421 => x"08",
          4422 => x"06",
          4423 => x"81",
          4424 => x"8a",
          4425 => x"05",
          4426 => x"06",
          4427 => x"a8",
          4428 => x"38",
          4429 => x"55",
          4430 => x"19",
          4431 => x"51",
          4432 => x"81",
          4433 => x"55",
          4434 => x"ff",
          4435 => x"ff",
          4436 => x"38",
          4437 => x"0c",
          4438 => x"52",
          4439 => x"cb",
          4440 => x"f0",
          4441 => x"ff",
          4442 => x"fe",
          4443 => x"7c",
          4444 => x"57",
          4445 => x"80",
          4446 => x"1a",
          4447 => x"22",
          4448 => x"75",
          4449 => x"38",
          4450 => x"58",
          4451 => x"53",
          4452 => x"1b",
          4453 => x"88",
          4454 => x"f0",
          4455 => x"38",
          4456 => x"33",
          4457 => x"80",
          4458 => x"b0",
          4459 => x"31",
          4460 => x"27",
          4461 => x"80",
          4462 => x"52",
          4463 => x"77",
          4464 => x"7d",
          4465 => x"e0",
          4466 => x"2b",
          4467 => x"76",
          4468 => x"94",
          4469 => x"ff",
          4470 => x"71",
          4471 => x"7b",
          4472 => x"38",
          4473 => x"19",
          4474 => x"51",
          4475 => x"81",
          4476 => x"fe",
          4477 => x"53",
          4478 => x"83",
          4479 => x"b4",
          4480 => x"51",
          4481 => x"7b",
          4482 => x"08",
          4483 => x"76",
          4484 => x"08",
          4485 => x"0c",
          4486 => x"f3",
          4487 => x"75",
          4488 => x"0c",
          4489 => x"04",
          4490 => x"60",
          4491 => x"40",
          4492 => x"80",
          4493 => x"3d",
          4494 => x"77",
          4495 => x"3f",
          4496 => x"08",
          4497 => x"f0",
          4498 => x"91",
          4499 => x"74",
          4500 => x"38",
          4501 => x"b8",
          4502 => x"33",
          4503 => x"70",
          4504 => x"56",
          4505 => x"74",
          4506 => x"a4",
          4507 => x"82",
          4508 => x"34",
          4509 => x"98",
          4510 => x"91",
          4511 => x"56",
          4512 => x"94",
          4513 => x"11",
          4514 => x"76",
          4515 => x"75",
          4516 => x"80",
          4517 => x"38",
          4518 => x"70",
          4519 => x"56",
          4520 => x"fd",
          4521 => x"11",
          4522 => x"77",
          4523 => x"5c",
          4524 => x"38",
          4525 => x"88",
          4526 => x"74",
          4527 => x"52",
          4528 => x"18",
          4529 => x"51",
          4530 => x"81",
          4531 => x"55",
          4532 => x"08",
          4533 => x"ab",
          4534 => x"2e",
          4535 => x"74",
          4536 => x"95",
          4537 => x"19",
          4538 => x"08",
          4539 => x"88",
          4540 => x"55",
          4541 => x"9c",
          4542 => x"09",
          4543 => x"38",
          4544 => x"c1",
          4545 => x"f0",
          4546 => x"38",
          4547 => x"52",
          4548 => x"97",
          4549 => x"f0",
          4550 => x"fe",
          4551 => x"fe",
          4552 => x"7c",
          4553 => x"57",
          4554 => x"80",
          4555 => x"1b",
          4556 => x"22",
          4557 => x"75",
          4558 => x"38",
          4559 => x"59",
          4560 => x"53",
          4561 => x"1a",
          4562 => x"be",
          4563 => x"f0",
          4564 => x"38",
          4565 => x"08",
          4566 => x"56",
          4567 => x"9b",
          4568 => x"53",
          4569 => x"77",
          4570 => x"7d",
          4571 => x"16",
          4572 => x"3f",
          4573 => x"0b",
          4574 => x"78",
          4575 => x"80",
          4576 => x"18",
          4577 => x"08",
          4578 => x"7e",
          4579 => x"3f",
          4580 => x"08",
          4581 => x"7e",
          4582 => x"0c",
          4583 => x"19",
          4584 => x"08",
          4585 => x"84",
          4586 => x"57",
          4587 => x"27",
          4588 => x"56",
          4589 => x"52",
          4590 => x"f9",
          4591 => x"f0",
          4592 => x"38",
          4593 => x"52",
          4594 => x"83",
          4595 => x"b4",
          4596 => x"d4",
          4597 => x"81",
          4598 => x"34",
          4599 => x"7e",
          4600 => x"0c",
          4601 => x"1a",
          4602 => x"94",
          4603 => x"1b",
          4604 => x"5e",
          4605 => x"27",
          4606 => x"55",
          4607 => x"0c",
          4608 => x"90",
          4609 => x"c0",
          4610 => x"90",
          4611 => x"56",
          4612 => x"f0",
          4613 => x"0d",
          4614 => x"0d",
          4615 => x"fc",
          4616 => x"52",
          4617 => x"3f",
          4618 => x"08",
          4619 => x"f0",
          4620 => x"38",
          4621 => x"70",
          4622 => x"81",
          4623 => x"55",
          4624 => x"80",
          4625 => x"16",
          4626 => x"51",
          4627 => x"81",
          4628 => x"57",
          4629 => x"08",
          4630 => x"a4",
          4631 => x"11",
          4632 => x"55",
          4633 => x"16",
          4634 => x"08",
          4635 => x"75",
          4636 => x"e8",
          4637 => x"08",
          4638 => x"51",
          4639 => x"82",
          4640 => x"52",
          4641 => x"c9",
          4642 => x"52",
          4643 => x"c9",
          4644 => x"54",
          4645 => x"15",
          4646 => x"cc",
          4647 => x"fe",
          4648 => x"17",
          4649 => x"06",
          4650 => x"90",
          4651 => x"81",
          4652 => x"8a",
          4653 => x"fc",
          4654 => x"70",
          4655 => x"d9",
          4656 => x"f0",
          4657 => x"fe",
          4658 => x"38",
          4659 => x"05",
          4660 => x"f1",
          4661 => x"fe",
          4662 => x"81",
          4663 => x"87",
          4664 => x"f0",
          4665 => x"72",
          4666 => x"0c",
          4667 => x"04",
          4668 => x"84",
          4669 => x"e4",
          4670 => x"80",
          4671 => x"f0",
          4672 => x"38",
          4673 => x"08",
          4674 => x"34",
          4675 => x"81",
          4676 => x"83",
          4677 => x"ef",
          4678 => x"53",
          4679 => x"05",
          4680 => x"51",
          4681 => x"81",
          4682 => x"55",
          4683 => x"08",
          4684 => x"76",
          4685 => x"93",
          4686 => x"51",
          4687 => x"81",
          4688 => x"55",
          4689 => x"08",
          4690 => x"80",
          4691 => x"70",
          4692 => x"56",
          4693 => x"89",
          4694 => x"94",
          4695 => x"b2",
          4696 => x"05",
          4697 => x"2a",
          4698 => x"51",
          4699 => x"80",
          4700 => x"76",
          4701 => x"52",
          4702 => x"3f",
          4703 => x"08",
          4704 => x"8e",
          4705 => x"f0",
          4706 => x"09",
          4707 => x"38",
          4708 => x"81",
          4709 => x"93",
          4710 => x"e4",
          4711 => x"6f",
          4712 => x"7a",
          4713 => x"9e",
          4714 => x"05",
          4715 => x"51",
          4716 => x"81",
          4717 => x"57",
          4718 => x"08",
          4719 => x"7b",
          4720 => x"94",
          4721 => x"55",
          4722 => x"73",
          4723 => x"ed",
          4724 => x"93",
          4725 => x"55",
          4726 => x"81",
          4727 => x"57",
          4728 => x"08",
          4729 => x"68",
          4730 => x"c9",
          4731 => x"fe",
          4732 => x"81",
          4733 => x"82",
          4734 => x"52",
          4735 => x"a3",
          4736 => x"f0",
          4737 => x"52",
          4738 => x"b8",
          4739 => x"f0",
          4740 => x"fe",
          4741 => x"a2",
          4742 => x"74",
          4743 => x"3f",
          4744 => x"08",
          4745 => x"f0",
          4746 => x"69",
          4747 => x"d9",
          4748 => x"81",
          4749 => x"2e",
          4750 => x"52",
          4751 => x"cf",
          4752 => x"f0",
          4753 => x"fe",
          4754 => x"2e",
          4755 => x"84",
          4756 => x"06",
          4757 => x"57",
          4758 => x"76",
          4759 => x"9e",
          4760 => x"05",
          4761 => x"dc",
          4762 => x"90",
          4763 => x"81",
          4764 => x"56",
          4765 => x"80",
          4766 => x"02",
          4767 => x"81",
          4768 => x"70",
          4769 => x"56",
          4770 => x"81",
          4771 => x"78",
          4772 => x"38",
          4773 => x"99",
          4774 => x"81",
          4775 => x"18",
          4776 => x"18",
          4777 => x"58",
          4778 => x"33",
          4779 => x"ee",
          4780 => x"6f",
          4781 => x"af",
          4782 => x"8d",
          4783 => x"2e",
          4784 => x"8a",
          4785 => x"6f",
          4786 => x"af",
          4787 => x"0b",
          4788 => x"33",
          4789 => x"81",
          4790 => x"70",
          4791 => x"52",
          4792 => x"56",
          4793 => x"8d",
          4794 => x"70",
          4795 => x"51",
          4796 => x"f5",
          4797 => x"54",
          4798 => x"a7",
          4799 => x"74",
          4800 => x"38",
          4801 => x"73",
          4802 => x"81",
          4803 => x"81",
          4804 => x"39",
          4805 => x"81",
          4806 => x"74",
          4807 => x"81",
          4808 => x"91",
          4809 => x"6e",
          4810 => x"59",
          4811 => x"7a",
          4812 => x"5c",
          4813 => x"26",
          4814 => x"7a",
          4815 => x"fe",
          4816 => x"3d",
          4817 => x"3d",
          4818 => x"8d",
          4819 => x"54",
          4820 => x"55",
          4821 => x"81",
          4822 => x"53",
          4823 => x"08",
          4824 => x"91",
          4825 => x"72",
          4826 => x"8c",
          4827 => x"73",
          4828 => x"38",
          4829 => x"70",
          4830 => x"81",
          4831 => x"57",
          4832 => x"73",
          4833 => x"08",
          4834 => x"94",
          4835 => x"75",
          4836 => x"97",
          4837 => x"11",
          4838 => x"2b",
          4839 => x"73",
          4840 => x"38",
          4841 => x"16",
          4842 => x"82",
          4843 => x"f0",
          4844 => x"78",
          4845 => x"55",
          4846 => x"f2",
          4847 => x"f0",
          4848 => x"96",
          4849 => x"70",
          4850 => x"94",
          4851 => x"71",
          4852 => x"08",
          4853 => x"53",
          4854 => x"15",
          4855 => x"a6",
          4856 => x"74",
          4857 => x"3f",
          4858 => x"08",
          4859 => x"f0",
          4860 => x"81",
          4861 => x"fe",
          4862 => x"2e",
          4863 => x"81",
          4864 => x"88",
          4865 => x"98",
          4866 => x"80",
          4867 => x"38",
          4868 => x"80",
          4869 => x"77",
          4870 => x"08",
          4871 => x"0c",
          4872 => x"70",
          4873 => x"81",
          4874 => x"5a",
          4875 => x"2e",
          4876 => x"52",
          4877 => x"f9",
          4878 => x"f0",
          4879 => x"fe",
          4880 => x"38",
          4881 => x"08",
          4882 => x"73",
          4883 => x"c7",
          4884 => x"fe",
          4885 => x"73",
          4886 => x"38",
          4887 => x"af",
          4888 => x"73",
          4889 => x"27",
          4890 => x"98",
          4891 => x"a0",
          4892 => x"08",
          4893 => x"0c",
          4894 => x"06",
          4895 => x"2e",
          4896 => x"52",
          4897 => x"a3",
          4898 => x"f0",
          4899 => x"82",
          4900 => x"34",
          4901 => x"c4",
          4902 => x"91",
          4903 => x"53",
          4904 => x"89",
          4905 => x"f0",
          4906 => x"94",
          4907 => x"8c",
          4908 => x"27",
          4909 => x"8c",
          4910 => x"15",
          4911 => x"07",
          4912 => x"16",
          4913 => x"ff",
          4914 => x"80",
          4915 => x"77",
          4916 => x"2e",
          4917 => x"9c",
          4918 => x"53",
          4919 => x"f0",
          4920 => x"0d",
          4921 => x"0d",
          4922 => x"54",
          4923 => x"81",
          4924 => x"53",
          4925 => x"05",
          4926 => x"84",
          4927 => x"e7",
          4928 => x"f0",
          4929 => x"fe",
          4930 => x"ea",
          4931 => x"0c",
          4932 => x"51",
          4933 => x"81",
          4934 => x"55",
          4935 => x"08",
          4936 => x"ab",
          4937 => x"98",
          4938 => x"80",
          4939 => x"38",
          4940 => x"70",
          4941 => x"81",
          4942 => x"57",
          4943 => x"ad",
          4944 => x"08",
          4945 => x"d3",
          4946 => x"fe",
          4947 => x"17",
          4948 => x"86",
          4949 => x"17",
          4950 => x"75",
          4951 => x"3f",
          4952 => x"08",
          4953 => x"2e",
          4954 => x"85",
          4955 => x"86",
          4956 => x"2e",
          4957 => x"76",
          4958 => x"73",
          4959 => x"0c",
          4960 => x"04",
          4961 => x"76",
          4962 => x"05",
          4963 => x"53",
          4964 => x"81",
          4965 => x"87",
          4966 => x"f0",
          4967 => x"86",
          4968 => x"fb",
          4969 => x"79",
          4970 => x"05",
          4971 => x"56",
          4972 => x"3f",
          4973 => x"08",
          4974 => x"f0",
          4975 => x"38",
          4976 => x"81",
          4977 => x"52",
          4978 => x"f8",
          4979 => x"f0",
          4980 => x"ca",
          4981 => x"f0",
          4982 => x"51",
          4983 => x"81",
          4984 => x"53",
          4985 => x"08",
          4986 => x"81",
          4987 => x"80",
          4988 => x"81",
          4989 => x"a6",
          4990 => x"73",
          4991 => x"3f",
          4992 => x"51",
          4993 => x"81",
          4994 => x"84",
          4995 => x"70",
          4996 => x"2c",
          4997 => x"f0",
          4998 => x"51",
          4999 => x"81",
          5000 => x"87",
          5001 => x"ee",
          5002 => x"57",
          5003 => x"3d",
          5004 => x"3d",
          5005 => x"af",
          5006 => x"f0",
          5007 => x"fe",
          5008 => x"38",
          5009 => x"51",
          5010 => x"81",
          5011 => x"55",
          5012 => x"08",
          5013 => x"80",
          5014 => x"70",
          5015 => x"58",
          5016 => x"85",
          5017 => x"8d",
          5018 => x"2e",
          5019 => x"52",
          5020 => x"be",
          5021 => x"fe",
          5022 => x"3d",
          5023 => x"3d",
          5024 => x"55",
          5025 => x"92",
          5026 => x"52",
          5027 => x"de",
          5028 => x"fe",
          5029 => x"81",
          5030 => x"82",
          5031 => x"74",
          5032 => x"98",
          5033 => x"11",
          5034 => x"59",
          5035 => x"75",
          5036 => x"38",
          5037 => x"81",
          5038 => x"5b",
          5039 => x"82",
          5040 => x"39",
          5041 => x"08",
          5042 => x"59",
          5043 => x"09",
          5044 => x"38",
          5045 => x"57",
          5046 => x"3d",
          5047 => x"c1",
          5048 => x"fe",
          5049 => x"2e",
          5050 => x"fe",
          5051 => x"2e",
          5052 => x"fe",
          5053 => x"70",
          5054 => x"08",
          5055 => x"7a",
          5056 => x"7f",
          5057 => x"54",
          5058 => x"77",
          5059 => x"80",
          5060 => x"15",
          5061 => x"f0",
          5062 => x"75",
          5063 => x"52",
          5064 => x"52",
          5065 => x"8d",
          5066 => x"f0",
          5067 => x"fe",
          5068 => x"d6",
          5069 => x"33",
          5070 => x"1a",
          5071 => x"54",
          5072 => x"09",
          5073 => x"38",
          5074 => x"ff",
          5075 => x"81",
          5076 => x"83",
          5077 => x"70",
          5078 => x"25",
          5079 => x"59",
          5080 => x"9b",
          5081 => x"51",
          5082 => x"3f",
          5083 => x"08",
          5084 => x"70",
          5085 => x"25",
          5086 => x"59",
          5087 => x"75",
          5088 => x"7a",
          5089 => x"ff",
          5090 => x"7c",
          5091 => x"90",
          5092 => x"11",
          5093 => x"56",
          5094 => x"15",
          5095 => x"fe",
          5096 => x"3d",
          5097 => x"3d",
          5098 => x"3d",
          5099 => x"70",
          5100 => x"dd",
          5101 => x"f0",
          5102 => x"fe",
          5103 => x"a8",
          5104 => x"33",
          5105 => x"a0",
          5106 => x"33",
          5107 => x"70",
          5108 => x"55",
          5109 => x"73",
          5110 => x"8e",
          5111 => x"08",
          5112 => x"18",
          5113 => x"80",
          5114 => x"38",
          5115 => x"08",
          5116 => x"08",
          5117 => x"c4",
          5118 => x"fe",
          5119 => x"88",
          5120 => x"80",
          5121 => x"17",
          5122 => x"51",
          5123 => x"3f",
          5124 => x"08",
          5125 => x"81",
          5126 => x"81",
          5127 => x"f0",
          5128 => x"09",
          5129 => x"38",
          5130 => x"39",
          5131 => x"77",
          5132 => x"f0",
          5133 => x"08",
          5134 => x"98",
          5135 => x"81",
          5136 => x"52",
          5137 => x"bd",
          5138 => x"f0",
          5139 => x"17",
          5140 => x"0c",
          5141 => x"80",
          5142 => x"73",
          5143 => x"75",
          5144 => x"38",
          5145 => x"34",
          5146 => x"81",
          5147 => x"89",
          5148 => x"e2",
          5149 => x"53",
          5150 => x"a4",
          5151 => x"3d",
          5152 => x"3f",
          5153 => x"08",
          5154 => x"f0",
          5155 => x"38",
          5156 => x"3d",
          5157 => x"3d",
          5158 => x"d1",
          5159 => x"fe",
          5160 => x"81",
          5161 => x"81",
          5162 => x"80",
          5163 => x"70",
          5164 => x"81",
          5165 => x"56",
          5166 => x"81",
          5167 => x"98",
          5168 => x"74",
          5169 => x"38",
          5170 => x"05",
          5171 => x"06",
          5172 => x"55",
          5173 => x"38",
          5174 => x"51",
          5175 => x"81",
          5176 => x"74",
          5177 => x"81",
          5178 => x"56",
          5179 => x"80",
          5180 => x"54",
          5181 => x"08",
          5182 => x"2e",
          5183 => x"73",
          5184 => x"f0",
          5185 => x"52",
          5186 => x"52",
          5187 => x"3f",
          5188 => x"08",
          5189 => x"f0",
          5190 => x"38",
          5191 => x"08",
          5192 => x"cc",
          5193 => x"fe",
          5194 => x"81",
          5195 => x"86",
          5196 => x"80",
          5197 => x"fe",
          5198 => x"2e",
          5199 => x"fe",
          5200 => x"c0",
          5201 => x"ce",
          5202 => x"fe",
          5203 => x"fe",
          5204 => x"70",
          5205 => x"08",
          5206 => x"51",
          5207 => x"80",
          5208 => x"73",
          5209 => x"38",
          5210 => x"52",
          5211 => x"95",
          5212 => x"f0",
          5213 => x"8c",
          5214 => x"ff",
          5215 => x"81",
          5216 => x"55",
          5217 => x"f0",
          5218 => x"0d",
          5219 => x"0d",
          5220 => x"3d",
          5221 => x"9a",
          5222 => x"cb",
          5223 => x"f0",
          5224 => x"fe",
          5225 => x"b0",
          5226 => x"69",
          5227 => x"70",
          5228 => x"97",
          5229 => x"f0",
          5230 => x"fe",
          5231 => x"38",
          5232 => x"94",
          5233 => x"f0",
          5234 => x"09",
          5235 => x"88",
          5236 => x"df",
          5237 => x"85",
          5238 => x"51",
          5239 => x"74",
          5240 => x"78",
          5241 => x"8a",
          5242 => x"57",
          5243 => x"81",
          5244 => x"75",
          5245 => x"fe",
          5246 => x"38",
          5247 => x"fe",
          5248 => x"2e",
          5249 => x"83",
          5250 => x"81",
          5251 => x"ff",
          5252 => x"06",
          5253 => x"54",
          5254 => x"73",
          5255 => x"81",
          5256 => x"52",
          5257 => x"a4",
          5258 => x"f0",
          5259 => x"fe",
          5260 => x"9a",
          5261 => x"a0",
          5262 => x"51",
          5263 => x"3f",
          5264 => x"0b",
          5265 => x"78",
          5266 => x"bf",
          5267 => x"88",
          5268 => x"80",
          5269 => x"ff",
          5270 => x"75",
          5271 => x"11",
          5272 => x"f8",
          5273 => x"78",
          5274 => x"80",
          5275 => x"ff",
          5276 => x"78",
          5277 => x"80",
          5278 => x"7f",
          5279 => x"d4",
          5280 => x"c9",
          5281 => x"54",
          5282 => x"15",
          5283 => x"cb",
          5284 => x"fe",
          5285 => x"81",
          5286 => x"b2",
          5287 => x"b2",
          5288 => x"96",
          5289 => x"b5",
          5290 => x"53",
          5291 => x"51",
          5292 => x"64",
          5293 => x"8b",
          5294 => x"54",
          5295 => x"15",
          5296 => x"ff",
          5297 => x"81",
          5298 => x"54",
          5299 => x"53",
          5300 => x"51",
          5301 => x"3f",
          5302 => x"f0",
          5303 => x"0d",
          5304 => x"0d",
          5305 => x"05",
          5306 => x"3f",
          5307 => x"3d",
          5308 => x"52",
          5309 => x"d5",
          5310 => x"fe",
          5311 => x"81",
          5312 => x"82",
          5313 => x"4d",
          5314 => x"52",
          5315 => x"52",
          5316 => x"3f",
          5317 => x"08",
          5318 => x"f0",
          5319 => x"38",
          5320 => x"05",
          5321 => x"06",
          5322 => x"73",
          5323 => x"a0",
          5324 => x"08",
          5325 => x"ff",
          5326 => x"ff",
          5327 => x"ac",
          5328 => x"92",
          5329 => x"54",
          5330 => x"3f",
          5331 => x"52",
          5332 => x"f7",
          5333 => x"f0",
          5334 => x"fe",
          5335 => x"38",
          5336 => x"09",
          5337 => x"38",
          5338 => x"08",
          5339 => x"88",
          5340 => x"39",
          5341 => x"08",
          5342 => x"81",
          5343 => x"38",
          5344 => x"b1",
          5345 => x"f0",
          5346 => x"fe",
          5347 => x"c8",
          5348 => x"93",
          5349 => x"ff",
          5350 => x"8d",
          5351 => x"b4",
          5352 => x"af",
          5353 => x"17",
          5354 => x"33",
          5355 => x"70",
          5356 => x"55",
          5357 => x"38",
          5358 => x"54",
          5359 => x"34",
          5360 => x"0b",
          5361 => x"8b",
          5362 => x"84",
          5363 => x"06",
          5364 => x"73",
          5365 => x"e5",
          5366 => x"2e",
          5367 => x"75",
          5368 => x"c6",
          5369 => x"fe",
          5370 => x"78",
          5371 => x"bb",
          5372 => x"81",
          5373 => x"80",
          5374 => x"38",
          5375 => x"08",
          5376 => x"ff",
          5377 => x"81",
          5378 => x"79",
          5379 => x"58",
          5380 => x"fe",
          5381 => x"c0",
          5382 => x"33",
          5383 => x"2e",
          5384 => x"99",
          5385 => x"75",
          5386 => x"c6",
          5387 => x"54",
          5388 => x"15",
          5389 => x"81",
          5390 => x"9c",
          5391 => x"c8",
          5392 => x"fe",
          5393 => x"81",
          5394 => x"8c",
          5395 => x"ff",
          5396 => x"81",
          5397 => x"55",
          5398 => x"f0",
          5399 => x"0d",
          5400 => x"0d",
          5401 => x"05",
          5402 => x"05",
          5403 => x"33",
          5404 => x"53",
          5405 => x"05",
          5406 => x"51",
          5407 => x"81",
          5408 => x"55",
          5409 => x"08",
          5410 => x"78",
          5411 => x"95",
          5412 => x"51",
          5413 => x"81",
          5414 => x"55",
          5415 => x"08",
          5416 => x"80",
          5417 => x"81",
          5418 => x"86",
          5419 => x"38",
          5420 => x"61",
          5421 => x"12",
          5422 => x"7a",
          5423 => x"51",
          5424 => x"74",
          5425 => x"78",
          5426 => x"83",
          5427 => x"51",
          5428 => x"3f",
          5429 => x"08",
          5430 => x"fe",
          5431 => x"3d",
          5432 => x"3d",
          5433 => x"82",
          5434 => x"d0",
          5435 => x"3d",
          5436 => x"3f",
          5437 => x"08",
          5438 => x"f0",
          5439 => x"38",
          5440 => x"52",
          5441 => x"05",
          5442 => x"3f",
          5443 => x"08",
          5444 => x"f0",
          5445 => x"02",
          5446 => x"33",
          5447 => x"54",
          5448 => x"a6",
          5449 => x"22",
          5450 => x"71",
          5451 => x"53",
          5452 => x"51",
          5453 => x"3f",
          5454 => x"0b",
          5455 => x"76",
          5456 => x"b8",
          5457 => x"f0",
          5458 => x"81",
          5459 => x"93",
          5460 => x"ea",
          5461 => x"6b",
          5462 => x"53",
          5463 => x"05",
          5464 => x"51",
          5465 => x"81",
          5466 => x"81",
          5467 => x"30",
          5468 => x"f0",
          5469 => x"25",
          5470 => x"79",
          5471 => x"85",
          5472 => x"75",
          5473 => x"73",
          5474 => x"f9",
          5475 => x"80",
          5476 => x"8d",
          5477 => x"54",
          5478 => x"3f",
          5479 => x"08",
          5480 => x"f0",
          5481 => x"38",
          5482 => x"51",
          5483 => x"81",
          5484 => x"57",
          5485 => x"08",
          5486 => x"fe",
          5487 => x"fe",
          5488 => x"5b",
          5489 => x"18",
          5490 => x"18",
          5491 => x"74",
          5492 => x"81",
          5493 => x"78",
          5494 => x"8b",
          5495 => x"54",
          5496 => x"75",
          5497 => x"38",
          5498 => x"1b",
          5499 => x"55",
          5500 => x"2e",
          5501 => x"39",
          5502 => x"09",
          5503 => x"38",
          5504 => x"80",
          5505 => x"70",
          5506 => x"25",
          5507 => x"80",
          5508 => x"38",
          5509 => x"bc",
          5510 => x"11",
          5511 => x"ff",
          5512 => x"81",
          5513 => x"57",
          5514 => x"08",
          5515 => x"70",
          5516 => x"80",
          5517 => x"83",
          5518 => x"80",
          5519 => x"84",
          5520 => x"a7",
          5521 => x"b4",
          5522 => x"ad",
          5523 => x"fe",
          5524 => x"0c",
          5525 => x"f0",
          5526 => x"0d",
          5527 => x"0d",
          5528 => x"3d",
          5529 => x"52",
          5530 => x"ce",
          5531 => x"fe",
          5532 => x"fe",
          5533 => x"54",
          5534 => x"08",
          5535 => x"8b",
          5536 => x"8b",
          5537 => x"59",
          5538 => x"3f",
          5539 => x"33",
          5540 => x"06",
          5541 => x"57",
          5542 => x"81",
          5543 => x"58",
          5544 => x"06",
          5545 => x"4e",
          5546 => x"ff",
          5547 => x"81",
          5548 => x"80",
          5549 => x"6c",
          5550 => x"53",
          5551 => x"ae",
          5552 => x"fe",
          5553 => x"2e",
          5554 => x"88",
          5555 => x"6d",
          5556 => x"55",
          5557 => x"fe",
          5558 => x"ff",
          5559 => x"83",
          5560 => x"51",
          5561 => x"26",
          5562 => x"15",
          5563 => x"ff",
          5564 => x"80",
          5565 => x"87",
          5566 => x"dc",
          5567 => x"74",
          5568 => x"38",
          5569 => x"ec",
          5570 => x"ae",
          5571 => x"fe",
          5572 => x"38",
          5573 => x"27",
          5574 => x"89",
          5575 => x"8b",
          5576 => x"27",
          5577 => x"55",
          5578 => x"81",
          5579 => x"8f",
          5580 => x"2a",
          5581 => x"70",
          5582 => x"34",
          5583 => x"74",
          5584 => x"05",
          5585 => x"17",
          5586 => x"70",
          5587 => x"52",
          5588 => x"73",
          5589 => x"c8",
          5590 => x"33",
          5591 => x"73",
          5592 => x"81",
          5593 => x"80",
          5594 => x"02",
          5595 => x"76",
          5596 => x"51",
          5597 => x"2e",
          5598 => x"87",
          5599 => x"57",
          5600 => x"79",
          5601 => x"80",
          5602 => x"70",
          5603 => x"ba",
          5604 => x"fe",
          5605 => x"81",
          5606 => x"80",
          5607 => x"52",
          5608 => x"bf",
          5609 => x"fe",
          5610 => x"81",
          5611 => x"8d",
          5612 => x"c4",
          5613 => x"e5",
          5614 => x"c6",
          5615 => x"f0",
          5616 => x"09",
          5617 => x"cc",
          5618 => x"76",
          5619 => x"c4",
          5620 => x"74",
          5621 => x"b0",
          5622 => x"f0",
          5623 => x"fe",
          5624 => x"38",
          5625 => x"fe",
          5626 => x"67",
          5627 => x"db",
          5628 => x"88",
          5629 => x"34",
          5630 => x"52",
          5631 => x"ab",
          5632 => x"54",
          5633 => x"15",
          5634 => x"ff",
          5635 => x"81",
          5636 => x"54",
          5637 => x"81",
          5638 => x"9c",
          5639 => x"f2",
          5640 => x"62",
          5641 => x"80",
          5642 => x"93",
          5643 => x"55",
          5644 => x"5e",
          5645 => x"3f",
          5646 => x"08",
          5647 => x"f0",
          5648 => x"38",
          5649 => x"58",
          5650 => x"38",
          5651 => x"97",
          5652 => x"08",
          5653 => x"38",
          5654 => x"70",
          5655 => x"81",
          5656 => x"55",
          5657 => x"87",
          5658 => x"39",
          5659 => x"90",
          5660 => x"82",
          5661 => x"8a",
          5662 => x"89",
          5663 => x"7f",
          5664 => x"56",
          5665 => x"3f",
          5666 => x"06",
          5667 => x"72",
          5668 => x"81",
          5669 => x"05",
          5670 => x"7c",
          5671 => x"55",
          5672 => x"27",
          5673 => x"16",
          5674 => x"83",
          5675 => x"76",
          5676 => x"80",
          5677 => x"79",
          5678 => x"99",
          5679 => x"7f",
          5680 => x"14",
          5681 => x"83",
          5682 => x"81",
          5683 => x"81",
          5684 => x"38",
          5685 => x"08",
          5686 => x"95",
          5687 => x"f0",
          5688 => x"81",
          5689 => x"7b",
          5690 => x"06",
          5691 => x"39",
          5692 => x"56",
          5693 => x"09",
          5694 => x"b9",
          5695 => x"80",
          5696 => x"80",
          5697 => x"78",
          5698 => x"7a",
          5699 => x"38",
          5700 => x"73",
          5701 => x"81",
          5702 => x"ff",
          5703 => x"74",
          5704 => x"ff",
          5705 => x"81",
          5706 => x"58",
          5707 => x"08",
          5708 => x"74",
          5709 => x"16",
          5710 => x"73",
          5711 => x"39",
          5712 => x"7e",
          5713 => x"0c",
          5714 => x"2e",
          5715 => x"88",
          5716 => x"8c",
          5717 => x"1a",
          5718 => x"07",
          5719 => x"1b",
          5720 => x"08",
          5721 => x"16",
          5722 => x"75",
          5723 => x"38",
          5724 => x"90",
          5725 => x"15",
          5726 => x"54",
          5727 => x"34",
          5728 => x"81",
          5729 => x"90",
          5730 => x"e9",
          5731 => x"6d",
          5732 => x"80",
          5733 => x"9d",
          5734 => x"5c",
          5735 => x"3f",
          5736 => x"0b",
          5737 => x"08",
          5738 => x"38",
          5739 => x"08",
          5740 => x"ff",
          5741 => x"08",
          5742 => x"80",
          5743 => x"80",
          5744 => x"fe",
          5745 => x"ff",
          5746 => x"52",
          5747 => x"a0",
          5748 => x"fe",
          5749 => x"ff",
          5750 => x"06",
          5751 => x"56",
          5752 => x"38",
          5753 => x"70",
          5754 => x"55",
          5755 => x"8b",
          5756 => x"3d",
          5757 => x"83",
          5758 => x"ff",
          5759 => x"81",
          5760 => x"99",
          5761 => x"74",
          5762 => x"38",
          5763 => x"80",
          5764 => x"ff",
          5765 => x"55",
          5766 => x"83",
          5767 => x"78",
          5768 => x"38",
          5769 => x"26",
          5770 => x"81",
          5771 => x"8b",
          5772 => x"79",
          5773 => x"80",
          5774 => x"93",
          5775 => x"39",
          5776 => x"6e",
          5777 => x"89",
          5778 => x"48",
          5779 => x"83",
          5780 => x"61",
          5781 => x"25",
          5782 => x"55",
          5783 => x"8a",
          5784 => x"3d",
          5785 => x"81",
          5786 => x"ff",
          5787 => x"81",
          5788 => x"f0",
          5789 => x"38",
          5790 => x"70",
          5791 => x"fe",
          5792 => x"56",
          5793 => x"38",
          5794 => x"55",
          5795 => x"75",
          5796 => x"38",
          5797 => x"70",
          5798 => x"ff",
          5799 => x"83",
          5800 => x"78",
          5801 => x"89",
          5802 => x"81",
          5803 => x"06",
          5804 => x"80",
          5805 => x"77",
          5806 => x"74",
          5807 => x"8d",
          5808 => x"06",
          5809 => x"2e",
          5810 => x"77",
          5811 => x"93",
          5812 => x"74",
          5813 => x"cb",
          5814 => x"7d",
          5815 => x"81",
          5816 => x"38",
          5817 => x"66",
          5818 => x"81",
          5819 => x"80",
          5820 => x"74",
          5821 => x"38",
          5822 => x"98",
          5823 => x"80",
          5824 => x"82",
          5825 => x"57",
          5826 => x"80",
          5827 => x"76",
          5828 => x"38",
          5829 => x"51",
          5830 => x"3f",
          5831 => x"08",
          5832 => x"87",
          5833 => x"2a",
          5834 => x"5c",
          5835 => x"fe",
          5836 => x"80",
          5837 => x"44",
          5838 => x"0a",
          5839 => x"ec",
          5840 => x"39",
          5841 => x"66",
          5842 => x"81",
          5843 => x"f0",
          5844 => x"74",
          5845 => x"38",
          5846 => x"98",
          5847 => x"f0",
          5848 => x"82",
          5849 => x"57",
          5850 => x"80",
          5851 => x"76",
          5852 => x"38",
          5853 => x"51",
          5854 => x"3f",
          5855 => x"08",
          5856 => x"57",
          5857 => x"08",
          5858 => x"96",
          5859 => x"81",
          5860 => x"10",
          5861 => x"08",
          5862 => x"72",
          5863 => x"59",
          5864 => x"ff",
          5865 => x"5d",
          5866 => x"44",
          5867 => x"11",
          5868 => x"70",
          5869 => x"71",
          5870 => x"06",
          5871 => x"52",
          5872 => x"40",
          5873 => x"09",
          5874 => x"38",
          5875 => x"18",
          5876 => x"39",
          5877 => x"79",
          5878 => x"70",
          5879 => x"58",
          5880 => x"76",
          5881 => x"38",
          5882 => x"7d",
          5883 => x"70",
          5884 => x"55",
          5885 => x"3f",
          5886 => x"08",
          5887 => x"2e",
          5888 => x"9b",
          5889 => x"f0",
          5890 => x"f5",
          5891 => x"38",
          5892 => x"38",
          5893 => x"59",
          5894 => x"38",
          5895 => x"7d",
          5896 => x"81",
          5897 => x"38",
          5898 => x"0b",
          5899 => x"08",
          5900 => x"78",
          5901 => x"1a",
          5902 => x"c0",
          5903 => x"74",
          5904 => x"39",
          5905 => x"55",
          5906 => x"8f",
          5907 => x"fd",
          5908 => x"fe",
          5909 => x"f5",
          5910 => x"78",
          5911 => x"79",
          5912 => x"80",
          5913 => x"f1",
          5914 => x"39",
          5915 => x"81",
          5916 => x"06",
          5917 => x"55",
          5918 => x"27",
          5919 => x"81",
          5920 => x"56",
          5921 => x"38",
          5922 => x"80",
          5923 => x"ff",
          5924 => x"8b",
          5925 => x"98",
          5926 => x"ff",
          5927 => x"84",
          5928 => x"1b",
          5929 => x"b3",
          5930 => x"1c",
          5931 => x"ff",
          5932 => x"8e",
          5933 => x"a1",
          5934 => x"0b",
          5935 => x"7d",
          5936 => x"30",
          5937 => x"84",
          5938 => x"51",
          5939 => x"51",
          5940 => x"3f",
          5941 => x"83",
          5942 => x"90",
          5943 => x"ff",
          5944 => x"93",
          5945 => x"a0",
          5946 => x"39",
          5947 => x"1b",
          5948 => x"85",
          5949 => x"95",
          5950 => x"52",
          5951 => x"ff",
          5952 => x"81",
          5953 => x"1b",
          5954 => x"cf",
          5955 => x"9c",
          5956 => x"a0",
          5957 => x"83",
          5958 => x"06",
          5959 => x"82",
          5960 => x"52",
          5961 => x"51",
          5962 => x"3f",
          5963 => x"1b",
          5964 => x"c5",
          5965 => x"ac",
          5966 => x"a0",
          5967 => x"52",
          5968 => x"ff",
          5969 => x"86",
          5970 => x"51",
          5971 => x"3f",
          5972 => x"80",
          5973 => x"a9",
          5974 => x"1c",
          5975 => x"81",
          5976 => x"80",
          5977 => x"ae",
          5978 => x"b2",
          5979 => x"1b",
          5980 => x"85",
          5981 => x"ff",
          5982 => x"96",
          5983 => x"9f",
          5984 => x"80",
          5985 => x"34",
          5986 => x"1c",
          5987 => x"81",
          5988 => x"ab",
          5989 => x"a0",
          5990 => x"d4",
          5991 => x"fe",
          5992 => x"59",
          5993 => x"3f",
          5994 => x"53",
          5995 => x"51",
          5996 => x"3f",
          5997 => x"fe",
          5998 => x"e7",
          5999 => x"2e",
          6000 => x"80",
          6001 => x"54",
          6002 => x"53",
          6003 => x"51",
          6004 => x"3f",
          6005 => x"80",
          6006 => x"ff",
          6007 => x"84",
          6008 => x"d2",
          6009 => x"ff",
          6010 => x"86",
          6011 => x"f2",
          6012 => x"1b",
          6013 => x"81",
          6014 => x"52",
          6015 => x"51",
          6016 => x"3f",
          6017 => x"ec",
          6018 => x"9e",
          6019 => x"d4",
          6020 => x"51",
          6021 => x"3f",
          6022 => x"87",
          6023 => x"52",
          6024 => x"9a",
          6025 => x"54",
          6026 => x"7a",
          6027 => x"ff",
          6028 => x"65",
          6029 => x"7a",
          6030 => x"8f",
          6031 => x"80",
          6032 => x"2e",
          6033 => x"9a",
          6034 => x"7a",
          6035 => x"a9",
          6036 => x"84",
          6037 => x"9e",
          6038 => x"0a",
          6039 => x"51",
          6040 => x"ff",
          6041 => x"7d",
          6042 => x"38",
          6043 => x"52",
          6044 => x"9e",
          6045 => x"55",
          6046 => x"62",
          6047 => x"74",
          6048 => x"75",
          6049 => x"7e",
          6050 => x"fe",
          6051 => x"f0",
          6052 => x"38",
          6053 => x"81",
          6054 => x"52",
          6055 => x"9e",
          6056 => x"16",
          6057 => x"56",
          6058 => x"38",
          6059 => x"77",
          6060 => x"8d",
          6061 => x"7d",
          6062 => x"38",
          6063 => x"57",
          6064 => x"83",
          6065 => x"76",
          6066 => x"7a",
          6067 => x"ff",
          6068 => x"81",
          6069 => x"81",
          6070 => x"16",
          6071 => x"56",
          6072 => x"38",
          6073 => x"83",
          6074 => x"86",
          6075 => x"ff",
          6076 => x"38",
          6077 => x"82",
          6078 => x"81",
          6079 => x"06",
          6080 => x"fe",
          6081 => x"53",
          6082 => x"51",
          6083 => x"3f",
          6084 => x"52",
          6085 => x"9c",
          6086 => x"be",
          6087 => x"75",
          6088 => x"81",
          6089 => x"0b",
          6090 => x"77",
          6091 => x"75",
          6092 => x"60",
          6093 => x"80",
          6094 => x"75",
          6095 => x"ee",
          6096 => x"85",
          6097 => x"fe",
          6098 => x"2a",
          6099 => x"75",
          6100 => x"81",
          6101 => x"87",
          6102 => x"52",
          6103 => x"51",
          6104 => x"3f",
          6105 => x"ca",
          6106 => x"9c",
          6107 => x"54",
          6108 => x"52",
          6109 => x"98",
          6110 => x"56",
          6111 => x"08",
          6112 => x"53",
          6113 => x"51",
          6114 => x"3f",
          6115 => x"fe",
          6116 => x"38",
          6117 => x"56",
          6118 => x"56",
          6119 => x"fe",
          6120 => x"75",
          6121 => x"0c",
          6122 => x"04",
          6123 => x"7d",
          6124 => x"80",
          6125 => x"05",
          6126 => x"76",
          6127 => x"38",
          6128 => x"11",
          6129 => x"53",
          6130 => x"79",
          6131 => x"3f",
          6132 => x"09",
          6133 => x"38",
          6134 => x"55",
          6135 => x"db",
          6136 => x"70",
          6137 => x"34",
          6138 => x"74",
          6139 => x"81",
          6140 => x"80",
          6141 => x"55",
          6142 => x"76",
          6143 => x"fe",
          6144 => x"3d",
          6145 => x"3d",
          6146 => x"84",
          6147 => x"33",
          6148 => x"8a",
          6149 => x"06",
          6150 => x"52",
          6151 => x"3f",
          6152 => x"56",
          6153 => x"be",
          6154 => x"08",
          6155 => x"05",
          6156 => x"75",
          6157 => x"56",
          6158 => x"a1",
          6159 => x"fc",
          6160 => x"53",
          6161 => x"76",
          6162 => x"dc",
          6163 => x"32",
          6164 => x"72",
          6165 => x"70",
          6166 => x"56",
          6167 => x"18",
          6168 => x"88",
          6169 => x"3d",
          6170 => x"3d",
          6171 => x"11",
          6172 => x"80",
          6173 => x"38",
          6174 => x"05",
          6175 => x"8c",
          6176 => x"08",
          6177 => x"3f",
          6178 => x"08",
          6179 => x"16",
          6180 => x"09",
          6181 => x"38",
          6182 => x"55",
          6183 => x"55",
          6184 => x"f0",
          6185 => x"0d",
          6186 => x"0d",
          6187 => x"cc",
          6188 => x"73",
          6189 => x"93",
          6190 => x"0c",
          6191 => x"04",
          6192 => x"02",
          6193 => x"33",
          6194 => x"3d",
          6195 => x"54",
          6196 => x"52",
          6197 => x"ae",
          6198 => x"ff",
          6199 => x"3d",
          6200 => x"3d",
          6201 => x"08",
          6202 => x"59",
          6203 => x"80",
          6204 => x"39",
          6205 => x"0c",
          6206 => x"54",
          6207 => x"74",
          6208 => x"a0",
          6209 => x"06",
          6210 => x"15",
          6211 => x"80",
          6212 => x"29",
          6213 => x"05",
          6214 => x"56",
          6215 => x"3f",
          6216 => x"08",
          6217 => x"08",
          6218 => x"76",
          6219 => x"fe",
          6220 => x"81",
          6221 => x"8b",
          6222 => x"33",
          6223 => x"2e",
          6224 => x"81",
          6225 => x"ff",
          6226 => x"98",
          6227 => x"38",
          6228 => x"81",
          6229 => x"8a",
          6230 => x"ff",
          6231 => x"52",
          6232 => x"81",
          6233 => x"84",
          6234 => x"84",
          6235 => x"08",
          6236 => x"b8",
          6237 => x"39",
          6238 => x"51",
          6239 => x"81",
          6240 => x"80",
          6241 => x"ee",
          6242 => x"eb",
          6243 => x"fc",
          6244 => x"39",
          6245 => x"51",
          6246 => x"81",
          6247 => x"80",
          6248 => x"ef",
          6249 => x"cf",
          6250 => x"c8",
          6251 => x"39",
          6252 => x"51",
          6253 => x"81",
          6254 => x"bb",
          6255 => x"94",
          6256 => x"81",
          6257 => x"af",
          6258 => x"d4",
          6259 => x"81",
          6260 => x"a3",
          6261 => x"88",
          6262 => x"81",
          6263 => x"97",
          6264 => x"b4",
          6265 => x"81",
          6266 => x"8b",
          6267 => x"e4",
          6268 => x"81",
          6269 => x"fe",
          6270 => x"83",
          6271 => x"fb",
          6272 => x"79",
          6273 => x"87",
          6274 => x"38",
          6275 => x"87",
          6276 => x"91",
          6277 => x"52",
          6278 => x"cf",
          6279 => x"fe",
          6280 => x"75",
          6281 => x"86",
          6282 => x"f0",
          6283 => x"53",
          6284 => x"f2",
          6285 => x"f7",
          6286 => x"3d",
          6287 => x"3d",
          6288 => x"84",
          6289 => x"05",
          6290 => x"80",
          6291 => x"70",
          6292 => x"25",
          6293 => x"59",
          6294 => x"87",
          6295 => x"38",
          6296 => x"76",
          6297 => x"ff",
          6298 => x"93",
          6299 => x"80",
          6300 => x"76",
          6301 => x"70",
          6302 => x"bf",
          6303 => x"fe",
          6304 => x"81",
          6305 => x"b8",
          6306 => x"f0",
          6307 => x"98",
          6308 => x"fe",
          6309 => x"96",
          6310 => x"54",
          6311 => x"77",
          6312 => x"c4",
          6313 => x"fe",
          6314 => x"81",
          6315 => x"90",
          6316 => x"74",
          6317 => x"38",
          6318 => x"19",
          6319 => x"39",
          6320 => x"05",
          6321 => x"3f",
          6322 => x"78",
          6323 => x"7b",
          6324 => x"2a",
          6325 => x"57",
          6326 => x"80",
          6327 => x"81",
          6328 => x"87",
          6329 => x"08",
          6330 => x"fe",
          6331 => x"56",
          6332 => x"f0",
          6333 => x"0d",
          6334 => x"0d",
          6335 => x"05",
          6336 => x"57",
          6337 => x"80",
          6338 => x"79",
          6339 => x"3f",
          6340 => x"08",
          6341 => x"80",
          6342 => x"75",
          6343 => x"38",
          6344 => x"55",
          6345 => x"fe",
          6346 => x"52",
          6347 => x"2d",
          6348 => x"08",
          6349 => x"77",
          6350 => x"fe",
          6351 => x"3d",
          6352 => x"3d",
          6353 => x"63",
          6354 => x"80",
          6355 => x"73",
          6356 => x"41",
          6357 => x"5e",
          6358 => x"52",
          6359 => x"51",
          6360 => x"3f",
          6361 => x"51",
          6362 => x"3f",
          6363 => x"79",
          6364 => x"38",
          6365 => x"89",
          6366 => x"2e",
          6367 => x"c6",
          6368 => x"53",
          6369 => x"8e",
          6370 => x"52",
          6371 => x"51",
          6372 => x"3f",
          6373 => x"f2",
          6374 => x"ef",
          6375 => x"15",
          6376 => x"39",
          6377 => x"72",
          6378 => x"38",
          6379 => x"81",
          6380 => x"fe",
          6381 => x"89",
          6382 => x"c0",
          6383 => x"e8",
          6384 => x"55",
          6385 => x"18",
          6386 => x"27",
          6387 => x"33",
          6388 => x"cc",
          6389 => x"b4",
          6390 => x"81",
          6391 => x"fe",
          6392 => x"81",
          6393 => x"51",
          6394 => x"3f",
          6395 => x"81",
          6396 => x"fe",
          6397 => x"80",
          6398 => x"27",
          6399 => x"18",
          6400 => x"53",
          6401 => x"7a",
          6402 => x"81",
          6403 => x"9f",
          6404 => x"38",
          6405 => x"73",
          6406 => x"ff",
          6407 => x"72",
          6408 => x"38",
          6409 => x"26",
          6410 => x"51",
          6411 => x"51",
          6412 => x"3f",
          6413 => x"c1",
          6414 => x"dc",
          6415 => x"e8",
          6416 => x"79",
          6417 => x"fe",
          6418 => x"81",
          6419 => x"98",
          6420 => x"2c",
          6421 => x"a0",
          6422 => x"06",
          6423 => x"dd",
          6424 => x"fe",
          6425 => x"2b",
          6426 => x"70",
          6427 => x"30",
          6428 => x"70",
          6429 => x"07",
          6430 => x"06",
          6431 => x"59",
          6432 => x"80",
          6433 => x"38",
          6434 => x"09",
          6435 => x"38",
          6436 => x"39",
          6437 => x"72",
          6438 => x"be",
          6439 => x"72",
          6440 => x"0c",
          6441 => x"04",
          6442 => x"02",
          6443 => x"81",
          6444 => x"81",
          6445 => x"55",
          6446 => x"3f",
          6447 => x"22",
          6448 => x"d7",
          6449 => x"f4",
          6450 => x"80",
          6451 => x"a1",
          6452 => x"f3",
          6453 => x"f2",
          6454 => x"80",
          6455 => x"fe",
          6456 => x"86",
          6457 => x"fe",
          6458 => x"c0",
          6459 => x"53",
          6460 => x"3f",
          6461 => x"d8",
          6462 => x"f3",
          6463 => x"da",
          6464 => x"51",
          6465 => x"3f",
          6466 => x"70",
          6467 => x"52",
          6468 => x"95",
          6469 => x"fe",
          6470 => x"81",
          6471 => x"fe",
          6472 => x"80",
          6473 => x"cc",
          6474 => x"2a",
          6475 => x"51",
          6476 => x"2e",
          6477 => x"51",
          6478 => x"3f",
          6479 => x"51",
          6480 => x"3f",
          6481 => x"d8",
          6482 => x"83",
          6483 => x"06",
          6484 => x"80",
          6485 => x"81",
          6486 => x"98",
          6487 => x"e4",
          6488 => x"90",
          6489 => x"fe",
          6490 => x"72",
          6491 => x"81",
          6492 => x"71",
          6493 => x"38",
          6494 => x"d7",
          6495 => x"f3",
          6496 => x"d9",
          6497 => x"51",
          6498 => x"3f",
          6499 => x"70",
          6500 => x"52",
          6501 => x"95",
          6502 => x"fe",
          6503 => x"81",
          6504 => x"fe",
          6505 => x"80",
          6506 => x"c8",
          6507 => x"2a",
          6508 => x"51",
          6509 => x"2e",
          6510 => x"51",
          6511 => x"3f",
          6512 => x"51",
          6513 => x"3f",
          6514 => x"d7",
          6515 => x"87",
          6516 => x"06",
          6517 => x"80",
          6518 => x"81",
          6519 => x"94",
          6520 => x"b4",
          6521 => x"8c",
          6522 => x"fe",
          6523 => x"72",
          6524 => x"81",
          6525 => x"71",
          6526 => x"38",
          6527 => x"d6",
          6528 => x"f4",
          6529 => x"d8",
          6530 => x"51",
          6531 => x"3f",
          6532 => x"3f",
          6533 => x"04",
          6534 => x"77",
          6535 => x"a3",
          6536 => x"55",
          6537 => x"52",
          6538 => x"ce",
          6539 => x"fb",
          6540 => x"73",
          6541 => x"53",
          6542 => x"52",
          6543 => x"51",
          6544 => x"3f",
          6545 => x"08",
          6546 => x"fe",
          6547 => x"80",
          6548 => x"31",
          6549 => x"73",
          6550 => x"34",
          6551 => x"33",
          6552 => x"2e",
          6553 => x"ac",
          6554 => x"88",
          6555 => x"75",
          6556 => x"3f",
          6557 => x"08",
          6558 => x"38",
          6559 => x"08",
          6560 => x"a4",
          6561 => x"82",
          6562 => x"c4",
          6563 => x"0b",
          6564 => x"34",
          6565 => x"33",
          6566 => x"2e",
          6567 => x"89",
          6568 => x"75",
          6569 => x"e4",
          6570 => x"81",
          6571 => x"87",
          6572 => x"ce",
          6573 => x"70",
          6574 => x"84",
          6575 => x"81",
          6576 => x"ff",
          6577 => x"81",
          6578 => x"81",
          6579 => x"78",
          6580 => x"81",
          6581 => x"81",
          6582 => x"96",
          6583 => x"59",
          6584 => x"3f",
          6585 => x"52",
          6586 => x"51",
          6587 => x"3f",
          6588 => x"08",
          6589 => x"38",
          6590 => x"51",
          6591 => x"81",
          6592 => x"81",
          6593 => x"fe",
          6594 => x"96",
          6595 => x"5a",
          6596 => x"79",
          6597 => x"3f",
          6598 => x"84",
          6599 => x"c2",
          6600 => x"f0",
          6601 => x"70",
          6602 => x"59",
          6603 => x"2e",
          6604 => x"78",
          6605 => x"80",
          6606 => x"ab",
          6607 => x"38",
          6608 => x"a4",
          6609 => x"2e",
          6610 => x"78",
          6611 => x"38",
          6612 => x"ff",
          6613 => x"a5",
          6614 => x"2e",
          6615 => x"78",
          6616 => x"b1",
          6617 => x"39",
          6618 => x"85",
          6619 => x"bd",
          6620 => x"78",
          6621 => x"af",
          6622 => x"2e",
          6623 => x"8e",
          6624 => x"bf",
          6625 => x"38",
          6626 => x"2e",
          6627 => x"8e",
          6628 => x"80",
          6629 => x"c2",
          6630 => x"d5",
          6631 => x"78",
          6632 => x"8c",
          6633 => x"80",
          6634 => x"38",
          6635 => x"2e",
          6636 => x"78",
          6637 => x"8b",
          6638 => x"c1",
          6639 => x"d1",
          6640 => x"38",
          6641 => x"2e",
          6642 => x"8e",
          6643 => x"81",
          6644 => x"86",
          6645 => x"82",
          6646 => x"78",
          6647 => x"8d",
          6648 => x"80",
          6649 => x"b4",
          6650 => x"39",
          6651 => x"2e",
          6652 => x"78",
          6653 => x"8d",
          6654 => x"81",
          6655 => x"ff",
          6656 => x"ff",
          6657 => x"fe",
          6658 => x"81",
          6659 => x"88",
          6660 => x"d8",
          6661 => x"39",
          6662 => x"fc",
          6663 => x"84",
          6664 => x"ed",
          6665 => x"fe",
          6666 => x"2e",
          6667 => x"63",
          6668 => x"80",
          6669 => x"cb",
          6670 => x"02",
          6671 => x"33",
          6672 => x"dd",
          6673 => x"f0",
          6674 => x"06",
          6675 => x"38",
          6676 => x"51",
          6677 => x"3f",
          6678 => x"a7",
          6679 => x"f8",
          6680 => x"39",
          6681 => x"80",
          6682 => x"84",
          6683 => x"ed",
          6684 => x"fe",
          6685 => x"2e",
          6686 => x"80",
          6687 => x"02",
          6688 => x"33",
          6689 => x"e6",
          6690 => x"f0",
          6691 => x"f6",
          6692 => x"bf",
          6693 => x"ff",
          6694 => x"ff",
          6695 => x"fe",
          6696 => x"81",
          6697 => x"80",
          6698 => x"63",
          6699 => x"d3",
          6700 => x"fe",
          6701 => x"ff",
          6702 => x"fe",
          6703 => x"81",
          6704 => x"86",
          6705 => x"f0",
          6706 => x"53",
          6707 => x"52",
          6708 => x"ea",
          6709 => x"80",
          6710 => x"53",
          6711 => x"84",
          6712 => x"80",
          6713 => x"ff",
          6714 => x"81",
          6715 => x"81",
          6716 => x"f5",
          6717 => x"e4",
          6718 => x"5d",
          6719 => x"b4",
          6720 => x"05",
          6721 => x"9d",
          6722 => x"f0",
          6723 => x"ff",
          6724 => x"5b",
          6725 => x"3f",
          6726 => x"fe",
          6727 => x"7a",
          6728 => x"3f",
          6729 => x"b4",
          6730 => x"05",
          6731 => x"f5",
          6732 => x"f0",
          6733 => x"ff",
          6734 => x"5b",
          6735 => x"3f",
          6736 => x"08",
          6737 => x"84",
          6738 => x"fe",
          6739 => x"81",
          6740 => x"b5",
          6741 => x"05",
          6742 => x"cd",
          6743 => x"f9",
          6744 => x"ff",
          6745 => x"56",
          6746 => x"fe",
          6747 => x"ff",
          6748 => x"53",
          6749 => x"51",
          6750 => x"81",
          6751 => x"80",
          6752 => x"38",
          6753 => x"08",
          6754 => x"3f",
          6755 => x"b4",
          6756 => x"11",
          6757 => x"05",
          6758 => x"e5",
          6759 => x"f0",
          6760 => x"fa",
          6761 => x"3d",
          6762 => x"53",
          6763 => x"51",
          6764 => x"3f",
          6765 => x"08",
          6766 => x"c7",
          6767 => x"fe",
          6768 => x"ff",
          6769 => x"fe",
          6770 => x"81",
          6771 => x"86",
          6772 => x"f0",
          6773 => x"f6",
          6774 => x"e2",
          6775 => x"63",
          6776 => x"7b",
          6777 => x"38",
          6778 => x"7a",
          6779 => x"5c",
          6780 => x"26",
          6781 => x"e1",
          6782 => x"ff",
          6783 => x"ff",
          6784 => x"fe",
          6785 => x"81",
          6786 => x"80",
          6787 => x"38",
          6788 => x"fc",
          6789 => x"84",
          6790 => x"e9",
          6791 => x"fe",
          6792 => x"2e",
          6793 => x"b4",
          6794 => x"11",
          6795 => x"05",
          6796 => x"cd",
          6797 => x"f0",
          6798 => x"f9",
          6799 => x"f6",
          6800 => x"e1",
          6801 => x"5a",
          6802 => x"81",
          6803 => x"59",
          6804 => x"05",
          6805 => x"34",
          6806 => x"42",
          6807 => x"3d",
          6808 => x"53",
          6809 => x"51",
          6810 => x"3f",
          6811 => x"08",
          6812 => x"8f",
          6813 => x"fe",
          6814 => x"ff",
          6815 => x"fe",
          6816 => x"81",
          6817 => x"80",
          6818 => x"38",
          6819 => x"f8",
          6820 => x"84",
          6821 => x"e8",
          6822 => x"fe",
          6823 => x"2e",
          6824 => x"81",
          6825 => x"fe",
          6826 => x"63",
          6827 => x"27",
          6828 => x"70",
          6829 => x"5e",
          6830 => x"7c",
          6831 => x"78",
          6832 => x"79",
          6833 => x"52",
          6834 => x"51",
          6835 => x"3f",
          6836 => x"81",
          6837 => x"d5",
          6838 => x"e4",
          6839 => x"39",
          6840 => x"80",
          6841 => x"84",
          6842 => x"e8",
          6843 => x"fe",
          6844 => x"df",
          6845 => x"b4",
          6846 => x"80",
          6847 => x"81",
          6848 => x"44",
          6849 => x"81",
          6850 => x"59",
          6851 => x"88",
          6852 => x"f4",
          6853 => x"39",
          6854 => x"33",
          6855 => x"2e",
          6856 => x"f9",
          6857 => x"ab",
          6858 => x"b7",
          6859 => x"80",
          6860 => x"81",
          6861 => x"44",
          6862 => x"fa",
          6863 => x"78",
          6864 => x"38",
          6865 => x"08",
          6866 => x"81",
          6867 => x"fc",
          6868 => x"b4",
          6869 => x"11",
          6870 => x"05",
          6871 => x"a1",
          6872 => x"f0",
          6873 => x"38",
          6874 => x"33",
          6875 => x"2e",
          6876 => x"f9",
          6877 => x"80",
          6878 => x"fa",
          6879 => x"78",
          6880 => x"38",
          6881 => x"08",
          6882 => x"81",
          6883 => x"59",
          6884 => x"88",
          6885 => x"80",
          6886 => x"39",
          6887 => x"33",
          6888 => x"2e",
          6889 => x"fa",
          6890 => x"99",
          6891 => x"b2",
          6892 => x"80",
          6893 => x"81",
          6894 => x"43",
          6895 => x"fa",
          6896 => x"05",
          6897 => x"fe",
          6898 => x"ff",
          6899 => x"fe",
          6900 => x"81",
          6901 => x"80",
          6902 => x"80",
          6903 => x"7a",
          6904 => x"38",
          6905 => x"90",
          6906 => x"70",
          6907 => x"2a",
          6908 => x"51",
          6909 => x"78",
          6910 => x"38",
          6911 => x"83",
          6912 => x"81",
          6913 => x"fe",
          6914 => x"a0",
          6915 => x"61",
          6916 => x"63",
          6917 => x"3f",
          6918 => x"51",
          6919 => x"3f",
          6920 => x"b4",
          6921 => x"11",
          6922 => x"05",
          6923 => x"d1",
          6924 => x"f0",
          6925 => x"f5",
          6926 => x"3d",
          6927 => x"53",
          6928 => x"51",
          6929 => x"3f",
          6930 => x"08",
          6931 => x"38",
          6932 => x"80",
          6933 => x"79",
          6934 => x"05",
          6935 => x"fe",
          6936 => x"ff",
          6937 => x"fe",
          6938 => x"81",
          6939 => x"e0",
          6940 => x"39",
          6941 => x"54",
          6942 => x"80",
          6943 => x"8c",
          6944 => x"52",
          6945 => x"e3",
          6946 => x"45",
          6947 => x"78",
          6948 => x"ef",
          6949 => x"27",
          6950 => x"3d",
          6951 => x"53",
          6952 => x"51",
          6953 => x"3f",
          6954 => x"08",
          6955 => x"38",
          6956 => x"80",
          6957 => x"79",
          6958 => x"05",
          6959 => x"39",
          6960 => x"51",
          6961 => x"3f",
          6962 => x"b4",
          6963 => x"11",
          6964 => x"05",
          6965 => x"9b",
          6966 => x"f0",
          6967 => x"f4",
          6968 => x"3d",
          6969 => x"53",
          6970 => x"51",
          6971 => x"3f",
          6972 => x"08",
          6973 => x"38",
          6974 => x"be",
          6975 => x"70",
          6976 => x"23",
          6977 => x"3d",
          6978 => x"53",
          6979 => x"51",
          6980 => x"3f",
          6981 => x"08",
          6982 => x"e7",
          6983 => x"22",
          6984 => x"f7",
          6985 => x"e1",
          6986 => x"f8",
          6987 => x"fe",
          6988 => x"79",
          6989 => x"59",
          6990 => x"f3",
          6991 => x"9f",
          6992 => x"60",
          6993 => x"d5",
          6994 => x"fe",
          6995 => x"ff",
          6996 => x"fe",
          6997 => x"81",
          6998 => x"80",
          6999 => x"60",
          7000 => x"05",
          7001 => x"82",
          7002 => x"78",
          7003 => x"39",
          7004 => x"51",
          7005 => x"3f",
          7006 => x"b4",
          7007 => x"11",
          7008 => x"05",
          7009 => x"eb",
          7010 => x"f0",
          7011 => x"f2",
          7012 => x"3d",
          7013 => x"53",
          7014 => x"51",
          7015 => x"3f",
          7016 => x"08",
          7017 => x"38",
          7018 => x"0c",
          7019 => x"05",
          7020 => x"fe",
          7021 => x"ff",
          7022 => x"fe",
          7023 => x"81",
          7024 => x"e4",
          7025 => x"39",
          7026 => x"54",
          7027 => x"a0",
          7028 => x"b8",
          7029 => x"52",
          7030 => x"e1",
          7031 => x"45",
          7032 => x"78",
          7033 => x"9b",
          7034 => x"27",
          7035 => x"3d",
          7036 => x"53",
          7037 => x"51",
          7038 => x"3f",
          7039 => x"08",
          7040 => x"38",
          7041 => x"0c",
          7042 => x"05",
          7043 => x"39",
          7044 => x"51",
          7045 => x"3f",
          7046 => x"81",
          7047 => x"fe",
          7048 => x"82",
          7049 => x"d7",
          7050 => x"39",
          7051 => x"51",
          7052 => x"3f",
          7053 => x"d4",
          7054 => x"c7",
          7055 => x"dc",
          7056 => x"e4",
          7057 => x"81",
          7058 => x"94",
          7059 => x"80",
          7060 => x"c0",
          7061 => x"f1",
          7062 => x"f7",
          7063 => x"d9",
          7064 => x"80",
          7065 => x"c0",
          7066 => x"8c",
          7067 => x"87",
          7068 => x"0c",
          7069 => x"b4",
          7070 => x"11",
          7071 => x"05",
          7072 => x"fd",
          7073 => x"f0",
          7074 => x"f0",
          7075 => x"52",
          7076 => x"51",
          7077 => x"3f",
          7078 => x"04",
          7079 => x"80",
          7080 => x"84",
          7081 => x"e0",
          7082 => x"fe",
          7083 => x"2e",
          7084 => x"63",
          7085 => x"a0",
          7086 => x"d0",
          7087 => x"78",
          7088 => x"f0",
          7089 => x"f0",
          7090 => x"fe",
          7091 => x"81",
          7092 => x"fe",
          7093 => x"f0",
          7094 => x"f8",
          7095 => x"d8",
          7096 => x"b5",
          7097 => x"9b",
          7098 => x"f4",
          7099 => x"b8",
          7100 => x"ff",
          7101 => x"ce",
          7102 => x"87",
          7103 => x"79",
          7104 => x"80",
          7105 => x"38",
          7106 => x"59",
          7107 => x"81",
          7108 => x"3d",
          7109 => x"51",
          7110 => x"3f",
          7111 => x"08",
          7112 => x"7b",
          7113 => x"38",
          7114 => x"89",
          7115 => x"2e",
          7116 => x"cd",
          7117 => x"2e",
          7118 => x"c5",
          7119 => x"88",
          7120 => x"81",
          7121 => x"80",
          7122 => x"90",
          7123 => x"ff",
          7124 => x"fe",
          7125 => x"bb",
          7126 => x"b0",
          7127 => x"ff",
          7128 => x"fe",
          7129 => x"ab",
          7130 => x"81",
          7131 => x"80",
          7132 => x"a0",
          7133 => x"ff",
          7134 => x"fe",
          7135 => x"93",
          7136 => x"80",
          7137 => x"ac",
          7138 => x"ff",
          7139 => x"fe",
          7140 => x"81",
          7141 => x"81",
          7142 => x"80",
          7143 => x"80",
          7144 => x"80",
          7145 => x"80",
          7146 => x"ff",
          7147 => x"e6",
          7148 => x"fe",
          7149 => x"fe",
          7150 => x"70",
          7151 => x"07",
          7152 => x"5b",
          7153 => x"5a",
          7154 => x"83",
          7155 => x"78",
          7156 => x"78",
          7157 => x"38",
          7158 => x"81",
          7159 => x"59",
          7160 => x"38",
          7161 => x"7d",
          7162 => x"59",
          7163 => x"7e",
          7164 => x"81",
          7165 => x"38",
          7166 => x"51",
          7167 => x"3f",
          7168 => x"fc",
          7169 => x"0b",
          7170 => x"34",
          7171 => x"8c",
          7172 => x"55",
          7173 => x"52",
          7174 => x"b3",
          7175 => x"fe",
          7176 => x"2b",
          7177 => x"53",
          7178 => x"52",
          7179 => x"b2",
          7180 => x"81",
          7181 => x"07",
          7182 => x"c0",
          7183 => x"08",
          7184 => x"84",
          7185 => x"51",
          7186 => x"3f",
          7187 => x"08",
          7188 => x"08",
          7189 => x"84",
          7190 => x"51",
          7191 => x"3f",
          7192 => x"f0",
          7193 => x"0c",
          7194 => x"0b",
          7195 => x"84",
          7196 => x"83",
          7197 => x"94",
          7198 => x"8b",
          7199 => x"84",
          7200 => x"0b",
          7201 => x"0c",
          7202 => x"3f",
          7203 => x"3f",
          7204 => x"51",
          7205 => x"3f",
          7206 => x"51",
          7207 => x"3f",
          7208 => x"51",
          7209 => x"3f",
          7210 => x"fc",
          7211 => x"3f",
          7212 => x"00",
          7213 => x"ff",
          7214 => x"ff",
          7215 => x"ff",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"25",
          7254 => x"64",
          7255 => x"20",
          7256 => x"25",
          7257 => x"64",
          7258 => x"25",
          7259 => x"53",
          7260 => x"43",
          7261 => x"69",
          7262 => x"61",
          7263 => x"6e",
          7264 => x"20",
          7265 => x"6f",
          7266 => x"6f",
          7267 => x"6f",
          7268 => x"67",
          7269 => x"3a",
          7270 => x"76",
          7271 => x"73",
          7272 => x"70",
          7273 => x"65",
          7274 => x"64",
          7275 => x"20",
          7276 => x"57",
          7277 => x"44",
          7278 => x"20",
          7279 => x"30",
          7280 => x"25",
          7281 => x"29",
          7282 => x"20",
          7283 => x"53",
          7284 => x"4d",
          7285 => x"20",
          7286 => x"30",
          7287 => x"25",
          7288 => x"29",
          7289 => x"20",
          7290 => x"49",
          7291 => x"20",
          7292 => x"4d",
          7293 => x"30",
          7294 => x"25",
          7295 => x"29",
          7296 => x"20",
          7297 => x"42",
          7298 => x"20",
          7299 => x"20",
          7300 => x"30",
          7301 => x"25",
          7302 => x"29",
          7303 => x"20",
          7304 => x"52",
          7305 => x"20",
          7306 => x"20",
          7307 => x"30",
          7308 => x"25",
          7309 => x"29",
          7310 => x"20",
          7311 => x"53",
          7312 => x"41",
          7313 => x"20",
          7314 => x"65",
          7315 => x"65",
          7316 => x"25",
          7317 => x"29",
          7318 => x"20",
          7319 => x"54",
          7320 => x"52",
          7321 => x"20",
          7322 => x"69",
          7323 => x"73",
          7324 => x"25",
          7325 => x"29",
          7326 => x"20",
          7327 => x"49",
          7328 => x"20",
          7329 => x"4c",
          7330 => x"68",
          7331 => x"65",
          7332 => x"25",
          7333 => x"29",
          7334 => x"20",
          7335 => x"57",
          7336 => x"42",
          7337 => x"20",
          7338 => x"0a",
          7339 => x"20",
          7340 => x"57",
          7341 => x"32",
          7342 => x"20",
          7343 => x"49",
          7344 => x"4c",
          7345 => x"20",
          7346 => x"50",
          7347 => x"00",
          7348 => x"20",
          7349 => x"53",
          7350 => x"00",
          7351 => x"41",
          7352 => x"65",
          7353 => x"73",
          7354 => x"20",
          7355 => x"43",
          7356 => x"52",
          7357 => x"74",
          7358 => x"63",
          7359 => x"20",
          7360 => x"72",
          7361 => x"20",
          7362 => x"30",
          7363 => x"00",
          7364 => x"20",
          7365 => x"43",
          7366 => x"4d",
          7367 => x"72",
          7368 => x"74",
          7369 => x"20",
          7370 => x"72",
          7371 => x"20",
          7372 => x"30",
          7373 => x"00",
          7374 => x"20",
          7375 => x"53",
          7376 => x"6b",
          7377 => x"61",
          7378 => x"41",
          7379 => x"65",
          7380 => x"20",
          7381 => x"20",
          7382 => x"30",
          7383 => x"00",
          7384 => x"4d",
          7385 => x"3a",
          7386 => x"20",
          7387 => x"5a",
          7388 => x"49",
          7389 => x"20",
          7390 => x"20",
          7391 => x"20",
          7392 => x"20",
          7393 => x"20",
          7394 => x"30",
          7395 => x"00",
          7396 => x"20",
          7397 => x"53",
          7398 => x"65",
          7399 => x"6c",
          7400 => x"20",
          7401 => x"71",
          7402 => x"20",
          7403 => x"20",
          7404 => x"64",
          7405 => x"34",
          7406 => x"7a",
          7407 => x"20",
          7408 => x"53",
          7409 => x"4d",
          7410 => x"6f",
          7411 => x"46",
          7412 => x"20",
          7413 => x"20",
          7414 => x"20",
          7415 => x"64",
          7416 => x"34",
          7417 => x"7a",
          7418 => x"20",
          7419 => x"57",
          7420 => x"62",
          7421 => x"20",
          7422 => x"41",
          7423 => x"6c",
          7424 => x"20",
          7425 => x"71",
          7426 => x"64",
          7427 => x"34",
          7428 => x"7a",
          7429 => x"53",
          7430 => x"6c",
          7431 => x"4d",
          7432 => x"75",
          7433 => x"46",
          7434 => x"00",
          7435 => x"45",
          7436 => x"45",
          7437 => x"69",
          7438 => x"55",
          7439 => x"6f",
          7440 => x"68",
          7441 => x"6f",
          7442 => x"74",
          7443 => x"68",
          7444 => x"6f",
          7445 => x"68",
          7446 => x"00",
          7447 => x"21",
          7448 => x"25",
          7449 => x"20",
          7450 => x"0a",
          7451 => x"46",
          7452 => x"65",
          7453 => x"6f",
          7454 => x"73",
          7455 => x"74",
          7456 => x"68",
          7457 => x"6f",
          7458 => x"66",
          7459 => x"20",
          7460 => x"45",
          7461 => x"0a",
          7462 => x"43",
          7463 => x"6f",
          7464 => x"70",
          7465 => x"63",
          7466 => x"74",
          7467 => x"69",
          7468 => x"72",
          7469 => x"69",
          7470 => x"20",
          7471 => x"61",
          7472 => x"6e",
          7473 => x"00",
          7474 => x"00",
          7475 => x"01",
          7476 => x"00",
          7477 => x"00",
          7478 => x"01",
          7479 => x"00",
          7480 => x"00",
          7481 => x"04",
          7482 => x"00",
          7483 => x"00",
          7484 => x"04",
          7485 => x"00",
          7486 => x"00",
          7487 => x"04",
          7488 => x"00",
          7489 => x"00",
          7490 => x"04",
          7491 => x"00",
          7492 => x"00",
          7493 => x"04",
          7494 => x"00",
          7495 => x"00",
          7496 => x"03",
          7497 => x"00",
          7498 => x"00",
          7499 => x"03",
          7500 => x"00",
          7501 => x"00",
          7502 => x"03",
          7503 => x"00",
          7504 => x"00",
          7505 => x"03",
          7506 => x"00",
          7507 => x"1b",
          7508 => x"1b",
          7509 => x"1b",
          7510 => x"1b",
          7511 => x"1b",
          7512 => x"1b",
          7513 => x"1b",
          7514 => x"1b",
          7515 => x"1b",
          7516 => x"0d",
          7517 => x"08",
          7518 => x"53",
          7519 => x"22",
          7520 => x"3a",
          7521 => x"3e",
          7522 => x"7c",
          7523 => x"46",
          7524 => x"46",
          7525 => x"32",
          7526 => x"eb",
          7527 => x"53",
          7528 => x"35",
          7529 => x"4e",
          7530 => x"41",
          7531 => x"20",
          7532 => x"41",
          7533 => x"20",
          7534 => x"4e",
          7535 => x"41",
          7536 => x"20",
          7537 => x"41",
          7538 => x"20",
          7539 => x"00",
          7540 => x"00",
          7541 => x"00",
          7542 => x"00",
          7543 => x"80",
          7544 => x"8e",
          7545 => x"45",
          7546 => x"49",
          7547 => x"90",
          7548 => x"99",
          7549 => x"59",
          7550 => x"9c",
          7551 => x"41",
          7552 => x"a5",
          7553 => x"a8",
          7554 => x"ac",
          7555 => x"b0",
          7556 => x"b4",
          7557 => x"b8",
          7558 => x"bc",
          7559 => x"c0",
          7560 => x"c4",
          7561 => x"c8",
          7562 => x"cc",
          7563 => x"d0",
          7564 => x"d4",
          7565 => x"d8",
          7566 => x"dc",
          7567 => x"e0",
          7568 => x"e4",
          7569 => x"e8",
          7570 => x"ec",
          7571 => x"f0",
          7572 => x"f4",
          7573 => x"f8",
          7574 => x"fc",
          7575 => x"2b",
          7576 => x"3d",
          7577 => x"5c",
          7578 => x"3c",
          7579 => x"7f",
          7580 => x"00",
          7581 => x"00",
          7582 => x"01",
          7583 => x"00",
          7584 => x"00",
          7585 => x"00",
          7586 => x"00",
          7587 => x"00",
          7588 => x"64",
          7589 => x"74",
          7590 => x"64",
          7591 => x"74",
          7592 => x"66",
          7593 => x"74",
          7594 => x"66",
          7595 => x"64",
          7596 => x"66",
          7597 => x"63",
          7598 => x"6d",
          7599 => x"61",
          7600 => x"6d",
          7601 => x"79",
          7602 => x"6d",
          7603 => x"66",
          7604 => x"6d",
          7605 => x"70",
          7606 => x"6d",
          7607 => x"6d",
          7608 => x"6d",
          7609 => x"68",
          7610 => x"68",
          7611 => x"68",
          7612 => x"68",
          7613 => x"63",
          7614 => x"00",
          7615 => x"6a",
          7616 => x"72",
          7617 => x"61",
          7618 => x"72",
          7619 => x"74",
          7620 => x"69",
          7621 => x"00",
          7622 => x"74",
          7623 => x"00",
          7624 => x"74",
          7625 => x"69",
          7626 => x"6d",
          7627 => x"69",
          7628 => x"6b",
          7629 => x"00",
          7630 => x"44",
          7631 => x"20",
          7632 => x"6f",
          7633 => x"49",
          7634 => x"72",
          7635 => x"20",
          7636 => x"6f",
          7637 => x"00",
          7638 => x"44",
          7639 => x"20",
          7640 => x"20",
          7641 => x"64",
          7642 => x"00",
          7643 => x"4e",
          7644 => x"69",
          7645 => x"66",
          7646 => x"64",
          7647 => x"4e",
          7648 => x"61",
          7649 => x"66",
          7650 => x"64",
          7651 => x"49",
          7652 => x"6c",
          7653 => x"66",
          7654 => x"6e",
          7655 => x"2e",
          7656 => x"41",
          7657 => x"73",
          7658 => x"65",
          7659 => x"64",
          7660 => x"46",
          7661 => x"20",
          7662 => x"65",
          7663 => x"20",
          7664 => x"73",
          7665 => x"0a",
          7666 => x"46",
          7667 => x"20",
          7668 => x"64",
          7669 => x"69",
          7670 => x"6c",
          7671 => x"0a",
          7672 => x"53",
          7673 => x"73",
          7674 => x"69",
          7675 => x"70",
          7676 => x"65",
          7677 => x"64",
          7678 => x"44",
          7679 => x"65",
          7680 => x"6d",
          7681 => x"20",
          7682 => x"69",
          7683 => x"6c",
          7684 => x"0a",
          7685 => x"44",
          7686 => x"20",
          7687 => x"20",
          7688 => x"62",
          7689 => x"2e",
          7690 => x"4e",
          7691 => x"6f",
          7692 => x"74",
          7693 => x"65",
          7694 => x"6c",
          7695 => x"73",
          7696 => x"20",
          7697 => x"6e",
          7698 => x"6e",
          7699 => x"73",
          7700 => x"00",
          7701 => x"46",
          7702 => x"61",
          7703 => x"62",
          7704 => x"65",
          7705 => x"00",
          7706 => x"54",
          7707 => x"6f",
          7708 => x"20",
          7709 => x"72",
          7710 => x"6f",
          7711 => x"61",
          7712 => x"6c",
          7713 => x"2e",
          7714 => x"46",
          7715 => x"20",
          7716 => x"6c",
          7717 => x"65",
          7718 => x"00",
          7719 => x"49",
          7720 => x"66",
          7721 => x"69",
          7722 => x"20",
          7723 => x"6f",
          7724 => x"0a",
          7725 => x"54",
          7726 => x"6d",
          7727 => x"20",
          7728 => x"6e",
          7729 => x"6c",
          7730 => x"0a",
          7731 => x"50",
          7732 => x"6d",
          7733 => x"72",
          7734 => x"6e",
          7735 => x"72",
          7736 => x"2e",
          7737 => x"53",
          7738 => x"65",
          7739 => x"0a",
          7740 => x"55",
          7741 => x"6f",
          7742 => x"65",
          7743 => x"72",
          7744 => x"0a",
          7745 => x"20",
          7746 => x"65",
          7747 => x"73",
          7748 => x"20",
          7749 => x"20",
          7750 => x"65",
          7751 => x"65",
          7752 => x"00",
          7753 => x"72",
          7754 => x"00",
          7755 => x"25",
          7756 => x"00",
          7757 => x"3a",
          7758 => x"25",
          7759 => x"00",
          7760 => x"20",
          7761 => x"20",
          7762 => x"00",
          7763 => x"25",
          7764 => x"00",
          7765 => x"20",
          7766 => x"20",
          7767 => x"7c",
          7768 => x"5a",
          7769 => x"41",
          7770 => x"0a",
          7771 => x"25",
          7772 => x"00",
          7773 => x"32",
          7774 => x"34",
          7775 => x"32",
          7776 => x"76",
          7777 => x"31",
          7778 => x"20",
          7779 => x"2c",
          7780 => x"76",
          7781 => x"32",
          7782 => x"25",
          7783 => x"73",
          7784 => x"0a",
          7785 => x"5a",
          7786 => x"41",
          7787 => x"74",
          7788 => x"75",
          7789 => x"48",
          7790 => x"6c",
          7791 => x"00",
          7792 => x"54",
          7793 => x"72",
          7794 => x"74",
          7795 => x"75",
          7796 => x"00",
          7797 => x"50",
          7798 => x"69",
          7799 => x"72",
          7800 => x"74",
          7801 => x"49",
          7802 => x"4c",
          7803 => x"20",
          7804 => x"65",
          7805 => x"70",
          7806 => x"49",
          7807 => x"4c",
          7808 => x"20",
          7809 => x"65",
          7810 => x"70",
          7811 => x"55",
          7812 => x"30",
          7813 => x"20",
          7814 => x"65",
          7815 => x"70",
          7816 => x"55",
          7817 => x"30",
          7818 => x"20",
          7819 => x"65",
          7820 => x"70",
          7821 => x"55",
          7822 => x"31",
          7823 => x"20",
          7824 => x"65",
          7825 => x"70",
          7826 => x"55",
          7827 => x"31",
          7828 => x"20",
          7829 => x"65",
          7830 => x"70",
          7831 => x"53",
          7832 => x"69",
          7833 => x"75",
          7834 => x"69",
          7835 => x"2e",
          7836 => x"00",
          7837 => x"45",
          7838 => x"6c",
          7839 => x"20",
          7840 => x"65",
          7841 => x"2e",
          7842 => x"61",
          7843 => x"65",
          7844 => x"2e",
          7845 => x"00",
          7846 => x"30",
          7847 => x"46",
          7848 => x"65",
          7849 => x"6f",
          7850 => x"69",
          7851 => x"6c",
          7852 => x"20",
          7853 => x"63",
          7854 => x"20",
          7855 => x"70",
          7856 => x"73",
          7857 => x"6e",
          7858 => x"6d",
          7859 => x"61",
          7860 => x"2e",
          7861 => x"2a",
          7862 => x"42",
          7863 => x"64",
          7864 => x"20",
          7865 => x"0a",
          7866 => x"49",
          7867 => x"69",
          7868 => x"73",
          7869 => x"0a",
          7870 => x"46",
          7871 => x"65",
          7872 => x"6f",
          7873 => x"69",
          7874 => x"6c",
          7875 => x"2e",
          7876 => x"72",
          7877 => x"64",
          7878 => x"25",
          7879 => x"43",
          7880 => x"72",
          7881 => x"2e",
          7882 => x"00",
          7883 => x"43",
          7884 => x"69",
          7885 => x"2e",
          7886 => x"43",
          7887 => x"61",
          7888 => x"67",
          7889 => x"00",
          7890 => x"25",
          7891 => x"78",
          7892 => x"38",
          7893 => x"3e",
          7894 => x"6c",
          7895 => x"30",
          7896 => x"0a",
          7897 => x"44",
          7898 => x"20",
          7899 => x"6f",
          7900 => x"00",
          7901 => x"0a",
          7902 => x"70",
          7903 => x"65",
          7904 => x"25",
          7905 => x"20",
          7906 => x"58",
          7907 => x"3f",
          7908 => x"00",
          7909 => x"25",
          7910 => x"20",
          7911 => x"58",
          7912 => x"25",
          7913 => x"20",
          7914 => x"58",
          7915 => x"44",
          7916 => x"62",
          7917 => x"67",
          7918 => x"74",
          7919 => x"75",
          7920 => x"0a",
          7921 => x"45",
          7922 => x"6c",
          7923 => x"20",
          7924 => x"65",
          7925 => x"70",
          7926 => x"00",
          7927 => x"44",
          7928 => x"62",
          7929 => x"20",
          7930 => x"74",
          7931 => x"66",
          7932 => x"45",
          7933 => x"6c",
          7934 => x"20",
          7935 => x"74",
          7936 => x"66",
          7937 => x"45",
          7938 => x"75",
          7939 => x"67",
          7940 => x"64",
          7941 => x"20",
          7942 => x"78",
          7943 => x"2e",
          7944 => x"43",
          7945 => x"69",
          7946 => x"63",
          7947 => x"20",
          7948 => x"30",
          7949 => x"2e",
          7950 => x"00",
          7951 => x"43",
          7952 => x"20",
          7953 => x"75",
          7954 => x"64",
          7955 => x"64",
          7956 => x"25",
          7957 => x"0a",
          7958 => x"52",
          7959 => x"61",
          7960 => x"6e",
          7961 => x"70",
          7962 => x"63",
          7963 => x"6f",
          7964 => x"2e",
          7965 => x"43",
          7966 => x"20",
          7967 => x"6f",
          7968 => x"6e",
          7969 => x"2e",
          7970 => x"5a",
          7971 => x"62",
          7972 => x"25",
          7973 => x"25",
          7974 => x"73",
          7975 => x"00",
          7976 => x"25",
          7977 => x"25",
          7978 => x"73",
          7979 => x"25",
          7980 => x"25",
          7981 => x"42",
          7982 => x"63",
          7983 => x"61",
          7984 => x"0a",
          7985 => x"52",
          7986 => x"69",
          7987 => x"2e",
          7988 => x"45",
          7989 => x"6c",
          7990 => x"20",
          7991 => x"65",
          7992 => x"70",
          7993 => x"2e",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"00",
          8000 => x"00",
          8001 => x"00",
          8002 => x"00",
          8003 => x"01",
          8004 => x"01",
          8005 => x"00",
          8006 => x"00",
          8007 => x"00",
          8008 => x"00",
          8009 => x"05",
          8010 => x"05",
          8011 => x"05",
          8012 => x"00",
          8013 => x"01",
          8014 => x"01",
          8015 => x"01",
          8016 => x"01",
          8017 => x"00",
          8018 => x"00",
          8019 => x"00",
          8020 => x"00",
          8021 => x"00",
          8022 => x"00",
          8023 => x"00",
          8024 => x"00",
          8025 => x"00",
          8026 => x"00",
          8027 => x"00",
          8028 => x"00",
          8029 => x"00",
          8030 => x"00",
          8031 => x"00",
          8032 => x"00",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"01",
          8050 => x"00",
          8051 => x"01",
          8052 => x"00",
          8053 => x"02",
          8054 => x"01",
          8055 => x"00",
          8056 => x"00",
          8057 => x"01",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"01",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"01",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"01",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"01",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"01",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"01",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"01",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"01",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"01",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"01",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"01",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"01",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"01",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"01",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"01",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"01",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"01",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"01",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"01",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"01",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"01",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"01",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"01",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"01",
          8154 => x"00",
          8155 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
