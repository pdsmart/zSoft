-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b83ff",
             1 => x"f80d0b0b",
             2 => x"0b93b904",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"9d040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b9380",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b82ac",
           162 => x"cc738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93850400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b80c5",
           171 => x"9f2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b80c7",
           179 => x"8b2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"95040b0b",
           269 => x"0b8ca404",
           270 => x"0b0b0b8c",
           271 => x"b3040b0b",
           272 => x"0b8cc204",
           273 => x"0b0b0b8c",
           274 => x"d1040b0b",
           275 => x"0b8ce004",
           276 => x"0b0b0b8c",
           277 => x"f0040b0b",
           278 => x"0b8d8004",
           279 => x"0b0b0b8d",
           280 => x"8f040b0b",
           281 => x"0b8d9e04",
           282 => x"0b0b0b8d",
           283 => x"ad040b0b",
           284 => x"0b8dbd04",
           285 => x"0b0b0b8d",
           286 => x"cd040b0b",
           287 => x"0b8ddd04",
           288 => x"0b0b0b8d",
           289 => x"ed040b0b",
           290 => x"0b8dfd04",
           291 => x"0b0b0b8e",
           292 => x"8d040b0b",
           293 => x"0b8e9d04",
           294 => x"0b0b0b8e",
           295 => x"ad040b0b",
           296 => x"0b8ebd04",
           297 => x"0b0b0b8e",
           298 => x"cd040b0b",
           299 => x"0b8edd04",
           300 => x"0b0b0b8e",
           301 => x"ed040b0b",
           302 => x"0b8efd04",
           303 => x"0b0b0b8f",
           304 => x"8d040b0b",
           305 => x"0b8f9d04",
           306 => x"0b0b0b8f",
           307 => x"ad040b0b",
           308 => x"0b8fbd04",
           309 => x"0b0b0b8f",
           310 => x"cd040b0b",
           311 => x"0b8fdd04",
           312 => x"0b0b0b8f",
           313 => x"ed040b0b",
           314 => x"0b8ffd04",
           315 => x"0b0b0b90",
           316 => x"8d040b0b",
           317 => x"0b909d04",
           318 => x"0b0b0b90",
           319 => x"ad040b0b",
           320 => x"0b90bd04",
           321 => x"0b0b0b90",
           322 => x"cd040b0b",
           323 => x"0b90dd04",
           324 => x"0b0b0b90",
           325 => x"ed040b0b",
           326 => x"0b90fd04",
           327 => x"0b0b0b91",
           328 => x"8d040b0b",
           329 => x"0b919d04",
           330 => x"0b0b0b91",
           331 => x"ad040b0b",
           332 => x"0b91bd04",
           333 => x"0b0b0b91",
           334 => x"cd040b0b",
           335 => x"0b91dd04",
           336 => x"0b0b0b91",
           337 => x"ed040b0b",
           338 => x"0b91fd04",
           339 => x"0b0b0b92",
           340 => x"8d040b0b",
           341 => x"0b929d04",
           342 => x"0b0b0b92",
           343 => x"ad040b0b",
           344 => x"0b92bd04",
           345 => x"0b0b0b92",
           346 => x"cd04ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0482d6e4",
           386 => x"0c80f7d4",
           387 => x"2d82d6e4",
           388 => x"08848090",
           389 => x"0482d6e4",
           390 => x"0cb3b22d",
           391 => x"82d6e408",
           392 => x"84809004",
           393 => x"82d6e40c",
           394 => x"afe32d82",
           395 => x"d6e40884",
           396 => x"80900482",
           397 => x"d6e40caf",
           398 => x"ad2d82d6",
           399 => x"e4088480",
           400 => x"900482d6",
           401 => x"e40c94ad",
           402 => x"2d82d6e4",
           403 => x"08848090",
           404 => x"0482d6e4",
           405 => x"0cb1c22d",
           406 => x"82d6e408",
           407 => x"84809004",
           408 => x"82d6e40c",
           409 => x"80d0f72d",
           410 => x"82d6e408",
           411 => x"84809004",
           412 => x"82d6e40c",
           413 => x"80cba62d",
           414 => x"82d6e408",
           415 => x"84809004",
           416 => x"82d6e40c",
           417 => x"93d82d82",
           418 => x"d6e40884",
           419 => x"80900482",
           420 => x"d6e40c96",
           421 => x"c02d82d6",
           422 => x"e4088480",
           423 => x"900482d6",
           424 => x"e40c97cd",
           425 => x"2d82d6e4",
           426 => x"08848090",
           427 => x"0482d6e4",
           428 => x"0c80f9fa",
           429 => x"2d82d6e4",
           430 => x"08848090",
           431 => x"0482d6e4",
           432 => x"0c80fac9",
           433 => x"2d82d6e4",
           434 => x"08848090",
           435 => x"0482d6e4",
           436 => x"0c80f399",
           437 => x"2d82d6e4",
           438 => x"08848090",
           439 => x"0482d6e4",
           440 => x"0c80f590",
           441 => x"2d82d6e4",
           442 => x"08848090",
           443 => x"0482d6e4",
           444 => x"0c80f6c3",
           445 => x"2d82d6e4",
           446 => x"08848090",
           447 => x"0482d6e4",
           448 => x"0c81ecad",
           449 => x"2d82d6e4",
           450 => x"08848090",
           451 => x"0482d6e4",
           452 => x"0c81f9ac",
           453 => x"2d82d6e4",
           454 => x"08848090",
           455 => x"0482d6e4",
           456 => x"0c81f192",
           457 => x"2d82d6e4",
           458 => x"08848090",
           459 => x"0482d6e4",
           460 => x"0c81f492",
           461 => x"2d82d6e4",
           462 => x"08848090",
           463 => x"0482d6e4",
           464 => x"0c81feea",
           465 => x"2d82d6e4",
           466 => x"08848090",
           467 => x"0482d6e4",
           468 => x"0c8287d3",
           469 => x"2d82d6e4",
           470 => x"08848090",
           471 => x"0482d6e4",
           472 => x"0c81f889",
           473 => x"2d82d6e4",
           474 => x"08848090",
           475 => x"0482d6e4",
           476 => x"0c82828d",
           477 => x"2d82d6e4",
           478 => x"08848090",
           479 => x"0482d6e4",
           480 => x"0c8283ad",
           481 => x"2d82d6e4",
           482 => x"08848090",
           483 => x"0482d6e4",
           484 => x"0c8283cc",
           485 => x"2d82d6e4",
           486 => x"08848090",
           487 => x"0482d6e4",
           488 => x"0c828bc0",
           489 => x"2d82d6e4",
           490 => x"08848090",
           491 => x"0482d6e4",
           492 => x"0c8289a2",
           493 => x"2d82d6e4",
           494 => x"08848090",
           495 => x"0482d6e4",
           496 => x"0c828e9c",
           497 => x"2d82d6e4",
           498 => x"08848090",
           499 => x"0482d6e4",
           500 => x"0c8284d2",
           501 => x"2d82d6e4",
           502 => x"08848090",
           503 => x"0482d6e4",
           504 => x"0c8291a1",
           505 => x"2d82d6e4",
           506 => x"08848090",
           507 => x"0482d6e4",
           508 => x"0c8292a2",
           509 => x"2d82d6e4",
           510 => x"08848090",
           511 => x"0482d6e4",
           512 => x"0c81fa8c",
           513 => x"2d82d6e4",
           514 => x"08848090",
           515 => x"0482d6e4",
           516 => x"0c81f9e5",
           517 => x"2d82d6e4",
           518 => x"08848090",
           519 => x"0482d6e4",
           520 => x"0c81fb90",
           521 => x"2d82d6e4",
           522 => x"08848090",
           523 => x"0482d6e4",
           524 => x"0c8285a9",
           525 => x"2d82d6e4",
           526 => x"08848090",
           527 => x"0482d6e4",
           528 => x"0c829393",
           529 => x"2d82d6e4",
           530 => x"08848090",
           531 => x"0482d6e4",
           532 => x"0c82959e",
           533 => x"2d82d6e4",
           534 => x"08848090",
           535 => x"0482d6e4",
           536 => x"0c8298a5",
           537 => x"2d82d6e4",
           538 => x"08848090",
           539 => x"0482d6e4",
           540 => x"0c81ebcc",
           541 => x"2d82d6e4",
           542 => x"08848090",
           543 => x"0482d6e4",
           544 => x"0c829b91",
           545 => x"2d82d6e4",
           546 => x"08848090",
           547 => x"0482d6e4",
           548 => x"0c82a9c6",
           549 => x"2d82d6e4",
           550 => x"08848090",
           551 => x"0482d6e4",
           552 => x"0c82a7b2",
           553 => x"2d82d6e4",
           554 => x"08848090",
           555 => x"0482d6e4",
           556 => x"0c81abd4",
           557 => x"2d82d6e4",
           558 => x"08848090",
           559 => x"0482d6e4",
           560 => x"0c81adbe",
           561 => x"2d82d6e4",
           562 => x"08848090",
           563 => x"0482d6e4",
           564 => x"0c81afa2",
           565 => x"2d82d6e4",
           566 => x"08848090",
           567 => x"0482d6e4",
           568 => x"0c80f3c2",
           569 => x"2d82d6e4",
           570 => x"08848090",
           571 => x"0482d6e4",
           572 => x"0c80f4e6",
           573 => x"2d82d6e4",
           574 => x"08848090",
           575 => x"0482d6e4",
           576 => x"0c80f8c9",
           577 => x"2d82d6e4",
           578 => x"08848090",
           579 => x"0482d6e4",
           580 => x"0c80d7bf",
           581 => x"2d82d6e4",
           582 => x"08848090",
           583 => x"0482d6e4",
           584 => x"0c81a5e8",
           585 => x"2d82d6e4",
           586 => x"08848090",
           587 => x"0482d6e4",
           588 => x"0c81a690",
           589 => x"2d82d6e4",
           590 => x"08848090",
           591 => x"0482d6e4",
           592 => x"0c81aa88",
           593 => x"2d82d6e4",
           594 => x"08848090",
           595 => x"0482d6e4",
           596 => x"0c81a2d2",
           597 => x"2d82d6e4",
           598 => x"08848090",
           599 => x"043c0400",
           600 => x"00101010",
           601 => x"10101010",
           602 => x"10101010",
           603 => x"10101010",
           604 => x"10101010",
           605 => x"10101010",
           606 => x"10101010",
           607 => x"10101010",
           608 => x"53510400",
           609 => x"007381ff",
           610 => x"06738306",
           611 => x"09810583",
           612 => x"05101010",
           613 => x"2b0772fc",
           614 => x"060c5151",
           615 => x"04727280",
           616 => x"728106ff",
           617 => x"05097206",
           618 => x"05711052",
           619 => x"720a100a",
           620 => x"5372ed38",
           621 => x"51515351",
           622 => x"0482d6d8",
           623 => x"7082f2c4",
           624 => x"278e3880",
           625 => x"71708405",
           626 => x"530c0b0b",
           627 => x"0b93bc04",
           628 => x"8c815180",
           629 => x"f0ec0400",
           630 => x"82d6e408",
           631 => x"0282d6e4",
           632 => x"0cfb3d0d",
           633 => x"82d6e408",
           634 => x"8c057082",
           635 => x"d6e408fc",
           636 => x"050c82d6",
           637 => x"e408fc05",
           638 => x"085482d6",
           639 => x"e4088805",
           640 => x"085382f2",
           641 => x"bc085254",
           642 => x"849a3f82",
           643 => x"d6d80870",
           644 => x"82d6e408",
           645 => x"f8050c82",
           646 => x"d6e408f8",
           647 => x"05087082",
           648 => x"d6d80c51",
           649 => x"54873d0d",
           650 => x"82d6e40c",
           651 => x"0482d6e4",
           652 => x"080282d6",
           653 => x"e40cfb3d",
           654 => x"0d82d6e4",
           655 => x"08900508",
           656 => x"85113370",
           657 => x"81327081",
           658 => x"06515151",
           659 => x"52718f38",
           660 => x"800b82d6",
           661 => x"e4088c05",
           662 => x"08258338",
           663 => x"8d39800b",
           664 => x"82d6e408",
           665 => x"f4050c81",
           666 => x"c43982d6",
           667 => x"e4088c05",
           668 => x"08ff0582",
           669 => x"d6e4088c",
           670 => x"050c800b",
           671 => x"82d6e408",
           672 => x"f8050c82",
           673 => x"d6e40888",
           674 => x"050882d6",
           675 => x"e408fc05",
           676 => x"0c82d6e4",
           677 => x"08f80508",
           678 => x"8a2e80f6",
           679 => x"38800b82",
           680 => x"d6e4088c",
           681 => x"05082580",
           682 => x"e93882d6",
           683 => x"e4089005",
           684 => x"0851a090",
           685 => x"3f82d6d8",
           686 => x"087082d6",
           687 => x"e408f805",
           688 => x"0c5282d6",
           689 => x"e408f805",
           690 => x"08ff2e09",
           691 => x"81068d38",
           692 => x"800b82d6",
           693 => x"e408f405",
           694 => x"0c80d239",
           695 => x"82d6e408",
           696 => x"fc050882",
           697 => x"d6e408f8",
           698 => x"05085353",
           699 => x"71733482",
           700 => x"d6e4088c",
           701 => x"0508ff05",
           702 => x"82d6e408",
           703 => x"8c050c82",
           704 => x"d6e408fc",
           705 => x"05088105",
           706 => x"82d6e408",
           707 => x"fc050cff",
           708 => x"803982d6",
           709 => x"e408fc05",
           710 => x"08528072",
           711 => x"3482d6e4",
           712 => x"08880508",
           713 => x"7082d6e4",
           714 => x"08f4050c",
           715 => x"5282d6e4",
           716 => x"08f40508",
           717 => x"82d6d80c",
           718 => x"873d0d82",
           719 => x"d6e40c04",
           720 => x"82d6e408",
           721 => x"0282d6e4",
           722 => x"0cf43d0d",
           723 => x"860b82d6",
           724 => x"e408e505",
           725 => x"3482d6e4",
           726 => x"08880508",
           727 => x"82d6e408",
           728 => x"e0050cfe",
           729 => x"0a0b82d6",
           730 => x"e408e805",
           731 => x"0c82d6e4",
           732 => x"08900570",
           733 => x"82d6e408",
           734 => x"fc050c82",
           735 => x"d6e408fc",
           736 => x"05085482",
           737 => x"d6e4088c",
           738 => x"05085382",
           739 => x"d6e408e0",
           740 => x"05705351",
           741 => x"54818d3f",
           742 => x"82d6d808",
           743 => x"7082d6e4",
           744 => x"08dc050c",
           745 => x"82d6e408",
           746 => x"ec050882",
           747 => x"d6e40888",
           748 => x"05080551",
           749 => x"54807434",
           750 => x"82d6e408",
           751 => x"dc050870",
           752 => x"82d6d80c",
           753 => x"548e3d0d",
           754 => x"82d6e40c",
           755 => x"0482d6e4",
           756 => x"080282d6",
           757 => x"e40cfb3d",
           758 => x"0d82d6e4",
           759 => x"08900570",
           760 => x"82d6e408",
           761 => x"fc050c82",
           762 => x"d6e408fc",
           763 => x"05085482",
           764 => x"d6e4088c",
           765 => x"05085382",
           766 => x"d6e40888",
           767 => x"05085254",
           768 => x"a33f82d6",
           769 => x"d8087082",
           770 => x"d6e408f8",
           771 => x"050c82d6",
           772 => x"e408f805",
           773 => x"087082d6",
           774 => x"d80c5154",
           775 => x"873d0d82",
           776 => x"d6e40c04",
           777 => x"82d6e408",
           778 => x"0282d6e4",
           779 => x"0ced3d0d",
           780 => x"800b82d6",
           781 => x"e408e405",
           782 => x"2382d6e4",
           783 => x"08880508",
           784 => x"53800b8c",
           785 => x"140c82d6",
           786 => x"e4088805",
           787 => x"08851133",
           788 => x"70812a70",
           789 => x"81327081",
           790 => x"06515151",
           791 => x"51537280",
           792 => x"2e8d38ff",
           793 => x"0b82d6e4",
           794 => x"08e0050c",
           795 => x"96ac3982",
           796 => x"d6e4088c",
           797 => x"05085372",
           798 => x"33537282",
           799 => x"d6e408f8",
           800 => x"05347281",
           801 => x"ff065372",
           802 => x"802e95fa",
           803 => x"3882d6e4",
           804 => x"088c0508",
           805 => x"810582d6",
           806 => x"e4088c05",
           807 => x"0c82d6e4",
           808 => x"08e40522",
           809 => x"70810651",
           810 => x"5372802e",
           811 => x"958b3882",
           812 => x"d6e408f8",
           813 => x"053353af",
           814 => x"732781fc",
           815 => x"3882d6e4",
           816 => x"08f80533",
           817 => x"5372b926",
           818 => x"81ee3882",
           819 => x"d6e408f8",
           820 => x"05335372",
           821 => x"b02e0981",
           822 => x"0680c538",
           823 => x"82d6e408",
           824 => x"e8053370",
           825 => x"982b7098",
           826 => x"2c515153",
           827 => x"72b23882",
           828 => x"d6e408e4",
           829 => x"05227083",
           830 => x"2a708132",
           831 => x"70810651",
           832 => x"51515372",
           833 => x"802e9938",
           834 => x"82d6e408",
           835 => x"e4052270",
           836 => x"82800751",
           837 => x"537282d6",
           838 => x"e408e405",
           839 => x"23fed039",
           840 => x"82d6e408",
           841 => x"e8053370",
           842 => x"982b7098",
           843 => x"2c707083",
           844 => x"2b721173",
           845 => x"11515151",
           846 => x"53515553",
           847 => x"7282d6e4",
           848 => x"08e80534",
           849 => x"82d6e408",
           850 => x"e8053354",
           851 => x"82d6e408",
           852 => x"f8053370",
           853 => x"15d01151",
           854 => x"51537282",
           855 => x"d6e408e8",
           856 => x"053482d6",
           857 => x"e408e805",
           858 => x"3370982b",
           859 => x"70982c51",
           860 => x"51537280",
           861 => x"258b3880",
           862 => x"ff0b82d6",
           863 => x"e408e805",
           864 => x"3482d6e4",
           865 => x"08e40522",
           866 => x"70832a70",
           867 => x"81065151",
           868 => x"5372fddb",
           869 => x"3882d6e4",
           870 => x"08e80533",
           871 => x"70882b70",
           872 => x"902b7090",
           873 => x"2c70882c",
           874 => x"51515151",
           875 => x"537282d6",
           876 => x"e408ec05",
           877 => x"23fdb839",
           878 => x"82d6e408",
           879 => x"e4052270",
           880 => x"832a7081",
           881 => x"06515153",
           882 => x"72802e9d",
           883 => x"3882d6e4",
           884 => x"08e80533",
           885 => x"70982b70",
           886 => x"982c5151",
           887 => x"53728a38",
           888 => x"810b82d6",
           889 => x"e408e805",
           890 => x"3482d6e4",
           891 => x"08f80533",
           892 => x"e01182d6",
           893 => x"e408c405",
           894 => x"0c5382d6",
           895 => x"e408c405",
           896 => x"0880d826",
           897 => x"92943882",
           898 => x"d6e408c4",
           899 => x"05087082",
           900 => x"2b82aebc",
           901 => x"11700851",
           902 => x"51515372",
           903 => x"0482d6e4",
           904 => x"08e40522",
           905 => x"70900751",
           906 => x"537282d6",
           907 => x"e408e405",
           908 => x"2382d6e4",
           909 => x"08e40522",
           910 => x"70a00751",
           911 => x"537282d6",
           912 => x"e408e405",
           913 => x"23fca839",
           914 => x"82d6e408",
           915 => x"e4052270",
           916 => x"81800751",
           917 => x"537282d6",
           918 => x"e408e405",
           919 => x"23fc9039",
           920 => x"82d6e408",
           921 => x"e4052270",
           922 => x"80c00751",
           923 => x"537282d6",
           924 => x"e408e405",
           925 => x"23fbf839",
           926 => x"82d6e408",
           927 => x"e4052270",
           928 => x"88075153",
           929 => x"7282d6e4",
           930 => x"08e40523",
           931 => x"800b82d6",
           932 => x"e408e805",
           933 => x"34fbd839",
           934 => x"82d6e408",
           935 => x"e4052270",
           936 => x"84075153",
           937 => x"7282d6e4",
           938 => x"08e40523",
           939 => x"fbc139bf",
           940 => x"0b82d6e4",
           941 => x"08fc0534",
           942 => x"82d6e408",
           943 => x"ec0522ff",
           944 => x"11515372",
           945 => x"82d6e408",
           946 => x"ec052380",
           947 => x"e30b82d6",
           948 => x"e408f805",
           949 => x"348da839",
           950 => x"82d6e408",
           951 => x"90050882",
           952 => x"d6e40890",
           953 => x"05088405",
           954 => x"82d6e408",
           955 => x"90050c70",
           956 => x"08515372",
           957 => x"82d6e408",
           958 => x"fc053482",
           959 => x"d6e408ec",
           960 => x"0522ff11",
           961 => x"51537282",
           962 => x"d6e408ec",
           963 => x"05238cef",
           964 => x"3982d6e4",
           965 => x"08900508",
           966 => x"82d6e408",
           967 => x"90050884",
           968 => x"0582d6e4",
           969 => x"0890050c",
           970 => x"700882d6",
           971 => x"e408fc05",
           972 => x"0c82d6e4",
           973 => x"08e40522",
           974 => x"70832a70",
           975 => x"81065151",
           976 => x"51537280",
           977 => x"2eab3882",
           978 => x"d6e408e8",
           979 => x"05337098",
           980 => x"2b537298",
           981 => x"2c5382d6",
           982 => x"e408fc05",
           983 => x"085253a4",
           984 => x"833f82d6",
           985 => x"d8085372",
           986 => x"82d6e408",
           987 => x"f4052399",
           988 => x"3982d6e4",
           989 => x"08fc0508",
           990 => x"519d8a3f",
           991 => x"82d6d808",
           992 => x"537282d6",
           993 => x"e408f405",
           994 => x"2382d6e4",
           995 => x"08ec0522",
           996 => x"5382d6e4",
           997 => x"08f40522",
           998 => x"73713154",
           999 => x"547282d6",
          1000 => x"e408ec05",
          1001 => x"238bd839",
          1002 => x"82d6e408",
          1003 => x"90050882",
          1004 => x"d6e40890",
          1005 => x"05088405",
          1006 => x"82d6e408",
          1007 => x"90050c70",
          1008 => x"0882d6e4",
          1009 => x"08fc050c",
          1010 => x"82d6e408",
          1011 => x"e4052270",
          1012 => x"832a7081",
          1013 => x"06515151",
          1014 => x"5372802e",
          1015 => x"ab3882d6",
          1016 => x"e408e805",
          1017 => x"3370982b",
          1018 => x"5372982c",
          1019 => x"5382d6e4",
          1020 => x"08fc0508",
          1021 => x"5253a2ec",
          1022 => x"3f82d6d8",
          1023 => x"08537282",
          1024 => x"d6e408f4",
          1025 => x"05239939",
          1026 => x"82d6e408",
          1027 => x"fc050851",
          1028 => x"9bf33f82",
          1029 => x"d6d80853",
          1030 => x"7282d6e4",
          1031 => x"08f40523",
          1032 => x"82d6e408",
          1033 => x"ec052253",
          1034 => x"82d6e408",
          1035 => x"f4052273",
          1036 => x"71315454",
          1037 => x"7282d6e4",
          1038 => x"08ec0523",
          1039 => x"8ac13982",
          1040 => x"d6e408e4",
          1041 => x"05227082",
          1042 => x"2a708106",
          1043 => x"51515372",
          1044 => x"802ea438",
          1045 => x"82d6e408",
          1046 => x"90050882",
          1047 => x"d6e40890",
          1048 => x"05088405",
          1049 => x"82d6e408",
          1050 => x"90050c70",
          1051 => x"0882d6e4",
          1052 => x"08dc050c",
          1053 => x"53a23982",
          1054 => x"d6e40890",
          1055 => x"050882d6",
          1056 => x"e4089005",
          1057 => x"08840582",
          1058 => x"d6e40890",
          1059 => x"050c7008",
          1060 => x"82d6e408",
          1061 => x"dc050c53",
          1062 => x"82d6e408",
          1063 => x"dc050882",
          1064 => x"d6e408fc",
          1065 => x"050c82d6",
          1066 => x"e408fc05",
          1067 => x"088025a4",
          1068 => x"3882d6e4",
          1069 => x"08e40522",
          1070 => x"70820751",
          1071 => x"537282d6",
          1072 => x"e408e405",
          1073 => x"2382d6e4",
          1074 => x"08fc0508",
          1075 => x"3082d6e4",
          1076 => x"08fc050c",
          1077 => x"82d6e408",
          1078 => x"e4052270",
          1079 => x"ffbf0651",
          1080 => x"537282d6",
          1081 => x"e408e405",
          1082 => x"2381af39",
          1083 => x"880b82d6",
          1084 => x"e408f405",
          1085 => x"23a93982",
          1086 => x"d6e408e4",
          1087 => x"05227080",
          1088 => x"c0075153",
          1089 => x"7282d6e4",
          1090 => x"08e40523",
          1091 => x"80f80b82",
          1092 => x"d6e408f8",
          1093 => x"0534900b",
          1094 => x"82d6e408",
          1095 => x"f4052382",
          1096 => x"d6e408e4",
          1097 => x"05227082",
          1098 => x"2a708106",
          1099 => x"51515372",
          1100 => x"802ea438",
          1101 => x"82d6e408",
          1102 => x"90050882",
          1103 => x"d6e40890",
          1104 => x"05088405",
          1105 => x"82d6e408",
          1106 => x"90050c70",
          1107 => x"0882d6e4",
          1108 => x"08d8050c",
          1109 => x"53a23982",
          1110 => x"d6e40890",
          1111 => x"050882d6",
          1112 => x"e4089005",
          1113 => x"08840582",
          1114 => x"d6e40890",
          1115 => x"050c7008",
          1116 => x"82d6e408",
          1117 => x"d8050c53",
          1118 => x"82d6e408",
          1119 => x"d8050882",
          1120 => x"d6e408fc",
          1121 => x"050c82d6",
          1122 => x"e408e405",
          1123 => x"2270cf06",
          1124 => x"51537282",
          1125 => x"d6e408e4",
          1126 => x"052382d6",
          1127 => x"e80b82d6",
          1128 => x"e408f005",
          1129 => x"0c82d6e4",
          1130 => x"08f00508",
          1131 => x"82d6e408",
          1132 => x"f4052282",
          1133 => x"d6e408fc",
          1134 => x"05087155",
          1135 => x"70545654",
          1136 => x"55a59e3f",
          1137 => x"82d6d808",
          1138 => x"53727534",
          1139 => x"82d6e408",
          1140 => x"f0050882",
          1141 => x"d6e408d4",
          1142 => x"050c82d6",
          1143 => x"e408f005",
          1144 => x"08703351",
          1145 => x"53897327",
          1146 => x"a43882d6",
          1147 => x"e408f005",
          1148 => x"08537233",
          1149 => x"5482d6e4",
          1150 => x"08f80533",
          1151 => x"7015df11",
          1152 => x"51515372",
          1153 => x"82d6e408",
          1154 => x"d0053497",
          1155 => x"3982d6e4",
          1156 => x"08f00508",
          1157 => x"537233b0",
          1158 => x"11515372",
          1159 => x"82d6e408",
          1160 => x"d0053482",
          1161 => x"d6e408d4",
          1162 => x"05085382",
          1163 => x"d6e408d0",
          1164 => x"05337334",
          1165 => x"82d6e408",
          1166 => x"f0050881",
          1167 => x"0582d6e4",
          1168 => x"08f0050c",
          1169 => x"82d6e408",
          1170 => x"f4052270",
          1171 => x"5382d6e4",
          1172 => x"08fc0508",
          1173 => x"5253a3d6",
          1174 => x"3f82d6d8",
          1175 => x"087082d6",
          1176 => x"e408fc05",
          1177 => x"0c5382d6",
          1178 => x"e408fc05",
          1179 => x"08802e84",
          1180 => x"38feb239",
          1181 => x"82d6e408",
          1182 => x"f0050882",
          1183 => x"d6e85455",
          1184 => x"72547470",
          1185 => x"75315153",
          1186 => x"7282d6e4",
          1187 => x"08fc0534",
          1188 => x"82d6e408",
          1189 => x"e4052270",
          1190 => x"b2065153",
          1191 => x"72802e94",
          1192 => x"3882d6e4",
          1193 => x"08ec0522",
          1194 => x"ff115153",
          1195 => x"7282d6e4",
          1196 => x"08ec0523",
          1197 => x"82d6e408",
          1198 => x"e4052270",
          1199 => x"862a7081",
          1200 => x"06515153",
          1201 => x"72802e80",
          1202 => x"e73882d6",
          1203 => x"e408ec05",
          1204 => x"2270902b",
          1205 => x"82d6e408",
          1206 => x"cc050c82",
          1207 => x"d6e408cc",
          1208 => x"0508902c",
          1209 => x"82d6e408",
          1210 => x"cc050c82",
          1211 => x"d6e408f4",
          1212 => x"05225153",
          1213 => x"72902e09",
          1214 => x"81069538",
          1215 => x"82d6e408",
          1216 => x"cc0508fe",
          1217 => x"05537282",
          1218 => x"d6e408c8",
          1219 => x"05239339",
          1220 => x"82d6e408",
          1221 => x"cc0508ff",
          1222 => x"05537282",
          1223 => x"d6e408c8",
          1224 => x"052382d6",
          1225 => x"e408c805",
          1226 => x"2282d6e4",
          1227 => x"08ec0523",
          1228 => x"82d6e408",
          1229 => x"e4052270",
          1230 => x"832a7081",
          1231 => x"06515153",
          1232 => x"72802e80",
          1233 => x"d03882d6",
          1234 => x"e408e805",
          1235 => x"3370982b",
          1236 => x"70982c82",
          1237 => x"d6e408fc",
          1238 => x"05335751",
          1239 => x"51537274",
          1240 => x"24973882",
          1241 => x"d6e408e4",
          1242 => x"052270f7",
          1243 => x"06515372",
          1244 => x"82d6e408",
          1245 => x"e405239d",
          1246 => x"3982d6e4",
          1247 => x"08e80533",
          1248 => x"5382d6e4",
          1249 => x"08fc0533",
          1250 => x"73713154",
          1251 => x"547282d6",
          1252 => x"e408e805",
          1253 => x"3482d6e4",
          1254 => x"08e40522",
          1255 => x"70832a70",
          1256 => x"81065151",
          1257 => x"5372802e",
          1258 => x"b13882d6",
          1259 => x"e408e805",
          1260 => x"3370882b",
          1261 => x"70902b70",
          1262 => x"902c7088",
          1263 => x"2c515151",
          1264 => x"51537254",
          1265 => x"82d6e408",
          1266 => x"ec052270",
          1267 => x"75315153",
          1268 => x"7282d6e4",
          1269 => x"08ec0523",
          1270 => x"af3982d6",
          1271 => x"e408fc05",
          1272 => x"3370882b",
          1273 => x"70902b70",
          1274 => x"902c7088",
          1275 => x"2c515151",
          1276 => x"51537254",
          1277 => x"82d6e408",
          1278 => x"ec052270",
          1279 => x"75315153",
          1280 => x"7282d6e4",
          1281 => x"08ec0523",
          1282 => x"82d6e408",
          1283 => x"e4052270",
          1284 => x"83800651",
          1285 => x"5372b038",
          1286 => x"82d6e408",
          1287 => x"ec0522ff",
          1288 => x"11545472",
          1289 => x"82d6e408",
          1290 => x"ec052373",
          1291 => x"902b7090",
          1292 => x"2c515380",
          1293 => x"73259038",
          1294 => x"82d6e408",
          1295 => x"88050852",
          1296 => x"a0518aee",
          1297 => x"3fd23982",
          1298 => x"d6e408e4",
          1299 => x"05227081",
          1300 => x"2a708106",
          1301 => x"51515372",
          1302 => x"802e9138",
          1303 => x"82d6e408",
          1304 => x"88050852",
          1305 => x"ad518aca",
          1306 => x"3f80c739",
          1307 => x"82d6e408",
          1308 => x"e4052270",
          1309 => x"842a7081",
          1310 => x"06515153",
          1311 => x"72802e90",
          1312 => x"3882d6e4",
          1313 => x"08880508",
          1314 => x"52ab518a",
          1315 => x"a53fa339",
          1316 => x"82d6e408",
          1317 => x"e4052270",
          1318 => x"852a7081",
          1319 => x"06515153",
          1320 => x"72802e8e",
          1321 => x"3882d6e4",
          1322 => x"08880508",
          1323 => x"52a0518a",
          1324 => x"813f82d6",
          1325 => x"e408e405",
          1326 => x"2270862a",
          1327 => x"70810651",
          1328 => x"51537280",
          1329 => x"2eb13882",
          1330 => x"d6e40888",
          1331 => x"050852b0",
          1332 => x"5189df3f",
          1333 => x"82d6e408",
          1334 => x"f4052253",
          1335 => x"72902e09",
          1336 => x"81069438",
          1337 => x"82d6e408",
          1338 => x"88050852",
          1339 => x"82d6e408",
          1340 => x"f8053351",
          1341 => x"89bc3f82",
          1342 => x"d6e408e4",
          1343 => x"05227088",
          1344 => x"2a708106",
          1345 => x"51515372",
          1346 => x"802eb038",
          1347 => x"82d6e408",
          1348 => x"ec0522ff",
          1349 => x"11545472",
          1350 => x"82d6e408",
          1351 => x"ec052373",
          1352 => x"902b7090",
          1353 => x"2c515380",
          1354 => x"73259038",
          1355 => x"82d6e408",
          1356 => x"88050852",
          1357 => x"b05188fa",
          1358 => x"3fd23982",
          1359 => x"d6e408e4",
          1360 => x"05227083",
          1361 => x"2a708106",
          1362 => x"51515372",
          1363 => x"802eb038",
          1364 => x"82d6e408",
          1365 => x"e80533ff",
          1366 => x"11545472",
          1367 => x"82d6e408",
          1368 => x"e8053473",
          1369 => x"982b7098",
          1370 => x"2c515380",
          1371 => x"73259038",
          1372 => x"82d6e408",
          1373 => x"88050852",
          1374 => x"b05188b6",
          1375 => x"3fd23982",
          1376 => x"d6e408e4",
          1377 => x"05227087",
          1378 => x"2a708106",
          1379 => x"51515372",
          1380 => x"b03882d6",
          1381 => x"e408ec05",
          1382 => x"22ff1154",
          1383 => x"547282d6",
          1384 => x"e408ec05",
          1385 => x"2373902b",
          1386 => x"70902c51",
          1387 => x"53807325",
          1388 => x"903882d6",
          1389 => x"e4088805",
          1390 => x"0852a051",
          1391 => x"87f43fd2",
          1392 => x"3982d6e4",
          1393 => x"08f80533",
          1394 => x"537280e3",
          1395 => x"2e098106",
          1396 => x"973882d6",
          1397 => x"e4088805",
          1398 => x"085282d6",
          1399 => x"e408fc05",
          1400 => x"335187ce",
          1401 => x"3f81ee39",
          1402 => x"82d6e408",
          1403 => x"f8053353",
          1404 => x"7280f32e",
          1405 => x"09810680",
          1406 => x"cb3882d6",
          1407 => x"e408f405",
          1408 => x"22ff1151",
          1409 => x"537282d6",
          1410 => x"e408f405",
          1411 => x"237283ff",
          1412 => x"ff065372",
          1413 => x"83ffff2e",
          1414 => x"81bb3882",
          1415 => x"d6e40888",
          1416 => x"05085282",
          1417 => x"d6e408fc",
          1418 => x"05087033",
          1419 => x"5282d6e4",
          1420 => x"08fc0508",
          1421 => x"810582d6",
          1422 => x"e408fc05",
          1423 => x"0c5386f2",
          1424 => x"3fffb739",
          1425 => x"82d6e408",
          1426 => x"f8053353",
          1427 => x"7280d32e",
          1428 => x"09810680",
          1429 => x"cb3882d6",
          1430 => x"e408f405",
          1431 => x"22ff1151",
          1432 => x"537282d6",
          1433 => x"e408f405",
          1434 => x"237283ff",
          1435 => x"ff065372",
          1436 => x"83ffff2e",
          1437 => x"80df3882",
          1438 => x"d6e40888",
          1439 => x"05085282",
          1440 => x"d6e408fc",
          1441 => x"05087033",
          1442 => x"525386a6",
          1443 => x"3f82d6e4",
          1444 => x"08fc0508",
          1445 => x"810582d6",
          1446 => x"e408fc05",
          1447 => x"0cffb739",
          1448 => x"82d6e408",
          1449 => x"f0050882",
          1450 => x"d6e82ea9",
          1451 => x"3882d6e4",
          1452 => x"08880508",
          1453 => x"5282d6e4",
          1454 => x"08f00508",
          1455 => x"ff0582d6",
          1456 => x"e408f005",
          1457 => x"0c82d6e4",
          1458 => x"08f00508",
          1459 => x"70335253",
          1460 => x"85e03fcc",
          1461 => x"3982d6e4",
          1462 => x"08e40522",
          1463 => x"70872a70",
          1464 => x"81065151",
          1465 => x"5372802e",
          1466 => x"80c33882",
          1467 => x"d6e408ec",
          1468 => x"0522ff11",
          1469 => x"54547282",
          1470 => x"d6e408ec",
          1471 => x"05237390",
          1472 => x"2b70902c",
          1473 => x"51538073",
          1474 => x"25a33882",
          1475 => x"d6e40888",
          1476 => x"050852a0",
          1477 => x"51859b3f",
          1478 => x"d23982d6",
          1479 => x"e4088805",
          1480 => x"085282d6",
          1481 => x"e408f805",
          1482 => x"33518586",
          1483 => x"3f800b82",
          1484 => x"d6e408e4",
          1485 => x"0523eab7",
          1486 => x"3982d6e4",
          1487 => x"08f80533",
          1488 => x"5372a52e",
          1489 => x"098106a8",
          1490 => x"38810b82",
          1491 => x"d6e408e4",
          1492 => x"0523800b",
          1493 => x"82d6e408",
          1494 => x"ec052380",
          1495 => x"0b82d6e4",
          1496 => x"08e80534",
          1497 => x"8a0b82d6",
          1498 => x"e408f405",
          1499 => x"23ea8039",
          1500 => x"82d6e408",
          1501 => x"88050852",
          1502 => x"82d6e408",
          1503 => x"f8053351",
          1504 => x"84b03fe9",
          1505 => x"ea3982d6",
          1506 => x"e4088805",
          1507 => x"088c1108",
          1508 => x"7082d6e4",
          1509 => x"08e0050c",
          1510 => x"515382d6",
          1511 => x"e408e005",
          1512 => x"0882d6d8",
          1513 => x"0c953d0d",
          1514 => x"82d6e40c",
          1515 => x"0482d6e4",
          1516 => x"080282d6",
          1517 => x"e40cfd3d",
          1518 => x"0d82f2b8",
          1519 => x"085382d6",
          1520 => x"e4088c05",
          1521 => x"085282d6",
          1522 => x"e4088805",
          1523 => x"0851e4dd",
          1524 => x"3f82d6d8",
          1525 => x"087082d6",
          1526 => x"d80c5485",
          1527 => x"3d0d82d6",
          1528 => x"e40c0482",
          1529 => x"d6e40802",
          1530 => x"82d6e40c",
          1531 => x"fb3d0d80",
          1532 => x"0b82d6e4",
          1533 => x"08f8050c",
          1534 => x"82f2bc08",
          1535 => x"85113370",
          1536 => x"812a7081",
          1537 => x"32708106",
          1538 => x"51515151",
          1539 => x"5372802e",
          1540 => x"8d38ff0b",
          1541 => x"82d6e408",
          1542 => x"f4050c81",
          1543 => x"923982d6",
          1544 => x"e4088805",
          1545 => x"08537233",
          1546 => x"82d6e408",
          1547 => x"88050881",
          1548 => x"0582d6e4",
          1549 => x"0888050c",
          1550 => x"537282d6",
          1551 => x"e408fc05",
          1552 => x"347281ff",
          1553 => x"06537280",
          1554 => x"2eb03882",
          1555 => x"f2bc0882",
          1556 => x"f2bc0853",
          1557 => x"82d6e408",
          1558 => x"fc053352",
          1559 => x"90110851",
          1560 => x"53722d82",
          1561 => x"d6d80853",
          1562 => x"72802eff",
          1563 => x"b138ff0b",
          1564 => x"82d6e408",
          1565 => x"f8050cff",
          1566 => x"a53982f2",
          1567 => x"bc0882f2",
          1568 => x"bc085353",
          1569 => x"8a519013",
          1570 => x"0853722d",
          1571 => x"82d6d808",
          1572 => x"5372802e",
          1573 => x"8a38ff0b",
          1574 => x"82d6e408",
          1575 => x"f8050c82",
          1576 => x"d6e408f8",
          1577 => x"05087082",
          1578 => x"d6e408f4",
          1579 => x"050c5382",
          1580 => x"d6e408f4",
          1581 => x"050882d6",
          1582 => x"d80c873d",
          1583 => x"0d82d6e4",
          1584 => x"0c0482d6",
          1585 => x"e4080282",
          1586 => x"d6e40cfb",
          1587 => x"3d0d800b",
          1588 => x"82d6e408",
          1589 => x"f8050c82",
          1590 => x"d6e4088c",
          1591 => x"05088511",
          1592 => x"3370812a",
          1593 => x"70813270",
          1594 => x"81065151",
          1595 => x"51515372",
          1596 => x"802e8d38",
          1597 => x"ff0b82d6",
          1598 => x"e408f405",
          1599 => x"0c80f339",
          1600 => x"82d6e408",
          1601 => x"88050853",
          1602 => x"723382d6",
          1603 => x"e4088805",
          1604 => x"08810582",
          1605 => x"d6e40888",
          1606 => x"050c5372",
          1607 => x"82d6e408",
          1608 => x"fc053472",
          1609 => x"81ff0653",
          1610 => x"72802eb6",
          1611 => x"3882d6e4",
          1612 => x"088c0508",
          1613 => x"82d6e408",
          1614 => x"8c050853",
          1615 => x"82d6e408",
          1616 => x"fc053352",
          1617 => x"90110851",
          1618 => x"53722d82",
          1619 => x"d6d80853",
          1620 => x"72802eff",
          1621 => x"ab38ff0b",
          1622 => x"82d6e408",
          1623 => x"f8050cff",
          1624 => x"9f3982d6",
          1625 => x"e408f805",
          1626 => x"087082d6",
          1627 => x"e408f405",
          1628 => x"0c5382d6",
          1629 => x"e408f405",
          1630 => x"0882d6d8",
          1631 => x"0c873d0d",
          1632 => x"82d6e40c",
          1633 => x"0482d6e4",
          1634 => x"080282d6",
          1635 => x"e40cfe3d",
          1636 => x"0d82f2bc",
          1637 => x"085282d6",
          1638 => x"e4088805",
          1639 => x"0851933f",
          1640 => x"82d6d808",
          1641 => x"7082d6d8",
          1642 => x"0c53843d",
          1643 => x"0d82d6e4",
          1644 => x"0c0482d6",
          1645 => x"e4080282",
          1646 => x"d6e40cfb",
          1647 => x"3d0d82d6",
          1648 => x"e4088c05",
          1649 => x"08851133",
          1650 => x"70812a70",
          1651 => x"81327081",
          1652 => x"06515151",
          1653 => x"51537280",
          1654 => x"2e8d38ff",
          1655 => x"0b82d6e4",
          1656 => x"08fc050c",
          1657 => x"81cb3982",
          1658 => x"d6e4088c",
          1659 => x"05088511",
          1660 => x"3370822a",
          1661 => x"70810651",
          1662 => x"51515372",
          1663 => x"802e80db",
          1664 => x"3882d6e4",
          1665 => x"088c0508",
          1666 => x"82d6e408",
          1667 => x"8c050854",
          1668 => x"548c1408",
          1669 => x"88140825",
          1670 => x"9f3882d6",
          1671 => x"e4088c05",
          1672 => x"08700870",
          1673 => x"82d6e408",
          1674 => x"88050852",
          1675 => x"57545472",
          1676 => x"75347308",
          1677 => x"8105740c",
          1678 => x"82d6e408",
          1679 => x"8c05088c",
          1680 => x"11088105",
          1681 => x"8c120c82",
          1682 => x"d6e40888",
          1683 => x"05087082",
          1684 => x"d6e408fc",
          1685 => x"050c5153",
          1686 => x"80d73982",
          1687 => x"d6e4088c",
          1688 => x"050882d6",
          1689 => x"e4088c05",
          1690 => x"085382d6",
          1691 => x"e4088805",
          1692 => x"087081ff",
          1693 => x"06539012",
          1694 => x"08515454",
          1695 => x"722d82d6",
          1696 => x"d8085372",
          1697 => x"a33882d6",
          1698 => x"e4088c05",
          1699 => x"088c1108",
          1700 => x"81058c12",
          1701 => x"0c82d6e4",
          1702 => x"08880508",
          1703 => x"7082d6e4",
          1704 => x"08fc050c",
          1705 => x"51538a39",
          1706 => x"ff0b82d6",
          1707 => x"e408fc05",
          1708 => x"0c82d6e4",
          1709 => x"08fc0508",
          1710 => x"82d6d80c",
          1711 => x"873d0d82",
          1712 => x"d6e40c04",
          1713 => x"82d6e408",
          1714 => x"0282d6e4",
          1715 => x"0cf93d0d",
          1716 => x"82d6e408",
          1717 => x"88050885",
          1718 => x"11337081",
          1719 => x"32708106",
          1720 => x"51515152",
          1721 => x"71802e8d",
          1722 => x"38ff0b82",
          1723 => x"d6e408f8",
          1724 => x"050c8394",
          1725 => x"3982d6e4",
          1726 => x"08880508",
          1727 => x"85113370",
          1728 => x"862a7081",
          1729 => x"06515151",
          1730 => x"5271802e",
          1731 => x"80c53882",
          1732 => x"d6e40888",
          1733 => x"050882d6",
          1734 => x"e4088805",
          1735 => x"08535385",
          1736 => x"123370ff",
          1737 => x"bf065152",
          1738 => x"71851434",
          1739 => x"82d6e408",
          1740 => x"8805088c",
          1741 => x"11088105",
          1742 => x"8c120c82",
          1743 => x"d6e40888",
          1744 => x"05088411",
          1745 => x"337082d6",
          1746 => x"e408f805",
          1747 => x"0c515152",
          1748 => x"82b63982",
          1749 => x"d6e40888",
          1750 => x"05088511",
          1751 => x"3370822a",
          1752 => x"70810651",
          1753 => x"51515271",
          1754 => x"802e80d7",
          1755 => x"3882d6e4",
          1756 => x"08880508",
          1757 => x"70087033",
          1758 => x"82d6e408",
          1759 => x"fc050c51",
          1760 => x"5282d6e4",
          1761 => x"08fc0508",
          1762 => x"a93882d6",
          1763 => x"e4088805",
          1764 => x"0882d6e4",
          1765 => x"08880508",
          1766 => x"53538512",
          1767 => x"3370a007",
          1768 => x"51527185",
          1769 => x"1434ff0b",
          1770 => x"82d6e408",
          1771 => x"f8050c81",
          1772 => x"d73982d6",
          1773 => x"e4088805",
          1774 => x"08700881",
          1775 => x"05710c52",
          1776 => x"81a13982",
          1777 => x"d6e40888",
          1778 => x"050882d6",
          1779 => x"e4088805",
          1780 => x"08529411",
          1781 => x"08515271",
          1782 => x"2d82d6d8",
          1783 => x"087082d6",
          1784 => x"e408fc05",
          1785 => x"0c5282d6",
          1786 => x"e408fc05",
          1787 => x"08802580",
          1788 => x"f23882d6",
          1789 => x"e4088805",
          1790 => x"0882d6e4",
          1791 => x"08f4050c",
          1792 => x"82d6e408",
          1793 => x"88050885",
          1794 => x"113382d6",
          1795 => x"e408f005",
          1796 => x"0c5282d6",
          1797 => x"e408fc05",
          1798 => x"08ff2e09",
          1799 => x"81069538",
          1800 => x"82d6e408",
          1801 => x"f0050890",
          1802 => x"07527182",
          1803 => x"d6e408ec",
          1804 => x"05349339",
          1805 => x"82d6e408",
          1806 => x"f00508a0",
          1807 => x"07527182",
          1808 => x"d6e408ec",
          1809 => x"053482d6",
          1810 => x"e408f405",
          1811 => x"085282d6",
          1812 => x"e408ec05",
          1813 => x"33851334",
          1814 => x"ff0b82d6",
          1815 => x"e408f805",
          1816 => x"0ca63982",
          1817 => x"d6e40888",
          1818 => x"05088c11",
          1819 => x"0881058c",
          1820 => x"120c82d6",
          1821 => x"e408fc05",
          1822 => x"087081ff",
          1823 => x"067082d6",
          1824 => x"e408f805",
          1825 => x"0c515152",
          1826 => x"82d6e408",
          1827 => x"f8050882",
          1828 => x"d6d80c89",
          1829 => x"3d0d82d6",
          1830 => x"e40c0482",
          1831 => x"d6e40802",
          1832 => x"82d6e40c",
          1833 => x"fd3d0d82",
          1834 => x"d6e40888",
          1835 => x"050882d6",
          1836 => x"e408fc05",
          1837 => x"0c82d6e4",
          1838 => x"088c0508",
          1839 => x"82d6e408",
          1840 => x"f8050c82",
          1841 => x"d6e40890",
          1842 => x"0508802e",
          1843 => x"82a23882",
          1844 => x"d6e408f8",
          1845 => x"050882d6",
          1846 => x"e408fc05",
          1847 => x"082681ac",
          1848 => x"3882d6e4",
          1849 => x"08f80508",
          1850 => x"82d6e408",
          1851 => x"90050805",
          1852 => x"5182d6e4",
          1853 => x"08fc0508",
          1854 => x"71278190",
          1855 => x"3882d6e4",
          1856 => x"08fc0508",
          1857 => x"82d6e408",
          1858 => x"90050805",
          1859 => x"82d6e408",
          1860 => x"fc050c82",
          1861 => x"d6e408f8",
          1862 => x"050882d6",
          1863 => x"e4089005",
          1864 => x"080582d6",
          1865 => x"e408f805",
          1866 => x"0c82d6e4",
          1867 => x"08900508",
          1868 => x"810582d6",
          1869 => x"e4089005",
          1870 => x"0c82d6e4",
          1871 => x"08900508",
          1872 => x"ff0582d6",
          1873 => x"e4089005",
          1874 => x"0c82d6e4",
          1875 => x"08900508",
          1876 => x"802e819c",
          1877 => x"3882d6e4",
          1878 => x"08fc0508",
          1879 => x"ff0582d6",
          1880 => x"e408fc05",
          1881 => x"0c82d6e4",
          1882 => x"08f80508",
          1883 => x"ff0582d6",
          1884 => x"e408f805",
          1885 => x"0c82d6e4",
          1886 => x"08fc0508",
          1887 => x"82d6e408",
          1888 => x"f8050853",
          1889 => x"51713371",
          1890 => x"34ffae39",
          1891 => x"82d6e408",
          1892 => x"90050881",
          1893 => x"0582d6e4",
          1894 => x"0890050c",
          1895 => x"82d6e408",
          1896 => x"900508ff",
          1897 => x"0582d6e4",
          1898 => x"0890050c",
          1899 => x"82d6e408",
          1900 => x"90050880",
          1901 => x"2eba3882",
          1902 => x"d6e408f8",
          1903 => x"05085170",
          1904 => x"3382d6e4",
          1905 => x"08f80508",
          1906 => x"810582d6",
          1907 => x"e408f805",
          1908 => x"0c82d6e4",
          1909 => x"08fc0508",
          1910 => x"52527171",
          1911 => x"3482d6e4",
          1912 => x"08fc0508",
          1913 => x"810582d6",
          1914 => x"e408fc05",
          1915 => x"0cffad39",
          1916 => x"82d6e408",
          1917 => x"88050870",
          1918 => x"82d6d80c",
          1919 => x"51853d0d",
          1920 => x"82d6e40c",
          1921 => x"0482d6e4",
          1922 => x"080282d6",
          1923 => x"e40cfe3d",
          1924 => x"0d82d6e4",
          1925 => x"08880508",
          1926 => x"82d6e408",
          1927 => x"fc050c82",
          1928 => x"d6e408fc",
          1929 => x"05085271",
          1930 => x"3382d6e4",
          1931 => x"08fc0508",
          1932 => x"810582d6",
          1933 => x"e408fc05",
          1934 => x"0c7081ff",
          1935 => x"06515170",
          1936 => x"802e8338",
          1937 => x"da3982d6",
          1938 => x"e408fc05",
          1939 => x"08ff0582",
          1940 => x"d6e408fc",
          1941 => x"050c82d6",
          1942 => x"e408fc05",
          1943 => x"0882d6e4",
          1944 => x"08880508",
          1945 => x"317082d6",
          1946 => x"d80c5184",
          1947 => x"3d0d82d6",
          1948 => x"e40c0482",
          1949 => x"d6e40802",
          1950 => x"82d6e40c",
          1951 => x"fe3d0d82",
          1952 => x"d6e40888",
          1953 => x"050882d6",
          1954 => x"e408fc05",
          1955 => x"0c82d6e4",
          1956 => x"088c0508",
          1957 => x"52713382",
          1958 => x"d6e4088c",
          1959 => x"05088105",
          1960 => x"82d6e408",
          1961 => x"8c050c82",
          1962 => x"d6e408fc",
          1963 => x"05085351",
          1964 => x"70723482",
          1965 => x"d6e408fc",
          1966 => x"05088105",
          1967 => x"82d6e408",
          1968 => x"fc050c70",
          1969 => x"81ff0651",
          1970 => x"70802e84",
          1971 => x"38ffbe39",
          1972 => x"82d6e408",
          1973 => x"88050870",
          1974 => x"82d6d80c",
          1975 => x"51843d0d",
          1976 => x"82d6e40c",
          1977 => x"0482d6e4",
          1978 => x"080282d6",
          1979 => x"e40cfd3d",
          1980 => x"0d82d6e4",
          1981 => x"08880508",
          1982 => x"82d6e408",
          1983 => x"fc050c82",
          1984 => x"d6e4088c",
          1985 => x"050882d6",
          1986 => x"e408f805",
          1987 => x"0c82d6e4",
          1988 => x"08900508",
          1989 => x"802e80e5",
          1990 => x"3882d6e4",
          1991 => x"08900508",
          1992 => x"810582d6",
          1993 => x"e4089005",
          1994 => x"0c82d6e4",
          1995 => x"08900508",
          1996 => x"ff0582d6",
          1997 => x"e4089005",
          1998 => x"0c82d6e4",
          1999 => x"08900508",
          2000 => x"802eba38",
          2001 => x"82d6e408",
          2002 => x"f8050851",
          2003 => x"703382d6",
          2004 => x"e408f805",
          2005 => x"08810582",
          2006 => x"d6e408f8",
          2007 => x"050c82d6",
          2008 => x"e408fc05",
          2009 => x"08525271",
          2010 => x"713482d6",
          2011 => x"e408fc05",
          2012 => x"08810582",
          2013 => x"d6e408fc",
          2014 => x"050cffad",
          2015 => x"3982d6e4",
          2016 => x"08880508",
          2017 => x"7082d6d8",
          2018 => x"0c51853d",
          2019 => x"0d82d6e4",
          2020 => x"0c0482d6",
          2021 => x"e4080282",
          2022 => x"d6e40cfd",
          2023 => x"3d0d82d6",
          2024 => x"e4089005",
          2025 => x"08802e81",
          2026 => x"f43882d6",
          2027 => x"e4088c05",
          2028 => x"08527133",
          2029 => x"82d6e408",
          2030 => x"8c050881",
          2031 => x"0582d6e4",
          2032 => x"088c050c",
          2033 => x"82d6e408",
          2034 => x"88050870",
          2035 => x"337281ff",
          2036 => x"06535454",
          2037 => x"5171712e",
          2038 => x"843880ce",
          2039 => x"3982d6e4",
          2040 => x"08880508",
          2041 => x"52713382",
          2042 => x"d6e40888",
          2043 => x"05088105",
          2044 => x"82d6e408",
          2045 => x"88050c70",
          2046 => x"81ff0651",
          2047 => x"51708d38",
          2048 => x"800b82d6",
          2049 => x"e408fc05",
          2050 => x"0c819b39",
          2051 => x"82d6e408",
          2052 => x"900508ff",
          2053 => x"0582d6e4",
          2054 => x"0890050c",
          2055 => x"82d6e408",
          2056 => x"90050880",
          2057 => x"2e8438ff",
          2058 => x"813982d6",
          2059 => x"e4089005",
          2060 => x"08802e80",
          2061 => x"e83882d6",
          2062 => x"e4088805",
          2063 => x"08703352",
          2064 => x"53708d38",
          2065 => x"ff0b82d6",
          2066 => x"e408fc05",
          2067 => x"0c80d739",
          2068 => x"82d6e408",
          2069 => x"8c0508ff",
          2070 => x"0582d6e4",
          2071 => x"088c050c",
          2072 => x"82d6e408",
          2073 => x"8c050870",
          2074 => x"33525270",
          2075 => x"8c38810b",
          2076 => x"82d6e408",
          2077 => x"fc050cae",
          2078 => x"3982d6e4",
          2079 => x"08880508",
          2080 => x"703382d6",
          2081 => x"e4088c05",
          2082 => x"08703372",
          2083 => x"71317082",
          2084 => x"d6e408fc",
          2085 => x"050c5355",
          2086 => x"5252538a",
          2087 => x"39800b82",
          2088 => x"d6e408fc",
          2089 => x"050c82d6",
          2090 => x"e408fc05",
          2091 => x"0882d6d8",
          2092 => x"0c853d0d",
          2093 => x"82d6e40c",
          2094 => x"0482d6e4",
          2095 => x"080282d6",
          2096 => x"e40cfa3d",
          2097 => x"0d82d6e4",
          2098 => x"088c0508",
          2099 => x"5282d6e4",
          2100 => x"08880508",
          2101 => x"51818d3f",
          2102 => x"82d6d808",
          2103 => x"7082d6e4",
          2104 => x"08f8050c",
          2105 => x"82d6e408",
          2106 => x"f8050881",
          2107 => x"05705351",
          2108 => x"5480e3f4",
          2109 => x"3f82d6d8",
          2110 => x"087082d6",
          2111 => x"e408fc05",
          2112 => x"0c5482d6",
          2113 => x"e408fc05",
          2114 => x"088c3880",
          2115 => x"0b82d6e4",
          2116 => x"08f4050c",
          2117 => x"bc3982d6",
          2118 => x"e408fc05",
          2119 => x"0882d6e4",
          2120 => x"08f80508",
          2121 => x"05548074",
          2122 => x"3482d6e4",
          2123 => x"08f80508",
          2124 => x"5382d6e4",
          2125 => x"08880508",
          2126 => x"5282d6e4",
          2127 => x"08fc0508",
          2128 => x"51fba23f",
          2129 => x"82d6d808",
          2130 => x"7082d6e4",
          2131 => x"08f4050c",
          2132 => x"5482d6e4",
          2133 => x"08f40508",
          2134 => x"82d6d80c",
          2135 => x"883d0d82",
          2136 => x"d6e40c04",
          2137 => x"82d6e408",
          2138 => x"0282d6e4",
          2139 => x"0cfd3d0d",
          2140 => x"82d6e408",
          2141 => x"88050882",
          2142 => x"d6e408f8",
          2143 => x"050c82d6",
          2144 => x"e4088c05",
          2145 => x"088d3880",
          2146 => x"0b82d6e4",
          2147 => x"08fc050c",
          2148 => x"80ec3982",
          2149 => x"d6e408f8",
          2150 => x"05085271",
          2151 => x"3382d6e4",
          2152 => x"08f80508",
          2153 => x"810582d6",
          2154 => x"e408f805",
          2155 => x"0c7081ff",
          2156 => x"06515170",
          2157 => x"802e9f38",
          2158 => x"82d6e408",
          2159 => x"8c0508ff",
          2160 => x"0582d6e4",
          2161 => x"088c050c",
          2162 => x"82d6e408",
          2163 => x"8c0508ff",
          2164 => x"2e8438ff",
          2165 => x"be3982d6",
          2166 => x"e408f805",
          2167 => x"08ff0582",
          2168 => x"d6e408f8",
          2169 => x"050c82d6",
          2170 => x"e408f805",
          2171 => x"0882d6e4",
          2172 => x"08880508",
          2173 => x"317082d6",
          2174 => x"e408fc05",
          2175 => x"0c5182d6",
          2176 => x"e408fc05",
          2177 => x"0882d6d8",
          2178 => x"0c853d0d",
          2179 => x"82d6e40c",
          2180 => x"0482d6e4",
          2181 => x"080282d6",
          2182 => x"e40cfe3d",
          2183 => x"0d82d6e4",
          2184 => x"08880508",
          2185 => x"82d6e408",
          2186 => x"fc050c82",
          2187 => x"d6e40890",
          2188 => x"0508802e",
          2189 => x"80d43882",
          2190 => x"d6e40890",
          2191 => x"05088105",
          2192 => x"82d6e408",
          2193 => x"90050c82",
          2194 => x"d6e40890",
          2195 => x"0508ff05",
          2196 => x"82d6e408",
          2197 => x"90050c82",
          2198 => x"d6e40890",
          2199 => x"0508802e",
          2200 => x"a93882d6",
          2201 => x"e4088c05",
          2202 => x"08517082",
          2203 => x"d6e408fc",
          2204 => x"05085252",
          2205 => x"71713482",
          2206 => x"d6e408fc",
          2207 => x"05088105",
          2208 => x"82d6e408",
          2209 => x"fc050cff",
          2210 => x"be3982d6",
          2211 => x"e4088805",
          2212 => x"087082d6",
          2213 => x"d80c5184",
          2214 => x"3d0d82d6",
          2215 => x"e40c0482",
          2216 => x"d6e40802",
          2217 => x"82d6e40c",
          2218 => x"f93d0d80",
          2219 => x"0b82d6e4",
          2220 => x"08fc050c",
          2221 => x"82d6e408",
          2222 => x"88050880",
          2223 => x"25b93882",
          2224 => x"d6e40888",
          2225 => x"05083082",
          2226 => x"d6e40888",
          2227 => x"050c800b",
          2228 => x"82d6e408",
          2229 => x"f4050c82",
          2230 => x"d6e408fc",
          2231 => x"05088a38",
          2232 => x"810b82d6",
          2233 => x"e408f405",
          2234 => x"0c82d6e4",
          2235 => x"08f40508",
          2236 => x"82d6e408",
          2237 => x"fc050c82",
          2238 => x"d6e4088c",
          2239 => x"05088025",
          2240 => x"b93882d6",
          2241 => x"e4088c05",
          2242 => x"083082d6",
          2243 => x"e4088c05",
          2244 => x"0c800b82",
          2245 => x"d6e408f0",
          2246 => x"050c82d6",
          2247 => x"e408fc05",
          2248 => x"088a3881",
          2249 => x"0b82d6e4",
          2250 => x"08f0050c",
          2251 => x"82d6e408",
          2252 => x"f0050882",
          2253 => x"d6e408fc",
          2254 => x"050c8053",
          2255 => x"82d6e408",
          2256 => x"8c050852",
          2257 => x"82d6e408",
          2258 => x"88050851",
          2259 => x"82c53f82",
          2260 => x"d6d80870",
          2261 => x"82d6e408",
          2262 => x"f8050c54",
          2263 => x"82d6e408",
          2264 => x"fc050880",
          2265 => x"2e903882",
          2266 => x"d6e408f8",
          2267 => x"05083082",
          2268 => x"d6e408f8",
          2269 => x"050c82d6",
          2270 => x"e408f805",
          2271 => x"087082d6",
          2272 => x"d80c5489",
          2273 => x"3d0d82d6",
          2274 => x"e40c0482",
          2275 => x"d6e40802",
          2276 => x"82d6e40c",
          2277 => x"fb3d0d80",
          2278 => x"0b82d6e4",
          2279 => x"08fc050c",
          2280 => x"82d6e408",
          2281 => x"88050880",
          2282 => x"25993882",
          2283 => x"d6e40888",
          2284 => x"05083082",
          2285 => x"d6e40888",
          2286 => x"050c810b",
          2287 => x"82d6e408",
          2288 => x"fc050c82",
          2289 => x"d6e4088c",
          2290 => x"05088025",
          2291 => x"903882d6",
          2292 => x"e4088c05",
          2293 => x"083082d6",
          2294 => x"e4088c05",
          2295 => x"0c815382",
          2296 => x"d6e4088c",
          2297 => x"05085282",
          2298 => x"d6e40888",
          2299 => x"05085181",
          2300 => x"a23f82d6",
          2301 => x"d8087082",
          2302 => x"d6e408f8",
          2303 => x"050c5482",
          2304 => x"d6e408fc",
          2305 => x"0508802e",
          2306 => x"903882d6",
          2307 => x"e408f805",
          2308 => x"083082d6",
          2309 => x"e408f805",
          2310 => x"0c82d6e4",
          2311 => x"08f80508",
          2312 => x"7082d6d8",
          2313 => x"0c54873d",
          2314 => x"0d82d6e4",
          2315 => x"0c0482d6",
          2316 => x"e4080282",
          2317 => x"d6e40cfd",
          2318 => x"3d0d8053",
          2319 => x"82d6e408",
          2320 => x"8c050852",
          2321 => x"82d6e408",
          2322 => x"88050851",
          2323 => x"80c53f82",
          2324 => x"d6d80870",
          2325 => x"82d6d80c",
          2326 => x"54853d0d",
          2327 => x"82d6e40c",
          2328 => x"0482d6e4",
          2329 => x"080282d6",
          2330 => x"e40cfd3d",
          2331 => x"0d815382",
          2332 => x"d6e4088c",
          2333 => x"05085282",
          2334 => x"d6e40888",
          2335 => x"05085193",
          2336 => x"3f82d6d8",
          2337 => x"087082d6",
          2338 => x"d80c5485",
          2339 => x"3d0d82d6",
          2340 => x"e40c0482",
          2341 => x"d6e40802",
          2342 => x"82d6e40c",
          2343 => x"fd3d0d81",
          2344 => x"0b82d6e4",
          2345 => x"08fc050c",
          2346 => x"800b82d6",
          2347 => x"e408f805",
          2348 => x"0c82d6e4",
          2349 => x"088c0508",
          2350 => x"82d6e408",
          2351 => x"88050827",
          2352 => x"b93882d6",
          2353 => x"e408fc05",
          2354 => x"08802eae",
          2355 => x"38800b82",
          2356 => x"d6e4088c",
          2357 => x"050824a2",
          2358 => x"3882d6e4",
          2359 => x"088c0508",
          2360 => x"1082d6e4",
          2361 => x"088c050c",
          2362 => x"82d6e408",
          2363 => x"fc050810",
          2364 => x"82d6e408",
          2365 => x"fc050cff",
          2366 => x"b83982d6",
          2367 => x"e408fc05",
          2368 => x"08802e80",
          2369 => x"e13882d6",
          2370 => x"e4088c05",
          2371 => x"0882d6e4",
          2372 => x"08880508",
          2373 => x"26ad3882",
          2374 => x"d6e40888",
          2375 => x"050882d6",
          2376 => x"e4088c05",
          2377 => x"083182d6",
          2378 => x"e4088805",
          2379 => x"0c82d6e4",
          2380 => x"08f80508",
          2381 => x"82d6e408",
          2382 => x"fc050807",
          2383 => x"82d6e408",
          2384 => x"f8050c82",
          2385 => x"d6e408fc",
          2386 => x"0508812a",
          2387 => x"82d6e408",
          2388 => x"fc050c82",
          2389 => x"d6e4088c",
          2390 => x"0508812a",
          2391 => x"82d6e408",
          2392 => x"8c050cff",
          2393 => x"953982d6",
          2394 => x"e4089005",
          2395 => x"08802e93",
          2396 => x"3882d6e4",
          2397 => x"08880508",
          2398 => x"7082d6e4",
          2399 => x"08f4050c",
          2400 => x"51913982",
          2401 => x"d6e408f8",
          2402 => x"05087082",
          2403 => x"d6e408f4",
          2404 => x"050c5182",
          2405 => x"d6e408f4",
          2406 => x"050882d6",
          2407 => x"d80c853d",
          2408 => x"0d82d6e4",
          2409 => x"0c0482d6",
          2410 => x"e4080282",
          2411 => x"d6e40cf7",
          2412 => x"3d0d800b",
          2413 => x"82d6e408",
          2414 => x"f0053482",
          2415 => x"d6e4088c",
          2416 => x"05085380",
          2417 => x"730c82d6",
          2418 => x"e4088805",
          2419 => x"08700851",
          2420 => x"53723353",
          2421 => x"7282d6e4",
          2422 => x"08f80534",
          2423 => x"7281ff06",
          2424 => x"5372a02e",
          2425 => x"09810691",
          2426 => x"3882d6e4",
          2427 => x"08880508",
          2428 => x"70088105",
          2429 => x"710c53ce",
          2430 => x"3982d6e4",
          2431 => x"08f80533",
          2432 => x"5372ad2e",
          2433 => x"098106a4",
          2434 => x"38810b82",
          2435 => x"d6e408f0",
          2436 => x"053482d6",
          2437 => x"e4088805",
          2438 => x"08700881",
          2439 => x"05710c70",
          2440 => x"08515372",
          2441 => x"3382d6e4",
          2442 => x"08f80534",
          2443 => x"82d6e408",
          2444 => x"f8053353",
          2445 => x"72b02e09",
          2446 => x"810681dc",
          2447 => x"3882d6e4",
          2448 => x"08880508",
          2449 => x"70088105",
          2450 => x"710c7008",
          2451 => x"51537233",
          2452 => x"82d6e408",
          2453 => x"f8053482",
          2454 => x"d6e408f8",
          2455 => x"053382d6",
          2456 => x"e408e805",
          2457 => x"0c82d6e4",
          2458 => x"08e80508",
          2459 => x"80e22eb6",
          2460 => x"3882d6e4",
          2461 => x"08e80508",
          2462 => x"80f82e84",
          2463 => x"3880cd39",
          2464 => x"900b82d6",
          2465 => x"e408f405",
          2466 => x"3482d6e4",
          2467 => x"08880508",
          2468 => x"70088105",
          2469 => x"710c7008",
          2470 => x"51537233",
          2471 => x"82d6e408",
          2472 => x"f8053481",
          2473 => x"a439820b",
          2474 => x"82d6e408",
          2475 => x"f4053482",
          2476 => x"d6e40888",
          2477 => x"05087008",
          2478 => x"8105710c",
          2479 => x"70085153",
          2480 => x"723382d6",
          2481 => x"e408f805",
          2482 => x"3480fe39",
          2483 => x"82d6e408",
          2484 => x"f8053353",
          2485 => x"72a0268d",
          2486 => x"38810b82",
          2487 => x"d6e408ec",
          2488 => x"050c8380",
          2489 => x"3982d6e4",
          2490 => x"08f80533",
          2491 => x"53af7327",
          2492 => x"903882d6",
          2493 => x"e408f805",
          2494 => x"335372b9",
          2495 => x"2683388d",
          2496 => x"39800b82",
          2497 => x"d6e408ec",
          2498 => x"050c82d8",
          2499 => x"39880b82",
          2500 => x"d6e408f4",
          2501 => x"0534b239",
          2502 => x"82d6e408",
          2503 => x"f8053353",
          2504 => x"af732790",
          2505 => x"3882d6e4",
          2506 => x"08f80533",
          2507 => x"5372b926",
          2508 => x"83388d39",
          2509 => x"800b82d6",
          2510 => x"e408ec05",
          2511 => x"0c82a539",
          2512 => x"8a0b82d6",
          2513 => x"e408f405",
          2514 => x"34800b82",
          2515 => x"d6e408fc",
          2516 => x"050c82d6",
          2517 => x"e408f805",
          2518 => x"3353a073",
          2519 => x"2781cf38",
          2520 => x"82d6e408",
          2521 => x"f8053353",
          2522 => x"80e07327",
          2523 => x"943882d6",
          2524 => x"e408f805",
          2525 => x"33e01151",
          2526 => x"537282d6",
          2527 => x"e408f805",
          2528 => x"3482d6e4",
          2529 => x"08f80533",
          2530 => x"d0115153",
          2531 => x"7282d6e4",
          2532 => x"08f80534",
          2533 => x"82d6e408",
          2534 => x"f8053353",
          2535 => x"907327ad",
          2536 => x"3882d6e4",
          2537 => x"08f80533",
          2538 => x"f9115153",
          2539 => x"7282d6e4",
          2540 => x"08f80534",
          2541 => x"82d6e408",
          2542 => x"f8053353",
          2543 => x"7289268d",
          2544 => x"38800b82",
          2545 => x"d6e408ec",
          2546 => x"050c8198",
          2547 => x"3982d6e4",
          2548 => x"08f80533",
          2549 => x"82d6e408",
          2550 => x"f4053354",
          2551 => x"54727426",
          2552 => x"8d38800b",
          2553 => x"82d6e408",
          2554 => x"ec050c80",
          2555 => x"f73982d6",
          2556 => x"e408f405",
          2557 => x"337082d6",
          2558 => x"e408fc05",
          2559 => x"082982d6",
          2560 => x"e408f805",
          2561 => x"33701282",
          2562 => x"d6e408fc",
          2563 => x"050c82d6",
          2564 => x"e4088805",
          2565 => x"08700881",
          2566 => x"05710c70",
          2567 => x"08515152",
          2568 => x"55537233",
          2569 => x"82d6e408",
          2570 => x"f80534fe",
          2571 => x"a53982d6",
          2572 => x"e408f005",
          2573 => x"33537280",
          2574 => x"2e903882",
          2575 => x"d6e408fc",
          2576 => x"05083082",
          2577 => x"d6e408fc",
          2578 => x"050c82d6",
          2579 => x"e4088c05",
          2580 => x"0882d6e4",
          2581 => x"08fc0508",
          2582 => x"710c5381",
          2583 => x"0b82d6e4",
          2584 => x"08ec050c",
          2585 => x"82d6e408",
          2586 => x"ec050882",
          2587 => x"d6d80c8b",
          2588 => x"3d0d82d6",
          2589 => x"e40c0482",
          2590 => x"d6e40802",
          2591 => x"82d6e40c",
          2592 => x"f73d0d80",
          2593 => x"0b82d6e4",
          2594 => x"08f00534",
          2595 => x"82d6e408",
          2596 => x"8c050853",
          2597 => x"80730c82",
          2598 => x"d6e40888",
          2599 => x"05087008",
          2600 => x"51537233",
          2601 => x"537282d6",
          2602 => x"e408f805",
          2603 => x"347281ff",
          2604 => x"065372a0",
          2605 => x"2e098106",
          2606 => x"913882d6",
          2607 => x"e4088805",
          2608 => x"08700881",
          2609 => x"05710c53",
          2610 => x"ce3982d6",
          2611 => x"e408f805",
          2612 => x"335372ad",
          2613 => x"2e098106",
          2614 => x"a438810b",
          2615 => x"82d6e408",
          2616 => x"f0053482",
          2617 => x"d6e40888",
          2618 => x"05087008",
          2619 => x"8105710c",
          2620 => x"70085153",
          2621 => x"723382d6",
          2622 => x"e408f805",
          2623 => x"3482d6e4",
          2624 => x"08f80533",
          2625 => x"5372b02e",
          2626 => x"09810681",
          2627 => x"dc3882d6",
          2628 => x"e4088805",
          2629 => x"08700881",
          2630 => x"05710c70",
          2631 => x"08515372",
          2632 => x"3382d6e4",
          2633 => x"08f80534",
          2634 => x"82d6e408",
          2635 => x"f8053382",
          2636 => x"d6e408e8",
          2637 => x"050c82d6",
          2638 => x"e408e805",
          2639 => x"0880e22e",
          2640 => x"b63882d6",
          2641 => x"e408e805",
          2642 => x"0880f82e",
          2643 => x"843880cd",
          2644 => x"39900b82",
          2645 => x"d6e408f4",
          2646 => x"053482d6",
          2647 => x"e4088805",
          2648 => x"08700881",
          2649 => x"05710c70",
          2650 => x"08515372",
          2651 => x"3382d6e4",
          2652 => x"08f80534",
          2653 => x"81a43982",
          2654 => x"0b82d6e4",
          2655 => x"08f40534",
          2656 => x"82d6e408",
          2657 => x"88050870",
          2658 => x"08810571",
          2659 => x"0c700851",
          2660 => x"53723382",
          2661 => x"d6e408f8",
          2662 => x"053480fe",
          2663 => x"3982d6e4",
          2664 => x"08f80533",
          2665 => x"5372a026",
          2666 => x"8d38810b",
          2667 => x"82d6e408",
          2668 => x"ec050c83",
          2669 => x"803982d6",
          2670 => x"e408f805",
          2671 => x"3353af73",
          2672 => x"27903882",
          2673 => x"d6e408f8",
          2674 => x"05335372",
          2675 => x"b9268338",
          2676 => x"8d39800b",
          2677 => x"82d6e408",
          2678 => x"ec050c82",
          2679 => x"d839880b",
          2680 => x"82d6e408",
          2681 => x"f40534b2",
          2682 => x"3982d6e4",
          2683 => x"08f80533",
          2684 => x"53af7327",
          2685 => x"903882d6",
          2686 => x"e408f805",
          2687 => x"335372b9",
          2688 => x"2683388d",
          2689 => x"39800b82",
          2690 => x"d6e408ec",
          2691 => x"050c82a5",
          2692 => x"398a0b82",
          2693 => x"d6e408f4",
          2694 => x"0534800b",
          2695 => x"82d6e408",
          2696 => x"fc050c82",
          2697 => x"d6e408f8",
          2698 => x"053353a0",
          2699 => x"732781cf",
          2700 => x"3882d6e4",
          2701 => x"08f80533",
          2702 => x"5380e073",
          2703 => x"27943882",
          2704 => x"d6e408f8",
          2705 => x"0533e011",
          2706 => x"51537282",
          2707 => x"d6e408f8",
          2708 => x"053482d6",
          2709 => x"e408f805",
          2710 => x"33d01151",
          2711 => x"537282d6",
          2712 => x"e408f805",
          2713 => x"3482d6e4",
          2714 => x"08f80533",
          2715 => x"53907327",
          2716 => x"ad3882d6",
          2717 => x"e408f805",
          2718 => x"33f91151",
          2719 => x"537282d6",
          2720 => x"e408f805",
          2721 => x"3482d6e4",
          2722 => x"08f80533",
          2723 => x"53728926",
          2724 => x"8d38800b",
          2725 => x"82d6e408",
          2726 => x"ec050c81",
          2727 => x"983982d6",
          2728 => x"e408f805",
          2729 => x"3382d6e4",
          2730 => x"08f40533",
          2731 => x"54547274",
          2732 => x"268d3880",
          2733 => x"0b82d6e4",
          2734 => x"08ec050c",
          2735 => x"80f73982",
          2736 => x"d6e408f4",
          2737 => x"05337082",
          2738 => x"d6e408fc",
          2739 => x"05082982",
          2740 => x"d6e408f8",
          2741 => x"05337012",
          2742 => x"82d6e408",
          2743 => x"fc050c82",
          2744 => x"d6e40888",
          2745 => x"05087008",
          2746 => x"8105710c",
          2747 => x"70085151",
          2748 => x"52555372",
          2749 => x"3382d6e4",
          2750 => x"08f80534",
          2751 => x"fea53982",
          2752 => x"d6e408f0",
          2753 => x"05335372",
          2754 => x"802e9038",
          2755 => x"82d6e408",
          2756 => x"fc050830",
          2757 => x"82d6e408",
          2758 => x"fc050c82",
          2759 => x"d6e4088c",
          2760 => x"050882d6",
          2761 => x"e408fc05",
          2762 => x"08710c53",
          2763 => x"810b82d6",
          2764 => x"e408ec05",
          2765 => x"0c82d6e4",
          2766 => x"08ec0508",
          2767 => x"82d6d80c",
          2768 => x"8b3d0d82",
          2769 => x"d6e40c04",
          2770 => x"f83d0d7a",
          2771 => x"70087056",
          2772 => x"56597480",
          2773 => x"2e80df38",
          2774 => x"8c397715",
          2775 => x"790c8516",
          2776 => x"335480d2",
          2777 => x"39743354",
          2778 => x"73a02e09",
          2779 => x"81068638",
          2780 => x"811555f1",
          2781 => x"39805776",
          2782 => x"902982d0",
          2783 => x"cc057008",
          2784 => x"5256e581",
          2785 => x"3f82d6d8",
          2786 => x"0882d6d8",
          2787 => x"08547553",
          2788 => x"76085258",
          2789 => x"e7fc3f82",
          2790 => x"d6d8088b",
          2791 => x"38841633",
          2792 => x"5473812e",
          2793 => x"ffb43881",
          2794 => x"177081ff",
          2795 => x"06585499",
          2796 => x"7727c438",
          2797 => x"ff547382",
          2798 => x"d6d80c8a",
          2799 => x"3d0d04ff",
          2800 => x"3d0d7352",
          2801 => x"71932681",
          2802 => x"8e387184",
          2803 => x"2982acdc",
          2804 => x"05527108",
          2805 => x"0482b2cc",
          2806 => x"51818039",
          2807 => x"82b2d851",
          2808 => x"80f93982",
          2809 => x"b2e85180",
          2810 => x"f23982b2",
          2811 => x"f85180eb",
          2812 => x"3982b388",
          2813 => x"5180e439",
          2814 => x"82b39851",
          2815 => x"80dd3982",
          2816 => x"b3ac5180",
          2817 => x"d63982b3",
          2818 => x"bc5180cf",
          2819 => x"3982b3d4",
          2820 => x"5180c839",
          2821 => x"82b3ec51",
          2822 => x"80c13982",
          2823 => x"b48451bb",
          2824 => x"3982b4a0",
          2825 => x"51b53982",
          2826 => x"b4b451af",
          2827 => x"3982b4dc",
          2828 => x"51a93982",
          2829 => x"b4ec51a3",
          2830 => x"3982b58c",
          2831 => x"519d3982",
          2832 => x"b59c5197",
          2833 => x"3982b5b4",
          2834 => x"51913982",
          2835 => x"b5cc518b",
          2836 => x"3982b5e4",
          2837 => x"51853982",
          2838 => x"b5f051d7",
          2839 => x"863f833d",
          2840 => x"0d04fb3d",
          2841 => x"0d777956",
          2842 => x"567487e7",
          2843 => x"268a3874",
          2844 => x"527587e8",
          2845 => x"29519039",
          2846 => x"87e85274",
          2847 => x"51efaf3f",
          2848 => x"82d6d808",
          2849 => x"527551ef",
          2850 => x"a53f82d6",
          2851 => x"d8085479",
          2852 => x"53755282",
          2853 => x"b68051ff",
          2854 => x"babe3f87",
          2855 => x"3d0d04ec",
          2856 => x"3d0d6602",
          2857 => x"840580e3",
          2858 => x"05335b57",
          2859 => x"80687830",
          2860 => x"707a0773",
          2861 => x"25515759",
          2862 => x"59785677",
          2863 => x"87ff2683",
          2864 => x"38815674",
          2865 => x"76077081",
          2866 => x"ff065155",
          2867 => x"93567481",
          2868 => x"82388153",
          2869 => x"76528c3d",
          2870 => x"70525681",
          2871 => x"92cf3f82",
          2872 => x"d6d80857",
          2873 => x"82d6d808",
          2874 => x"b93882d6",
          2875 => x"d80887c0",
          2876 => x"98880c82",
          2877 => x"d6d80859",
          2878 => x"963dd405",
          2879 => x"54848053",
          2880 => x"77527551",
          2881 => x"81978b3f",
          2882 => x"82d6d808",
          2883 => x"5782d6d8",
          2884 => x"0890387a",
          2885 => x"5574802e",
          2886 => x"89387419",
          2887 => x"75195959",
          2888 => x"d739963d",
          2889 => x"d8055181",
          2890 => x"9f823f76",
          2891 => x"30707807",
          2892 => x"80257b30",
          2893 => x"709f2a72",
          2894 => x"06515751",
          2895 => x"5674802e",
          2896 => x"903882b6",
          2897 => x"a45387c0",
          2898 => x"98880852",
          2899 => x"7851fe92",
          2900 => x"3f765675",
          2901 => x"82d6d80c",
          2902 => x"963d0d04",
          2903 => x"f73d0d7d",
          2904 => x"028405bb",
          2905 => x"0533595a",
          2906 => x"ff598053",
          2907 => x"7c527b51",
          2908 => x"fead3f82",
          2909 => x"d6d80880",
          2910 => x"cb387780",
          2911 => x"2e883877",
          2912 => x"812ebf38",
          2913 => x"bf3982f2",
          2914 => x"b85782f2",
          2915 => x"b85682f2",
          2916 => x"b85582f2",
          2917 => x"c0085482",
          2918 => x"f2bc0853",
          2919 => x"82f2b808",
          2920 => x"5282b6ac",
          2921 => x"51ffb8b0",
          2922 => x"3f82f2b8",
          2923 => x"56625561",
          2924 => x"5482d6d8",
          2925 => x"5360527f",
          2926 => x"51792d82",
          2927 => x"d6d80859",
          2928 => x"83397904",
          2929 => x"7882d6d8",
          2930 => x"0c8b3d0d",
          2931 => x"04f33d0d",
          2932 => x"7f616302",
          2933 => x"8c0580cf",
          2934 => x"05337373",
          2935 => x"1568415f",
          2936 => x"5c5c5e5e",
          2937 => x"5e7a5282",
          2938 => x"b6e051ff",
          2939 => x"b7ea3f82",
          2940 => x"b6e851ff",
          2941 => x"b7e23f80",
          2942 => x"55747927",
          2943 => x"8180387b",
          2944 => x"902e8938",
          2945 => x"7ba02ea7",
          2946 => x"3880c639",
          2947 => x"74185372",
          2948 => x"7a278e38",
          2949 => x"72225282",
          2950 => x"b6ec51ff",
          2951 => x"b7ba3f89",
          2952 => x"3982b6f8",
          2953 => x"51ffb7b0",
          2954 => x"3f821555",
          2955 => x"80c33974",
          2956 => x"1853727a",
          2957 => x"278e3872",
          2958 => x"085282b6",
          2959 => x"e051ffb7",
          2960 => x"973f8939",
          2961 => x"82b6f451",
          2962 => x"ffb78d3f",
          2963 => x"841555a1",
          2964 => x"39741853",
          2965 => x"727a278e",
          2966 => x"38723352",
          2967 => x"82b78051",
          2968 => x"ffb6f53f",
          2969 => x"893982b7",
          2970 => x"8851ffb6",
          2971 => x"eb3f8115",
          2972 => x"5582f2bc",
          2973 => x"0852a051",
          2974 => x"d6b83ffe",
          2975 => x"fc3982b7",
          2976 => x"8c51ffb6",
          2977 => x"d33f8055",
          2978 => x"74792780",
          2979 => x"c6387418",
          2980 => x"70335553",
          2981 => x"8056727a",
          2982 => x"27833881",
          2983 => x"5680539f",
          2984 => x"74278338",
          2985 => x"81537573",
          2986 => x"067081ff",
          2987 => x"06515372",
          2988 => x"802e9038",
          2989 => x"7380fe26",
          2990 => x"8a3882f2",
          2991 => x"bc085273",
          2992 => x"51883982",
          2993 => x"f2bc0852",
          2994 => x"a051d5e6",
          2995 => x"3f811555",
          2996 => x"ffb63982",
          2997 => x"b79051d2",
          2998 => x"8a3f7818",
          2999 => x"791c5c58",
          3000 => x"9ce73f82",
          3001 => x"d6d80898",
          3002 => x"2b70982c",
          3003 => x"515776a0",
          3004 => x"2e098106",
          3005 => x"aa389cd1",
          3006 => x"3f82d6d8",
          3007 => x"08982b70",
          3008 => x"982c70a0",
          3009 => x"32703072",
          3010 => x"9b327030",
          3011 => x"70720773",
          3012 => x"75070651",
          3013 => x"58585957",
          3014 => x"51578073",
          3015 => x"24d83876",
          3016 => x"9b2e0981",
          3017 => x"06853880",
          3018 => x"538c397c",
          3019 => x"1e537278",
          3020 => x"26fdb238",
          3021 => x"ff537282",
          3022 => x"d6d80c8f",
          3023 => x"3d0d04fc",
          3024 => x"3d0d029b",
          3025 => x"053382b7",
          3026 => x"945382b7",
          3027 => x"985255ff",
          3028 => x"b5863f82",
          3029 => x"d4a42251",
          3030 => x"a5c03f82",
          3031 => x"b7a45482",
          3032 => x"b7b05382",
          3033 => x"d4a53352",
          3034 => x"82b7b851",
          3035 => x"ffb4e93f",
          3036 => x"74802e84",
          3037 => x"38a0f43f",
          3038 => x"863d0d04",
          3039 => x"fe3d0d87",
          3040 => x"c0968008",
          3041 => x"53a5dc3f",
          3042 => x"815199bd",
          3043 => x"3f82b7d4",
          3044 => x"5199ce3f",
          3045 => x"805199b1",
          3046 => x"3f72812a",
          3047 => x"70810651",
          3048 => x"5271802e",
          3049 => x"92388151",
          3050 => x"999f3f82",
          3051 => x"b7ec5199",
          3052 => x"b03f8051",
          3053 => x"99933f72",
          3054 => x"822a7081",
          3055 => x"06515271",
          3056 => x"802e9238",
          3057 => x"81519981",
          3058 => x"3f82b7fc",
          3059 => x"5199923f",
          3060 => x"805198f5",
          3061 => x"3f72832a",
          3062 => x"70810651",
          3063 => x"5271802e",
          3064 => x"92388151",
          3065 => x"98e33f82",
          3066 => x"b88c5198",
          3067 => x"f43f8051",
          3068 => x"98d73f72",
          3069 => x"842a7081",
          3070 => x"06515271",
          3071 => x"802e9238",
          3072 => x"815198c5",
          3073 => x"3f82b8a0",
          3074 => x"5198d63f",
          3075 => x"805198b9",
          3076 => x"3f72852a",
          3077 => x"70810651",
          3078 => x"5271802e",
          3079 => x"92388151",
          3080 => x"98a73f82",
          3081 => x"b8b45198",
          3082 => x"b83f8051",
          3083 => x"989b3f72",
          3084 => x"862a7081",
          3085 => x"06515271",
          3086 => x"802e9238",
          3087 => x"81519889",
          3088 => x"3f82b8c8",
          3089 => x"51989a3f",
          3090 => x"805197fd",
          3091 => x"3f72872a",
          3092 => x"70810651",
          3093 => x"5271802e",
          3094 => x"92388151",
          3095 => x"97eb3f82",
          3096 => x"b8dc5197",
          3097 => x"fc3f8051",
          3098 => x"97df3f72",
          3099 => x"882a7081",
          3100 => x"06515271",
          3101 => x"802e9238",
          3102 => x"815197cd",
          3103 => x"3f82b8f0",
          3104 => x"5197de3f",
          3105 => x"805197c1",
          3106 => x"3fa3e03f",
          3107 => x"843d0d04",
          3108 => x"fb3d0d77",
          3109 => x"028405a3",
          3110 => x"05337055",
          3111 => x"56568052",
          3112 => x"7551e2ed",
          3113 => x"3f0b0b82",
          3114 => x"d0c83354",
          3115 => x"73a93881",
          3116 => x"5382b9ac",
          3117 => x"5282ede8",
          3118 => x"51818af1",
          3119 => x"3f82d6d8",
          3120 => x"08307082",
          3121 => x"d6d80807",
          3122 => x"80258271",
          3123 => x"31515154",
          3124 => x"730b0b82",
          3125 => x"d0c8340b",
          3126 => x"0b82d0c8",
          3127 => x"33547381",
          3128 => x"2e098106",
          3129 => x"af3882ed",
          3130 => x"e8537452",
          3131 => x"755181c5",
          3132 => x"c13f82d6",
          3133 => x"d808802e",
          3134 => x"8b3882d6",
          3135 => x"d80851cd",
          3136 => x"e23f9139",
          3137 => x"82ede851",
          3138 => x"8197a13f",
          3139 => x"820b0b0b",
          3140 => x"82d0c834",
          3141 => x"0b0b82d0",
          3142 => x"c8335473",
          3143 => x"822e0981",
          3144 => x"068c3882",
          3145 => x"b9bc5374",
          3146 => x"527551a9",
          3147 => x"d83f800b",
          3148 => x"82d6d80c",
          3149 => x"873d0d04",
          3150 => x"cd3d0d80",
          3151 => x"70415eff",
          3152 => x"7e82ede4",
          3153 => x"0c5f8152",
          3154 => x"7d5180c8",
          3155 => x"883f82d6",
          3156 => x"d80881ff",
          3157 => x"0659787e",
          3158 => x"2e098106",
          3159 => x"a338973d",
          3160 => x"59835382",
          3161 => x"b9c45278",
          3162 => x"51dafa3f",
          3163 => x"7d537852",
          3164 => x"82d88451",
          3165 => x"8188d53f",
          3166 => x"82d6d808",
          3167 => x"7e2e8838",
          3168 => x"82b9c851",
          3169 => x"8ddf3981",
          3170 => x"70415e82",
          3171 => x"ba8051ff",
          3172 => x"b0c63f97",
          3173 => x"3d70475a",
          3174 => x"80f85279",
          3175 => x"51fdf13f",
          3176 => x"b53dff84",
          3177 => x"0551f3a0",
          3178 => x"3f82d6d8",
          3179 => x"08902b70",
          3180 => x"902c5159",
          3181 => x"7880c22e",
          3182 => x"87a33878",
          3183 => x"80c224b2",
          3184 => x"3878bd2e",
          3185 => x"81d23878",
          3186 => x"bd249038",
          3187 => x"78802eff",
          3188 => x"ba3878bc",
          3189 => x"2e80da38",
          3190 => x"8ad63978",
          3191 => x"80c02e83",
          3192 => x"99387880",
          3193 => x"c02485cd",
          3194 => x"3878bf2e",
          3195 => x"828c388a",
          3196 => x"bf397880",
          3197 => x"f92e89db",
          3198 => x"387880f9",
          3199 => x"24923878",
          3200 => x"80c32e88",
          3201 => x"8a387880",
          3202 => x"f82e89a3",
          3203 => x"388aa139",
          3204 => x"7881832e",
          3205 => x"8a883878",
          3206 => x"8183248b",
          3207 => x"38788182",
          3208 => x"2e89ed38",
          3209 => x"8a8a3978",
          3210 => x"81852e89",
          3211 => x"fd388a80",
          3212 => x"39b53dff",
          3213 => x"801153ff",
          3214 => x"840551ec",
          3215 => x"ba3f82d6",
          3216 => x"d808802e",
          3217 => x"fec538b5",
          3218 => x"3dfefc11",
          3219 => x"53ff8405",
          3220 => x"51eca43f",
          3221 => x"82d6d808",
          3222 => x"802efeaf",
          3223 => x"38b53dfe",
          3224 => x"f81153ff",
          3225 => x"840551ec",
          3226 => x"8e3f82d6",
          3227 => x"d8088638",
          3228 => x"82d6d808",
          3229 => x"4382ba84",
          3230 => x"51ffaedc",
          3231 => x"3f64645c",
          3232 => x"5a797b27",
          3233 => x"81ec3862",
          3234 => x"59787a70",
          3235 => x"84055c0c",
          3236 => x"7a7a26f5",
          3237 => x"3881db39",
          3238 => x"b53dff80",
          3239 => x"1153ff84",
          3240 => x"0551ebd3",
          3241 => x"3f82d6d8",
          3242 => x"08802efd",
          3243 => x"de38b53d",
          3244 => x"fefc1153",
          3245 => x"ff840551",
          3246 => x"ebbd3f82",
          3247 => x"d6d80880",
          3248 => x"2efdc838",
          3249 => x"b53dfef8",
          3250 => x"1153ff84",
          3251 => x"0551eba7",
          3252 => x"3f82d6d8",
          3253 => x"08802efd",
          3254 => x"b23882ba",
          3255 => x"9451ffad",
          3256 => x"f73f645a",
          3257 => x"79642781",
          3258 => x"89386259",
          3259 => x"79708105",
          3260 => x"5b337934",
          3261 => x"62810543",
          3262 => x"eb39b53d",
          3263 => x"ff801153",
          3264 => x"ff840551",
          3265 => x"eaf13f82",
          3266 => x"d6d80880",
          3267 => x"2efcfc38",
          3268 => x"b53dfefc",
          3269 => x"1153ff84",
          3270 => x"0551eadb",
          3271 => x"3f82d6d8",
          3272 => x"08802efc",
          3273 => x"e638b53d",
          3274 => x"fef81153",
          3275 => x"ff840551",
          3276 => x"eac53f82",
          3277 => x"d6d80880",
          3278 => x"2efcd038",
          3279 => x"82baa051",
          3280 => x"ffad953f",
          3281 => x"645a7964",
          3282 => x"27a83862",
          3283 => x"70337b33",
          3284 => x"5e5a5b78",
          3285 => x"7c2e9238",
          3286 => x"78557a54",
          3287 => x"79335379",
          3288 => x"5282bab0",
          3289 => x"51ffacf0",
          3290 => x"3f811a63",
          3291 => x"8105445a",
          3292 => x"d5398a51",
          3293 => x"cc8f3ffc",
          3294 => x"9239b53d",
          3295 => x"ff801153",
          3296 => x"ff840551",
          3297 => x"e9f13f82",
          3298 => x"d6d80880",
          3299 => x"df3882d4",
          3300 => x"b8335978",
          3301 => x"802e8938",
          3302 => x"82d3f008",
          3303 => x"4580cd39",
          3304 => x"82d4b933",
          3305 => x"5978802e",
          3306 => x"883882d3",
          3307 => x"f80845bc",
          3308 => x"3982d4ba",
          3309 => x"33597880",
          3310 => x"2e883882",
          3311 => x"d4800845",
          3312 => x"ab3982d4",
          3313 => x"bb335978",
          3314 => x"802e8838",
          3315 => x"82d48808",
          3316 => x"459a3982",
          3317 => x"d4b63359",
          3318 => x"78802e88",
          3319 => x"3882d490",
          3320 => x"08458939",
          3321 => x"82d4a008",
          3322 => x"fc800545",
          3323 => x"b53dfefc",
          3324 => x"1153ff84",
          3325 => x"0551e8ff",
          3326 => x"3f82d6d8",
          3327 => x"0880de38",
          3328 => x"82d4b833",
          3329 => x"5978802e",
          3330 => x"893882d3",
          3331 => x"f4084480",
          3332 => x"cc3982d4",
          3333 => x"b9335978",
          3334 => x"802e8838",
          3335 => x"82d3fc08",
          3336 => x"44bb3982",
          3337 => x"d4ba3359",
          3338 => x"78802e88",
          3339 => x"3882d484",
          3340 => x"0844aa39",
          3341 => x"82d4bb33",
          3342 => x"5978802e",
          3343 => x"883882d4",
          3344 => x"8c084499",
          3345 => x"3982d4b6",
          3346 => x"33597880",
          3347 => x"2e883882",
          3348 => x"d4940844",
          3349 => x"883982d4",
          3350 => x"a0088805",
          3351 => x"44b53dfe",
          3352 => x"f81153ff",
          3353 => x"840551e8",
          3354 => x"8e3f82d6",
          3355 => x"d808802e",
          3356 => x"a7388063",
          3357 => x"5c5c7a88",
          3358 => x"2e833881",
          3359 => x"5c7a9032",
          3360 => x"70307072",
          3361 => x"079f2a70",
          3362 => x"7f065151",
          3363 => x"5a5a7880",
          3364 => x"2e88387a",
          3365 => x"a02e8338",
          3366 => x"884382ba",
          3367 => x"cc51c6c3",
          3368 => x"3fa05564",
          3369 => x"54625363",
          3370 => x"526451f2",
          3371 => x"a03f82ba",
          3372 => x"d85187b1",
          3373 => x"39b53dff",
          3374 => x"801153ff",
          3375 => x"840551e7",
          3376 => x"b63f82d6",
          3377 => x"d808802e",
          3378 => x"f9c138b5",
          3379 => x"3dfefc11",
          3380 => x"53ff8405",
          3381 => x"51e7a03f",
          3382 => x"82d6d808",
          3383 => x"802ea438",
          3384 => x"64590280",
          3385 => x"cf053379",
          3386 => x"34648105",
          3387 => x"45b53dfe",
          3388 => x"fc1153ff",
          3389 => x"840551e6",
          3390 => x"fe3f82d6",
          3391 => x"d808e138",
          3392 => x"f9893964",
          3393 => x"70335452",
          3394 => x"82bae451",
          3395 => x"ffa9c93f",
          3396 => x"82f2b808",
          3397 => x"5380f852",
          3398 => x"7951ffaa",
          3399 => x"903f7946",
          3400 => x"79335978",
          3401 => x"ae2ef8e3",
          3402 => x"389f7927",
          3403 => x"9f38b53d",
          3404 => x"fefc1153",
          3405 => x"ff840551",
          3406 => x"e6bd3f82",
          3407 => x"d6d80880",
          3408 => x"2e913864",
          3409 => x"590280cf",
          3410 => x"05337934",
          3411 => x"64810545",
          3412 => x"ffb13982",
          3413 => x"baf051c5",
          3414 => x"8a3fffa7",
          3415 => x"39b53dfe",
          3416 => x"f41153ff",
          3417 => x"840551e0",
          3418 => x"bd3f82d6",
          3419 => x"d808802e",
          3420 => x"f89938b5",
          3421 => x"3dfef011",
          3422 => x"53ff8405",
          3423 => x"51e0a73f",
          3424 => x"82d6d808",
          3425 => x"802ea638",
          3426 => x"61590280",
          3427 => x"c2052279",
          3428 => x"7082055b",
          3429 => x"237842b5",
          3430 => x"3dfef011",
          3431 => x"53ff8405",
          3432 => x"51e0833f",
          3433 => x"82d6d808",
          3434 => x"df38f7df",
          3435 => x"39617022",
          3436 => x"545282ba",
          3437 => x"f451ffa8",
          3438 => x"9f3f82f2",
          3439 => x"b8085380",
          3440 => x"f8527951",
          3441 => x"ffa8e63f",
          3442 => x"79467933",
          3443 => x"5978ae2e",
          3444 => x"f7b93878",
          3445 => x"9f268738",
          3446 => x"61820542",
          3447 => x"d039b53d",
          3448 => x"fef01153",
          3449 => x"ff840551",
          3450 => x"dfbc3f82",
          3451 => x"d6d80880",
          3452 => x"2e933861",
          3453 => x"590280c2",
          3454 => x"05227970",
          3455 => x"82055b23",
          3456 => x"7842ffa9",
          3457 => x"3982baf0",
          3458 => x"51c3d83f",
          3459 => x"ff9f39b5",
          3460 => x"3dfef411",
          3461 => x"53ff8405",
          3462 => x"51df8b3f",
          3463 => x"82d6d808",
          3464 => x"802ef6e7",
          3465 => x"38b53dfe",
          3466 => x"f01153ff",
          3467 => x"840551de",
          3468 => x"f53f82d6",
          3469 => x"d808802e",
          3470 => x"a0386161",
          3471 => x"710c5961",
          3472 => x"840542b5",
          3473 => x"3dfef011",
          3474 => x"53ff8405",
          3475 => x"51ded73f",
          3476 => x"82d6d808",
          3477 => x"e538f6b3",
          3478 => x"39617008",
          3479 => x"545282bb",
          3480 => x"8051ffa6",
          3481 => x"f33f82f2",
          3482 => x"b8085380",
          3483 => x"f8527951",
          3484 => x"ffa7ba3f",
          3485 => x"79467933",
          3486 => x"5978ae2e",
          3487 => x"f68d389f",
          3488 => x"79279b38",
          3489 => x"b53dfef0",
          3490 => x"1153ff84",
          3491 => x"0551de96",
          3492 => x"3f82d6d8",
          3493 => x"08802e8d",
          3494 => x"38616171",
          3495 => x"0c596184",
          3496 => x"0542ffb5",
          3497 => x"3982baf0",
          3498 => x"51c2b83f",
          3499 => x"ffab39b5",
          3500 => x"3dff8011",
          3501 => x"53ff8405",
          3502 => x"51e3bc3f",
          3503 => x"82d6d808",
          3504 => x"802ef5c7",
          3505 => x"38645282",
          3506 => x"bb9051ff",
          3507 => x"a68a3f64",
          3508 => x"597804b5",
          3509 => x"3dff8011",
          3510 => x"53ff8405",
          3511 => x"51e3983f",
          3512 => x"82d6d808",
          3513 => x"802ef5a3",
          3514 => x"38645282",
          3515 => x"bbac51ff",
          3516 => x"a5e63f64",
          3517 => x"59782d82",
          3518 => x"d6d80880",
          3519 => x"2ef58c38",
          3520 => x"82d6d808",
          3521 => x"5282bbc8",
          3522 => x"51ffa5cc",
          3523 => x"3ff4fc39",
          3524 => x"82bbe451",
          3525 => x"c1cd3fff",
          3526 => x"a59f3ff4",
          3527 => x"ee3982bc",
          3528 => x"8051c1bf",
          3529 => x"3f8059ff",
          3530 => x"a83991bf",
          3531 => x"3ff4dc39",
          3532 => x"973d3359",
          3533 => x"78802ef4",
          3534 => x"d23880f8",
          3535 => x"527951d2",
          3536 => x"f83f82d6",
          3537 => x"d8085d82",
          3538 => x"d6d80880",
          3539 => x"2e829238",
          3540 => x"82d6d808",
          3541 => x"46b53dff",
          3542 => x"84055184",
          3543 => x"e53f82d6",
          3544 => x"d808607f",
          3545 => x"065a5c78",
          3546 => x"802e81d2",
          3547 => x"3882d6d8",
          3548 => x"0851cd91",
          3549 => x"3f82d6d8",
          3550 => x"088f2681",
          3551 => x"c138815b",
          3552 => x"7a822eb2",
          3553 => x"387a8224",
          3554 => x"89387a81",
          3555 => x"2e8c3880",
          3556 => x"ca397a83",
          3557 => x"2ead3880",
          3558 => x"c23982bc",
          3559 => x"94567b55",
          3560 => x"82bc9854",
          3561 => x"805382bc",
          3562 => x"9c52b53d",
          3563 => x"ffb00551",
          3564 => x"ffa78d3f",
          3565 => x"b8397b52",
          3566 => x"b53dffb0",
          3567 => x"0551cdb3",
          3568 => x"3fab397b",
          3569 => x"5582bc98",
          3570 => x"54805382",
          3571 => x"bcac52b5",
          3572 => x"3dffb005",
          3573 => x"51ffa6e8",
          3574 => x"3f93397b",
          3575 => x"54805382",
          3576 => x"bcb852b5",
          3577 => x"3dffb005",
          3578 => x"51ffa6d4",
          3579 => x"3f82d3f0",
          3580 => x"5882d788",
          3581 => x"577c5665",
          3582 => x"55805484",
          3583 => x"80805384",
          3584 => x"808052b5",
          3585 => x"3dffb005",
          3586 => x"51ead13f",
          3587 => x"82d6d808",
          3588 => x"82d6d808",
          3589 => x"09703070",
          3590 => x"72078025",
          3591 => x"515b5b5f",
          3592 => x"805a7a83",
          3593 => x"26833881",
          3594 => x"5a787a06",
          3595 => x"5978802e",
          3596 => x"8d38811b",
          3597 => x"7081ff06",
          3598 => x"5c597afe",
          3599 => x"c3387f81",
          3600 => x"327e8132",
          3601 => x"07597889",
          3602 => x"387eff2e",
          3603 => x"09810689",
          3604 => x"3882bcc0",
          3605 => x"51ffbf8b",
          3606 => x"3f7c51b1",
          3607 => x"f53ff2ab",
          3608 => x"3982bcd0",
          3609 => x"51ffbefb",
          3610 => x"3ff2a039",
          3611 => x"f63d0d80",
          3612 => x"0b82d788",
          3613 => x"3487c094",
          3614 => x"8c085387",
          3615 => x"84805272",
          3616 => x"51d7ab3f",
          3617 => x"82d6d808",
          3618 => x"902b87c0",
          3619 => x"948c0855",
          3620 => x"53878480",
          3621 => x"527351d7",
          3622 => x"953f7282",
          3623 => x"d6d80807",
          3624 => x"87c0948c",
          3625 => x"0c87c094",
          3626 => x"9c085387",
          3627 => x"84805272",
          3628 => x"51d6fb3f",
          3629 => x"82d6d808",
          3630 => x"902b87c0",
          3631 => x"949c0855",
          3632 => x"53878480",
          3633 => x"527351d6",
          3634 => x"e53f7282",
          3635 => x"d6d80807",
          3636 => x"87c0949c",
          3637 => x"0c8c8083",
          3638 => x"0b87c094",
          3639 => x"840c8c80",
          3640 => x"830b87c0",
          3641 => x"94940c87",
          3642 => x"a0a08053",
          3643 => x"80737084",
          3644 => x"05550c87",
          3645 => x"a0affe73",
          3646 => x"27f23887",
          3647 => x"a0b08053",
          3648 => x"878bc5e2",
          3649 => x"f1737084",
          3650 => x"05550c87",
          3651 => x"a0bffe73",
          3652 => x"27ee3880",
          3653 => x"5280c851",
          3654 => x"a79e3f80",
          3655 => x"5280c551",
          3656 => x"a7963f80",
          3657 => x"5280cc51",
          3658 => x"a78e3f80",
          3659 => x"5280cc51",
          3660 => x"a7863f80",
          3661 => x"5280cf51",
          3662 => x"a6fe3f80",
          3663 => x"528a51a6",
          3664 => x"f73f8052",
          3665 => x"be51a6f0",
          3666 => x"3f8199b8",
          3667 => x"59819aca",
          3668 => x"5a830284",
          3669 => x"05950534",
          3670 => x"805b853d",
          3671 => x"7082f2c0",
          3672 => x"0c7082f2",
          3673 => x"b80c82f2",
          3674 => x"bc0c82bc",
          3675 => x"fc51ffbc",
          3676 => x"f23f88ab",
          3677 => x"3f91ec3f",
          3678 => x"82bd8c51",
          3679 => x"ffbce43f",
          3680 => x"82bd9851",
          3681 => x"ffbcdc3f",
          3682 => x"80defc51",
          3683 => x"91d03f81",
          3684 => x"51ebac3f",
          3685 => x"efa23f80",
          3686 => x"04fe3d0d",
          3687 => x"80528353",
          3688 => x"71882b52",
          3689 => x"86d43f82",
          3690 => x"d6d80881",
          3691 => x"ff067207",
          3692 => x"ff145452",
          3693 => x"728025e8",
          3694 => x"387182d6",
          3695 => x"d80c843d",
          3696 => x"0d04fc3d",
          3697 => x"0d767008",
          3698 => x"54558073",
          3699 => x"52547274",
          3700 => x"2e818a38",
          3701 => x"72335170",
          3702 => x"a02e0981",
          3703 => x"06863881",
          3704 => x"1353f139",
          3705 => x"72335170",
          3706 => x"a22e0981",
          3707 => x"06863881",
          3708 => x"13538154",
          3709 => x"72527381",
          3710 => x"2e098106",
          3711 => x"9f388439",
          3712 => x"81125280",
          3713 => x"72335254",
          3714 => x"70a22e83",
          3715 => x"38815470",
          3716 => x"802e9d38",
          3717 => x"73ea3898",
          3718 => x"39811252",
          3719 => x"80723352",
          3720 => x"5470a02e",
          3721 => x"83388154",
          3722 => x"70802e84",
          3723 => x"3873ea38",
          3724 => x"80723352",
          3725 => x"5470a02e",
          3726 => x"09810683",
          3727 => x"38815470",
          3728 => x"a2327030",
          3729 => x"70802576",
          3730 => x"07515151",
          3731 => x"70802e88",
          3732 => x"38807270",
          3733 => x"81055434",
          3734 => x"71750c72",
          3735 => x"517082d6",
          3736 => x"d80c863d",
          3737 => x"0d04fc3d",
          3738 => x"0d765372",
          3739 => x"08802e91",
          3740 => x"38863dfc",
          3741 => x"05527251",
          3742 => x"d6ac3f82",
          3743 => x"d6d80885",
          3744 => x"38805383",
          3745 => x"39745372",
          3746 => x"82d6d80c",
          3747 => x"863d0d04",
          3748 => x"fc3d0d76",
          3749 => x"821133ff",
          3750 => x"05525381",
          3751 => x"52708b26",
          3752 => x"81983883",
          3753 => x"1333ff05",
          3754 => x"51825270",
          3755 => x"9e26818a",
          3756 => x"38841333",
          3757 => x"51835270",
          3758 => x"972680fe",
          3759 => x"38851333",
          3760 => x"51845270",
          3761 => x"bb2680f2",
          3762 => x"38861333",
          3763 => x"51855270",
          3764 => x"bb2680e6",
          3765 => x"38881322",
          3766 => x"55865274",
          3767 => x"87e72680",
          3768 => x"d9388a13",
          3769 => x"22548752",
          3770 => x"7387e726",
          3771 => x"80cc3881",
          3772 => x"0b87c098",
          3773 => x"9c0c7222",
          3774 => x"87c098bc",
          3775 => x"0c821333",
          3776 => x"87c098b8",
          3777 => x"0c831333",
          3778 => x"87c098b4",
          3779 => x"0c841333",
          3780 => x"87c098b0",
          3781 => x"0c851333",
          3782 => x"87c098ac",
          3783 => x"0c861333",
          3784 => x"87c098a8",
          3785 => x"0c7487c0",
          3786 => x"98a40c73",
          3787 => x"87c098a0",
          3788 => x"0c800b87",
          3789 => x"c0989c0c",
          3790 => x"80527182",
          3791 => x"d6d80c86",
          3792 => x"3d0d04f3",
          3793 => x"3d0d7f5b",
          3794 => x"87c0989c",
          3795 => x"5d817d0c",
          3796 => x"87c098bc",
          3797 => x"085e7d7b",
          3798 => x"2387c098",
          3799 => x"b8085a79",
          3800 => x"821c3487",
          3801 => x"c098b408",
          3802 => x"5a79831c",
          3803 => x"3487c098",
          3804 => x"b0085a79",
          3805 => x"841c3487",
          3806 => x"c098ac08",
          3807 => x"5a79851c",
          3808 => x"3487c098",
          3809 => x"a8085a79",
          3810 => x"861c3487",
          3811 => x"c098a408",
          3812 => x"5c7b881c",
          3813 => x"2387c098",
          3814 => x"a0085a79",
          3815 => x"8a1c2380",
          3816 => x"7d0c7983",
          3817 => x"ffff0659",
          3818 => x"7b83ffff",
          3819 => x"0658861b",
          3820 => x"3357851b",
          3821 => x"3356841b",
          3822 => x"3355831b",
          3823 => x"3354821b",
          3824 => x"33537d83",
          3825 => x"ffff0652",
          3826 => x"82bdb051",
          3827 => x"ff9c893f",
          3828 => x"8f3d0d04",
          3829 => x"fb3d0d02",
          3830 => x"9f053382",
          3831 => x"d3ec3370",
          3832 => x"81ff0658",
          3833 => x"555587c0",
          3834 => x"94845175",
          3835 => x"802e8638",
          3836 => x"87c09494",
          3837 => x"51700870",
          3838 => x"962a7081",
          3839 => x"06535452",
          3840 => x"70802e8c",
          3841 => x"3871912a",
          3842 => x"70810651",
          3843 => x"5170d738",
          3844 => x"72813270",
          3845 => x"81065151",
          3846 => x"70802e8d",
          3847 => x"3871932a",
          3848 => x"70810651",
          3849 => x"5170ffbe",
          3850 => x"387381ff",
          3851 => x"065187c0",
          3852 => x"94805270",
          3853 => x"802e8638",
          3854 => x"87c09490",
          3855 => x"5274720c",
          3856 => x"7482d6d8",
          3857 => x"0c873d0d",
          3858 => x"04ff3d0d",
          3859 => x"028f0533",
          3860 => x"7030709f",
          3861 => x"2a515252",
          3862 => x"7082d3ec",
          3863 => x"34833d0d",
          3864 => x"04f93d0d",
          3865 => x"79548074",
          3866 => x"337081ff",
          3867 => x"06535357",
          3868 => x"70772e80",
          3869 => x"fc387181",
          3870 => x"ff068115",
          3871 => x"82d3ec33",
          3872 => x"7081ff06",
          3873 => x"59575558",
          3874 => x"87c09484",
          3875 => x"5175802e",
          3876 => x"863887c0",
          3877 => x"94945170",
          3878 => x"0870962a",
          3879 => x"70810653",
          3880 => x"54527080",
          3881 => x"2e8c3871",
          3882 => x"912a7081",
          3883 => x"06515170",
          3884 => x"d7387281",
          3885 => x"32708106",
          3886 => x"51517080",
          3887 => x"2e8d3871",
          3888 => x"932a7081",
          3889 => x"06515170",
          3890 => x"ffbe3874",
          3891 => x"81ff0651",
          3892 => x"87c09480",
          3893 => x"5270802e",
          3894 => x"863887c0",
          3895 => x"94905277",
          3896 => x"720c8117",
          3897 => x"74337081",
          3898 => x"ff065353",
          3899 => x"5770ff86",
          3900 => x"387682d6",
          3901 => x"d80c893d",
          3902 => x"0d04fe3d",
          3903 => x"0d82d3ec",
          3904 => x"337081ff",
          3905 => x"06545287",
          3906 => x"c0948451",
          3907 => x"72802e86",
          3908 => x"3887c094",
          3909 => x"94517008",
          3910 => x"70822a70",
          3911 => x"81065151",
          3912 => x"5170802e",
          3913 => x"e2387181",
          3914 => x"ff065187",
          3915 => x"c0948052",
          3916 => x"70802e86",
          3917 => x"3887c094",
          3918 => x"90527108",
          3919 => x"7081ff06",
          3920 => x"82d6d80c",
          3921 => x"51843d0d",
          3922 => x"04fe3d0d",
          3923 => x"82d3ec33",
          3924 => x"7081ff06",
          3925 => x"525387c0",
          3926 => x"94845270",
          3927 => x"802e8638",
          3928 => x"87c09494",
          3929 => x"52710870",
          3930 => x"822a7081",
          3931 => x"06515151",
          3932 => x"ff527080",
          3933 => x"2ea03872",
          3934 => x"81ff0651",
          3935 => x"87c09480",
          3936 => x"5270802e",
          3937 => x"863887c0",
          3938 => x"94905271",
          3939 => x"0870982b",
          3940 => x"70982c51",
          3941 => x"53517182",
          3942 => x"d6d80c84",
          3943 => x"3d0d04ff",
          3944 => x"3d0d87c0",
          3945 => x"9e800870",
          3946 => x"9c2a8a06",
          3947 => x"51517080",
          3948 => x"2e84b438",
          3949 => x"87c09ea4",
          3950 => x"0882d3f0",
          3951 => x"0c87c09e",
          3952 => x"a80882d3",
          3953 => x"f40c87c0",
          3954 => x"9e940882",
          3955 => x"d3f80c87",
          3956 => x"c09e9808",
          3957 => x"82d3fc0c",
          3958 => x"87c09e9c",
          3959 => x"0882d480",
          3960 => x"0c87c09e",
          3961 => x"a00882d4",
          3962 => x"840c87c0",
          3963 => x"9eac0882",
          3964 => x"d4880c87",
          3965 => x"c09eb008",
          3966 => x"82d48c0c",
          3967 => x"87c09eb4",
          3968 => x"0882d490",
          3969 => x"0c87c09e",
          3970 => x"b80882d4",
          3971 => x"940c87c0",
          3972 => x"9ebc0882",
          3973 => x"d4980c87",
          3974 => x"c09ec008",
          3975 => x"82d49c0c",
          3976 => x"87c09ec4",
          3977 => x"0882d4a0",
          3978 => x"0c87c09e",
          3979 => x"80085170",
          3980 => x"82d4a423",
          3981 => x"87c09e84",
          3982 => x"0882d4a8",
          3983 => x"0c87c09e",
          3984 => x"880882d4",
          3985 => x"ac0c87c0",
          3986 => x"9e8c0882",
          3987 => x"d4b00c81",
          3988 => x"0b82d4b4",
          3989 => x"34800b87",
          3990 => x"c09e9008",
          3991 => x"7084800a",
          3992 => x"06515252",
          3993 => x"70802e83",
          3994 => x"38815271",
          3995 => x"82d4b534",
          3996 => x"800b87c0",
          3997 => x"9e900870",
          3998 => x"88800a06",
          3999 => x"51525270",
          4000 => x"802e8338",
          4001 => x"81527182",
          4002 => x"d4b63480",
          4003 => x"0b87c09e",
          4004 => x"90087090",
          4005 => x"800a0651",
          4006 => x"52527080",
          4007 => x"2e833881",
          4008 => x"527182d4",
          4009 => x"b734800b",
          4010 => x"87c09e90",
          4011 => x"08708880",
          4012 => x"80065152",
          4013 => x"5270802e",
          4014 => x"83388152",
          4015 => x"7182d4b8",
          4016 => x"34800b87",
          4017 => x"c09e9008",
          4018 => x"70a08080",
          4019 => x"06515252",
          4020 => x"70802e83",
          4021 => x"38815271",
          4022 => x"82d4b934",
          4023 => x"800b87c0",
          4024 => x"9e900870",
          4025 => x"90808006",
          4026 => x"51525270",
          4027 => x"802e8338",
          4028 => x"81527182",
          4029 => x"d4ba3480",
          4030 => x"0b87c09e",
          4031 => x"90087084",
          4032 => x"80800651",
          4033 => x"52527080",
          4034 => x"2e833881",
          4035 => x"527182d4",
          4036 => x"bb34800b",
          4037 => x"87c09e90",
          4038 => x"08708280",
          4039 => x"80065152",
          4040 => x"5270802e",
          4041 => x"83388152",
          4042 => x"7182d4bc",
          4043 => x"34800b87",
          4044 => x"c09e9008",
          4045 => x"70818080",
          4046 => x"06515252",
          4047 => x"70802e83",
          4048 => x"38815271",
          4049 => x"82d4bd34",
          4050 => x"800b87c0",
          4051 => x"9e900870",
          4052 => x"80c08006",
          4053 => x"51525270",
          4054 => x"802e8338",
          4055 => x"81527182",
          4056 => x"d4be3480",
          4057 => x"0b87c09e",
          4058 => x"900870a0",
          4059 => x"80065152",
          4060 => x"5270802e",
          4061 => x"83388152",
          4062 => x"7182d4bf",
          4063 => x"3487c09e",
          4064 => x"90087098",
          4065 => x"8006708a",
          4066 => x"2a515151",
          4067 => x"7082d4c0",
          4068 => x"34800b87",
          4069 => x"c09e9008",
          4070 => x"70848006",
          4071 => x"51525270",
          4072 => x"802e8338",
          4073 => x"81527182",
          4074 => x"d4c13487",
          4075 => x"c09e9008",
          4076 => x"7083f006",
          4077 => x"70842a51",
          4078 => x"51517082",
          4079 => x"d4c23480",
          4080 => x"0b87c09e",
          4081 => x"90087088",
          4082 => x"06515252",
          4083 => x"70802e83",
          4084 => x"38815271",
          4085 => x"82d4c334",
          4086 => x"87c09e90",
          4087 => x"08708706",
          4088 => x"51517082",
          4089 => x"d4c43483",
          4090 => x"3d0d04fb",
          4091 => x"3d0d82bd",
          4092 => x"c851ff93",
          4093 => x"e33f82d4",
          4094 => x"b4335473",
          4095 => x"802e8938",
          4096 => x"82bddc51",
          4097 => x"ff93d13f",
          4098 => x"82bdf051",
          4099 => x"ffafd43f",
          4100 => x"82d4b633",
          4101 => x"5473802e",
          4102 => x"943882d4",
          4103 => x"900882d4",
          4104 => x"94081154",
          4105 => x"5282be88",
          4106 => x"51ff93ac",
          4107 => x"3f82d4bb",
          4108 => x"33547380",
          4109 => x"2e943882",
          4110 => x"d4880882",
          4111 => x"d48c0811",
          4112 => x"545282be",
          4113 => x"a451ff93",
          4114 => x"8f3f82d4",
          4115 => x"b8335473",
          4116 => x"802e9438",
          4117 => x"82d3f008",
          4118 => x"82d3f408",
          4119 => x"11545282",
          4120 => x"bec051ff",
          4121 => x"92f23f82",
          4122 => x"d4b93354",
          4123 => x"73802e94",
          4124 => x"3882d3f8",
          4125 => x"0882d3fc",
          4126 => x"08115452",
          4127 => x"82bedc51",
          4128 => x"ff92d53f",
          4129 => x"82d4ba33",
          4130 => x"5473802e",
          4131 => x"943882d4",
          4132 => x"800882d4",
          4133 => x"84081154",
          4134 => x"5282bef8",
          4135 => x"51ff92b8",
          4136 => x"3f82d4bf",
          4137 => x"33547380",
          4138 => x"2e8e3882",
          4139 => x"d4c03352",
          4140 => x"82bf9451",
          4141 => x"ff92a13f",
          4142 => x"82d4c333",
          4143 => x"5473802e",
          4144 => x"8e3882d4",
          4145 => x"c4335282",
          4146 => x"bfb451ff",
          4147 => x"928a3f82",
          4148 => x"d4c13354",
          4149 => x"73802e8e",
          4150 => x"3882d4c2",
          4151 => x"335282bf",
          4152 => x"d451ff91",
          4153 => x"f33f82d4",
          4154 => x"b5335473",
          4155 => x"802e8938",
          4156 => x"82bff451",
          4157 => x"ffadec3f",
          4158 => x"82d4b733",
          4159 => x"5473802e",
          4160 => x"893882c0",
          4161 => x"8851ffad",
          4162 => x"da3f82d4",
          4163 => x"bc335473",
          4164 => x"802e8938",
          4165 => x"82c09451",
          4166 => x"ffadc83f",
          4167 => x"82d4bd33",
          4168 => x"5473802e",
          4169 => x"893882c0",
          4170 => x"a051ffad",
          4171 => x"b63f82d4",
          4172 => x"be335473",
          4173 => x"802e8938",
          4174 => x"82c0a851",
          4175 => x"ffada43f",
          4176 => x"82c0b051",
          4177 => x"ffad9c3f",
          4178 => x"82d49808",
          4179 => x"5282c0bc",
          4180 => x"51ff9184",
          4181 => x"3f82d49c",
          4182 => x"085282c0",
          4183 => x"e451ff90",
          4184 => x"f73f82d4",
          4185 => x"a0085282",
          4186 => x"c18c51ff",
          4187 => x"90ea3f82",
          4188 => x"c1b451ff",
          4189 => x"aced3f82",
          4190 => x"d4a42252",
          4191 => x"82c1bc51",
          4192 => x"ff90d53f",
          4193 => x"82d4a808",
          4194 => x"56bd84c0",
          4195 => x"527551c5",
          4196 => x"9d3f82d6",
          4197 => x"d808bd84",
          4198 => x"c0297671",
          4199 => x"31545482",
          4200 => x"d6d80852",
          4201 => x"82c1e451",
          4202 => x"ff90ad3f",
          4203 => x"82d4bb33",
          4204 => x"5473802e",
          4205 => x"a93882d4",
          4206 => x"ac0856bd",
          4207 => x"84c05275",
          4208 => x"51c4eb3f",
          4209 => x"82d6d808",
          4210 => x"bd84c029",
          4211 => x"76713154",
          4212 => x"5482d6d8",
          4213 => x"085282c2",
          4214 => x"9051ff8f",
          4215 => x"fb3f82d4",
          4216 => x"b6335473",
          4217 => x"802ea938",
          4218 => x"82d4b008",
          4219 => x"56bd84c0",
          4220 => x"527551c4",
          4221 => x"b93f82d6",
          4222 => x"d808bd84",
          4223 => x"c0297671",
          4224 => x"31545482",
          4225 => x"d6d80852",
          4226 => x"82c2bc51",
          4227 => x"ff8fc93f",
          4228 => x"8a51ffae",
          4229 => x"f03f873d",
          4230 => x"0d04fe3d",
          4231 => x"0d029205",
          4232 => x"33ff0552",
          4233 => x"718426aa",
          4234 => x"38718429",
          4235 => x"82adac05",
          4236 => x"52710804",
          4237 => x"82c2e851",
          4238 => x"9d3982c2",
          4239 => x"f0519739",
          4240 => x"82c2f851",
          4241 => x"913982c3",
          4242 => x"80518b39",
          4243 => x"82c38451",
          4244 => x"853982c3",
          4245 => x"8c51ff8e",
          4246 => x"ff3f843d",
          4247 => x"0d047188",
          4248 => x"800c0480",
          4249 => x"0b87c096",
          4250 => x"840c0482",
          4251 => x"d4c80887",
          4252 => x"c096840c",
          4253 => x"04fd3d0d",
          4254 => x"76982b70",
          4255 => x"982c7998",
          4256 => x"2b70982c",
          4257 => x"72101370",
          4258 => x"822b5153",
          4259 => x"51545151",
          4260 => x"800b82c3",
          4261 => x"98123355",
          4262 => x"53717425",
          4263 => x"9c3882c3",
          4264 => x"94110812",
          4265 => x"02840597",
          4266 => x"05337133",
          4267 => x"52525270",
          4268 => x"722e0981",
          4269 => x"06833881",
          4270 => x"537282d6",
          4271 => x"d80c853d",
          4272 => x"0d04fb3d",
          4273 => x"0d790284",
          4274 => x"05a30533",
          4275 => x"71335556",
          4276 => x"5472802e",
          4277 => x"b13882f2",
          4278 => x"bc085288",
          4279 => x"51ffadd2",
          4280 => x"3f82f2bc",
          4281 => x"0852a051",
          4282 => x"ffadc73f",
          4283 => x"82f2bc08",
          4284 => x"528851ff",
          4285 => x"adbc3f73",
          4286 => x"33ff0553",
          4287 => x"72743472",
          4288 => x"81ff0653",
          4289 => x"cc397751",
          4290 => x"ff8dcd3f",
          4291 => x"74743487",
          4292 => x"3d0d04f6",
          4293 => x"3d0d7c02",
          4294 => x"8405b705",
          4295 => x"33028805",
          4296 => x"bb053382",
          4297 => x"d5a43370",
          4298 => x"842982d4",
          4299 => x"cc057008",
          4300 => x"5159595a",
          4301 => x"58597480",
          4302 => x"2e863874",
          4303 => x"519c933f",
          4304 => x"82d5a433",
          4305 => x"70842982",
          4306 => x"d4cc0581",
          4307 => x"19705458",
          4308 => x"565a9f94",
          4309 => x"3f82d6d8",
          4310 => x"08750c82",
          4311 => x"d5a43370",
          4312 => x"842982d4",
          4313 => x"cc057008",
          4314 => x"51565a74",
          4315 => x"802ea738",
          4316 => x"75537852",
          4317 => x"7451ffb6",
          4318 => x"ec3f82d5",
          4319 => x"a4338105",
          4320 => x"557482d5",
          4321 => x"a4347481",
          4322 => x"ff065593",
          4323 => x"75278738",
          4324 => x"800b82d5",
          4325 => x"a4347780",
          4326 => x"2eb63882",
          4327 => x"d5a00856",
          4328 => x"75802eac",
          4329 => x"3882d59c",
          4330 => x"335574a4",
          4331 => x"388c3dfc",
          4332 => x"05547653",
          4333 => x"78527551",
          4334 => x"80ecd73f",
          4335 => x"82d5a008",
          4336 => x"528a5181",
          4337 => x"a2803f82",
          4338 => x"d5a00851",
          4339 => x"80f0ba3f",
          4340 => x"8c3d0d04",
          4341 => x"fd3d0d82",
          4342 => x"d4cc5393",
          4343 => x"54720852",
          4344 => x"71802e89",
          4345 => x"3871519a",
          4346 => x"e93f8073",
          4347 => x"0cff1484",
          4348 => x"14545473",
          4349 => x"8025e638",
          4350 => x"800b82d5",
          4351 => x"a43482d5",
          4352 => x"a0085271",
          4353 => x"802e9538",
          4354 => x"715180f1",
          4355 => x"9f3f82d5",
          4356 => x"a008519a",
          4357 => x"bd3f800b",
          4358 => x"82d5a00c",
          4359 => x"853d0d04",
          4360 => x"dc3d0d81",
          4361 => x"57805282",
          4362 => x"d5a00851",
          4363 => x"80f6bb3f",
          4364 => x"82d6d808",
          4365 => x"80d33882",
          4366 => x"d5a00853",
          4367 => x"80f85288",
          4368 => x"3d705256",
          4369 => x"819eeb3f",
          4370 => x"82d6d808",
          4371 => x"802eba38",
          4372 => x"7551ffb3",
          4373 => x"b03f82d6",
          4374 => x"d8085580",
          4375 => x"0b82d6d8",
          4376 => x"08259d38",
          4377 => x"82d6d808",
          4378 => x"ff057017",
          4379 => x"55558074",
          4380 => x"34755376",
          4381 => x"52811782",
          4382 => x"c6885257",
          4383 => x"ff8ad93f",
          4384 => x"74ff2e09",
          4385 => x"8106ffaf",
          4386 => x"38a63d0d",
          4387 => x"04d93d0d",
          4388 => x"aa3d08ad",
          4389 => x"3d085a5a",
          4390 => x"81705858",
          4391 => x"805282d5",
          4392 => x"a0085180",
          4393 => x"f5c43f82",
          4394 => x"d6d80881",
          4395 => x"9538ff0b",
          4396 => x"82d5a008",
          4397 => x"545580f8",
          4398 => x"528b3d70",
          4399 => x"5256819d",
          4400 => x"f13f82d6",
          4401 => x"d808802e",
          4402 => x"a5387551",
          4403 => x"ffb2b63f",
          4404 => x"82d6d808",
          4405 => x"81185855",
          4406 => x"800b82d6",
          4407 => x"d808258e",
          4408 => x"3882d6d8",
          4409 => x"08ff0570",
          4410 => x"17555580",
          4411 => x"74347409",
          4412 => x"70307072",
          4413 => x"079f2a51",
          4414 => x"55557877",
          4415 => x"2e853873",
          4416 => x"ffac3882",
          4417 => x"d5a0088c",
          4418 => x"11085351",
          4419 => x"80f4db3f",
          4420 => x"82d6d808",
          4421 => x"802e8938",
          4422 => x"82c69451",
          4423 => x"ff89b93f",
          4424 => x"78772e09",
          4425 => x"81069b38",
          4426 => x"75527951",
          4427 => x"ffb2c43f",
          4428 => x"7951ffb1",
          4429 => x"d03fab3d",
          4430 => x"085482d6",
          4431 => x"d8087434",
          4432 => x"80587782",
          4433 => x"d6d80ca9",
          4434 => x"3d0d04f6",
          4435 => x"3d0d7c7e",
          4436 => x"715c7172",
          4437 => x"3357595a",
          4438 => x"5873a02e",
          4439 => x"098106a2",
          4440 => x"38783378",
          4441 => x"05567776",
          4442 => x"27983881",
          4443 => x"17705b70",
          4444 => x"71335658",
          4445 => x"5573a02e",
          4446 => x"09810686",
          4447 => x"38757526",
          4448 => x"ea388054",
          4449 => x"73882982",
          4450 => x"d5a80570",
          4451 => x"085255ff",
          4452 => x"b0f33f82",
          4453 => x"d6d80853",
          4454 => x"79527408",
          4455 => x"51ffb3f2",
          4456 => x"3f82d6d8",
          4457 => x"0880c538",
          4458 => x"84153355",
          4459 => x"74812e88",
          4460 => x"3874822e",
          4461 => x"8838b539",
          4462 => x"fce63fac",
          4463 => x"39811a5a",
          4464 => x"8c3dfc11",
          4465 => x"53f80551",
          4466 => x"c5ad3f82",
          4467 => x"d6d80880",
          4468 => x"2e9a38ff",
          4469 => x"1b537852",
          4470 => x"7751fdb1",
          4471 => x"3f82d6d8",
          4472 => x"0881ff06",
          4473 => x"55748538",
          4474 => x"74549139",
          4475 => x"81147081",
          4476 => x"ff065154",
          4477 => x"827427ff",
          4478 => x"8b388054",
          4479 => x"7382d6d8",
          4480 => x"0c8c3d0d",
          4481 => x"04d33d0d",
          4482 => x"b03d08b2",
          4483 => x"3d08b43d",
          4484 => x"08595f5a",
          4485 => x"800baf3d",
          4486 => x"3482d5a4",
          4487 => x"3382d5a0",
          4488 => x"08555b73",
          4489 => x"81cb3873",
          4490 => x"82d59c33",
          4491 => x"55557383",
          4492 => x"38815576",
          4493 => x"802e81bc",
          4494 => x"38817076",
          4495 => x"06555673",
          4496 => x"802e81ad",
          4497 => x"38a85199",
          4498 => x"9f3f82d6",
          4499 => x"d80882d5",
          4500 => x"a00c82d6",
          4501 => x"d808802e",
          4502 => x"81923893",
          4503 => x"53765282",
          4504 => x"d6d80851",
          4505 => x"80dfc63f",
          4506 => x"82d6d808",
          4507 => x"802e8c38",
          4508 => x"82c6c051",
          4509 => x"ffa2ec3f",
          4510 => x"80f73982",
          4511 => x"d6d8085b",
          4512 => x"82d5a008",
          4513 => x"5380f852",
          4514 => x"903d7052",
          4515 => x"54819aa2",
          4516 => x"3f82d6d8",
          4517 => x"085682d6",
          4518 => x"d808742e",
          4519 => x"09810680",
          4520 => x"d03882d6",
          4521 => x"d80851ff",
          4522 => x"aedb3f82",
          4523 => x"d6d80855",
          4524 => x"800b82d6",
          4525 => x"d80825a9",
          4526 => x"3882d6d8",
          4527 => x"08ff0570",
          4528 => x"17555580",
          4529 => x"74348053",
          4530 => x"7481ff06",
          4531 => x"527551f8",
          4532 => x"c23f811b",
          4533 => x"7081ff06",
          4534 => x"5c54937b",
          4535 => x"27833880",
          4536 => x"5b74ff2e",
          4537 => x"098106ff",
          4538 => x"97388639",
          4539 => x"7582d59c",
          4540 => x"34768c38",
          4541 => x"82d5a008",
          4542 => x"802e8438",
          4543 => x"f9d63f8f",
          4544 => x"3d5decc5",
          4545 => x"3f82d6d8",
          4546 => x"08982b70",
          4547 => x"982c5159",
          4548 => x"78ff2eee",
          4549 => x"387881ff",
          4550 => x"0682ee94",
          4551 => x"3370982b",
          4552 => x"70982c82",
          4553 => x"ee903370",
          4554 => x"982b7097",
          4555 => x"2c71982c",
          4556 => x"05708429",
          4557 => x"82c39405",
          4558 => x"70081570",
          4559 => x"33515151",
          4560 => x"51595951",
          4561 => x"595d5881",
          4562 => x"5673782e",
          4563 => x"80e93877",
          4564 => x"7427b438",
          4565 => x"7481800a",
          4566 => x"2981ff0a",
          4567 => x"0570982c",
          4568 => x"51558075",
          4569 => x"2480ce38",
          4570 => x"76537452",
          4571 => x"7751f685",
          4572 => x"3f82d6d8",
          4573 => x"0881ff06",
          4574 => x"5473802e",
          4575 => x"d7387482",
          4576 => x"ee903481",
          4577 => x"56b13974",
          4578 => x"81800a29",
          4579 => x"81800a05",
          4580 => x"70982c70",
          4581 => x"81ff0656",
          4582 => x"51557395",
          4583 => x"26973876",
          4584 => x"53745277",
          4585 => x"51f5ce3f",
          4586 => x"82d6d808",
          4587 => x"81ff0654",
          4588 => x"73cc38d3",
          4589 => x"39805675",
          4590 => x"802e80ca",
          4591 => x"38811c55",
          4592 => x"7482ee94",
          4593 => x"3474982b",
          4594 => x"70982c82",
          4595 => x"ee903370",
          4596 => x"982b7098",
          4597 => x"2c701011",
          4598 => x"70822b82",
          4599 => x"c3981133",
          4600 => x"5e515151",
          4601 => x"57585155",
          4602 => x"74772e09",
          4603 => x"8106fe92",
          4604 => x"3882c39c",
          4605 => x"14087d0c",
          4606 => x"800b82ee",
          4607 => x"9434800b",
          4608 => x"82ee9034",
          4609 => x"92397582",
          4610 => x"ee943475",
          4611 => x"82ee9034",
          4612 => x"78af3d34",
          4613 => x"757d0c7e",
          4614 => x"54739526",
          4615 => x"fde13873",
          4616 => x"842982ad",
          4617 => x"c0055473",
          4618 => x"080482ee",
          4619 => x"9c335473",
          4620 => x"7e2efdcb",
          4621 => x"3882ee98",
          4622 => x"33557375",
          4623 => x"27ab3874",
          4624 => x"982b7098",
          4625 => x"2c515573",
          4626 => x"75249e38",
          4627 => x"741a5473",
          4628 => x"33811534",
          4629 => x"7481800a",
          4630 => x"2981ff0a",
          4631 => x"0570982c",
          4632 => x"82ee9c33",
          4633 => x"565155df",
          4634 => x"3982ee9c",
          4635 => x"33811156",
          4636 => x"547482ee",
          4637 => x"9c34731a",
          4638 => x"54ae3d33",
          4639 => x"743482ee",
          4640 => x"98335473",
          4641 => x"7e258938",
          4642 => x"81145473",
          4643 => x"82ee9834",
          4644 => x"82ee9c33",
          4645 => x"7081800a",
          4646 => x"2981ff0a",
          4647 => x"0570982c",
          4648 => x"82ee9833",
          4649 => x"5a515656",
          4650 => x"747725a8",
          4651 => x"3882f2bc",
          4652 => x"0852741a",
          4653 => x"70335254",
          4654 => x"ffa1f73f",
          4655 => x"7481800a",
          4656 => x"2981800a",
          4657 => x"0570982c",
          4658 => x"82ee9833",
          4659 => x"56515573",
          4660 => x"7524da38",
          4661 => x"82ee9c33",
          4662 => x"70982b70",
          4663 => x"982c82ee",
          4664 => x"98335a51",
          4665 => x"56567477",
          4666 => x"25fc9438",
          4667 => x"82f2bc08",
          4668 => x"528851ff",
          4669 => x"a1bc3f74",
          4670 => x"81800a29",
          4671 => x"81800a05",
          4672 => x"70982c82",
          4673 => x"ee983356",
          4674 => x"51557375",
          4675 => x"24de38fb",
          4676 => x"ee39837a",
          4677 => x"34800b81",
          4678 => x"1b3482ee",
          4679 => x"9c538052",
          4680 => x"82b6a051",
          4681 => x"f39c3f81",
          4682 => x"fd3982ee",
          4683 => x"9c337081",
          4684 => x"ff065555",
          4685 => x"73802efb",
          4686 => x"c63882ee",
          4687 => x"9833ff05",
          4688 => x"547382ee",
          4689 => x"9834ff15",
          4690 => x"547382ee",
          4691 => x"9c3482f2",
          4692 => x"bc085288",
          4693 => x"51ffa0da",
          4694 => x"3f82ee9c",
          4695 => x"3370982b",
          4696 => x"70982c82",
          4697 => x"ee983357",
          4698 => x"51565774",
          4699 => x"7425ad38",
          4700 => x"741a5481",
          4701 => x"14337434",
          4702 => x"82f2bc08",
          4703 => x"52733351",
          4704 => x"ffa0af3f",
          4705 => x"7481800a",
          4706 => x"2981800a",
          4707 => x"0570982c",
          4708 => x"82ee9833",
          4709 => x"58515575",
          4710 => x"7524d538",
          4711 => x"82f2bc08",
          4712 => x"52a051ff",
          4713 => x"a08c3f82",
          4714 => x"ee9c3370",
          4715 => x"982b7098",
          4716 => x"2c82ee98",
          4717 => x"33575156",
          4718 => x"57747424",
          4719 => x"fac13882",
          4720 => x"f2bc0852",
          4721 => x"8851ff9f",
          4722 => x"e93f7481",
          4723 => x"800a2981",
          4724 => x"800a0570",
          4725 => x"982c82ee",
          4726 => x"98335851",
          4727 => x"55757525",
          4728 => x"de38fa9b",
          4729 => x"3982ee98",
          4730 => x"337a0554",
          4731 => x"80743482",
          4732 => x"f2bc0852",
          4733 => x"8a51ff9f",
          4734 => x"b93f82ee",
          4735 => x"98527951",
          4736 => x"f6c93f82",
          4737 => x"d6d80881",
          4738 => x"ff065473",
          4739 => x"963882ee",
          4740 => x"98335473",
          4741 => x"802e8f38",
          4742 => x"81537352",
          4743 => x"7951f1f3",
          4744 => x"3f843980",
          4745 => x"7a34800b",
          4746 => x"82ee9c34",
          4747 => x"800b82ee",
          4748 => x"98347982",
          4749 => x"d6d80caf",
          4750 => x"3d0d0482",
          4751 => x"ee9c3354",
          4752 => x"73802ef9",
          4753 => x"ba3882f2",
          4754 => x"bc085288",
          4755 => x"51ff9ee2",
          4756 => x"3f82ee9c",
          4757 => x"33ff0554",
          4758 => x"7382ee9c",
          4759 => x"347381ff",
          4760 => x"0654dd39",
          4761 => x"82ee9c33",
          4762 => x"82ee9833",
          4763 => x"55557375",
          4764 => x"2ef98c38",
          4765 => x"ff145473",
          4766 => x"82ee9834",
          4767 => x"74982b70",
          4768 => x"982c7581",
          4769 => x"ff065651",
          4770 => x"55747425",
          4771 => x"ad38741a",
          4772 => x"54811433",
          4773 => x"743482f2",
          4774 => x"bc085273",
          4775 => x"3351ff9e",
          4776 => x"913f7481",
          4777 => x"800a2981",
          4778 => x"800a0570",
          4779 => x"982c82ee",
          4780 => x"98335851",
          4781 => x"55757524",
          4782 => x"d53882f2",
          4783 => x"bc0852a0",
          4784 => x"51ff9dee",
          4785 => x"3f82ee9c",
          4786 => x"3370982b",
          4787 => x"70982c82",
          4788 => x"ee983357",
          4789 => x"51565774",
          4790 => x"7424f8a3",
          4791 => x"3882f2bc",
          4792 => x"08528851",
          4793 => x"ff9dcb3f",
          4794 => x"7481800a",
          4795 => x"2981800a",
          4796 => x"0570982c",
          4797 => x"82ee9833",
          4798 => x"58515575",
          4799 => x"7525de38",
          4800 => x"f7fd3982",
          4801 => x"ee9c3370",
          4802 => x"81ff0682",
          4803 => x"ee983359",
          4804 => x"56547477",
          4805 => x"27f7e838",
          4806 => x"82f2bc08",
          4807 => x"52811454",
          4808 => x"7382ee9c",
          4809 => x"34741a70",
          4810 => x"335254ff",
          4811 => x"9d843f82",
          4812 => x"ee9c3370",
          4813 => x"81ff0682",
          4814 => x"ee983358",
          4815 => x"56547575",
          4816 => x"26d638f7",
          4817 => x"ba3982ee",
          4818 => x"9c538052",
          4819 => x"82b6a051",
          4820 => x"eef03f80",
          4821 => x"0b82ee9c",
          4822 => x"34800b82",
          4823 => x"ee9834f7",
          4824 => x"9e397ab0",
          4825 => x"3882d598",
          4826 => x"08557480",
          4827 => x"2ea63874",
          4828 => x"51ffa591",
          4829 => x"3f82d6d8",
          4830 => x"0882ee98",
          4831 => x"3482d6d8",
          4832 => x"0881ff06",
          4833 => x"81055374",
          4834 => x"527951ff",
          4835 => x"a6d73f93",
          4836 => x"5b81c039",
          4837 => x"7a842982",
          4838 => x"d4cc05fc",
          4839 => x"11085654",
          4840 => x"74802ea7",
          4841 => x"387451ff",
          4842 => x"a4db3f82",
          4843 => x"d6d80882",
          4844 => x"ee983482",
          4845 => x"d6d80881",
          4846 => x"ff068105",
          4847 => x"53745279",
          4848 => x"51ffa6a1",
          4849 => x"3fff1b54",
          4850 => x"80fa3973",
          4851 => x"08557480",
          4852 => x"2ef6ac38",
          4853 => x"7451ffa4",
          4854 => x"ac3f9939",
          4855 => x"7a932e09",
          4856 => x"8106ae38",
          4857 => x"82d4cc08",
          4858 => x"5574802e",
          4859 => x"a4387451",
          4860 => x"ffa4923f",
          4861 => x"82d6d808",
          4862 => x"82ee9834",
          4863 => x"82d6d808",
          4864 => x"81ff0681",
          4865 => x"05537452",
          4866 => x"7951ffa5",
          4867 => x"d83f80c3",
          4868 => x"397a8429",
          4869 => x"82d4d005",
          4870 => x"70085654",
          4871 => x"74802eab",
          4872 => x"387451ff",
          4873 => x"a3df3f82",
          4874 => x"d6d80882",
          4875 => x"ee983482",
          4876 => x"d6d80881",
          4877 => x"ff068105",
          4878 => x"53745279",
          4879 => x"51ffa5a5",
          4880 => x"3f811b54",
          4881 => x"7381ff06",
          4882 => x"5b893974",
          4883 => x"82ee9834",
          4884 => x"747a3482",
          4885 => x"ee9c5382",
          4886 => x"ee983352",
          4887 => x"7951ece2",
          4888 => x"3ff59c39",
          4889 => x"82ee9c33",
          4890 => x"7081ff06",
          4891 => x"82ee9833",
          4892 => x"59565474",
          4893 => x"7727f587",
          4894 => x"3882f2bc",
          4895 => x"08528114",
          4896 => x"547382ee",
          4897 => x"9c34741a",
          4898 => x"70335254",
          4899 => x"ff9aa33f",
          4900 => x"f4ed3982",
          4901 => x"ee9c3354",
          4902 => x"73802ef4",
          4903 => x"e23882f2",
          4904 => x"bc085288",
          4905 => x"51ff9a8a",
          4906 => x"3f82ee9c",
          4907 => x"33ff0554",
          4908 => x"7382ee9c",
          4909 => x"34f4c839",
          4910 => x"ff3d0d02",
          4911 => x"8f053352",
          4912 => x"718a2e09",
          4913 => x"8106a038",
          4914 => x"82d6c408",
          4915 => x"810582d6",
          4916 => x"c40c980b",
          4917 => x"82d6c408",
          4918 => x"25873898",
          4919 => x"0b82d6c4",
          4920 => x"0c800b82",
          4921 => x"d6c80c82",
          4922 => x"d6c40884",
          4923 => x"2982d6c4",
          4924 => x"08057088",
          4925 => x"2982d6c8",
          4926 => x"080587a0",
          4927 => x"a0801170",
          4928 => x"82d6c00c",
          4929 => x"51515182",
          4930 => x"d5c01233",
          4931 => x"713482d6",
          4932 => x"c8088105",
          4933 => x"82d6c80c",
          4934 => x"a70b82d6",
          4935 => x"c80825a0",
          4936 => x"3882d6c4",
          4937 => x"08810582",
          4938 => x"d6c40c98",
          4939 => x"0b82d6c4",
          4940 => x"08258738",
          4941 => x"980b82d6",
          4942 => x"c40c800b",
          4943 => x"82d6c80c",
          4944 => x"800b82d6",
          4945 => x"d80c833d",
          4946 => x"0d04ff0b",
          4947 => x"82d6d80c",
          4948 => x"04f93d0d",
          4949 => x"83bff40b",
          4950 => x"82d6d00c",
          4951 => x"84800b82",
          4952 => x"d6cc23a0",
          4953 => x"80538052",
          4954 => x"83bff451",
          4955 => x"ffa9a23f",
          4956 => x"82d6d008",
          4957 => x"54805877",
          4958 => x"74348157",
          4959 => x"76811534",
          4960 => x"82d6d008",
          4961 => x"54778415",
          4962 => x"34768515",
          4963 => x"3482d6d0",
          4964 => x"08547786",
          4965 => x"15347687",
          4966 => x"153482d6",
          4967 => x"d00882d6",
          4968 => x"cc22ff05",
          4969 => x"fe808007",
          4970 => x"7083ffff",
          4971 => x"0670882a",
          4972 => x"58515556",
          4973 => x"74881734",
          4974 => x"73891734",
          4975 => x"82d6cc22",
          4976 => x"70882982",
          4977 => x"d6d00805",
          4978 => x"f8115155",
          4979 => x"55778215",
          4980 => x"34768315",
          4981 => x"34893d0d",
          4982 => x"04ff3d0d",
          4983 => x"73528151",
          4984 => x"8472278f",
          4985 => x"38fb1283",
          4986 => x"2a821170",
          4987 => x"83ffff06",
          4988 => x"51515170",
          4989 => x"82d6d80c",
          4990 => x"833d0d04",
          4991 => x"f93d0d02",
          4992 => x"a6052202",
          4993 => x"8405aa05",
          4994 => x"22710582",
          4995 => x"d6d00871",
          4996 => x"832b7111",
          4997 => x"74832b73",
          4998 => x"11703381",
          4999 => x"12337188",
          5000 => x"2b0702a4",
          5001 => x"05ae0522",
          5002 => x"7181ffff",
          5003 => x"06077088",
          5004 => x"2a535152",
          5005 => x"59545b5b",
          5006 => x"57535455",
          5007 => x"71773470",
          5008 => x"81183482",
          5009 => x"d6d00814",
          5010 => x"75882a52",
          5011 => x"54708215",
          5012 => x"34748315",
          5013 => x"3482d6d0",
          5014 => x"08701770",
          5015 => x"33811233",
          5016 => x"71882b07",
          5017 => x"70832b8f",
          5018 => x"fff80651",
          5019 => x"52565271",
          5020 => x"057383ff",
          5021 => x"ff067088",
          5022 => x"2a545451",
          5023 => x"71821234",
          5024 => x"7281ff06",
          5025 => x"53728312",
          5026 => x"3482d6d0",
          5027 => x"08165671",
          5028 => x"76347281",
          5029 => x"1734893d",
          5030 => x"0d04fb3d",
          5031 => x"0d82d6d0",
          5032 => x"08028405",
          5033 => x"9e052270",
          5034 => x"832b7211",
          5035 => x"86113387",
          5036 => x"1233718b",
          5037 => x"2b71832b",
          5038 => x"07585b59",
          5039 => x"52555272",
          5040 => x"05841233",
          5041 => x"85133371",
          5042 => x"882b0770",
          5043 => x"882a5456",
          5044 => x"56527084",
          5045 => x"13347385",
          5046 => x"133482d6",
          5047 => x"d0087014",
          5048 => x"84113385",
          5049 => x"1233718b",
          5050 => x"2b71832b",
          5051 => x"07565957",
          5052 => x"52720586",
          5053 => x"12338713",
          5054 => x"3371882b",
          5055 => x"0770882a",
          5056 => x"54565652",
          5057 => x"70861334",
          5058 => x"73871334",
          5059 => x"82d6d008",
          5060 => x"13703381",
          5061 => x"12337188",
          5062 => x"2b077081",
          5063 => x"ffff0670",
          5064 => x"882a5351",
          5065 => x"53535371",
          5066 => x"73347081",
          5067 => x"1434873d",
          5068 => x"0d04fa3d",
          5069 => x"0d02a205",
          5070 => x"2282d6d0",
          5071 => x"0871832b",
          5072 => x"71117033",
          5073 => x"81123371",
          5074 => x"882b0770",
          5075 => x"88291570",
          5076 => x"33811233",
          5077 => x"71982b71",
          5078 => x"902b0753",
          5079 => x"5f535552",
          5080 => x"5a565753",
          5081 => x"54718025",
          5082 => x"80f63872",
          5083 => x"51feab3f",
          5084 => x"82d6d008",
          5085 => x"70167033",
          5086 => x"81123371",
          5087 => x"8b2b7183",
          5088 => x"2b077411",
          5089 => x"70338112",
          5090 => x"3371882b",
          5091 => x"0770832b",
          5092 => x"8ffff806",
          5093 => x"51525451",
          5094 => x"535a5853",
          5095 => x"72057488",
          5096 => x"2a545272",
          5097 => x"82133473",
          5098 => x"83133482",
          5099 => x"d6d00870",
          5100 => x"16703381",
          5101 => x"1233718b",
          5102 => x"2b71832b",
          5103 => x"07565957",
          5104 => x"55720570",
          5105 => x"33811233",
          5106 => x"71882b07",
          5107 => x"7081ffff",
          5108 => x"0670882a",
          5109 => x"57515258",
          5110 => x"52727434",
          5111 => x"71811534",
          5112 => x"883d0d04",
          5113 => x"fb3d0d82",
          5114 => x"d6d00802",
          5115 => x"84059e05",
          5116 => x"2270832b",
          5117 => x"72118211",
          5118 => x"33831233",
          5119 => x"718b2b71",
          5120 => x"832b0759",
          5121 => x"5b595256",
          5122 => x"52730571",
          5123 => x"33811333",
          5124 => x"71882b07",
          5125 => x"028c05a2",
          5126 => x"05227107",
          5127 => x"70882a53",
          5128 => x"51535353",
          5129 => x"71733470",
          5130 => x"81143482",
          5131 => x"d6d00870",
          5132 => x"15703381",
          5133 => x"1233718b",
          5134 => x"2b71832b",
          5135 => x"07565957",
          5136 => x"52720582",
          5137 => x"12338313",
          5138 => x"3371882b",
          5139 => x"0770882a",
          5140 => x"54555652",
          5141 => x"70821334",
          5142 => x"72831334",
          5143 => x"82d6d008",
          5144 => x"14821133",
          5145 => x"83123371",
          5146 => x"882b0782",
          5147 => x"d6d80c52",
          5148 => x"54873d0d",
          5149 => x"04f73d0d",
          5150 => x"7b82d6d0",
          5151 => x"0831832a",
          5152 => x"7083ffff",
          5153 => x"06705357",
          5154 => x"53fda73f",
          5155 => x"82d6d008",
          5156 => x"76832b71",
          5157 => x"11821133",
          5158 => x"83123371",
          5159 => x"8b2b7183",
          5160 => x"2b077511",
          5161 => x"70338112",
          5162 => x"3371982b",
          5163 => x"71902b07",
          5164 => x"53424051",
          5165 => x"535b5855",
          5166 => x"59547280",
          5167 => x"258d3882",
          5168 => x"80805275",
          5169 => x"51fe9d3f",
          5170 => x"81843984",
          5171 => x"14338515",
          5172 => x"33718b2b",
          5173 => x"71832b07",
          5174 => x"76117988",
          5175 => x"2a535155",
          5176 => x"58557686",
          5177 => x"14347581",
          5178 => x"ff065675",
          5179 => x"87143482",
          5180 => x"d6d00870",
          5181 => x"19841233",
          5182 => x"85133371",
          5183 => x"882b0770",
          5184 => x"882a5457",
          5185 => x"5b565372",
          5186 => x"84163473",
          5187 => x"85163482",
          5188 => x"d6d00818",
          5189 => x"53800b86",
          5190 => x"1434800b",
          5191 => x"87143482",
          5192 => x"d6d00853",
          5193 => x"76841434",
          5194 => x"75851434",
          5195 => x"82d6d008",
          5196 => x"18703381",
          5197 => x"12337188",
          5198 => x"2b077082",
          5199 => x"80800770",
          5200 => x"882a5351",
          5201 => x"55565474",
          5202 => x"74347281",
          5203 => x"15348b3d",
          5204 => x"0d04ff3d",
          5205 => x"0d735282",
          5206 => x"d6d00884",
          5207 => x"38f7f23f",
          5208 => x"71802e86",
          5209 => x"387151fe",
          5210 => x"8c3f833d",
          5211 => x"0d04f53d",
          5212 => x"0d807e52",
          5213 => x"58f8e23f",
          5214 => x"82d6d808",
          5215 => x"83ffff06",
          5216 => x"82d6d008",
          5217 => x"84113385",
          5218 => x"12337188",
          5219 => x"2b07705f",
          5220 => x"5956585a",
          5221 => x"81ffff59",
          5222 => x"75782e80",
          5223 => x"cb387588",
          5224 => x"29177033",
          5225 => x"81123371",
          5226 => x"882b0770",
          5227 => x"81ffff06",
          5228 => x"79317083",
          5229 => x"ffff0670",
          5230 => x"7f275253",
          5231 => x"51565955",
          5232 => x"7779278a",
          5233 => x"3873802e",
          5234 => x"85387578",
          5235 => x"5a5b8415",
          5236 => x"33851633",
          5237 => x"71882b07",
          5238 => x"575475c2",
          5239 => x"387881ff",
          5240 => x"ff2e8538",
          5241 => x"7a795956",
          5242 => x"8076832b",
          5243 => x"82d6d008",
          5244 => x"11703381",
          5245 => x"12337188",
          5246 => x"2b077081",
          5247 => x"ffff0651",
          5248 => x"525a565c",
          5249 => x"5573752e",
          5250 => x"83388155",
          5251 => x"80547978",
          5252 => x"2681cc38",
          5253 => x"74547480",
          5254 => x"2e81c438",
          5255 => x"777a2e09",
          5256 => x"81068938",
          5257 => x"7551f8f2",
          5258 => x"3f81ac39",
          5259 => x"82808053",
          5260 => x"79527551",
          5261 => x"f7c63f82",
          5262 => x"d6d00870",
          5263 => x"1c861133",
          5264 => x"87123371",
          5265 => x"8b2b7183",
          5266 => x"2b07535a",
          5267 => x"5e557405",
          5268 => x"7a177083",
          5269 => x"ffff0670",
          5270 => x"882a5c59",
          5271 => x"56547884",
          5272 => x"15347681",
          5273 => x"ff065776",
          5274 => x"85153482",
          5275 => x"d6d00875",
          5276 => x"832b7111",
          5277 => x"721e8611",
          5278 => x"33871233",
          5279 => x"71882b07",
          5280 => x"70882a53",
          5281 => x"5b5e535a",
          5282 => x"56547386",
          5283 => x"19347587",
          5284 => x"193482d6",
          5285 => x"d008701c",
          5286 => x"84113385",
          5287 => x"1233718b",
          5288 => x"2b71832b",
          5289 => x"07535d5a",
          5290 => x"55740554",
          5291 => x"78861534",
          5292 => x"76871534",
          5293 => x"82d6d008",
          5294 => x"7016711d",
          5295 => x"84113385",
          5296 => x"12337188",
          5297 => x"2b077088",
          5298 => x"2a535a5f",
          5299 => x"52565473",
          5300 => x"84163475",
          5301 => x"85163482",
          5302 => x"d6d0081b",
          5303 => x"84055473",
          5304 => x"82d6d80c",
          5305 => x"8d3d0d04",
          5306 => x"fe3d0d74",
          5307 => x"5282d6d0",
          5308 => x"088438f4",
          5309 => x"dc3f7153",
          5310 => x"71802e8b",
          5311 => x"387151fc",
          5312 => x"ed3f82d6",
          5313 => x"d8085372",
          5314 => x"82d6d80c",
          5315 => x"843d0d04",
          5316 => x"ee3d0d64",
          5317 => x"66405c80",
          5318 => x"70424082",
          5319 => x"d6d00860",
          5320 => x"2e098106",
          5321 => x"8438f4a9",
          5322 => x"3f7b8e38",
          5323 => x"7e51ffb8",
          5324 => x"3f82d6d8",
          5325 => x"085483c7",
          5326 => x"397e8b38",
          5327 => x"7b51fc92",
          5328 => x"3f7e5483",
          5329 => x"ba397e51",
          5330 => x"f58f3f82",
          5331 => x"d6d80883",
          5332 => x"ffff0682",
          5333 => x"d6d0087d",
          5334 => x"7131832a",
          5335 => x"7083ffff",
          5336 => x"0670832b",
          5337 => x"73117033",
          5338 => x"81123371",
          5339 => x"882b0770",
          5340 => x"75317083",
          5341 => x"ffff0670",
          5342 => x"8829fc05",
          5343 => x"7388291a",
          5344 => x"70338112",
          5345 => x"3371882b",
          5346 => x"0770902b",
          5347 => x"53444e53",
          5348 => x"4841525c",
          5349 => x"545b415c",
          5350 => x"565b5b73",
          5351 => x"80258f38",
          5352 => x"7681ffff",
          5353 => x"06753170",
          5354 => x"83ffff06",
          5355 => x"42548216",
          5356 => x"33831733",
          5357 => x"71882b07",
          5358 => x"7088291c",
          5359 => x"70338112",
          5360 => x"3371982b",
          5361 => x"71902b07",
          5362 => x"53474552",
          5363 => x"56547380",
          5364 => x"258b3878",
          5365 => x"75317083",
          5366 => x"ffff0641",
          5367 => x"54777b27",
          5368 => x"81fe3860",
          5369 => x"1854737b",
          5370 => x"2e098106",
          5371 => x"8f387851",
          5372 => x"f6c03f7a",
          5373 => x"83ffff06",
          5374 => x"5881e539",
          5375 => x"7f8e387a",
          5376 => x"74248938",
          5377 => x"7851f6aa",
          5378 => x"3f81a539",
          5379 => x"7f18557a",
          5380 => x"752480c8",
          5381 => x"38791d82",
          5382 => x"11338312",
          5383 => x"3371882b",
          5384 => x"07535754",
          5385 => x"f4f43f80",
          5386 => x"527851f7",
          5387 => x"b73f82d6",
          5388 => x"d80883ff",
          5389 => x"ff067e54",
          5390 => x"7c537083",
          5391 => x"2b82d6d0",
          5392 => x"08118405",
          5393 => x"535559ff",
          5394 => x"90d13f82",
          5395 => x"d6d00814",
          5396 => x"84057583",
          5397 => x"ffff0659",
          5398 => x"5c818539",
          5399 => x"6015547a",
          5400 => x"742480d4",
          5401 => x"387851f5",
          5402 => x"c93f82d6",
          5403 => x"d0081d82",
          5404 => x"11338312",
          5405 => x"3371882b",
          5406 => x"07534354",
          5407 => x"f49c3f80",
          5408 => x"527851f6",
          5409 => x"df3f82d6",
          5410 => x"d80883ff",
          5411 => x"ff067e54",
          5412 => x"7c537083",
          5413 => x"2b82d6d0",
          5414 => x"08118405",
          5415 => x"535559ff",
          5416 => x"8ff93f82",
          5417 => x"d6d00814",
          5418 => x"84056062",
          5419 => x"0519555c",
          5420 => x"7383ffff",
          5421 => x"0658a939",
          5422 => x"7b7f5254",
          5423 => x"f9b03f82",
          5424 => x"d6d8085c",
          5425 => x"82d6d808",
          5426 => x"802e9338",
          5427 => x"7d537352",
          5428 => x"82d6d808",
          5429 => x"51ff948d",
          5430 => x"3f7351f7",
          5431 => x"983f7a58",
          5432 => x"7a782799",
          5433 => x"3880537a",
          5434 => x"527851f2",
          5435 => x"8f3f7a19",
          5436 => x"832b82d6",
          5437 => x"d0080584",
          5438 => x"0551f6f9",
          5439 => x"3f7b5473",
          5440 => x"82d6d80c",
          5441 => x"943d0d04",
          5442 => x"fc3d0d77",
          5443 => x"77297052",
          5444 => x"54fbd53f",
          5445 => x"82d6d808",
          5446 => x"5582d6d8",
          5447 => x"08802e8e",
          5448 => x"38735380",
          5449 => x"5282d6d8",
          5450 => x"0851ff99",
          5451 => x"e43f7482",
          5452 => x"d6d80c86",
          5453 => x"3d0d04ff",
          5454 => x"3d0d028f",
          5455 => x"05335181",
          5456 => x"52707226",
          5457 => x"873882d6",
          5458 => x"d4113352",
          5459 => x"7182d6d8",
          5460 => x"0c833d0d",
          5461 => x"04fc3d0d",
          5462 => x"029b0533",
          5463 => x"0284059f",
          5464 => x"05335653",
          5465 => x"83517281",
          5466 => x"2680e038",
          5467 => x"72842b87",
          5468 => x"c0928c11",
          5469 => x"53518854",
          5470 => x"74802e84",
          5471 => x"38818854",
          5472 => x"73720c87",
          5473 => x"c0928c11",
          5474 => x"5181710c",
          5475 => x"850b87c0",
          5476 => x"988c0c70",
          5477 => x"52710870",
          5478 => x"82065151",
          5479 => x"70802e8a",
          5480 => x"3887c098",
          5481 => x"8c085170",
          5482 => x"ec387108",
          5483 => x"fc808006",
          5484 => x"52719238",
          5485 => x"87c0988c",
          5486 => x"08517080",
          5487 => x"2e873871",
          5488 => x"82d6d414",
          5489 => x"3482d6d4",
          5490 => x"13335170",
          5491 => x"82d6d80c",
          5492 => x"863d0d04",
          5493 => x"f33d0d60",
          5494 => x"6264028c",
          5495 => x"05bf0533",
          5496 => x"5740585b",
          5497 => x"8374525a",
          5498 => x"fecd3f82",
          5499 => x"d6d80881",
          5500 => x"067a5452",
          5501 => x"7181be38",
          5502 => x"71727584",
          5503 => x"2b87c092",
          5504 => x"801187c0",
          5505 => x"928c1287",
          5506 => x"c0928413",
          5507 => x"415a4057",
          5508 => x"5a58850b",
          5509 => x"87c0988c",
          5510 => x"0c767d0c",
          5511 => x"84760c75",
          5512 => x"0870852a",
          5513 => x"70810651",
          5514 => x"53547180",
          5515 => x"2e8e387b",
          5516 => x"0852717b",
          5517 => x"7081055d",
          5518 => x"34811959",
          5519 => x"8074a206",
          5520 => x"53537173",
          5521 => x"2e833881",
          5522 => x"537883ff",
          5523 => x"268f3872",
          5524 => x"802e8a38",
          5525 => x"87c0988c",
          5526 => x"085271c3",
          5527 => x"3887c098",
          5528 => x"8c085271",
          5529 => x"802e8738",
          5530 => x"7884802e",
          5531 => x"99388176",
          5532 => x"0c87c092",
          5533 => x"8c155372",
          5534 => x"08708206",
          5535 => x"515271f7",
          5536 => x"38ff1a5a",
          5537 => x"8d398480",
          5538 => x"17811970",
          5539 => x"81ff065a",
          5540 => x"53577980",
          5541 => x"2e903873",
          5542 => x"fc808006",
          5543 => x"52718738",
          5544 => x"7d7826fe",
          5545 => x"ed3873fc",
          5546 => x"80800652",
          5547 => x"71802e83",
          5548 => x"38815271",
          5549 => x"537282d6",
          5550 => x"d80c8f3d",
          5551 => x"0d04f33d",
          5552 => x"0d606264",
          5553 => x"028c05bf",
          5554 => x"05335740",
          5555 => x"585b8359",
          5556 => x"80745258",
          5557 => x"fce13f82",
          5558 => x"d6d80881",
          5559 => x"06795452",
          5560 => x"71782e09",
          5561 => x"810681b1",
          5562 => x"38777484",
          5563 => x"2b87c092",
          5564 => x"801187c0",
          5565 => x"928c1287",
          5566 => x"c0928413",
          5567 => x"40595f56",
          5568 => x"5a850b87",
          5569 => x"c0988c0c",
          5570 => x"767d0c82",
          5571 => x"760c8058",
          5572 => x"75087084",
          5573 => x"2a708106",
          5574 => x"51535471",
          5575 => x"802e8c38",
          5576 => x"7a708105",
          5577 => x"5c337c0c",
          5578 => x"81185873",
          5579 => x"812a7081",
          5580 => x"06515271",
          5581 => x"802e8a38",
          5582 => x"87c0988c",
          5583 => x"085271d0",
          5584 => x"3887c098",
          5585 => x"8c085271",
          5586 => x"802e8738",
          5587 => x"7784802e",
          5588 => x"99388176",
          5589 => x"0c87c092",
          5590 => x"8c155372",
          5591 => x"08708206",
          5592 => x"515271f7",
          5593 => x"38ff1959",
          5594 => x"8d39811a",
          5595 => x"7081ff06",
          5596 => x"84801959",
          5597 => x"5b527880",
          5598 => x"2e903873",
          5599 => x"fc808006",
          5600 => x"52718738",
          5601 => x"7d7a26fe",
          5602 => x"f83873fc",
          5603 => x"80800652",
          5604 => x"71802e83",
          5605 => x"38815271",
          5606 => x"537282d6",
          5607 => x"d80c8f3d",
          5608 => x"0d04fa3d",
          5609 => x"0d7a0284",
          5610 => x"05a30533",
          5611 => x"028805a7",
          5612 => x"05337154",
          5613 => x"545657fa",
          5614 => x"fe3f82d6",
          5615 => x"d8088106",
          5616 => x"53835472",
          5617 => x"80fe3885",
          5618 => x"0b87c098",
          5619 => x"8c0c8156",
          5620 => x"71762e80",
          5621 => x"dc387176",
          5622 => x"24933874",
          5623 => x"842b87c0",
          5624 => x"928c1154",
          5625 => x"5471802e",
          5626 => x"8d3880d4",
          5627 => x"3971832e",
          5628 => x"80c63880",
          5629 => x"cb397208",
          5630 => x"70812a70",
          5631 => x"81065151",
          5632 => x"5271802e",
          5633 => x"8a3887c0",
          5634 => x"988c0852",
          5635 => x"71e83887",
          5636 => x"c0988c08",
          5637 => x"52719638",
          5638 => x"81730c87",
          5639 => x"c0928c14",
          5640 => x"53720870",
          5641 => x"82065152",
          5642 => x"71f73896",
          5643 => x"39805692",
          5644 => x"3988800a",
          5645 => x"770c8539",
          5646 => x"8180770c",
          5647 => x"72568339",
          5648 => x"84567554",
          5649 => x"7382d6d8",
          5650 => x"0c883d0d",
          5651 => x"04fe3d0d",
          5652 => x"74811133",
          5653 => x"71337188",
          5654 => x"2b0782d6",
          5655 => x"d80c5351",
          5656 => x"843d0d04",
          5657 => x"fd3d0d75",
          5658 => x"83113382",
          5659 => x"12337190",
          5660 => x"2b71882b",
          5661 => x"07811433",
          5662 => x"70720788",
          5663 => x"2b753371",
          5664 => x"0782d6d8",
          5665 => x"0c525354",
          5666 => x"56545285",
          5667 => x"3d0d04ff",
          5668 => x"3d0d7302",
          5669 => x"84059205",
          5670 => x"22525270",
          5671 => x"72708105",
          5672 => x"54347088",
          5673 => x"2a517072",
          5674 => x"34833d0d",
          5675 => x"04ff3d0d",
          5676 => x"73755252",
          5677 => x"70727081",
          5678 => x"05543470",
          5679 => x"882a5170",
          5680 => x"72708105",
          5681 => x"54347088",
          5682 => x"2a517072",
          5683 => x"70810554",
          5684 => x"3470882a",
          5685 => x"51707234",
          5686 => x"833d0d04",
          5687 => x"fe3d0d76",
          5688 => x"75775454",
          5689 => x"5170802e",
          5690 => x"92387170",
          5691 => x"81055333",
          5692 => x"73708105",
          5693 => x"5534ff11",
          5694 => x"51eb3984",
          5695 => x"3d0d04fe",
          5696 => x"3d0d7577",
          5697 => x"76545253",
          5698 => x"72727081",
          5699 => x"055434ff",
          5700 => x"115170f4",
          5701 => x"38843d0d",
          5702 => x"04fc3d0d",
          5703 => x"78777956",
          5704 => x"56537470",
          5705 => x"81055633",
          5706 => x"74708105",
          5707 => x"56337171",
          5708 => x"31ff1656",
          5709 => x"52525272",
          5710 => x"802e8638",
          5711 => x"71802ee2",
          5712 => x"387182d6",
          5713 => x"d80c863d",
          5714 => x"0d04fe3d",
          5715 => x"0d747654",
          5716 => x"51893971",
          5717 => x"732e8a38",
          5718 => x"81115170",
          5719 => x"335271f3",
          5720 => x"38703382",
          5721 => x"d6d80c84",
          5722 => x"3d0d0480",
          5723 => x"0b82d6d8",
          5724 => x"0c04fb3d",
          5725 => x"0d777008",
          5726 => x"70708105",
          5727 => x"52337054",
          5728 => x"555556e7",
          5729 => x"3fff5582",
          5730 => x"d6d808a2",
          5731 => x"3872802e",
          5732 => x"983883b5",
          5733 => x"52725180",
          5734 => x"f7b63f82",
          5735 => x"d6d80883",
          5736 => x"ffff0653",
          5737 => x"72802e86",
          5738 => x"3873760c",
          5739 => x"72557482",
          5740 => x"d6d80c87",
          5741 => x"3d0d04f7",
          5742 => x"3d0d7b56",
          5743 => x"800b8317",
          5744 => x"33565a74",
          5745 => x"7a2e80d6",
          5746 => x"388154b4",
          5747 => x"160853b8",
          5748 => x"16705381",
          5749 => x"17335259",
          5750 => x"f9e43f82",
          5751 => x"d6d8087a",
          5752 => x"2e098106",
          5753 => x"b73882d6",
          5754 => x"d8088317",
          5755 => x"34b41608",
          5756 => x"70a81808",
          5757 => x"31a01808",
          5758 => x"59565874",
          5759 => x"77279f38",
          5760 => x"82163355",
          5761 => x"74822e09",
          5762 => x"81069338",
          5763 => x"81547618",
          5764 => x"53785281",
          5765 => x"163351f9",
          5766 => x"a53f8339",
          5767 => x"815a7982",
          5768 => x"d6d80c8b",
          5769 => x"3d0d04fa",
          5770 => x"3d0d787a",
          5771 => x"56568057",
          5772 => x"74b41708",
          5773 => x"2eaf3875",
          5774 => x"51fefc3f",
          5775 => x"82d6d808",
          5776 => x"5782d6d8",
          5777 => x"089f3881",
          5778 => x"547453b8",
          5779 => x"16528116",
          5780 => x"3351f780",
          5781 => x"3f82d6d8",
          5782 => x"08802e85",
          5783 => x"38ff5581",
          5784 => x"5774b417",
          5785 => x"0c7682d6",
          5786 => x"d80c883d",
          5787 => x"0d04f83d",
          5788 => x"0d7a7052",
          5789 => x"57fec03f",
          5790 => x"82d6d808",
          5791 => x"5882d6d8",
          5792 => x"08819138",
          5793 => x"76335574",
          5794 => x"832e0981",
          5795 => x"0680f038",
          5796 => x"84173359",
          5797 => x"78812e09",
          5798 => x"810680e3",
          5799 => x"38848053",
          5800 => x"82d6d808",
          5801 => x"52b81770",
          5802 => x"5256fcd3",
          5803 => x"3f82d4d5",
          5804 => x"5284b617",
          5805 => x"51fbd83f",
          5806 => x"848b85a4",
          5807 => x"d2527551",
          5808 => x"fbeb3f86",
          5809 => x"8a85e4f2",
          5810 => x"52849c17",
          5811 => x"51fbde3f",
          5812 => x"94170852",
          5813 => x"84a01751",
          5814 => x"fbd33f90",
          5815 => x"17085284",
          5816 => x"a41751fb",
          5817 => x"c83fa417",
          5818 => x"08810570",
          5819 => x"b4190c79",
          5820 => x"55537552",
          5821 => x"81173351",
          5822 => x"f7c43f77",
          5823 => x"84183480",
          5824 => x"53805281",
          5825 => x"173351f9",
          5826 => x"993f82d6",
          5827 => x"d808802e",
          5828 => x"83388158",
          5829 => x"7782d6d8",
          5830 => x"0c8a3d0d",
          5831 => x"04fb3d0d",
          5832 => x"77fe1a9c",
          5833 => x"1208fe05",
          5834 => x"55565480",
          5835 => x"56747327",
          5836 => x"8d388a14",
          5837 => x"22757129",
          5838 => x"b0160805",
          5839 => x"57537582",
          5840 => x"d6d80c87",
          5841 => x"3d0d04f9",
          5842 => x"3d0d7a7a",
          5843 => x"70085654",
          5844 => x"57817727",
          5845 => x"81df3876",
          5846 => x"9c150827",
          5847 => x"81d738ff",
          5848 => x"74335458",
          5849 => x"72822e80",
          5850 => x"f5387282",
          5851 => x"24893872",
          5852 => x"812e8d38",
          5853 => x"81bf3972",
          5854 => x"832e818e",
          5855 => x"3881b639",
          5856 => x"76812a17",
          5857 => x"70892aa8",
          5858 => x"16080553",
          5859 => x"745255fd",
          5860 => x"963f82d6",
          5861 => x"d808819f",
          5862 => x"387483ff",
          5863 => x"0614b811",
          5864 => x"33811770",
          5865 => x"892aa818",
          5866 => x"08055576",
          5867 => x"54575753",
          5868 => x"fcf53f82",
          5869 => x"d6d80880",
          5870 => x"fe387483",
          5871 => x"ff0614b8",
          5872 => x"11337088",
          5873 => x"2b780779",
          5874 => x"81067184",
          5875 => x"2a5c5258",
          5876 => x"51537280",
          5877 => x"e238759f",
          5878 => x"ff065880",
          5879 => x"da397688",
          5880 => x"2aa81508",
          5881 => x"05527351",
          5882 => x"fcbd3f82",
          5883 => x"d6d80880",
          5884 => x"c6387610",
          5885 => x"83fe0674",
          5886 => x"05b80551",
          5887 => x"f8cf3f82",
          5888 => x"d6d80883",
          5889 => x"ffff0658",
          5890 => x"ae397687",
          5891 => x"2aa81508",
          5892 => x"05527351",
          5893 => x"fc913f82",
          5894 => x"d6d8089b",
          5895 => x"3876822b",
          5896 => x"83fc0674",
          5897 => x"05b80551",
          5898 => x"f8ba3f82",
          5899 => x"d6d808f0",
          5900 => x"0a065883",
          5901 => x"39815877",
          5902 => x"82d6d80c",
          5903 => x"893d0d04",
          5904 => x"f83d0d7a",
          5905 => x"7c7e5a58",
          5906 => x"56825981",
          5907 => x"7727829e",
          5908 => x"38769c17",
          5909 => x"08278296",
          5910 => x"38753353",
          5911 => x"72792e81",
          5912 => x"9d387279",
          5913 => x"24893872",
          5914 => x"812e8d38",
          5915 => x"82803972",
          5916 => x"832e81b8",
          5917 => x"3881f739",
          5918 => x"76812a17",
          5919 => x"70892aa8",
          5920 => x"18080553",
          5921 => x"765255fb",
          5922 => x"9e3f82d6",
          5923 => x"d8085982",
          5924 => x"d6d80881",
          5925 => x"d9387483",
          5926 => x"ff0616b8",
          5927 => x"05811678",
          5928 => x"81065956",
          5929 => x"54775376",
          5930 => x"802e8f38",
          5931 => x"77842b9f",
          5932 => x"f0067433",
          5933 => x"8f067107",
          5934 => x"51537274",
          5935 => x"34810b83",
          5936 => x"17347489",
          5937 => x"2aa81708",
          5938 => x"05527551",
          5939 => x"fad93f82",
          5940 => x"d6d80859",
          5941 => x"82d6d808",
          5942 => x"81943874",
          5943 => x"83ff0616",
          5944 => x"b8057884",
          5945 => x"2a545476",
          5946 => x"8f387788",
          5947 => x"2a743381",
          5948 => x"f006718f",
          5949 => x"06075153",
          5950 => x"72743480",
          5951 => x"ec397688",
          5952 => x"2aa81708",
          5953 => x"05527551",
          5954 => x"fa9d3f82",
          5955 => x"d6d80859",
          5956 => x"82d6d808",
          5957 => x"80d83877",
          5958 => x"83ffff06",
          5959 => x"52761083",
          5960 => x"fe067605",
          5961 => x"b80551f6",
          5962 => x"e63fbe39",
          5963 => x"76872aa8",
          5964 => x"17080552",
          5965 => x"7551f9ef",
          5966 => x"3f82d6d8",
          5967 => x"085982d6",
          5968 => x"d808ab38",
          5969 => x"77f00a06",
          5970 => x"77822b83",
          5971 => x"fc067018",
          5972 => x"b8057054",
          5973 => x"515454f6",
          5974 => x"8b3f82d6",
          5975 => x"d8088f0a",
          5976 => x"06740752",
          5977 => x"7251f6c5",
          5978 => x"3f810b83",
          5979 => x"17347882",
          5980 => x"d6d80c8a",
          5981 => x"3d0d04f8",
          5982 => x"3d0d7a7c",
          5983 => x"7e720859",
          5984 => x"56565981",
          5985 => x"7527a438",
          5986 => x"749c1708",
          5987 => x"279d3873",
          5988 => x"802eaa38",
          5989 => x"ff537352",
          5990 => x"7551fda4",
          5991 => x"3f82d6d8",
          5992 => x"085482d6",
          5993 => x"d80880f2",
          5994 => x"38933982",
          5995 => x"5480eb39",
          5996 => x"815480e6",
          5997 => x"3982d6d8",
          5998 => x"085480de",
          5999 => x"39745278",
          6000 => x"51fb843f",
          6001 => x"82d6d808",
          6002 => x"5882d6d8",
          6003 => x"08802e80",
          6004 => x"c73882d6",
          6005 => x"d808812e",
          6006 => x"d23882d6",
          6007 => x"d808ff2e",
          6008 => x"cf388053",
          6009 => x"74527551",
          6010 => x"fcd63f82",
          6011 => x"d6d808c5",
          6012 => x"389c1608",
          6013 => x"fe119418",
          6014 => x"08575557",
          6015 => x"74742790",
          6016 => x"38811594",
          6017 => x"170c8416",
          6018 => x"33810754",
          6019 => x"73841734",
          6020 => x"77557678",
          6021 => x"26ffa638",
          6022 => x"80547382",
          6023 => x"d6d80c8a",
          6024 => x"3d0d04f6",
          6025 => x"3d0d7c7e",
          6026 => x"7108595b",
          6027 => x"5b799538",
          6028 => x"90170858",
          6029 => x"77802e88",
          6030 => x"389c1708",
          6031 => x"7826b238",
          6032 => x"8158ae39",
          6033 => x"79527a51",
          6034 => x"f9fd3f81",
          6035 => x"557482d6",
          6036 => x"d8082782",
          6037 => x"e03882d6",
          6038 => x"d8085582",
          6039 => x"d6d808ff",
          6040 => x"2e82d238",
          6041 => x"9c170882",
          6042 => x"d6d80826",
          6043 => x"82c73879",
          6044 => x"58941708",
          6045 => x"70565473",
          6046 => x"802e82b9",
          6047 => x"38777a2e",
          6048 => x"09810680",
          6049 => x"e238811a",
          6050 => x"569c1708",
          6051 => x"76268338",
          6052 => x"82567552",
          6053 => x"7a51f9af",
          6054 => x"3f805982",
          6055 => x"d6d80881",
          6056 => x"2e098106",
          6057 => x"863882d6",
          6058 => x"d8085982",
          6059 => x"d6d80809",
          6060 => x"70307072",
          6061 => x"07802570",
          6062 => x"7c0782d6",
          6063 => x"d8085451",
          6064 => x"51555573",
          6065 => x"81ef3882",
          6066 => x"d6d80880",
          6067 => x"2e953890",
          6068 => x"17085481",
          6069 => x"74279038",
          6070 => x"739c1808",
          6071 => x"27893873",
          6072 => x"58853975",
          6073 => x"80db3877",
          6074 => x"56811656",
          6075 => x"9c170876",
          6076 => x"26893882",
          6077 => x"56757826",
          6078 => x"81ac3875",
          6079 => x"527a51f8",
          6080 => x"c63f82d6",
          6081 => x"d808802e",
          6082 => x"b8388059",
          6083 => x"82d6d808",
          6084 => x"812e0981",
          6085 => x"06863882",
          6086 => x"d6d80859",
          6087 => x"82d6d808",
          6088 => x"09703070",
          6089 => x"72078025",
          6090 => x"707c0751",
          6091 => x"51555573",
          6092 => x"80f83875",
          6093 => x"782e0981",
          6094 => x"06ffae38",
          6095 => x"735580f5",
          6096 => x"39ff5375",
          6097 => x"527651f9",
          6098 => x"f73f82d6",
          6099 => x"d80882d6",
          6100 => x"d8083070",
          6101 => x"82d6d808",
          6102 => x"07802551",
          6103 => x"55557980",
          6104 => x"2e943873",
          6105 => x"802e8f38",
          6106 => x"75537952",
          6107 => x"7651f9d0",
          6108 => x"3f82d6d8",
          6109 => x"085574a5",
          6110 => x"38759018",
          6111 => x"0c9c1708",
          6112 => x"fe059418",
          6113 => x"08565474",
          6114 => x"74268638",
          6115 => x"ff159418",
          6116 => x"0c841733",
          6117 => x"81075473",
          6118 => x"84183497",
          6119 => x"39ff5674",
          6120 => x"812e9038",
          6121 => x"8c398055",
          6122 => x"8c3982d6",
          6123 => x"d8085585",
          6124 => x"39815675",
          6125 => x"557482d6",
          6126 => x"d80c8c3d",
          6127 => x"0d04f83d",
          6128 => x"0d7a7052",
          6129 => x"55f3f03f",
          6130 => x"82d6d808",
          6131 => x"58815682",
          6132 => x"d6d80880",
          6133 => x"d8387b52",
          6134 => x"7451f6c1",
          6135 => x"3f82d6d8",
          6136 => x"0882d6d8",
          6137 => x"08b4170c",
          6138 => x"59848053",
          6139 => x"7752b815",
          6140 => x"705257f2",
          6141 => x"8a3f7756",
          6142 => x"84398116",
          6143 => x"568a1522",
          6144 => x"58757827",
          6145 => x"97388154",
          6146 => x"75195376",
          6147 => x"52811533",
          6148 => x"51edab3f",
          6149 => x"82d6d808",
          6150 => x"802edf38",
          6151 => x"8a152276",
          6152 => x"32703070",
          6153 => x"7207709f",
          6154 => x"2a535156",
          6155 => x"567582d6",
          6156 => x"d80c8a3d",
          6157 => x"0d04f83d",
          6158 => x"0d7a7c71",
          6159 => x"08585657",
          6160 => x"74f0800a",
          6161 => x"2680f138",
          6162 => x"749f0653",
          6163 => x"7280e938",
          6164 => x"7490180c",
          6165 => x"88170854",
          6166 => x"73aa3875",
          6167 => x"33538273",
          6168 => x"278838ac",
          6169 => x"16085473",
          6170 => x"9b387485",
          6171 => x"2a53820b",
          6172 => x"8817225a",
          6173 => x"58727927",
          6174 => x"80fe38ac",
          6175 => x"16089818",
          6176 => x"0c80cd39",
          6177 => x"8a162270",
          6178 => x"892b5458",
          6179 => x"727526b2",
          6180 => x"38735276",
          6181 => x"51f5b03f",
          6182 => x"82d6d808",
          6183 => x"5482d6d8",
          6184 => x"08ff2ebd",
          6185 => x"38810b82",
          6186 => x"d6d80827",
          6187 => x"8b389c16",
          6188 => x"0882d6d8",
          6189 => x"08268538",
          6190 => x"8258bd39",
          6191 => x"74733155",
          6192 => x"cb397352",
          6193 => x"7551f4d5",
          6194 => x"3f82d6d8",
          6195 => x"0898180c",
          6196 => x"7394180c",
          6197 => x"98170853",
          6198 => x"82587280",
          6199 => x"2e9a3885",
          6200 => x"39815894",
          6201 => x"3974892a",
          6202 => x"1398180c",
          6203 => x"7483ff06",
          6204 => x"16b8059c",
          6205 => x"180c8058",
          6206 => x"7782d6d8",
          6207 => x"0c8a3d0d",
          6208 => x"04f83d0d",
          6209 => x"7a700890",
          6210 => x"1208a005",
          6211 => x"595754f0",
          6212 => x"800a7727",
          6213 => x"8638800b",
          6214 => x"98150c98",
          6215 => x"14085384",
          6216 => x"5572802e",
          6217 => x"81cb3876",
          6218 => x"83ff0658",
          6219 => x"7781b538",
          6220 => x"81139815",
          6221 => x"0c941408",
          6222 => x"55749238",
          6223 => x"76852a88",
          6224 => x"17225653",
          6225 => x"74732681",
          6226 => x"9b3880c0",
          6227 => x"398a1622",
          6228 => x"ff057789",
          6229 => x"2a065372",
          6230 => x"818a3874",
          6231 => x"527351f3",
          6232 => x"e63f82d6",
          6233 => x"d8085382",
          6234 => x"55810b82",
          6235 => x"d6d80827",
          6236 => x"80ff3881",
          6237 => x"5582d6d8",
          6238 => x"08ff2e80",
          6239 => x"f4389c16",
          6240 => x"0882d6d8",
          6241 => x"082680ca",
          6242 => x"387b8a38",
          6243 => x"7798150c",
          6244 => x"845580dd",
          6245 => x"39941408",
          6246 => x"527351f9",
          6247 => x"863f82d6",
          6248 => x"d8085387",
          6249 => x"5582d6d8",
          6250 => x"08802e80",
          6251 => x"c4388255",
          6252 => x"82d6d808",
          6253 => x"812eba38",
          6254 => x"815582d6",
          6255 => x"d808ff2e",
          6256 => x"b03882d6",
          6257 => x"d8085275",
          6258 => x"51fbf33f",
          6259 => x"82d6d808",
          6260 => x"a0387294",
          6261 => x"150c7252",
          6262 => x"7551f2c1",
          6263 => x"3f82d6d8",
          6264 => x"0898150c",
          6265 => x"7690150c",
          6266 => x"7716b805",
          6267 => x"9c150c80",
          6268 => x"557482d6",
          6269 => x"d80c8a3d",
          6270 => x"0d04f73d",
          6271 => x"0d7b7d71",
          6272 => x"085b5b57",
          6273 => x"80527651",
          6274 => x"fcac3f82",
          6275 => x"d6d80854",
          6276 => x"82d6d808",
          6277 => x"80ec3882",
          6278 => x"d6d80856",
          6279 => x"98170852",
          6280 => x"7851f083",
          6281 => x"3f82d6d8",
          6282 => x"085482d6",
          6283 => x"d80880d2",
          6284 => x"3882d6d8",
          6285 => x"089c1808",
          6286 => x"70335154",
          6287 => x"587281e5",
          6288 => x"2e098106",
          6289 => x"83388158",
          6290 => x"82d6d808",
          6291 => x"55728338",
          6292 => x"81557775",
          6293 => x"07537280",
          6294 => x"2e8e3881",
          6295 => x"1656757a",
          6296 => x"2e098106",
          6297 => x"8838a539",
          6298 => x"82d6d808",
          6299 => x"56815276",
          6300 => x"51fd8e3f",
          6301 => x"82d6d808",
          6302 => x"5482d6d8",
          6303 => x"08802eff",
          6304 => x"9b387384",
          6305 => x"2e098106",
          6306 => x"83388754",
          6307 => x"7382d6d8",
          6308 => x"0c8b3d0d",
          6309 => x"04fd3d0d",
          6310 => x"769a1152",
          6311 => x"54ebae3f",
          6312 => x"82d6d808",
          6313 => x"83ffff06",
          6314 => x"76703351",
          6315 => x"53537183",
          6316 => x"2e098106",
          6317 => x"90389414",
          6318 => x"51eb923f",
          6319 => x"82d6d808",
          6320 => x"902b7307",
          6321 => x"537282d6",
          6322 => x"d80c853d",
          6323 => x"0d04fc3d",
          6324 => x"0d777970",
          6325 => x"83ffff06",
          6326 => x"549a1253",
          6327 => x"5555ebaf",
          6328 => x"3f767033",
          6329 => x"51537283",
          6330 => x"2e098106",
          6331 => x"8b387390",
          6332 => x"2a529415",
          6333 => x"51eb983f",
          6334 => x"863d0d04",
          6335 => x"fd3d0d75",
          6336 => x"5480518b",
          6337 => x"5370812a",
          6338 => x"71818029",
          6339 => x"05747081",
          6340 => x"05563371",
          6341 => x"057081ff",
          6342 => x"06ff1656",
          6343 => x"51515172",
          6344 => x"e4387082",
          6345 => x"d6d80c85",
          6346 => x"3d0d04f2",
          6347 => x"3d0d6062",
          6348 => x"40598479",
          6349 => x"085f5b81",
          6350 => x"ff705d5d",
          6351 => x"98190880",
          6352 => x"2e838038",
          6353 => x"98190852",
          6354 => x"7d51eddb",
          6355 => x"3f82d6d8",
          6356 => x"085b82d6",
          6357 => x"d80882eb",
          6358 => x"389c1908",
          6359 => x"70335555",
          6360 => x"73863884",
          6361 => x"5b82dc39",
          6362 => x"8b1533bf",
          6363 => x"067081ff",
          6364 => x"06585372",
          6365 => x"861a3482",
          6366 => x"d6d80856",
          6367 => x"7381e52e",
          6368 => x"09810683",
          6369 => x"38815682",
          6370 => x"d6d80853",
          6371 => x"73ae2e09",
          6372 => x"81068338",
          6373 => x"81537573",
          6374 => x"07537299",
          6375 => x"3882d6d8",
          6376 => x"0877df06",
          6377 => x"54567288",
          6378 => x"2e098106",
          6379 => x"83388156",
          6380 => x"757f2e87",
          6381 => x"3881ff5c",
          6382 => x"81ef3976",
          6383 => x"8f2e0981",
          6384 => x"0681ca38",
          6385 => x"73862a70",
          6386 => x"81065153",
          6387 => x"72802e92",
          6388 => x"388d1533",
          6389 => x"7481bf06",
          6390 => x"70901c08",
          6391 => x"ac1d0c56",
          6392 => x"5d5d737c",
          6393 => x"2e098106",
          6394 => x"819c388d",
          6395 => x"1533537c",
          6396 => x"732e0981",
          6397 => x"06818f38",
          6398 => x"8c1e089a",
          6399 => x"16525ae8",
          6400 => x"cc3f82d6",
          6401 => x"d80883ff",
          6402 => x"ff065372",
          6403 => x"80f83874",
          6404 => x"337081bf",
          6405 => x"068d29f3",
          6406 => x"05515481",
          6407 => x"7b585882",
          6408 => x"c7d41733",
          6409 => x"750551e8",
          6410 => x"a43f82d6",
          6411 => x"d80883ff",
          6412 => x"ff065677",
          6413 => x"802e9638",
          6414 => x"7381fe26",
          6415 => x"80c83873",
          6416 => x"101a7659",
          6417 => x"53757323",
          6418 => x"8114548b",
          6419 => x"397583ff",
          6420 => x"ff2e0981",
          6421 => x"06b03881",
          6422 => x"17578c77",
          6423 => x"27c13874",
          6424 => x"3370862a",
          6425 => x"70810651",
          6426 => x"54557280",
          6427 => x"2e8e3873",
          6428 => x"81fe2692",
          6429 => x"3873101a",
          6430 => x"53807323",
          6431 => x"ff1c7081",
          6432 => x"ff065153",
          6433 => x"843981ff",
          6434 => x"53725c9d",
          6435 => x"397b9338",
          6436 => x"7451fce8",
          6437 => x"3f82d6d8",
          6438 => x"0881ff06",
          6439 => x"53727d2e",
          6440 => x"a738ff0b",
          6441 => x"ac1a0ca0",
          6442 => x"39805278",
          6443 => x"51f8d23f",
          6444 => x"82d6d808",
          6445 => x"5b82d6d8",
          6446 => x"08893898",
          6447 => x"1908fd84",
          6448 => x"38863980",
          6449 => x"0b981a0c",
          6450 => x"7a82d6d8",
          6451 => x"0c903d0d",
          6452 => x"04f23d0d",
          6453 => x"60700840",
          6454 => x"59805278",
          6455 => x"51f6d73f",
          6456 => x"82d6d808",
          6457 => x"5882d6d8",
          6458 => x"0883a438",
          6459 => x"81ff705f",
          6460 => x"5cff0bac",
          6461 => x"1a0c9819",
          6462 => x"08527e51",
          6463 => x"eaa93f82",
          6464 => x"d6d80858",
          6465 => x"82d6d808",
          6466 => x"8385389c",
          6467 => x"19087033",
          6468 => x"57577586",
          6469 => x"38845882",
          6470 => x"f6398b17",
          6471 => x"33bf0670",
          6472 => x"81ff0656",
          6473 => x"5473861a",
          6474 => x"347581e5",
          6475 => x"2e82c338",
          6476 => x"74832a70",
          6477 => x"81065154",
          6478 => x"748f2e8e",
          6479 => x"387382b2",
          6480 => x"38748f2e",
          6481 => x"09810681",
          6482 => x"f738ab19",
          6483 => x"3370862a",
          6484 => x"70810651",
          6485 => x"55557382",
          6486 => x"a1387586",
          6487 => x"2a708106",
          6488 => x"51547380",
          6489 => x"2e92388d",
          6490 => x"17337681",
          6491 => x"bf067090",
          6492 => x"1c08ac1d",
          6493 => x"0c585d5e",
          6494 => x"757c2e09",
          6495 => x"810681b9",
          6496 => x"388d1733",
          6497 => x"567d762e",
          6498 => x"09810681",
          6499 => x"ac388c1f",
          6500 => x"089a1852",
          6501 => x"5de5b63f",
          6502 => x"82d6d808",
          6503 => x"83ffff06",
          6504 => x"55748195",
          6505 => x"38763370",
          6506 => x"bf068d29",
          6507 => x"f3055956",
          6508 => x"81755c5a",
          6509 => x"82c7d41b",
          6510 => x"33770551",
          6511 => x"e58f3f82",
          6512 => x"d6d80883",
          6513 => x"ffff0656",
          6514 => x"79802eb1",
          6515 => x"387781fe",
          6516 => x"2680e638",
          6517 => x"755180df",
          6518 => x"b43f82d6",
          6519 => x"d8087810",
          6520 => x"1e702253",
          6521 => x"55811959",
          6522 => x"5580dfa1",
          6523 => x"3f7482d6",
          6524 => x"d8082e09",
          6525 => x"810680c1",
          6526 => x"38755a8b",
          6527 => x"397583ff",
          6528 => x"ff2e0981",
          6529 => x"06b33881",
          6530 => x"1b5b8c7b",
          6531 => x"27ffa538",
          6532 => x"76337086",
          6533 => x"2a708106",
          6534 => x"51555779",
          6535 => x"802e9038",
          6536 => x"73802e8b",
          6537 => x"3877101d",
          6538 => x"70225154",
          6539 => x"738b38ff",
          6540 => x"1c7081ff",
          6541 => x"06515484",
          6542 => x"3981ff54",
          6543 => x"735cbb39",
          6544 => x"7b933876",
          6545 => x"51f9b53f",
          6546 => x"82d6d808",
          6547 => x"81ff0654",
          6548 => x"737e2ebb",
          6549 => x"38ab1933",
          6550 => x"81065473",
          6551 => x"95388b53",
          6552 => x"a019529c",
          6553 => x"190851e5",
          6554 => x"b03f82d6",
          6555 => x"d808802e",
          6556 => x"9e3881ff",
          6557 => x"5cff0bac",
          6558 => x"1a0c8052",
          6559 => x"7851f581",
          6560 => x"3f82d6d8",
          6561 => x"085882d6",
          6562 => x"d808802e",
          6563 => x"fce83877",
          6564 => x"82d6d80c",
          6565 => x"903d0d04",
          6566 => x"ee3d0d64",
          6567 => x"7008ab12",
          6568 => x"3381a006",
          6569 => x"565d5a86",
          6570 => x"557385b5",
          6571 => x"38738c1d",
          6572 => x"08702256",
          6573 => x"565d7380",
          6574 => x"2e8d3881",
          6575 => x"1d701016",
          6576 => x"70225155",
          6577 => x"5df0398c",
          6578 => x"53a01a70",
          6579 => x"53923d70",
          6580 => x"535f59e4",
          6581 => x"873f0280",
          6582 => x"cb053381",
          6583 => x"06547380",
          6584 => x"2e82a838",
          6585 => x"80c00bab",
          6586 => x"1b34815b",
          6587 => x"8c1c087b",
          6588 => x"56588b53",
          6589 => x"7d527851",
          6590 => x"e3e23f85",
          6591 => x"7b2780c6",
          6592 => x"387a5677",
          6593 => x"227083ff",
          6594 => x"ff065555",
          6595 => x"73802eb4",
          6596 => x"387483ff",
          6597 => x"ff068219",
          6598 => x"59558f57",
          6599 => x"74810676",
          6600 => x"10077581",
          6601 => x"2a71902a",
          6602 => x"70810651",
          6603 => x"56565673",
          6604 => x"802e8738",
          6605 => x"7584a0a1",
          6606 => x"3256ff17",
          6607 => x"57768025",
          6608 => x"db38c039",
          6609 => x"75558702",
          6610 => x"8405bf05",
          6611 => x"575774b0",
          6612 => x"07bf0654",
          6613 => x"b9742784",
          6614 => x"38871454",
          6615 => x"737634ff",
          6616 => x"16ff1876",
          6617 => x"842a5758",
          6618 => x"5674e338",
          6619 => x"943dec05",
          6620 => x"175480fe",
          6621 => x"74348077",
          6622 => x"27b53878",
          6623 => x"335473a0",
          6624 => x"2ead3874",
          6625 => x"19703352",
          6626 => x"54e3e03f",
          6627 => x"82d6d808",
          6628 => x"802e8c38",
          6629 => x"ff175474",
          6630 => x"742e9438",
          6631 => x"81155581",
          6632 => x"15557477",
          6633 => x"27893874",
          6634 => x"19703351",
          6635 => x"54d03994",
          6636 => x"3d7705eb",
          6637 => x"05547815",
          6638 => x"81165658",
          6639 => x"a0567687",
          6640 => x"268a3881",
          6641 => x"17811570",
          6642 => x"33585557",
          6643 => x"75783487",
          6644 => x"7527e338",
          6645 => x"7951f9f9",
          6646 => x"3f82d6d8",
          6647 => x"088b3881",
          6648 => x"1b5b80e3",
          6649 => x"7b27fe84",
          6650 => x"3887557a",
          6651 => x"80e42e82",
          6652 => x"f03882d6",
          6653 => x"d8085582",
          6654 => x"d6d80884",
          6655 => x"2e098106",
          6656 => x"82df3802",
          6657 => x"80cb0533",
          6658 => x"ab1b3402",
          6659 => x"80cb0533",
          6660 => x"70812a70",
          6661 => x"81065155",
          6662 => x"5e815973",
          6663 => x"802e9038",
          6664 => x"8d528c1d",
          6665 => x"51fef886",
          6666 => x"3f82d6d8",
          6667 => x"08195978",
          6668 => x"527951f3",
          6669 => x"c53f82d6",
          6670 => x"d8085782",
          6671 => x"d6d80882",
          6672 => x"9e38ff19",
          6673 => x"5978802e",
          6674 => x"81d43878",
          6675 => x"852b901b",
          6676 => x"08713153",
          6677 => x"547951ef",
          6678 => x"dd3f82d6",
          6679 => x"d8085782",
          6680 => x"d6d80881",
          6681 => x"fa38a01a",
          6682 => x"51f5913f",
          6683 => x"82d6d808",
          6684 => x"81ff065d",
          6685 => x"981a0852",
          6686 => x"7b51e3ab",
          6687 => x"3f82d6d8",
          6688 => x"085782d6",
          6689 => x"d80881d7",
          6690 => x"388c1c08",
          6691 => x"9c1b087a",
          6692 => x"81ff065a",
          6693 => x"575b7c8d",
          6694 => x"17348f0b",
          6695 => x"8b173482",
          6696 => x"d6d8088c",
          6697 => x"173482d6",
          6698 => x"d808529a",
          6699 => x"1651dfdf",
          6700 => x"3f778d29",
          6701 => x"f3057755",
          6702 => x"557383ff",
          6703 => x"ff2e8b38",
          6704 => x"74101b70",
          6705 => x"22811757",
          6706 => x"51547352",
          6707 => x"82c7d417",
          6708 => x"33760551",
          6709 => x"dfb93f73",
          6710 => x"853883ff",
          6711 => x"ff548117",
          6712 => x"578c7727",
          6713 => x"d4387383",
          6714 => x"ffff2e8b",
          6715 => x"3874101b",
          6716 => x"70225154",
          6717 => x"73863877",
          6718 => x"80c00758",
          6719 => x"77763481",
          6720 => x"0b831d34",
          6721 => x"80527951",
          6722 => x"eff73f82",
          6723 => x"d6d80857",
          6724 => x"82d6d808",
          6725 => x"80c938ff",
          6726 => x"195978fe",
          6727 => x"d738981a",
          6728 => x"08527b51",
          6729 => x"e2813f82",
          6730 => x"d6d80857",
          6731 => x"82d6d808",
          6732 => x"ae38a053",
          6733 => x"82d6d808",
          6734 => x"529c1a08",
          6735 => x"51dfc03f",
          6736 => x"8b53a01a",
          6737 => x"529c1a08",
          6738 => x"51df913f",
          6739 => x"9c1a08ab",
          6740 => x"1b339806",
          6741 => x"5555738c",
          6742 => x"1634810b",
          6743 => x"831d3476",
          6744 => x"557482d6",
          6745 => x"d80c943d",
          6746 => x"0d04fa3d",
          6747 => x"0d787008",
          6748 => x"901208ac",
          6749 => x"13085659",
          6750 => x"575572ff",
          6751 => x"2e943872",
          6752 => x"527451ed",
          6753 => x"b13f82d6",
          6754 => x"d8085482",
          6755 => x"d6d80880",
          6756 => x"c9389815",
          6757 => x"08527551",
          6758 => x"e18d3f82",
          6759 => x"d6d80854",
          6760 => x"82d6d808",
          6761 => x"ab389c15",
          6762 => x"0853e573",
          6763 => x"34810b83",
          6764 => x"17349015",
          6765 => x"087727a2",
          6766 => x"3882d6d8",
          6767 => x"08527451",
          6768 => x"eebf3f82",
          6769 => x"d6d80854",
          6770 => x"82d6d808",
          6771 => x"802ec338",
          6772 => x"73842e09",
          6773 => x"81068338",
          6774 => x"82547382",
          6775 => x"d6d80c88",
          6776 => x"3d0d04f4",
          6777 => x"3d0d7e60",
          6778 => x"71085f59",
          6779 => x"5c800b96",
          6780 => x"1934981c",
          6781 => x"08802e83",
          6782 => x"e238ac1c",
          6783 => x"08ff2e81",
          6784 => x"bb388070",
          6785 => x"717f8c05",
          6786 => x"08702257",
          6787 => x"575b5c57",
          6788 => x"72772e81",
          6789 => x"9d387810",
          6790 => x"14702281",
          6791 => x"1b5b5653",
          6792 => x"7a973880",
          6793 => x"d0801570",
          6794 => x"83ffff06",
          6795 => x"5153728f",
          6796 => x"ff268638",
          6797 => x"745b80df",
          6798 => x"39761896",
          6799 => x"1181ff79",
          6800 => x"31585b54",
          6801 => x"83b5527a",
          6802 => x"902b7507",
          6803 => x"5180d598",
          6804 => x"3f82d6d8",
          6805 => x"0883ffff",
          6806 => x"065581ff",
          6807 => x"75279538",
          6808 => x"817627a5",
          6809 => x"3874882a",
          6810 => x"53727a34",
          6811 => x"74971534",
          6812 => x"82559f39",
          6813 => x"74307630",
          6814 => x"70780780",
          6815 => x"25728025",
          6816 => x"07525454",
          6817 => x"73802e85",
          6818 => x"3880579a",
          6819 => x"39747a34",
          6820 => x"81557417",
          6821 => x"57805b8c",
          6822 => x"1d087910",
          6823 => x"11702251",
          6824 => x"545472fe",
          6825 => x"f1387a30",
          6826 => x"70802570",
          6827 => x"30790659",
          6828 => x"51537717",
          6829 => x"94055380",
          6830 => x"0b821434",
          6831 => x"8070891a",
          6832 => x"585a579c",
          6833 => x"1c081970",
          6834 => x"33811b5b",
          6835 => x"565374a0",
          6836 => x"2eb73874",
          6837 => x"852e0981",
          6838 => x"06843881",
          6839 => x"e5557889",
          6840 => x"32703070",
          6841 => x"72078025",
          6842 => x"51545476",
          6843 => x"8b269038",
          6844 => x"72802e8b",
          6845 => x"38ae7670",
          6846 => x"81055834",
          6847 => x"81175774",
          6848 => x"76708105",
          6849 => x"58348117",
          6850 => x"578a7927",
          6851 => x"ffb53877",
          6852 => x"17880553",
          6853 => x"800b8114",
          6854 => x"34961833",
          6855 => x"53728187",
          6856 => x"38768b38",
          6857 => x"bf0b9619",
          6858 => x"34815780",
          6859 => x"e1397273",
          6860 => x"891a3355",
          6861 => x"5a577280",
          6862 => x"2e80d338",
          6863 => x"96188919",
          6864 => x"55567333",
          6865 => x"ffbf1154",
          6866 => x"55729926",
          6867 => x"aa389c1c",
          6868 => x"088c1133",
          6869 => x"51538879",
          6870 => x"27873872",
          6871 => x"842a5385",
          6872 => x"3972832a",
          6873 => x"53728106",
          6874 => x"5372802e",
          6875 => x"8a38a015",
          6876 => x"7083ffff",
          6877 => x"06565374",
          6878 => x"76708105",
          6879 => x"58348119",
          6880 => x"81158119",
          6881 => x"71335659",
          6882 => x"555972ff",
          6883 => x"b5387717",
          6884 => x"94055380",
          6885 => x"0b821434",
          6886 => x"9c1c088c",
          6887 => x"11335153",
          6888 => x"72853872",
          6889 => x"8919349c",
          6890 => x"1c08538b",
          6891 => x"13338819",
          6892 => x"349c1c08",
          6893 => x"9c115253",
          6894 => x"d9aa3f82",
          6895 => x"d6d80878",
          6896 => x"0c961351",
          6897 => x"d9873f82",
          6898 => x"d6d80886",
          6899 => x"19239813",
          6900 => x"51d8fa3f",
          6901 => x"82d6d808",
          6902 => x"8419238e",
          6903 => x"3d0d04f0",
          6904 => x"3d0d6270",
          6905 => x"08415e80",
          6906 => x"64703351",
          6907 => x"555573af",
          6908 => x"2e833881",
          6909 => x"557380dc",
          6910 => x"2e923874",
          6911 => x"802e8d38",
          6912 => x"7f980508",
          6913 => x"881f0caa",
          6914 => x"39811544",
          6915 => x"80647033",
          6916 => x"56565673",
          6917 => x"af2e0981",
          6918 => x"06833881",
          6919 => x"567380dc",
          6920 => x"32703070",
          6921 => x"80257807",
          6922 => x"51515473",
          6923 => x"dc387388",
          6924 => x"1f0c6370",
          6925 => x"33515473",
          6926 => x"9f269638",
          6927 => x"ff800bab",
          6928 => x"1f348052",
          6929 => x"7d51e7ee",
          6930 => x"3f82d6d8",
          6931 => x"085687e1",
          6932 => x"3963417d",
          6933 => x"088c1108",
          6934 => x"5b548059",
          6935 => x"923dfc05",
          6936 => x"51da8f3f",
          6937 => x"82d6d808",
          6938 => x"ff2e82b1",
          6939 => x"3883ffff",
          6940 => x"0b82d6d8",
          6941 => x"08279238",
          6942 => x"78101a82",
          6943 => x"d6d80890",
          6944 => x"2a555573",
          6945 => x"75238119",
          6946 => x"5982d6d8",
          6947 => x"0883ffff",
          6948 => x"0670af32",
          6949 => x"70309f73",
          6950 => x"27718025",
          6951 => x"07515155",
          6952 => x"5673b438",
          6953 => x"7580dc2e",
          6954 => x"ae387580",
          6955 => x"ff269138",
          6956 => x"755282c6",
          6957 => x"f051d992",
          6958 => x"3f82d6d8",
          6959 => x"0881de38",
          6960 => x"7881fe26",
          6961 => x"81d73878",
          6962 => x"101a5475",
          6963 => x"74238119",
          6964 => x"59ff8939",
          6965 => x"81154180",
          6966 => x"61703356",
          6967 => x"565773af",
          6968 => x"2e098106",
          6969 => x"83388157",
          6970 => x"7380dc32",
          6971 => x"70307080",
          6972 => x"25790751",
          6973 => x"515473dc",
          6974 => x"3874449f",
          6975 => x"7627822b",
          6976 => x"5778812e",
          6977 => x"0981068c",
          6978 => x"38792254",
          6979 => x"73ae2ea5",
          6980 => x"3880d239",
          6981 => x"78822e09",
          6982 => x"810680c9",
          6983 => x"38821a22",
          6984 => x"5473ae2e",
          6985 => x"09810680",
          6986 => x"c1387922",
          6987 => x"5473ae2e",
          6988 => x"098106b6",
          6989 => x"3878101a",
          6990 => x"54807423",
          6991 => x"800ba01f",
          6992 => x"5658ae54",
          6993 => x"78782683",
          6994 => x"38a05473",
          6995 => x"75708105",
          6996 => x"57348118",
          6997 => x"588a7827",
          6998 => x"e93876a0",
          6999 => x"075473ab",
          7000 => x"1f3484c4",
          7001 => x"3978802e",
          7002 => x"a8387810",
          7003 => x"1afe0555",
          7004 => x"7422fe16",
          7005 => x"7172a032",
          7006 => x"7030709f",
          7007 => x"2a515153",
          7008 => x"58565475",
          7009 => x"ae2e8438",
          7010 => x"738738ff",
          7011 => x"195978e0",
          7012 => x"3878197a",
          7013 => x"11555680",
          7014 => x"7423788d",
          7015 => x"38865685",
          7016 => x"90397683",
          7017 => x"07578399",
          7018 => x"39807a22",
          7019 => x"7083ffff",
          7020 => x"0656565d",
          7021 => x"73a02e09",
          7022 => x"81069338",
          7023 => x"811d7010",
          7024 => x"1b702251",
          7025 => x"555d73a0",
          7026 => x"2ef2387c",
          7027 => x"8f387483",
          7028 => x"ffff0654",
          7029 => x"73ae2e09",
          7030 => x"81068538",
          7031 => x"76830757",
          7032 => x"78802eaa",
          7033 => x"387916fe",
          7034 => x"05702251",
          7035 => x"5473ae2e",
          7036 => x"9d387810",
          7037 => x"1afe0555",
          7038 => x"ff195978",
          7039 => x"802e8f38",
          7040 => x"fe157022",
          7041 => x"555573ae",
          7042 => x"2e098106",
          7043 => x"eb388b53",
          7044 => x"a052a01e",
          7045 => x"51d5e83f",
          7046 => x"8070595c",
          7047 => x"885f7c10",
          7048 => x"1a702281",
          7049 => x"1f5f5754",
          7050 => x"75802e82",
          7051 => x"943875a0",
          7052 => x"2e963875",
          7053 => x"ae327030",
          7054 => x"70802551",
          7055 => x"51547c79",
          7056 => x"2e8c3873",
          7057 => x"802e8938",
          7058 => x"76830757",
          7059 => x"d1398054",
          7060 => x"735b7e78",
          7061 => x"26833881",
          7062 => x"5b7c7932",
          7063 => x"70307072",
          7064 => x"07802570",
          7065 => x"7e075151",
          7066 => x"55557380",
          7067 => x"2ea6387e",
          7068 => x"8b2efeae",
          7069 => x"387c792e",
          7070 => x"8b387683",
          7071 => x"07577c79",
          7072 => x"2681be38",
          7073 => x"785d8858",
          7074 => x"8b7c822b",
          7075 => x"81fc065d",
          7076 => x"5fff8b39",
          7077 => x"80ff7627",
          7078 => x"af387682",
          7079 => x"075783b5",
          7080 => x"52755180",
          7081 => x"ccc23f82",
          7082 => x"d6d80883",
          7083 => x"ffff0670",
          7084 => x"872a7081",
          7085 => x"06515556",
          7086 => x"73802e8c",
          7087 => x"387580ff",
          7088 => x"0682c7e4",
          7089 => x"11335754",
          7090 => x"81ff7627",
          7091 => x"a438ff1f",
          7092 => x"54737826",
          7093 => x"8a387683",
          7094 => x"077f5957",
          7095 => x"fec0397d",
          7096 => x"18a00576",
          7097 => x"882a5555",
          7098 => x"73753481",
          7099 => x"185880c3",
          7100 => x"3975802e",
          7101 => x"92387552",
          7102 => x"82c6fc51",
          7103 => x"d4cc3f82",
          7104 => x"d6d80880",
          7105 => x"2e8a3880",
          7106 => x"df778307",
          7107 => x"5856a439",
          7108 => x"ffbf1654",
          7109 => x"73992685",
          7110 => x"387b8207",
          7111 => x"5cff9f16",
          7112 => x"54739926",
          7113 => x"8e387b81",
          7114 => x"07e01770",
          7115 => x"83ffff06",
          7116 => x"58555c7d",
          7117 => x"18a00554",
          7118 => x"75743481",
          7119 => x"1858fdde",
          7120 => x"39a01e33",
          7121 => x"547381e5",
          7122 => x"2e098106",
          7123 => x"8638850b",
          7124 => x"a01f347e",
          7125 => x"882e0981",
          7126 => x"0688387b",
          7127 => x"822b81fc",
          7128 => x"065c7b8c",
          7129 => x"0654738c",
          7130 => x"2e8d387b",
          7131 => x"83065473",
          7132 => x"832e0981",
          7133 => x"06853876",
          7134 => x"82075776",
          7135 => x"812a7081",
          7136 => x"06515473",
          7137 => x"9f387b81",
          7138 => x"06547380",
          7139 => x"2e853876",
          7140 => x"9007577b",
          7141 => x"822a7081",
          7142 => x"06515473",
          7143 => x"802e8538",
          7144 => x"76880757",
          7145 => x"76ab1f34",
          7146 => x"7d51eaa5",
          7147 => x"3f82d6d8",
          7148 => x"08ab1f33",
          7149 => x"565682d6",
          7150 => x"d808802e",
          7151 => x"be3882d6",
          7152 => x"d808842e",
          7153 => x"09810680",
          7154 => x"e8387485",
          7155 => x"2a708106",
          7156 => x"76822a57",
          7157 => x"51547380",
          7158 => x"2e963874",
          7159 => x"81065473",
          7160 => x"802ef8ed",
          7161 => x"38ff800b",
          7162 => x"ab1f3480",
          7163 => x"5680c239",
          7164 => x"74810654",
          7165 => x"73bb3885",
          7166 => x"56b73974",
          7167 => x"822a7081",
          7168 => x"06515473",
          7169 => x"ac38861e",
          7170 => x"3370842a",
          7171 => x"70810651",
          7172 => x"55557380",
          7173 => x"2ee13890",
          7174 => x"1e0883ff",
          7175 => x"066005b8",
          7176 => x"05527f51",
          7177 => x"e4ef3f82",
          7178 => x"d6d80888",
          7179 => x"1f0cf8a1",
          7180 => x"397582d6",
          7181 => x"d80c923d",
          7182 => x"0d04f63d",
          7183 => x"0d7c5bff",
          7184 => x"7b087071",
          7185 => x"7355595c",
          7186 => x"55597380",
          7187 => x"2e81c638",
          7188 => x"75708105",
          7189 => x"5733709f",
          7190 => x"26525271",
          7191 => x"ba2e8d38",
          7192 => x"70ee3871",
          7193 => x"ba2e0981",
          7194 => x"0681a538",
          7195 => x"7333d011",
          7196 => x"7081ff06",
          7197 => x"51525370",
          7198 => x"89269138",
          7199 => x"82147381",
          7200 => x"ff06d005",
          7201 => x"56527176",
          7202 => x"2e80f738",
          7203 => x"800b82c7",
          7204 => x"c4595577",
          7205 => x"087a5557",
          7206 => x"76708105",
          7207 => x"58337470",
          7208 => x"81055633",
          7209 => x"ff9f1253",
          7210 => x"53537099",
          7211 => x"268938e0",
          7212 => x"137081ff",
          7213 => x"065451ff",
          7214 => x"9f125170",
          7215 => x"99268938",
          7216 => x"e0127081",
          7217 => x"ff065351",
          7218 => x"7230709f",
          7219 => x"2a515172",
          7220 => x"722e0981",
          7221 => x"06853870",
          7222 => x"ffbe3872",
          7223 => x"30747732",
          7224 => x"70307072",
          7225 => x"079f2a73",
          7226 => x"9f2a0753",
          7227 => x"54545170",
          7228 => x"802e8f38",
          7229 => x"81158419",
          7230 => x"59558375",
          7231 => x"25ff9438",
          7232 => x"8b397483",
          7233 => x"24863874",
          7234 => x"767c0c59",
          7235 => x"78518639",
          7236 => x"82eeb433",
          7237 => x"517082d6",
          7238 => x"d80c8c3d",
          7239 => x"0d04fa3d",
          7240 => x"0d785680",
          7241 => x"0b831734",
          7242 => x"ff0bb417",
          7243 => x"0c795275",
          7244 => x"51d1f43f",
          7245 => x"845582d6",
          7246 => x"d8088180",
          7247 => x"3884b616",
          7248 => x"51ce8a3f",
          7249 => x"82d6d808",
          7250 => x"83ffff06",
          7251 => x"54835573",
          7252 => x"82d4d52e",
          7253 => x"09810680",
          7254 => x"e338800b",
          7255 => x"b8173356",
          7256 => x"577481e9",
          7257 => x"2e098106",
          7258 => x"83388157",
          7259 => x"7481eb32",
          7260 => x"70307080",
          7261 => x"25790751",
          7262 => x"5154738a",
          7263 => x"387481e8",
          7264 => x"2e098106",
          7265 => x"b5388353",
          7266 => x"82c78452",
          7267 => x"80ee1651",
          7268 => x"cf873f82",
          7269 => x"d6d80855",
          7270 => x"82d6d808",
          7271 => x"802e9d38",
          7272 => x"855382c7",
          7273 => x"8852818a",
          7274 => x"1651ceed",
          7275 => x"3f82d6d8",
          7276 => x"085582d6",
          7277 => x"d808802e",
          7278 => x"83388255",
          7279 => x"7482d6d8",
          7280 => x"0c883d0d",
          7281 => x"04f23d0d",
          7282 => x"61028405",
          7283 => x"80cb0533",
          7284 => x"58558075",
          7285 => x"0c6051fc",
          7286 => x"e13f82d6",
          7287 => x"d808588b",
          7288 => x"56800b82",
          7289 => x"d6d80824",
          7290 => x"87843882",
          7291 => x"d6d80884",
          7292 => x"2982eea0",
          7293 => x"05700855",
          7294 => x"538c5673",
          7295 => x"802e86ee",
          7296 => x"3873750c",
          7297 => x"7681fe06",
          7298 => x"74335457",
          7299 => x"72802eae",
          7300 => x"38811433",
          7301 => x"51c6a03f",
          7302 => x"82d6d808",
          7303 => x"81ff0670",
          7304 => x"81065455",
          7305 => x"72983876",
          7306 => x"802e86c0",
          7307 => x"3874822a",
          7308 => x"70810651",
          7309 => x"538a5672",
          7310 => x"86b43886",
          7311 => x"af398074",
          7312 => x"34778115",
          7313 => x"34815281",
          7314 => x"143351c6",
          7315 => x"883f82d6",
          7316 => x"d80881ff",
          7317 => x"06708106",
          7318 => x"54558356",
          7319 => x"72868f38",
          7320 => x"76802e8f",
          7321 => x"3874822a",
          7322 => x"70810651",
          7323 => x"538a5672",
          7324 => x"85fc3880",
          7325 => x"70537452",
          7326 => x"5bfda33f",
          7327 => x"82d6d808",
          7328 => x"81ff0657",
          7329 => x"76822e09",
          7330 => x"810680e2",
          7331 => x"388c3d74",
          7332 => x"56588356",
          7333 => x"83fa1533",
          7334 => x"70585372",
          7335 => x"802e8d38",
          7336 => x"83fe1551",
          7337 => x"cbbe3f82",
          7338 => x"d6d80857",
          7339 => x"76787084",
          7340 => x"055a0cff",
          7341 => x"16901656",
          7342 => x"56758025",
          7343 => x"d738800b",
          7344 => x"8d3d5456",
          7345 => x"72708405",
          7346 => x"54085b83",
          7347 => x"577a802e",
          7348 => x"95387a52",
          7349 => x"7351fcc6",
          7350 => x"3f82d6d8",
          7351 => x"0881ff06",
          7352 => x"57817727",
          7353 => x"89388116",
          7354 => x"56837627",
          7355 => x"d7388156",
          7356 => x"76842e84",
          7357 => x"f9388d56",
          7358 => x"76812684",
          7359 => x"f13880c3",
          7360 => x"1451cac9",
          7361 => x"3f82d6d8",
          7362 => x"0883ffff",
          7363 => x"06537284",
          7364 => x"802e0981",
          7365 => x"0684d738",
          7366 => x"80ce1451",
          7367 => x"caaf3f82",
          7368 => x"d6d80883",
          7369 => x"ffff0658",
          7370 => x"778d3880",
          7371 => x"dc1451ca",
          7372 => x"b33f82d6",
          7373 => x"d8085877",
          7374 => x"a0150c80",
          7375 => x"c8143382",
          7376 => x"153480c8",
          7377 => x"1433ff11",
          7378 => x"7081ff06",
          7379 => x"5154558d",
          7380 => x"56728126",
          7381 => x"84983874",
          7382 => x"81ff0678",
          7383 => x"712980c5",
          7384 => x"16335259",
          7385 => x"53728a15",
          7386 => x"2372802e",
          7387 => x"8b38ff13",
          7388 => x"73065372",
          7389 => x"802e8638",
          7390 => x"8d5683f2",
          7391 => x"3980c914",
          7392 => x"51c9ca3f",
          7393 => x"82d6d808",
          7394 => x"5382d6d8",
          7395 => x"08881523",
          7396 => x"728f0657",
          7397 => x"8d567683",
          7398 => x"d53880cb",
          7399 => x"1451c9ad",
          7400 => x"3f82d6d8",
          7401 => x"0883ffff",
          7402 => x"0655748d",
          7403 => x"3880d814",
          7404 => x"51c9b13f",
          7405 => x"82d6d808",
          7406 => x"5580c614",
          7407 => x"51c98e3f",
          7408 => x"82d6d808",
          7409 => x"83ffff06",
          7410 => x"538d5672",
          7411 => x"802e839e",
          7412 => x"38881422",
          7413 => x"78147184",
          7414 => x"2a055a5a",
          7415 => x"78752683",
          7416 => x"8d388a14",
          7417 => x"22527479",
          7418 => x"3151fee0",
          7419 => x"c13f82d6",
          7420 => x"d8085582",
          7421 => x"d6d80880",
          7422 => x"2e82f338",
          7423 => x"82d6d808",
          7424 => x"80ffffff",
          7425 => x"f5268338",
          7426 => x"83577483",
          7427 => x"fff52683",
          7428 => x"38825774",
          7429 => x"9ff52685",
          7430 => x"38815789",
          7431 => x"398d5676",
          7432 => x"802e82ca",
          7433 => x"38821570",
          7434 => x"9c160c7b",
          7435 => x"a4160c73",
          7436 => x"1c70a817",
          7437 => x"0c7a1db0",
          7438 => x"170c5455",
          7439 => x"76832e09",
          7440 => x"8106af38",
          7441 => x"80e21451",
          7442 => x"c8833f82",
          7443 => x"d6d80883",
          7444 => x"ffff0653",
          7445 => x"8d567282",
          7446 => x"95387982",
          7447 => x"913880e4",
          7448 => x"1451c880",
          7449 => x"3f82d6d8",
          7450 => x"08ac150c",
          7451 => x"74822b53",
          7452 => x"a2398d56",
          7453 => x"79802e81",
          7454 => x"f5387713",
          7455 => x"ac150c74",
          7456 => x"15537682",
          7457 => x"2e8d3874",
          7458 => x"10157081",
          7459 => x"2a768106",
          7460 => x"05515383",
          7461 => x"ff13892a",
          7462 => x"538d5672",
          7463 => x"a0150826",
          7464 => x"81cc38ff",
          7465 => x"0b94150c",
          7466 => x"ff0b9015",
          7467 => x"0cff800b",
          7468 => x"84153476",
          7469 => x"832e0981",
          7470 => x"06819238",
          7471 => x"80e81451",
          7472 => x"c78b3f82",
          7473 => x"d6d80883",
          7474 => x"ffff0653",
          7475 => x"72812e09",
          7476 => x"810680f9",
          7477 => x"38811b52",
          7478 => x"7351cacb",
          7479 => x"3f82d6d8",
          7480 => x"0880ea38",
          7481 => x"82d6d808",
          7482 => x"84153484",
          7483 => x"b61451c6",
          7484 => x"dc3f82d6",
          7485 => x"d80883ff",
          7486 => x"ff065372",
          7487 => x"82d4d52e",
          7488 => x"09810680",
          7489 => x"c838b814",
          7490 => x"51c6d93f",
          7491 => x"82d6d808",
          7492 => x"848b85a4",
          7493 => x"d22e0981",
          7494 => x"06b33884",
          7495 => x"9c1451c6",
          7496 => x"c33f82d6",
          7497 => x"d808868a",
          7498 => x"85e4f22e",
          7499 => x"0981069d",
          7500 => x"3884a014",
          7501 => x"51c6ad3f",
          7502 => x"82d6d808",
          7503 => x"94150c84",
          7504 => x"a41451c6",
          7505 => x"9f3f82d6",
          7506 => x"d8089015",
          7507 => x"0c767434",
          7508 => x"82eeb022",
          7509 => x"81055372",
          7510 => x"82eeb023",
          7511 => x"72861523",
          7512 => x"82eeb80b",
          7513 => x"8c150c80",
          7514 => x"0b98150c",
          7515 => x"80567582",
          7516 => x"d6d80c90",
          7517 => x"3d0d04fb",
          7518 => x"3d0d7754",
          7519 => x"89557380",
          7520 => x"2eba3873",
          7521 => x"08537280",
          7522 => x"2eb23872",
          7523 => x"33527180",
          7524 => x"2eaa3886",
          7525 => x"13228415",
          7526 => x"22575271",
          7527 => x"762e0981",
          7528 => x"069a3881",
          7529 => x"133351ff",
          7530 => x"bf8d3f82",
          7531 => x"d6d80881",
          7532 => x"06527188",
          7533 => x"38717408",
          7534 => x"54558339",
          7535 => x"80537873",
          7536 => x"710c5274",
          7537 => x"82d6d80c",
          7538 => x"873d0d04",
          7539 => x"fa3d0d02",
          7540 => x"ab05337a",
          7541 => x"58893dfc",
          7542 => x"055256f4",
          7543 => x"dd3f8b54",
          7544 => x"800b82d6",
          7545 => x"d80824bc",
          7546 => x"3882d6d8",
          7547 => x"08842982",
          7548 => x"eea00570",
          7549 => x"08555573",
          7550 => x"802e8438",
          7551 => x"80743478",
          7552 => x"5473802e",
          7553 => x"84388074",
          7554 => x"3478750c",
          7555 => x"75547580",
          7556 => x"2e923880",
          7557 => x"53893d70",
          7558 => x"53840551",
          7559 => x"f7a73f82",
          7560 => x"d6d80854",
          7561 => x"7382d6d8",
          7562 => x"0c883d0d",
          7563 => x"04ea3d0d",
          7564 => x"68028405",
          7565 => x"80eb0533",
          7566 => x"59598954",
          7567 => x"78802e84",
          7568 => x"c83877bf",
          7569 => x"06705499",
          7570 => x"3dcc0553",
          7571 => x"9a3d8405",
          7572 => x"5258f6f1",
          7573 => x"3f82d6d8",
          7574 => x"085582d6",
          7575 => x"d80884a4",
          7576 => x"387a5c69",
          7577 => x"528c3d70",
          7578 => x"5256eaf3",
          7579 => x"3f82d6d8",
          7580 => x"085582d6",
          7581 => x"d8089238",
          7582 => x"0280d705",
          7583 => x"3370982b",
          7584 => x"55577380",
          7585 => x"25833886",
          7586 => x"55779c06",
          7587 => x"5473802e",
          7588 => x"81ab3874",
          7589 => x"802e9538",
          7590 => x"74842e09",
          7591 => x"8106aa38",
          7592 => x"7551dff4",
          7593 => x"3f82d6d8",
          7594 => x"08559e39",
          7595 => x"02b20533",
          7596 => x"91065473",
          7597 => x"81b83877",
          7598 => x"822a7081",
          7599 => x"06515473",
          7600 => x"802e8e38",
          7601 => x"885583bc",
          7602 => x"39778807",
          7603 => x"587483b4",
          7604 => x"3877832a",
          7605 => x"70810651",
          7606 => x"5473802e",
          7607 => x"81af3862",
          7608 => x"527a51d7",
          7609 => x"b03f82d6",
          7610 => x"d8085682",
          7611 => x"88b20a52",
          7612 => x"628e0551",
          7613 => x"c3b73f62",
          7614 => x"54a00b8b",
          7615 => x"15348053",
          7616 => x"62527a51",
          7617 => x"d7c83f80",
          7618 => x"52629c05",
          7619 => x"51c39e3f",
          7620 => x"7a54810b",
          7621 => x"83153475",
          7622 => x"802e80f1",
          7623 => x"387ab411",
          7624 => x"08515480",
          7625 => x"53755298",
          7626 => x"3dd00551",
          7627 => x"ccc93f82",
          7628 => x"d6d80855",
          7629 => x"82d6d808",
          7630 => x"82ca38b7",
          7631 => x"397482c4",
          7632 => x"3802b205",
          7633 => x"3370842a",
          7634 => x"70810651",
          7635 => x"55567380",
          7636 => x"2e863884",
          7637 => x"5582ad39",
          7638 => x"77812a70",
          7639 => x"81065154",
          7640 => x"73802ea9",
          7641 => x"38758106",
          7642 => x"5473802e",
          7643 => x"a0388755",
          7644 => x"82923973",
          7645 => x"527a51c5",
          7646 => x"ae3f82d6",
          7647 => x"d8087bff",
          7648 => x"1890120c",
          7649 => x"555582d6",
          7650 => x"d80881f8",
          7651 => x"3877832a",
          7652 => x"70810651",
          7653 => x"5473802e",
          7654 => x"86387780",
          7655 => x"c007587a",
          7656 => x"b41108a0",
          7657 => x"1b0c63a4",
          7658 => x"1b0c6353",
          7659 => x"705257d5",
          7660 => x"e43f82d6",
          7661 => x"d80882d6",
          7662 => x"d808881b",
          7663 => x"0c639c05",
          7664 => x"525ac1a0",
          7665 => x"3f82d6d8",
          7666 => x"0882d6d8",
          7667 => x"088c1b0c",
          7668 => x"777a0c56",
          7669 => x"86172284",
          7670 => x"1a237790",
          7671 => x"1a34800b",
          7672 => x"911a3480",
          7673 => x"0b9c1a0c",
          7674 => x"800b941a",
          7675 => x"0c77852a",
          7676 => x"70810651",
          7677 => x"5473802e",
          7678 => x"818d3882",
          7679 => x"d6d80880",
          7680 => x"2e818438",
          7681 => x"82d6d808",
          7682 => x"941a0c8a",
          7683 => x"17227089",
          7684 => x"2b7b5259",
          7685 => x"57a83976",
          7686 => x"527851c6",
          7687 => x"aa3f82d6",
          7688 => x"d8085782",
          7689 => x"d6d80881",
          7690 => x"26833882",
          7691 => x"5582d6d8",
          7692 => x"08ff2e09",
          7693 => x"81068338",
          7694 => x"79557578",
          7695 => x"31567430",
          7696 => x"70760780",
          7697 => x"25515477",
          7698 => x"76278a38",
          7699 => x"81707506",
          7700 => x"555a73c3",
          7701 => x"3876981a",
          7702 => x"0c74a938",
          7703 => x"7583ff06",
          7704 => x"5473802e",
          7705 => x"a2387652",
          7706 => x"7a51c5b1",
          7707 => x"3f82d6d8",
          7708 => x"08853882",
          7709 => x"558e3975",
          7710 => x"892a82d6",
          7711 => x"d808059c",
          7712 => x"1a0c8439",
          7713 => x"80790c74",
          7714 => x"547382d6",
          7715 => x"d80c983d",
          7716 => x"0d04f23d",
          7717 => x"0d606365",
          7718 => x"6440405d",
          7719 => x"59807e0c",
          7720 => x"903dfc05",
          7721 => x"527851f9",
          7722 => x"ce3f82d6",
          7723 => x"d8085582",
          7724 => x"d6d8088a",
          7725 => x"38911933",
          7726 => x"5574802e",
          7727 => x"86387456",
          7728 => x"82c73990",
          7729 => x"19338106",
          7730 => x"55875674",
          7731 => x"802e82b9",
          7732 => x"38953982",
          7733 => x"0b911a34",
          7734 => x"825682ad",
          7735 => x"39810b91",
          7736 => x"1a348156",
          7737 => x"82a3398c",
          7738 => x"1908941a",
          7739 => x"08315574",
          7740 => x"7c278338",
          7741 => x"745c7b80",
          7742 => x"2e828c38",
          7743 => x"94190870",
          7744 => x"83ff0656",
          7745 => x"567481b4",
          7746 => x"387e8a11",
          7747 => x"22ff0577",
          7748 => x"892a065b",
          7749 => x"5579a838",
          7750 => x"75873888",
          7751 => x"1908558f",
          7752 => x"39981908",
          7753 => x"527851c4",
          7754 => x"9e3f82d6",
          7755 => x"d8085581",
          7756 => x"7527ff9f",
          7757 => x"3874ff2e",
          7758 => x"ffa33874",
          7759 => x"981a0c98",
          7760 => x"1908527e",
          7761 => x"51c3d63f",
          7762 => x"82d6d808",
          7763 => x"802eff83",
          7764 => x"3882d6d8",
          7765 => x"081a7c89",
          7766 => x"2a595777",
          7767 => x"802e80d8",
          7768 => x"38771a7f",
          7769 => x"8a112258",
          7770 => x"5c557575",
          7771 => x"27853875",
          7772 => x"7a315877",
          7773 => x"5476537c",
          7774 => x"52811b33",
          7775 => x"51ffb8d4",
          7776 => x"3f82d6d8",
          7777 => x"08fed638",
          7778 => x"7e831133",
          7779 => x"56567480",
          7780 => x"2ea038b4",
          7781 => x"16087731",
          7782 => x"55747827",
          7783 => x"95388480",
          7784 => x"53b81652",
          7785 => x"b4160877",
          7786 => x"31892b7d",
          7787 => x"0551ffbe",
          7788 => x"ab3f7789",
          7789 => x"2b56ba39",
          7790 => x"769c1a0c",
          7791 => x"94190883",
          7792 => x"ff068480",
          7793 => x"71315755",
          7794 => x"7b762783",
          7795 => x"387b569c",
          7796 => x"1908527e",
          7797 => x"51c0d03f",
          7798 => x"82d6d808",
          7799 => x"fdff3875",
          7800 => x"53941908",
          7801 => x"83ff061f",
          7802 => x"b805527c",
          7803 => x"51ffbdec",
          7804 => x"3f7b7631",
          7805 => x"7e08177f",
          7806 => x"0c761e94",
          7807 => x"1b081894",
          7808 => x"1c0c5e5c",
          7809 => x"fdf03980",
          7810 => x"567582d6",
          7811 => x"d80c903d",
          7812 => x"0d04f23d",
          7813 => x"0d606365",
          7814 => x"6440405d",
          7815 => x"58807e0c",
          7816 => x"903dfc05",
          7817 => x"527751f6",
          7818 => x"ce3f82d6",
          7819 => x"d8085582",
          7820 => x"d6d8088a",
          7821 => x"38911833",
          7822 => x"5574802e",
          7823 => x"86387456",
          7824 => x"83be3990",
          7825 => x"18337081",
          7826 => x"2a708106",
          7827 => x"51565687",
          7828 => x"5674802e",
          7829 => x"83aa3895",
          7830 => x"39820b91",
          7831 => x"19348256",
          7832 => x"839e3981",
          7833 => x"0b911934",
          7834 => x"81568394",
          7835 => x"39941808",
          7836 => x"7c115656",
          7837 => x"74762784",
          7838 => x"3875095c",
          7839 => x"7b802e82",
          7840 => x"f2389418",
          7841 => x"087083ff",
          7842 => x"06565674",
          7843 => x"8281387e",
          7844 => x"8a1122ff",
          7845 => x"0577892a",
          7846 => x"065c557a",
          7847 => x"bf38758c",
          7848 => x"38881808",
          7849 => x"55749c38",
          7850 => x"7a528539",
          7851 => x"98180852",
          7852 => x"7751c6ef",
          7853 => x"3f82d6d8",
          7854 => x"085582d6",
          7855 => x"d808802e",
          7856 => x"82b13874",
          7857 => x"812eff91",
          7858 => x"3874ff2e",
          7859 => x"ff953874",
          7860 => x"98190c88",
          7861 => x"18088538",
          7862 => x"7488190c",
          7863 => x"7e55b415",
          7864 => x"089c1908",
          7865 => x"2e098106",
          7866 => x"8e387451",
          7867 => x"ffbdc83f",
          7868 => x"82d6d808",
          7869 => x"feed3898",
          7870 => x"1808527e",
          7871 => x"51c09e3f",
          7872 => x"82d6d808",
          7873 => x"802efed1",
          7874 => x"3882d6d8",
          7875 => x"081b7c89",
          7876 => x"2a5a5778",
          7877 => x"802e80d7",
          7878 => x"38781b7f",
          7879 => x"8a112258",
          7880 => x"5b557575",
          7881 => x"27853875",
          7882 => x"7b315978",
          7883 => x"5476537c",
          7884 => x"52811a33",
          7885 => x"51ffb786",
          7886 => x"3f82d6d8",
          7887 => x"08fea438",
          7888 => x"7eb41108",
          7889 => x"78315656",
          7890 => x"7479279c",
          7891 => x"38848053",
          7892 => x"b4160877",
          7893 => x"31892b7d",
          7894 => x"0552b816",
          7895 => x"51ffbafc",
          7896 => x"3f7e5580",
          7897 => x"0b831634",
          7898 => x"78892b56",
          7899 => x"80de398c",
          7900 => x"18089419",
          7901 => x"08269438",
          7902 => x"7e51ffbc",
          7903 => x"ba3f82d6",
          7904 => x"d808fddf",
          7905 => x"387e77b4",
          7906 => x"120c5576",
          7907 => x"9c190c94",
          7908 => x"180883ff",
          7909 => x"06848071",
          7910 => x"3157557b",
          7911 => x"76278338",
          7912 => x"7b569c18",
          7913 => x"08527e51",
          7914 => x"ffbcfc3f",
          7915 => x"82d6d808",
          7916 => x"fdb13875",
          7917 => x"537c5294",
          7918 => x"180883ff",
          7919 => x"061fb805",
          7920 => x"51ffba98",
          7921 => x"3f7e5581",
          7922 => x"0b831634",
          7923 => x"7b76317e",
          7924 => x"08177f0c",
          7925 => x"761e941a",
          7926 => x"08187094",
          7927 => x"1c0c8c1b",
          7928 => x"0858585e",
          7929 => x"5c747627",
          7930 => x"83387555",
          7931 => x"748c190c",
          7932 => x"fd8a3990",
          7933 => x"183380c0",
          7934 => x"07557490",
          7935 => x"19348056",
          7936 => x"7582d6d8",
          7937 => x"0c903d0d",
          7938 => x"04f83d0d",
          7939 => x"7a8b3dfc",
          7940 => x"05537052",
          7941 => x"56f2e03f",
          7942 => x"82d6d808",
          7943 => x"5782d6d8",
          7944 => x"08818038",
          7945 => x"90163370",
          7946 => x"862a7081",
          7947 => x"06515555",
          7948 => x"73802e80",
          7949 => x"ee38a016",
          7950 => x"08527851",
          7951 => x"ffbbe83f",
          7952 => x"82d6d808",
          7953 => x"5782d6d8",
          7954 => x"0880d838",
          7955 => x"a416088b",
          7956 => x"1133a007",
          7957 => x"5555738b",
          7958 => x"16348816",
          7959 => x"08537452",
          7960 => x"750851cc",
          7961 => x"e93f8c16",
          7962 => x"08529c15",
          7963 => x"51ffb8bd",
          7964 => x"3f8288b2",
          7965 => x"0a529615",
          7966 => x"51ffb8b1",
          7967 => x"3f765292",
          7968 => x"1551ffb8",
          7969 => x"8a3f7854",
          7970 => x"810b8315",
          7971 => x"347851ff",
          7972 => x"bbdc3f82",
          7973 => x"d6d80890",
          7974 => x"173381bf",
          7975 => x"06555773",
          7976 => x"90173476",
          7977 => x"82d6d80c",
          7978 => x"8a3d0d04",
          7979 => x"fc3d0d76",
          7980 => x"705254fe",
          7981 => x"d43f82d6",
          7982 => x"d8085382",
          7983 => x"d6d8089c",
          7984 => x"38863dfc",
          7985 => x"05527351",
          7986 => x"f1ad3f82",
          7987 => x"d6d80853",
          7988 => x"82d6d808",
          7989 => x"873882d6",
          7990 => x"d808740c",
          7991 => x"7282d6d8",
          7992 => x"0c863d0d",
          7993 => x"04ff3d0d",
          7994 => x"843d51e6",
          7995 => x"cd3f8b52",
          7996 => x"800b82d6",
          7997 => x"d808248b",
          7998 => x"3882d6d8",
          7999 => x"0882eeb4",
          8000 => x"34805271",
          8001 => x"82d6d80c",
          8002 => x"833d0d04",
          8003 => x"ee3d0d80",
          8004 => x"53943dcc",
          8005 => x"0552953d",
          8006 => x"51e9aa3f",
          8007 => x"82d6d808",
          8008 => x"5582d6d8",
          8009 => x"0880e038",
          8010 => x"76586452",
          8011 => x"943dd005",
          8012 => x"51ddac3f",
          8013 => x"82d6d808",
          8014 => x"5582d6d8",
          8015 => x"08bc3802",
          8016 => x"80c70533",
          8017 => x"70982b55",
          8018 => x"56738025",
          8019 => x"8938767a",
          8020 => x"98120c54",
          8021 => x"b23902a2",
          8022 => x"05337084",
          8023 => x"2a708106",
          8024 => x"51555673",
          8025 => x"802e9e38",
          8026 => x"767f5370",
          8027 => x"5254caa5",
          8028 => x"3f82d6d8",
          8029 => x"0898150c",
          8030 => x"8e3982d6",
          8031 => x"d808842e",
          8032 => x"09810683",
          8033 => x"38855574",
          8034 => x"82d6d80c",
          8035 => x"943d0d04",
          8036 => x"ffa33d0d",
          8037 => x"80e13d08",
          8038 => x"80e13d08",
          8039 => x"5b5b807a",
          8040 => x"34805380",
          8041 => x"df3dfdb4",
          8042 => x"055280e0",
          8043 => x"3d51e895",
          8044 => x"3f82d6d8",
          8045 => x"085782d6",
          8046 => x"d80883a1",
          8047 => x"387b80d4",
          8048 => x"3d0c7a7c",
          8049 => x"98110880",
          8050 => x"d83d0c55",
          8051 => x"5880d53d",
          8052 => x"08547380",
          8053 => x"2e828338",
          8054 => x"a05280d3",
          8055 => x"3d705255",
          8056 => x"c4d43f82",
          8057 => x"d6d80857",
          8058 => x"82d6d808",
          8059 => x"82ef3880",
          8060 => x"d93d0852",
          8061 => x"7b51ffb8",
          8062 => x"ae3f82d6",
          8063 => x"d8085782",
          8064 => x"d6d80882",
          8065 => x"d83880da",
          8066 => x"3d08527b",
          8067 => x"51c9863f",
          8068 => x"82d6d808",
          8069 => x"80d63d0c",
          8070 => x"76527451",
          8071 => x"c4983f82",
          8072 => x"d6d80857",
          8073 => x"82d6d808",
          8074 => x"82b33880",
          8075 => x"527451c9",
          8076 => x"fa3f82d6",
          8077 => x"d8085782",
          8078 => x"d6d808a7",
          8079 => x"3880da3d",
          8080 => x"08527b51",
          8081 => x"c8cf3f73",
          8082 => x"82d6d808",
          8083 => x"2ea63876",
          8084 => x"527451c5",
          8085 => x"ac3f82d6",
          8086 => x"d8085782",
          8087 => x"d6d80880",
          8088 => x"2ec93876",
          8089 => x"842e0981",
          8090 => x"06863882",
          8091 => x"5781ee39",
          8092 => x"7681ea38",
          8093 => x"80df3dfd",
          8094 => x"b8055274",
          8095 => x"51d6e43f",
          8096 => x"76933d78",
          8097 => x"11821133",
          8098 => x"51565a56",
          8099 => x"73802e92",
          8100 => x"380280c6",
          8101 => x"05558116",
          8102 => x"81167033",
          8103 => x"56565673",
          8104 => x"f5388116",
          8105 => x"54737826",
          8106 => x"81993875",
          8107 => x"802e9c38",
          8108 => x"78168205",
          8109 => x"55ff1880",
          8110 => x"e13d0811",
          8111 => x"ff18ff18",
          8112 => x"58585558",
          8113 => x"74337434",
          8114 => x"75eb38ff",
          8115 => x"1880e13d",
          8116 => x"08115558",
          8117 => x"af7434fd",
          8118 => x"f439777b",
          8119 => x"2e098106",
          8120 => x"8d38ff18",
          8121 => x"80e13d08",
          8122 => x"115558af",
          8123 => x"7434800b",
          8124 => x"82eeb433",
          8125 => x"70842982",
          8126 => x"c7c40570",
          8127 => x"08703352",
          8128 => x"5c565656",
          8129 => x"73762e8d",
          8130 => x"38811670",
          8131 => x"1a703351",
          8132 => x"555673f5",
          8133 => x"38821654",
          8134 => x"737826a7",
          8135 => x"38805574",
          8136 => x"76279138",
          8137 => x"74195473",
          8138 => x"337a7081",
          8139 => x"055c3481",
          8140 => x"1555ec39",
          8141 => x"ba7a7081",
          8142 => x"055c3474",
          8143 => x"ff2e0981",
          8144 => x"06853891",
          8145 => x"57973980",
          8146 => x"e03d0818",
          8147 => x"81195954",
          8148 => x"73337a70",
          8149 => x"81055c34",
          8150 => x"7a7826eb",
          8151 => x"38807a34",
          8152 => x"7682d6d8",
          8153 => x"0c80df3d",
          8154 => x"0d04f73d",
          8155 => x"0d7b7d8d",
          8156 => x"3dfc0554",
          8157 => x"71535755",
          8158 => x"ebfd3f82",
          8159 => x"d6d80853",
          8160 => x"82d6d808",
          8161 => x"82fe3891",
          8162 => x"15335372",
          8163 => x"82f6388c",
          8164 => x"15085473",
          8165 => x"76279238",
          8166 => x"90153370",
          8167 => x"812a7081",
          8168 => x"06515457",
          8169 => x"72833873",
          8170 => x"56941508",
          8171 => x"54807094",
          8172 => x"170c5875",
          8173 => x"782e829b",
          8174 => x"38798a11",
          8175 => x"2270892b",
          8176 => x"59515373",
          8177 => x"782eb738",
          8178 => x"7652ff16",
          8179 => x"51fec8de",
          8180 => x"3f82d6d8",
          8181 => x"08ff1578",
          8182 => x"54705355",
          8183 => x"53fec8ce",
          8184 => x"3f82d6d8",
          8185 => x"08732696",
          8186 => x"38763070",
          8187 => x"75067094",
          8188 => x"180c7771",
          8189 => x"31981808",
          8190 => x"57585153",
          8191 => x"b2398815",
          8192 => x"085473a7",
          8193 => x"38735274",
          8194 => x"51ffbc97",
          8195 => x"3f82d6d8",
          8196 => x"085482d6",
          8197 => x"d808812e",
          8198 => x"819d3882",
          8199 => x"d6d808ff",
          8200 => x"2e819e38",
          8201 => x"82d6d808",
          8202 => x"88160c73",
          8203 => x"98160c73",
          8204 => x"802e819f",
          8205 => x"38767627",
          8206 => x"80de3875",
          8207 => x"77319416",
          8208 => x"08189417",
          8209 => x"0c901633",
          8210 => x"70812a70",
          8211 => x"81065155",
          8212 => x"5a567280",
          8213 => x"2e9b3873",
          8214 => x"527451ff",
          8215 => x"bbc53f82",
          8216 => x"d6d80854",
          8217 => x"82d6d808",
          8218 => x"953882d6",
          8219 => x"d80856a8",
          8220 => x"39735274",
          8221 => x"51ffb5cf",
          8222 => x"3f82d6d8",
          8223 => x"085473ff",
          8224 => x"2ebf3881",
          8225 => x"7427b038",
          8226 => x"7953739c",
          8227 => x"140827a7",
          8228 => x"38739816",
          8229 => x"0cff9e39",
          8230 => x"94150816",
          8231 => x"94160c75",
          8232 => x"83ff0653",
          8233 => x"72802eab",
          8234 => x"38735279",
          8235 => x"51ffb4ed",
          8236 => x"3f82d6d8",
          8237 => x"08943882",
          8238 => x"0b911634",
          8239 => x"825380c4",
          8240 => x"39810b91",
          8241 => x"16348153",
          8242 => x"bb397589",
          8243 => x"2a82d6d8",
          8244 => x"08055894",
          8245 => x"1508548c",
          8246 => x"15087427",
          8247 => x"9038738c",
          8248 => x"160c9015",
          8249 => x"3380c007",
          8250 => x"53729016",
          8251 => x"347383ff",
          8252 => x"06537280",
          8253 => x"2e8c3877",
          8254 => x"9c16082e",
          8255 => x"8538779c",
          8256 => x"160c8053",
          8257 => x"7282d6d8",
          8258 => x"0c8b3d0d",
          8259 => x"04f93d0d",
          8260 => x"79568954",
          8261 => x"75802e81",
          8262 => x"8b388053",
          8263 => x"893dfc05",
          8264 => x"528a3d84",
          8265 => x"0551e19d",
          8266 => x"3f82d6d8",
          8267 => x"085582d6",
          8268 => x"d80880eb",
          8269 => x"3877760c",
          8270 => x"7a527551",
          8271 => x"d5a13f82",
          8272 => x"d6d80855",
          8273 => x"82d6d808",
          8274 => x"80c438ab",
          8275 => x"16337098",
          8276 => x"2b555780",
          8277 => x"7424a238",
          8278 => x"86163370",
          8279 => x"842a7081",
          8280 => x"06515557",
          8281 => x"73802eae",
          8282 => x"389c1608",
          8283 => x"527751c2",
          8284 => x"a43f82d6",
          8285 => x"d8088817",
          8286 => x"0c775486",
          8287 => x"14228417",
          8288 => x"23745275",
          8289 => x"51ffbdae",
          8290 => x"3f82d6d8",
          8291 => x"08557484",
          8292 => x"2e098106",
          8293 => x"85388555",
          8294 => x"86397480",
          8295 => x"2e843880",
          8296 => x"760c7454",
          8297 => x"7382d6d8",
          8298 => x"0c893d0d",
          8299 => x"04fc3d0d",
          8300 => x"76873dfc",
          8301 => x"05537052",
          8302 => x"53e7bc3f",
          8303 => x"82d6d808",
          8304 => x"873882d6",
          8305 => x"d808730c",
          8306 => x"863d0d04",
          8307 => x"fb3d0d77",
          8308 => x"79893dfc",
          8309 => x"05547153",
          8310 => x"5654e79b",
          8311 => x"3f82d6d8",
          8312 => x"085382d6",
          8313 => x"d80880e1",
          8314 => x"38749438",
          8315 => x"82d6d808",
          8316 => x"527351ff",
          8317 => x"bcc03f82",
          8318 => x"d6d80853",
          8319 => x"80cb3982",
          8320 => x"d6d80852",
          8321 => x"7351c2a3",
          8322 => x"3f82d6d8",
          8323 => x"085382d6",
          8324 => x"d808842e",
          8325 => x"09810685",
          8326 => x"38805387",
          8327 => x"3982d6d8",
          8328 => x"08a73874",
          8329 => x"527351cf",
          8330 => x"ba3f7252",
          8331 => x"7351ffbd",
          8332 => x"d03f82d6",
          8333 => x"d8088432",
          8334 => x"70307072",
          8335 => x"079f2c70",
          8336 => x"82d6d808",
          8337 => x"06515154",
          8338 => x"547282d6",
          8339 => x"d80c873d",
          8340 => x"0d04ed3d",
          8341 => x"0d665780",
          8342 => x"53893d70",
          8343 => x"53973d52",
          8344 => x"56dee23f",
          8345 => x"82d6d808",
          8346 => x"5582d6d8",
          8347 => x"08b23865",
          8348 => x"527551d2",
          8349 => x"ea3f82d6",
          8350 => x"d8085582",
          8351 => x"d6d808a0",
          8352 => x"380280cb",
          8353 => x"05337098",
          8354 => x"2b555873",
          8355 => x"80258538",
          8356 => x"86558d39",
          8357 => x"76802e88",
          8358 => x"38765275",
          8359 => x"51cec43f",
          8360 => x"7482d6d8",
          8361 => x"0c953d0d",
          8362 => x"04f03d0d",
          8363 => x"6365555c",
          8364 => x"8053923d",
          8365 => x"ec055293",
          8366 => x"3d51de89",
          8367 => x"3f82d6d8",
          8368 => x"085b82d6",
          8369 => x"d8088282",
          8370 => x"387c740c",
          8371 => x"73089c11",
          8372 => x"08fe1194",
          8373 => x"13085956",
          8374 => x"58557574",
          8375 => x"26913875",
          8376 => x"7c0c81e6",
          8377 => x"39815b81",
          8378 => x"ce39825b",
          8379 => x"81c93982",
          8380 => x"d6d80875",
          8381 => x"33555973",
          8382 => x"812e0981",
          8383 => x"0680c038",
          8384 => x"82755f57",
          8385 => x"7652923d",
          8386 => x"f00551ff",
          8387 => x"b0b93f82",
          8388 => x"d6d808ff",
          8389 => x"2ecf3882",
          8390 => x"d6d80881",
          8391 => x"2ecc3882",
          8392 => x"d6d80830",
          8393 => x"7082d6d8",
          8394 => x"08078025",
          8395 => x"7a058119",
          8396 => x"7f53595a",
          8397 => x"549c1408",
          8398 => x"7726c938",
          8399 => x"80f939a8",
          8400 => x"150882d6",
          8401 => x"d8085758",
          8402 => x"75983877",
          8403 => x"5281187d",
          8404 => x"5258ffad",
          8405 => x"d23f82d6",
          8406 => x"d8085b82",
          8407 => x"d6d80880",
          8408 => x"d6387c70",
          8409 => x"337712ff",
          8410 => x"1a5d5256",
          8411 => x"5474822e",
          8412 => x"0981069e",
          8413 => x"38b81451",
          8414 => x"ffa9d23f",
          8415 => x"82d6d808",
          8416 => x"83ffff06",
          8417 => x"70307080",
          8418 => x"251b8219",
          8419 => x"595b5154",
          8420 => x"9b39b814",
          8421 => x"51ffa9cc",
          8422 => x"3f82d6d8",
          8423 => x"08f00a06",
          8424 => x"70307080",
          8425 => x"251b8419",
          8426 => x"595b5154",
          8427 => x"7583ff06",
          8428 => x"7a585679",
          8429 => x"ff923878",
          8430 => x"7c0c7c79",
          8431 => x"94120c84",
          8432 => x"11338107",
          8433 => x"56547484",
          8434 => x"15347a82",
          8435 => x"d6d80c92",
          8436 => x"3d0d04f9",
          8437 => x"3d0d798a",
          8438 => x"3dfc0553",
          8439 => x"705257e3",
          8440 => x"963f82d6",
          8441 => x"d8085682",
          8442 => x"d6d80881",
          8443 => x"aa389117",
          8444 => x"33567581",
          8445 => x"a2389017",
          8446 => x"3370812a",
          8447 => x"70810651",
          8448 => x"55558755",
          8449 => x"73802e81",
          8450 => x"90389417",
          8451 => x"0854738c",
          8452 => x"18082781",
          8453 => x"8238739c",
          8454 => x"3882d6d8",
          8455 => x"08538817",
          8456 => x"08527651",
          8457 => x"ffb2d03f",
          8458 => x"82d6d808",
          8459 => x"7488190c",
          8460 => x"5680ca39",
          8461 => x"98170852",
          8462 => x"7651ffae",
          8463 => x"8a3f82d6",
          8464 => x"d808ff2e",
          8465 => x"09810683",
          8466 => x"38815682",
          8467 => x"d6d80881",
          8468 => x"2e098106",
          8469 => x"85388256",
          8470 => x"a43975a1",
          8471 => x"38775482",
          8472 => x"d6d8089c",
          8473 => x"15082795",
          8474 => x"38981708",
          8475 => x"5382d6d8",
          8476 => x"08527651",
          8477 => x"ffb2803f",
          8478 => x"82d6d808",
          8479 => x"56941708",
          8480 => x"8c180c90",
          8481 => x"173380c0",
          8482 => x"07547390",
          8483 => x"18347580",
          8484 => x"2e853875",
          8485 => x"91183475",
          8486 => x"557482d6",
          8487 => x"d80c893d",
          8488 => x"0d04e03d",
          8489 => x"0d8253a2",
          8490 => x"3dff9c05",
          8491 => x"52a33d51",
          8492 => x"da933f82",
          8493 => x"d6d80855",
          8494 => x"82d6d808",
          8495 => x"81f93878",
          8496 => x"46a33d08",
          8497 => x"52963d70",
          8498 => x"5258ce93",
          8499 => x"3f82d6d8",
          8500 => x"085582d6",
          8501 => x"d80881df",
          8502 => x"380280ff",
          8503 => x"05337085",
          8504 => x"2a708106",
          8505 => x"51555686",
          8506 => x"557381cb",
          8507 => x"3875982b",
          8508 => x"54807424",
          8509 => x"81c13802",
          8510 => x"80da0533",
          8511 => x"70810658",
          8512 => x"54875576",
          8513 => x"81b1386c",
          8514 => x"527851ff",
          8515 => x"bb873f82",
          8516 => x"d6d80874",
          8517 => x"842a7081",
          8518 => x"06515556",
          8519 => x"73802e80",
          8520 => x"d6387854",
          8521 => x"82d6d808",
          8522 => x"9815082e",
          8523 => x"81893873",
          8524 => x"5a82d6d8",
          8525 => x"085c7652",
          8526 => x"8a3d7052",
          8527 => x"54ffb5f6",
          8528 => x"3f82d6d8",
          8529 => x"085582d6",
          8530 => x"d80880eb",
          8531 => x"3882d6d8",
          8532 => x"08527351",
          8533 => x"ffbbd43f",
          8534 => x"82d6d808",
          8535 => x"5582d6d8",
          8536 => x"08863887",
          8537 => x"5580d039",
          8538 => x"82d6d808",
          8539 => x"842e8838",
          8540 => x"82d6d808",
          8541 => x"80c13877",
          8542 => x"51c7ef3f",
          8543 => x"82d6d808",
          8544 => x"82d6d808",
          8545 => x"307082d6",
          8546 => x"d8080780",
          8547 => x"25515555",
          8548 => x"75802e95",
          8549 => x"3873802e",
          8550 => x"90388053",
          8551 => x"75527751",
          8552 => x"ffafd43f",
          8553 => x"82d6d808",
          8554 => x"55748c38",
          8555 => x"7851ffa9",
          8556 => x"bd3f82d6",
          8557 => x"d8085574",
          8558 => x"82d6d80c",
          8559 => x"a23d0d04",
          8560 => x"e83d0d82",
          8561 => x"539a3dff",
          8562 => x"bc05529b",
          8563 => x"3d51d7f5",
          8564 => x"3f82d6d8",
          8565 => x"085482d6",
          8566 => x"d80882b7",
          8567 => x"38785e6a",
          8568 => x"528e3d70",
          8569 => x"5258cbf7",
          8570 => x"3f82d6d8",
          8571 => x"085482d6",
          8572 => x"d8088638",
          8573 => x"8854829b",
          8574 => x"3982d6d8",
          8575 => x"08842e09",
          8576 => x"8106828f",
          8577 => x"380280df",
          8578 => x"05337085",
          8579 => x"2a810651",
          8580 => x"55865474",
          8581 => x"81fd3878",
          8582 => x"5a74528a",
          8583 => x"3d705257",
          8584 => x"ffb0803f",
          8585 => x"82d6d808",
          8586 => x"75555682",
          8587 => x"d6d80883",
          8588 => x"38875482",
          8589 => x"d6d80881",
          8590 => x"2e098106",
          8591 => x"83388254",
          8592 => x"82d6d808",
          8593 => x"ff2e0981",
          8594 => x"06863881",
          8595 => x"5481ba39",
          8596 => x"7381b638",
          8597 => x"82d6d808",
          8598 => x"527851ff",
          8599 => x"b2e03f82",
          8600 => x"d6d80854",
          8601 => x"82d6d808",
          8602 => x"819f388b",
          8603 => x"53a052b8",
          8604 => x"1951ffa5",
          8605 => x"8a3f7854",
          8606 => x"ae0bb815",
          8607 => x"34785490",
          8608 => x"0b80c315",
          8609 => x"348288b2",
          8610 => x"0a5280ce",
          8611 => x"1951ffa4",
          8612 => x"9c3f7553",
          8613 => x"78b81153",
          8614 => x"51ffb8b2",
          8615 => x"3fa05378",
          8616 => x"b8115380",
          8617 => x"d80551ff",
          8618 => x"a4b23f78",
          8619 => x"54ae0b80",
          8620 => x"d915347f",
          8621 => x"537880d8",
          8622 => x"115351ff",
          8623 => x"b8903f78",
          8624 => x"54810b83",
          8625 => x"15347751",
          8626 => x"ffbfcd3f",
          8627 => x"82d6d808",
          8628 => x"5482d6d8",
          8629 => x"08b33882",
          8630 => x"88b20a52",
          8631 => x"64960551",
          8632 => x"ffa3ca3f",
          8633 => x"75536452",
          8634 => x"7851ffb7",
          8635 => x"e13f6454",
          8636 => x"900b8b15",
          8637 => x"34785481",
          8638 => x"0b831534",
          8639 => x"7851ffa6",
          8640 => x"ed3f82d6",
          8641 => x"d808548b",
          8642 => x"39805375",
          8643 => x"527651ff",
          8644 => x"ace53f73",
          8645 => x"82d6d80c",
          8646 => x"9a3d0d04",
          8647 => x"d83d0dab",
          8648 => x"3d840551",
          8649 => x"d2943f82",
          8650 => x"53aa3dfe",
          8651 => x"fc0552ab",
          8652 => x"3d51d591",
          8653 => x"3f82d6d8",
          8654 => x"085582d6",
          8655 => x"d80882d8",
          8656 => x"38784eab",
          8657 => x"3d08529e",
          8658 => x"3d705258",
          8659 => x"c9913f82",
          8660 => x"d6d80855",
          8661 => x"82d6d808",
          8662 => x"82be3802",
          8663 => x"819f0533",
          8664 => x"81a00654",
          8665 => x"86557382",
          8666 => x"af38a053",
          8667 => x"a53d0852",
          8668 => x"aa3dff80",
          8669 => x"0551ffa2",
          8670 => x"e33fb053",
          8671 => x"7752923d",
          8672 => x"705254ff",
          8673 => x"a2d63fac",
          8674 => x"3d085273",
          8675 => x"51c8d03f",
          8676 => x"82d6d808",
          8677 => x"5582d6d8",
          8678 => x"08973863",
          8679 => x"a13d082e",
          8680 => x"09810688",
          8681 => x"3865a33d",
          8682 => x"082e9238",
          8683 => x"885581e8",
          8684 => x"3982d6d8",
          8685 => x"08842e09",
          8686 => x"810681bb",
          8687 => x"387351ff",
          8688 => x"bdd63f82",
          8689 => x"d6d80855",
          8690 => x"82d6d808",
          8691 => x"81ca3868",
          8692 => x"569353aa",
          8693 => x"3dff8d05",
          8694 => x"528d1651",
          8695 => x"ffa1fd3f",
          8696 => x"02af0533",
          8697 => x"8b17348b",
          8698 => x"16337084",
          8699 => x"2a708106",
          8700 => x"51555573",
          8701 => x"893874a0",
          8702 => x"0754738b",
          8703 => x"17347854",
          8704 => x"810b8315",
          8705 => x"348b1633",
          8706 => x"70842a70",
          8707 => x"81065155",
          8708 => x"5573802e",
          8709 => x"80e7386f",
          8710 => x"642e80e1",
          8711 => x"38755278",
          8712 => x"51ffb4f1",
          8713 => x"3f82d6d8",
          8714 => x"08527851",
          8715 => x"ffa5ee3f",
          8716 => x"825582d6",
          8717 => x"d808802e",
          8718 => x"80de3882",
          8719 => x"d6d80852",
          8720 => x"7851ffa3",
          8721 => x"e23f82d6",
          8722 => x"d8087980",
          8723 => x"d8115858",
          8724 => x"5582d6d8",
          8725 => x"0880c138",
          8726 => x"81163354",
          8727 => x"73ae2e09",
          8728 => x"81069a38",
          8729 => x"63537552",
          8730 => x"7651ffb4",
          8731 => x"e13f7854",
          8732 => x"810b8315",
          8733 => x"34873982",
          8734 => x"d6d8089c",
          8735 => x"387751c1",
          8736 => x"e93f82d6",
          8737 => x"d8085582",
          8738 => x"d6d8088c",
          8739 => x"387851ff",
          8740 => x"a3dc3f82",
          8741 => x"d6d80855",
          8742 => x"7482d6d8",
          8743 => x"0caa3d0d",
          8744 => x"04ec3d0d",
          8745 => x"0280df05",
          8746 => x"33028405",
          8747 => x"80e30533",
          8748 => x"57578253",
          8749 => x"963dcc05",
          8750 => x"52973d51",
          8751 => x"d2873f82",
          8752 => x"d6d80855",
          8753 => x"82d6d808",
          8754 => x"80cf3878",
          8755 => x"5a665296",
          8756 => x"3dd00551",
          8757 => x"c6893f82",
          8758 => x"d6d80855",
          8759 => x"82d6d808",
          8760 => x"b8380280",
          8761 => x"cf053381",
          8762 => x"a0065486",
          8763 => x"5573aa38",
          8764 => x"75a70661",
          8765 => x"71098b12",
          8766 => x"3371067a",
          8767 => x"74060751",
          8768 => x"57555674",
          8769 => x"8b153478",
          8770 => x"54810b83",
          8771 => x"15347851",
          8772 => x"ffa2db3f",
          8773 => x"82d6d808",
          8774 => x"557482d6",
          8775 => x"d80c963d",
          8776 => x"0d04ee3d",
          8777 => x"0d655682",
          8778 => x"53943dcc",
          8779 => x"0552953d",
          8780 => x"51d1923f",
          8781 => x"82d6d808",
          8782 => x"5582d6d8",
          8783 => x"0880cb38",
          8784 => x"76586452",
          8785 => x"943dd005",
          8786 => x"51c5943f",
          8787 => x"82d6d808",
          8788 => x"5582d6d8",
          8789 => x"08b43802",
          8790 => x"80c70533",
          8791 => x"81a00654",
          8792 => x"865573a6",
          8793 => x"38841622",
          8794 => x"86172271",
          8795 => x"902b0753",
          8796 => x"54961f51",
          8797 => x"ff9eb63f",
          8798 => x"7654810b",
          8799 => x"83153476",
          8800 => x"51ffa1ea",
          8801 => x"3f82d6d8",
          8802 => x"08557482",
          8803 => x"d6d80c94",
          8804 => x"3d0d04e9",
          8805 => x"3d0d6a6c",
          8806 => x"5c5a8053",
          8807 => x"993dcc05",
          8808 => x"529a3d51",
          8809 => x"d09f3f82",
          8810 => x"d6d80882",
          8811 => x"d6d80830",
          8812 => x"7082d6d8",
          8813 => x"08078025",
          8814 => x"51555779",
          8815 => x"802e8186",
          8816 => x"38817075",
          8817 => x"06555573",
          8818 => x"802e80fa",
          8819 => x"387b5d80",
          8820 => x"5f80528d",
          8821 => x"3d705254",
          8822 => x"ffacdb3f",
          8823 => x"82d6d808",
          8824 => x"5782d6d8",
          8825 => x"0880d238",
          8826 => x"74527351",
          8827 => x"ffb2bc3f",
          8828 => x"82d6d808",
          8829 => x"5782d6d8",
          8830 => x"08bf3882",
          8831 => x"d6d80882",
          8832 => x"d6d80865",
          8833 => x"5b595678",
          8834 => x"1881197b",
          8835 => x"18565955",
          8836 => x"74337434",
          8837 => x"8116568a",
          8838 => x"7827ec38",
          8839 => x"8b56751a",
          8840 => x"54807434",
          8841 => x"75802e9e",
          8842 => x"38ff1670",
          8843 => x"1b703351",
          8844 => x"555673a0",
          8845 => x"2ee8388e",
          8846 => x"3976842e",
          8847 => x"09810686",
          8848 => x"38807a34",
          8849 => x"80577630",
          8850 => x"70780780",
          8851 => x"2551547a",
          8852 => x"802e80c1",
          8853 => x"3873802e",
          8854 => x"bc387ba4",
          8855 => x"11085351",
          8856 => x"ff9fc43f",
          8857 => x"82d6d808",
          8858 => x"5782d6d8",
          8859 => x"08a7387b",
          8860 => x"70335555",
          8861 => x"80c35673",
          8862 => x"832e8b38",
          8863 => x"80e45673",
          8864 => x"842e8338",
          8865 => x"a7567515",
          8866 => x"b80551ff",
          8867 => x"9bd63f82",
          8868 => x"d6d8087b",
          8869 => x"0c7682d6",
          8870 => x"d80c993d",
          8871 => x"0d04e63d",
          8872 => x"0d82539c",
          8873 => x"3dffb405",
          8874 => x"529d3d51",
          8875 => x"ce973f82",
          8876 => x"d6d80882",
          8877 => x"d6d80856",
          8878 => x"5482d6d8",
          8879 => x"0882dd38",
          8880 => x"8b53a052",
          8881 => x"8a3d7052",
          8882 => x"58ff9cb3",
          8883 => x"3f736d70",
          8884 => x"33515556",
          8885 => x"9f742781",
          8886 => x"86387757",
          8887 => x"9d3d51ff",
          8888 => x"9d903f82",
          8889 => x"d6d80883",
          8890 => x"ffff2680",
          8891 => x"c43882d6",
          8892 => x"d8085195",
          8893 => x"983f83b5",
          8894 => x"5282d6d8",
          8895 => x"085193e8",
          8896 => x"3f82d6d8",
          8897 => x"0883ffff",
          8898 => x"06557480",
          8899 => x"2ea33874",
          8900 => x"5282c8e4",
          8901 => x"51ff9cb2",
          8902 => x"3f82d6d8",
          8903 => x"08933881",
          8904 => x"ff752788",
          8905 => x"38758926",
          8906 => x"88388b39",
          8907 => x"8a762786",
          8908 => x"38865581",
          8909 => x"e73981ff",
          8910 => x"75278f38",
          8911 => x"74882a54",
          8912 => x"73777081",
          8913 => x"05593481",
          8914 => x"16567477",
          8915 => x"70810559",
          8916 => x"3481166d",
          8917 => x"70335155",
          8918 => x"56739f26",
          8919 => x"fefe388a",
          8920 => x"3d335486",
          8921 => x"557381e5",
          8922 => x"2e81b138",
          8923 => x"75802e99",
          8924 => x"3802a305",
          8925 => x"55751570",
          8926 => x"33515473",
          8927 => x"a02e0981",
          8928 => x"068738ff",
          8929 => x"165675ed",
          8930 => x"38784080",
          8931 => x"42805290",
          8932 => x"3d705255",
          8933 => x"ffa99f3f",
          8934 => x"82d6d808",
          8935 => x"5482d6d8",
          8936 => x"0880f738",
          8937 => x"81527451",
          8938 => x"ffaf803f",
          8939 => x"82d6d808",
          8940 => x"5482d6d8",
          8941 => x"088d3875",
          8942 => x"80c43866",
          8943 => x"54e57434",
          8944 => x"80c63982",
          8945 => x"d6d80884",
          8946 => x"2e098106",
          8947 => x"80cc3880",
          8948 => x"5475742e",
          8949 => x"80c43881",
          8950 => x"527451ff",
          8951 => x"ac9c3f82",
          8952 => x"d6d80854",
          8953 => x"82d6d808",
          8954 => x"b138a053",
          8955 => x"82d6d808",
          8956 => x"526651ff",
          8957 => x"9a893f66",
          8958 => x"54880b8b",
          8959 => x"15348b53",
          8960 => x"77526651",
          8961 => x"ff99d53f",
          8962 => x"7854810b",
          8963 => x"83153478",
          8964 => x"51ff9cda",
          8965 => x"3f82d6d8",
          8966 => x"08547355",
          8967 => x"7482d6d8",
          8968 => x"0c9c3d0d",
          8969 => x"04f23d0d",
          8970 => x"60620288",
          8971 => x"0580cb05",
          8972 => x"33933dfc",
          8973 => x"05557254",
          8974 => x"405e5ad2",
          8975 => x"ba3f82d6",
          8976 => x"d8085882",
          8977 => x"d6d80882",
          8978 => x"bd38911a",
          8979 => x"33587782",
          8980 => x"b5387c80",
          8981 => x"2e97388c",
          8982 => x"1a085978",
          8983 => x"9038901a",
          8984 => x"3370812a",
          8985 => x"70810651",
          8986 => x"55557390",
          8987 => x"38875482",
          8988 => x"97398258",
          8989 => x"82903981",
          8990 => x"58828b39",
          8991 => x"7e8a1122",
          8992 => x"70892b70",
          8993 => x"557f5456",
          8994 => x"5656feaf",
          8995 => x"a13fff14",
          8996 => x"7d067030",
          8997 => x"7072079f",
          8998 => x"2a82d6d8",
          8999 => x"08059019",
          9000 => x"087c405a",
          9001 => x"5d555581",
          9002 => x"77278838",
          9003 => x"9c160877",
          9004 => x"26833882",
          9005 => x"57767756",
          9006 => x"59805674",
          9007 => x"527951ff",
          9008 => x"9d853f81",
          9009 => x"157f5555",
          9010 => x"9c140875",
          9011 => x"26833882",
          9012 => x"5582d6d8",
          9013 => x"08812eff",
          9014 => x"993882d6",
          9015 => x"d808ff2e",
          9016 => x"ff953882",
          9017 => x"d6d8088e",
          9018 => x"38811656",
          9019 => x"757b2e09",
          9020 => x"81068738",
          9021 => x"93397459",
          9022 => x"80567477",
          9023 => x"2e098106",
          9024 => x"ffb93887",
          9025 => x"5880ff39",
          9026 => x"7d802eba",
          9027 => x"38787b55",
          9028 => x"557a802e",
          9029 => x"b4388115",
          9030 => x"5673812e",
          9031 => x"09810683",
          9032 => x"38ff5675",
          9033 => x"5374527e",
          9034 => x"51ff9e94",
          9035 => x"3f82d6d8",
          9036 => x"085882d6",
          9037 => x"d80880ce",
          9038 => x"38748116",
          9039 => x"ff165656",
          9040 => x"5c73d338",
          9041 => x"8439ff19",
          9042 => x"5c7e7c90",
          9043 => x"120c557d",
          9044 => x"802eb338",
          9045 => x"78881b0c",
          9046 => x"7c8c1b0c",
          9047 => x"901a3380",
          9048 => x"c0075473",
          9049 => x"901b349c",
          9050 => x"1508fe05",
          9051 => x"94160857",
          9052 => x"54757426",
          9053 => x"9138757b",
          9054 => x"3194160c",
          9055 => x"84153381",
          9056 => x"07547384",
          9057 => x"16347754",
          9058 => x"7382d6d8",
          9059 => x"0c903d0d",
          9060 => x"04e93d0d",
          9061 => x"6b6d0288",
          9062 => x"0580eb05",
          9063 => x"339d3d54",
          9064 => x"5a5c59c5",
          9065 => x"953f8b56",
          9066 => x"800b82d6",
          9067 => x"d808248b",
          9068 => x"f83882d6",
          9069 => x"d8088429",
          9070 => x"82eea005",
          9071 => x"70085155",
          9072 => x"74802e84",
          9073 => x"38807534",
          9074 => x"82d6d808",
          9075 => x"81ff065f",
          9076 => x"81527e51",
          9077 => x"ff8efe3f",
          9078 => x"82d6d808",
          9079 => x"81ff0670",
          9080 => x"81065657",
          9081 => x"8356748b",
          9082 => x"c0387682",
          9083 => x"2a708106",
          9084 => x"51558a56",
          9085 => x"748bb238",
          9086 => x"993dfc05",
          9087 => x"5383527e",
          9088 => x"51ff939e",
          9089 => x"3f82d6d8",
          9090 => x"08993867",
          9091 => x"5574802e",
          9092 => x"92387482",
          9093 => x"8080268b",
          9094 => x"38ff1575",
          9095 => x"06557480",
          9096 => x"2e833881",
          9097 => x"4878802e",
          9098 => x"87388480",
          9099 => x"79269238",
          9100 => x"7881800a",
          9101 => x"268b38ff",
          9102 => x"19790655",
          9103 => x"74802e86",
          9104 => x"3893568a",
          9105 => x"e4397889",
          9106 => x"2a6e892a",
          9107 => x"70892b77",
          9108 => x"59484359",
          9109 => x"7a833881",
          9110 => x"56613070",
          9111 => x"80257707",
          9112 => x"51559156",
          9113 => x"748ac238",
          9114 => x"993df805",
          9115 => x"5381527e",
          9116 => x"51ff92ae",
          9117 => x"3f815682",
          9118 => x"d6d8088a",
          9119 => x"ac387783",
          9120 => x"2a707706",
          9121 => x"82d6d808",
          9122 => x"43564574",
          9123 => x"8338bf41",
          9124 => x"66558e56",
          9125 => x"6075268a",
          9126 => x"90387461",
          9127 => x"31704855",
          9128 => x"80ff7527",
          9129 => x"8a833893",
          9130 => x"56788180",
          9131 => x"2689fa38",
          9132 => x"77812a70",
          9133 => x"81065643",
          9134 => x"74802e95",
          9135 => x"38778706",
          9136 => x"5574822e",
          9137 => x"838d3877",
          9138 => x"81065574",
          9139 => x"802e8383",
          9140 => x"38778106",
          9141 => x"55935682",
          9142 => x"5e74802e",
          9143 => x"89cb3878",
          9144 => x"5a7d832e",
          9145 => x"09810680",
          9146 => x"e13878ae",
          9147 => x"3866912a",
          9148 => x"57810b82",
          9149 => x"c9882256",
          9150 => x"5a74802e",
          9151 => x"9d387477",
          9152 => x"26983882",
          9153 => x"c9885679",
          9154 => x"10821770",
          9155 => x"2257575a",
          9156 => x"74802e86",
          9157 => x"38767527",
          9158 => x"ee387952",
          9159 => x"6651feaa",
          9160 => x"8d3f82d6",
          9161 => x"d8088429",
          9162 => x"84870570",
          9163 => x"892a5e55",
          9164 => x"a05c800b",
          9165 => x"82d6d808",
          9166 => x"fc808a05",
          9167 => x"5644fdff",
          9168 => x"f00a7527",
          9169 => x"80ec3888",
          9170 => x"d33978ae",
          9171 => x"38668c2a",
          9172 => x"57810b82",
          9173 => x"c8f82256",
          9174 => x"5a74802e",
          9175 => x"9d387477",
          9176 => x"26983882",
          9177 => x"c8f85679",
          9178 => x"10821770",
          9179 => x"2257575a",
          9180 => x"74802e86",
          9181 => x"38767527",
          9182 => x"ee387952",
          9183 => x"6651fea9",
          9184 => x"ad3f82d6",
          9185 => x"d8081084",
          9186 => x"055782d6",
          9187 => x"d8089ff5",
          9188 => x"26963881",
          9189 => x"0b82d6d8",
          9190 => x"081082d6",
          9191 => x"d8080571",
          9192 => x"11722a83",
          9193 => x"0559565e",
          9194 => x"83ff1789",
          9195 => x"2a5d815c",
          9196 => x"a044601c",
          9197 => x"7d116505",
          9198 => x"697012ff",
          9199 => x"05713070",
          9200 => x"72067431",
          9201 => x"5c525957",
          9202 => x"59407d83",
          9203 => x"2e098106",
          9204 => x"8938761c",
          9205 => x"6018415c",
          9206 => x"8439761d",
          9207 => x"5d799029",
          9208 => x"18706231",
          9209 => x"68585155",
          9210 => x"74762687",
          9211 => x"af38757c",
          9212 => x"317d317a",
          9213 => x"53706531",
          9214 => x"5255fea8",
          9215 => x"b13f82d6",
          9216 => x"d808587d",
          9217 => x"832e0981",
          9218 => x"069b3882",
          9219 => x"d6d80883",
          9220 => x"fff52680",
          9221 => x"dd387887",
          9222 => x"83387981",
          9223 => x"2a5978fd",
          9224 => x"be3886f8",
          9225 => x"397d822e",
          9226 => x"09810680",
          9227 => x"c53883ff",
          9228 => x"f50b82d6",
          9229 => x"d80827a0",
          9230 => x"38788f38",
          9231 => x"791a5574",
          9232 => x"80c02686",
          9233 => x"387459fd",
          9234 => x"96396281",
          9235 => x"06557480",
          9236 => x"2e8f3883",
          9237 => x"5efd8839",
          9238 => x"82d6d808",
          9239 => x"9ff52692",
          9240 => x"387886b8",
          9241 => x"38791a59",
          9242 => x"81807927",
          9243 => x"fcf13886",
          9244 => x"ab398055",
          9245 => x"7d812e09",
          9246 => x"81068338",
          9247 => x"7d559ff5",
          9248 => x"78278b38",
          9249 => x"74810655",
          9250 => x"8e567486",
          9251 => x"9c388480",
          9252 => x"5380527a",
          9253 => x"51ff90e7",
          9254 => x"3f8b5382",
          9255 => x"c790527a",
          9256 => x"51ff90b8",
          9257 => x"3f848052",
          9258 => x"8b1b51ff",
          9259 => x"8fe13f79",
          9260 => x"8d1c347b",
          9261 => x"83ffff06",
          9262 => x"528e1b51",
          9263 => x"ff8fd03f",
          9264 => x"810b901c",
          9265 => x"347d8332",
          9266 => x"70307096",
          9267 => x"2a848006",
          9268 => x"54515591",
          9269 => x"1b51ff8f",
          9270 => x"b63f6655",
          9271 => x"7483ffff",
          9272 => x"26903874",
          9273 => x"83ffff06",
          9274 => x"52931b51",
          9275 => x"ff8fa03f",
          9276 => x"8a397452",
          9277 => x"a01b51ff",
          9278 => x"8fb33ff8",
          9279 => x"0b951c34",
          9280 => x"bf52981b",
          9281 => x"51ff8f87",
          9282 => x"3f81ff52",
          9283 => x"9a1b51ff",
          9284 => x"8efd3f60",
          9285 => x"529c1b51",
          9286 => x"ff8f923f",
          9287 => x"7d832e09",
          9288 => x"810680cb",
          9289 => x"388288b2",
          9290 => x"0a5280c3",
          9291 => x"1b51ff8e",
          9292 => x"fc3f7c52",
          9293 => x"a41b51ff",
          9294 => x"8ef33f82",
          9295 => x"52ac1b51",
          9296 => x"ff8eea3f",
          9297 => x"8152b01b",
          9298 => x"51ff8ec3",
          9299 => x"3f8652b2",
          9300 => x"1b51ff8e",
          9301 => x"ba3fff80",
          9302 => x"0b80c01c",
          9303 => x"34a90b80",
          9304 => x"c21c3493",
          9305 => x"5382c79c",
          9306 => x"5280c71b",
          9307 => x"51ae3982",
          9308 => x"88b20a52",
          9309 => x"a71b51ff",
          9310 => x"8eb33f7c",
          9311 => x"83ffff06",
          9312 => x"52961b51",
          9313 => x"ff8e883f",
          9314 => x"ff800ba4",
          9315 => x"1c34a90b",
          9316 => x"a61c3493",
          9317 => x"5382c7b0",
          9318 => x"52ab1b51",
          9319 => x"ff8ebd3f",
          9320 => x"82d4d552",
          9321 => x"83fe1b70",
          9322 => x"5259ff8d",
          9323 => x"e23f8154",
          9324 => x"60537a52",
          9325 => x"7e51ff8a",
          9326 => x"853f8156",
          9327 => x"82d6d808",
          9328 => x"83e7387d",
          9329 => x"832e0981",
          9330 => x"0680ee38",
          9331 => x"75546086",
          9332 => x"05537a52",
          9333 => x"7e51ff89",
          9334 => x"e53f8480",
          9335 => x"5380527a",
          9336 => x"51ff8e9b",
          9337 => x"3f848b85",
          9338 => x"a4d2527a",
          9339 => x"51ff8dbd",
          9340 => x"3f868a85",
          9341 => x"e4f25283",
          9342 => x"e41b51ff",
          9343 => x"8daf3fff",
          9344 => x"185283e8",
          9345 => x"1b51ff8d",
          9346 => x"a43f8252",
          9347 => x"83ec1b51",
          9348 => x"ff8d9a3f",
          9349 => x"82d4d552",
          9350 => x"7851ff8c",
          9351 => x"f23f7554",
          9352 => x"60870553",
          9353 => x"7a527e51",
          9354 => x"ff89933f",
          9355 => x"75546016",
          9356 => x"537a527e",
          9357 => x"51ff8986",
          9358 => x"3f655380",
          9359 => x"527a51ff",
          9360 => x"8dbd3f7f",
          9361 => x"5680587d",
          9362 => x"832e0981",
          9363 => x"069a38f8",
          9364 => x"527a51ff",
          9365 => x"8cd73fff",
          9366 => x"52841b51",
          9367 => x"ff8cce3f",
          9368 => x"f00a5288",
          9369 => x"1b519139",
          9370 => x"87fffff8",
          9371 => x"557d812e",
          9372 => x"8338f855",
          9373 => x"74527a51",
          9374 => x"ff8cb23f",
          9375 => x"7c556157",
          9376 => x"74622683",
          9377 => x"38745776",
          9378 => x"5475537a",
          9379 => x"527e51ff",
          9380 => x"88ac3f82",
          9381 => x"d6d80882",
          9382 => x"87388480",
          9383 => x"5382d6d8",
          9384 => x"08527a51",
          9385 => x"ff8cd83f",
          9386 => x"76167578",
          9387 => x"31565674",
          9388 => x"cd388118",
          9389 => x"5877802e",
          9390 => x"ff8d3879",
          9391 => x"557d832e",
          9392 => x"83386355",
          9393 => x"61577462",
          9394 => x"26833874",
          9395 => x"57765475",
          9396 => x"537a527e",
          9397 => x"51ff87e6",
          9398 => x"3f82d6d8",
          9399 => x"0881c138",
          9400 => x"76167578",
          9401 => x"31565674",
          9402 => x"db388c56",
          9403 => x"7d832e93",
          9404 => x"38865666",
          9405 => x"83ffff26",
          9406 => x"8a388456",
          9407 => x"7d822e83",
          9408 => x"38815664",
          9409 => x"81065877",
          9410 => x"80fe3884",
          9411 => x"80537752",
          9412 => x"7a51ff8b",
          9413 => x"ea3f82d4",
          9414 => x"d5527851",
          9415 => x"ff8af03f",
          9416 => x"83be1b55",
          9417 => x"77753481",
          9418 => x"0b811634",
          9419 => x"810b8216",
          9420 => x"34778316",
          9421 => x"34758416",
          9422 => x"34606705",
          9423 => x"5680fdc1",
          9424 => x"527551fe",
          9425 => x"a1e83ffe",
          9426 => x"0b851634",
          9427 => x"82d6d808",
          9428 => x"822abf07",
          9429 => x"56758616",
          9430 => x"3482d6d8",
          9431 => x"08871634",
          9432 => x"605283c6",
          9433 => x"1b51ff8a",
          9434 => x"c43f6652",
          9435 => x"83ca1b51",
          9436 => x"ff8aba3f",
          9437 => x"81547753",
          9438 => x"7a527e51",
          9439 => x"ff86bf3f",
          9440 => x"815682d6",
          9441 => x"d808a238",
          9442 => x"80538052",
          9443 => x"7e51ff88",
          9444 => x"913f8156",
          9445 => x"82d6d808",
          9446 => x"90388939",
          9447 => x"8e568a39",
          9448 => x"81568639",
          9449 => x"82d6d808",
          9450 => x"567582d6",
          9451 => x"d80c993d",
          9452 => x"0d04f53d",
          9453 => x"0d7d605b",
          9454 => x"59807960",
          9455 => x"ff055a57",
          9456 => x"57767825",
          9457 => x"b4388d3d",
          9458 => x"f8115555",
          9459 => x"8153fc15",
          9460 => x"527951c9",
          9461 => x"bd3f7a81",
          9462 => x"2e098106",
          9463 => x"9c388c3d",
          9464 => x"3355748d",
          9465 => x"2edb3874",
          9466 => x"76708105",
          9467 => x"58348117",
          9468 => x"57748a2e",
          9469 => x"098106c9",
          9470 => x"38807634",
          9471 => x"78557683",
          9472 => x"38765574",
          9473 => x"82d6d80c",
          9474 => x"8d3d0d04",
          9475 => x"f73d0d7b",
          9476 => x"028405b3",
          9477 => x"05335957",
          9478 => x"778a2e09",
          9479 => x"81068738",
          9480 => x"8d527651",
          9481 => x"e73f8417",
          9482 => x"08568076",
          9483 => x"24be3888",
          9484 => x"17087717",
          9485 => x"8c055659",
          9486 => x"77753481",
          9487 => x"1656bb76",
          9488 => x"25a1388b",
          9489 => x"3dfc0554",
          9490 => x"75538c17",
          9491 => x"52760851",
          9492 => x"cbc03f79",
          9493 => x"76327030",
          9494 => x"7072079f",
          9495 => x"2a703053",
          9496 => x"51565675",
          9497 => x"84180c81",
          9498 => x"1988180c",
          9499 => x"8b3d0d04",
          9500 => x"f93d0d79",
          9501 => x"84110856",
          9502 => x"56807524",
          9503 => x"a738893d",
          9504 => x"fc055474",
          9505 => x"538c1652",
          9506 => x"750851cb",
          9507 => x"853f82d6",
          9508 => x"d8089138",
          9509 => x"84160878",
          9510 => x"2e098106",
          9511 => x"87388816",
          9512 => x"08558339",
          9513 => x"ff557482",
          9514 => x"d6d80c89",
          9515 => x"3d0d04fd",
          9516 => x"3d0d7554",
          9517 => x"80cc5380",
          9518 => x"527351ff",
          9519 => x"88c13f76",
          9520 => x"740c853d",
          9521 => x"0d04ea3d",
          9522 => x"0d0280e3",
          9523 => x"05336a53",
          9524 => x"863d7053",
          9525 => x"5454d83f",
          9526 => x"73527251",
          9527 => x"feae3f72",
          9528 => x"51ff8d3f",
          9529 => x"983d0d04",
          9530 => x"fd3d0d75",
          9531 => x"0284059a",
          9532 => x"05225553",
          9533 => x"80527280",
          9534 => x"ff268a38",
          9535 => x"7283ffff",
          9536 => x"065280c3",
          9537 => x"3983ffff",
          9538 => x"73275173",
          9539 => x"83b52e09",
          9540 => x"8106b438",
          9541 => x"70802eaf",
          9542 => x"3882c998",
          9543 => x"22517271",
          9544 => x"2e9c3881",
          9545 => x"127083ff",
          9546 => x"ff065351",
          9547 => x"7180ff26",
          9548 => x"8d387110",
          9549 => x"82c99805",
          9550 => x"70225151",
          9551 => x"e1398180",
          9552 => x"127081ff",
          9553 => x"06535171",
          9554 => x"82d6d80c",
          9555 => x"853d0d04",
          9556 => x"fe3d0d02",
          9557 => x"92052202",
          9558 => x"84059605",
          9559 => x"22535180",
          9560 => x"537080ff",
          9561 => x"26853870",
          9562 => x"539a3971",
          9563 => x"83b52e09",
          9564 => x"81069138",
          9565 => x"7081ff26",
          9566 => x"8b387010",
          9567 => x"82c79805",
          9568 => x"70225451",
          9569 => x"7282d6d8",
          9570 => x"0c843d0d",
          9571 => x"04fb3d0d",
          9572 => x"77517083",
          9573 => x"ffff2681",
          9574 => x"a7387083",
          9575 => x"ffff0682",
          9576 => x"cb985752",
          9577 => x"9fff7227",
          9578 => x"853882cf",
          9579 => x"8c567570",
          9580 => x"82055722",
          9581 => x"70307080",
          9582 => x"25727526",
          9583 => x"07515255",
          9584 => x"7080fb38",
          9585 => x"75708205",
          9586 => x"57227088",
          9587 => x"2a7181ff",
          9588 => x"06701854",
          9589 => x"52555371",
          9590 => x"712580d7",
          9591 => x"38738826",
          9592 => x"80dc3873",
          9593 => x"842982ae",
          9594 => x"98055170",
          9595 => x"08047175",
          9596 => x"31107611",
          9597 => x"70225451",
          9598 => x"5180c339",
          9599 => x"71753181",
          9600 => x"06727131",
          9601 => x"5151a439",
          9602 => x"f012519f",
          9603 => x"39e01251",
          9604 => x"9a39d012",
          9605 => x"519539e6",
          9606 => x"12519039",
          9607 => x"8812518b",
          9608 => x"39ffb012",
          9609 => x"518539c7",
          9610 => x"a0125170",
          9611 => x"83ffff06",
          9612 => x"528c3973",
          9613 => x"fef83872",
          9614 => x"101656fe",
          9615 => x"f1397151",
          9616 => x"7082d6d8",
          9617 => x"0c873d0d",
          9618 => x"04000000",
          9619 => x"00ffffff",
          9620 => x"ff00ffff",
          9621 => x"ffff00ff",
          9622 => x"ffffff00",
          9623 => x"00002c51",
          9624 => x"00002bd5",
          9625 => x"00002bdc",
          9626 => x"00002be3",
          9627 => x"00002bea",
          9628 => x"00002bf1",
          9629 => x"00002bf8",
          9630 => x"00002bff",
          9631 => x"00002c06",
          9632 => x"00002c0d",
          9633 => x"00002c14",
          9634 => x"00002c1b",
          9635 => x"00002c21",
          9636 => x"00002c27",
          9637 => x"00002c2d",
          9638 => x"00002c33",
          9639 => x"00002c39",
          9640 => x"00002c3f",
          9641 => x"00002c45",
          9642 => x"00002c4b",
          9643 => x"00004234",
          9644 => x"0000423a",
          9645 => x"00004240",
          9646 => x"00004246",
          9647 => x"0000424c",
          9648 => x"0000482a",
          9649 => x"0000492a",
          9650 => x"00004a3b",
          9651 => x"00004c93",
          9652 => x"00004912",
          9653 => x"000046ff",
          9654 => x"00004b03",
          9655 => x"00004c64",
          9656 => x"00004b46",
          9657 => x"00004bdc",
          9658 => x"00004b62",
          9659 => x"000049e5",
          9660 => x"000046ff",
          9661 => x"00004a3b",
          9662 => x"00004a64",
          9663 => x"00004b03",
          9664 => x"000046ff",
          9665 => x"000046ff",
          9666 => x"00004b62",
          9667 => x"00004bdc",
          9668 => x"00004c64",
          9669 => x"00004c93",
          9670 => x"000095ee",
          9671 => x"000095fc",
          9672 => x"00009608",
          9673 => x"0000960d",
          9674 => x"00009612",
          9675 => x"00009617",
          9676 => x"0000961c",
          9677 => x"00009621",
          9678 => x"00009627",
          9679 => x"00000e31",
          9680 => x"0000171a",
          9681 => x"0000171a",
          9682 => x"00000e60",
          9683 => x"0000171a",
          9684 => x"0000171a",
          9685 => x"0000171a",
          9686 => x"0000171a",
          9687 => x"0000171a",
          9688 => x"0000171a",
          9689 => x"0000171a",
          9690 => x"00000e1d",
          9691 => x"0000171a",
          9692 => x"00000e48",
          9693 => x"00000e78",
          9694 => x"0000171a",
          9695 => x"0000171a",
          9696 => x"0000171a",
          9697 => x"0000171a",
          9698 => x"0000171a",
          9699 => x"0000171a",
          9700 => x"0000171a",
          9701 => x"0000171a",
          9702 => x"0000171a",
          9703 => x"0000171a",
          9704 => x"0000171a",
          9705 => x"0000171a",
          9706 => x"0000171a",
          9707 => x"0000171a",
          9708 => x"0000171a",
          9709 => x"0000171a",
          9710 => x"0000171a",
          9711 => x"0000171a",
          9712 => x"0000171a",
          9713 => x"0000171a",
          9714 => x"0000171a",
          9715 => x"0000171a",
          9716 => x"0000171a",
          9717 => x"0000171a",
          9718 => x"0000171a",
          9719 => x"0000171a",
          9720 => x"0000171a",
          9721 => x"0000171a",
          9722 => x"0000171a",
          9723 => x"0000171a",
          9724 => x"0000171a",
          9725 => x"0000171a",
          9726 => x"0000171a",
          9727 => x"0000171a",
          9728 => x"0000171a",
          9729 => x"0000171a",
          9730 => x"00000fa8",
          9731 => x"0000171a",
          9732 => x"0000171a",
          9733 => x"0000171a",
          9734 => x"0000171a",
          9735 => x"00001116",
          9736 => x"0000171a",
          9737 => x"0000171a",
          9738 => x"0000171a",
          9739 => x"0000171a",
          9740 => x"0000171a",
          9741 => x"0000171a",
          9742 => x"0000171a",
          9743 => x"0000171a",
          9744 => x"0000171a",
          9745 => x"0000171a",
          9746 => x"00000ed8",
          9747 => x"0000103f",
          9748 => x"00000eaf",
          9749 => x"00000eaf",
          9750 => x"00000eaf",
          9751 => x"0000171a",
          9752 => x"0000103f",
          9753 => x"0000171a",
          9754 => x"0000171a",
          9755 => x"00000e98",
          9756 => x"0000171a",
          9757 => x"0000171a",
          9758 => x"000010ec",
          9759 => x"000010f7",
          9760 => x"0000171a",
          9761 => x"0000171a",
          9762 => x"00000f11",
          9763 => x"0000171a",
          9764 => x"0000111f",
          9765 => x"0000171a",
          9766 => x"0000171a",
          9767 => x"00001116",
          9768 => x"64696e69",
          9769 => x"74000000",
          9770 => x"64696f63",
          9771 => x"746c0000",
          9772 => x"66696e69",
          9773 => x"74000000",
          9774 => x"666c6f61",
          9775 => x"64000000",
          9776 => x"66657865",
          9777 => x"63000000",
          9778 => x"6d636c65",
          9779 => x"61720000",
          9780 => x"6d636f70",
          9781 => x"79000000",
          9782 => x"6d646966",
          9783 => x"66000000",
          9784 => x"6d64756d",
          9785 => x"70000000",
          9786 => x"6d656200",
          9787 => x"6d656800",
          9788 => x"6d657700",
          9789 => x"68696400",
          9790 => x"68696500",
          9791 => x"68666400",
          9792 => x"68666500",
          9793 => x"63616c6c",
          9794 => x"00000000",
          9795 => x"6a6d7000",
          9796 => x"72657374",
          9797 => x"61727400",
          9798 => x"72657365",
          9799 => x"74000000",
          9800 => x"696e666f",
          9801 => x"00000000",
          9802 => x"74657374",
          9803 => x"00000000",
          9804 => x"74626173",
          9805 => x"69630000",
          9806 => x"6d626173",
          9807 => x"69630000",
          9808 => x"6b696c6f",
          9809 => x"00000000",
          9810 => x"65640000",
          9811 => x"4469736b",
          9812 => x"20457272",
          9813 => x"6f720000",
          9814 => x"496e7465",
          9815 => x"726e616c",
          9816 => x"20657272",
          9817 => x"6f722e00",
          9818 => x"4469736b",
          9819 => x"206e6f74",
          9820 => x"20726561",
          9821 => x"64792e00",
          9822 => x"4e6f2066",
          9823 => x"696c6520",
          9824 => x"666f756e",
          9825 => x"642e0000",
          9826 => x"4e6f2070",
          9827 => x"61746820",
          9828 => x"666f756e",
          9829 => x"642e0000",
          9830 => x"496e7661",
          9831 => x"6c696420",
          9832 => x"66696c65",
          9833 => x"6e616d65",
          9834 => x"2e000000",
          9835 => x"41636365",
          9836 => x"73732064",
          9837 => x"656e6965",
          9838 => x"642e0000",
          9839 => x"46696c65",
          9840 => x"20616c72",
          9841 => x"65616479",
          9842 => x"20657869",
          9843 => x"7374732e",
          9844 => x"00000000",
          9845 => x"46696c65",
          9846 => x"2068616e",
          9847 => x"646c6520",
          9848 => x"696e7661",
          9849 => x"6c69642e",
          9850 => x"00000000",
          9851 => x"53442069",
          9852 => x"73207772",
          9853 => x"69746520",
          9854 => x"70726f74",
          9855 => x"65637465",
          9856 => x"642e0000",
          9857 => x"44726976",
          9858 => x"65206e75",
          9859 => x"6d626572",
          9860 => x"20697320",
          9861 => x"696e7661",
          9862 => x"6c69642e",
          9863 => x"00000000",
          9864 => x"4469736b",
          9865 => x"206e6f74",
          9866 => x"20656e61",
          9867 => x"626c6564",
          9868 => x"2e000000",
          9869 => x"4e6f2063",
          9870 => x"6f6d7061",
          9871 => x"7469626c",
          9872 => x"65206669",
          9873 => x"6c657379",
          9874 => x"7374656d",
          9875 => x"20666f75",
          9876 => x"6e64206f",
          9877 => x"6e206469",
          9878 => x"736b2e00",
          9879 => x"466f726d",
          9880 => x"61742061",
          9881 => x"626f7274",
          9882 => x"65642e00",
          9883 => x"54696d65",
          9884 => x"6f75742c",
          9885 => x"206f7065",
          9886 => x"72617469",
          9887 => x"6f6e2063",
          9888 => x"616e6365",
          9889 => x"6c6c6564",
          9890 => x"2e000000",
          9891 => x"46696c65",
          9892 => x"20697320",
          9893 => x"6c6f636b",
          9894 => x"65642e00",
          9895 => x"496e7375",
          9896 => x"66666963",
          9897 => x"69656e74",
          9898 => x"206d656d",
          9899 => x"6f72792e",
          9900 => x"00000000",
          9901 => x"546f6f20",
          9902 => x"6d616e79",
          9903 => x"206f7065",
          9904 => x"6e206669",
          9905 => x"6c65732e",
          9906 => x"00000000",
          9907 => x"50617261",
          9908 => x"6d657465",
          9909 => x"72732069",
          9910 => x"6e636f72",
          9911 => x"72656374",
          9912 => x"2e000000",
          9913 => x"53756363",
          9914 => x"6573732e",
          9915 => x"00000000",
          9916 => x"556e6b6e",
          9917 => x"6f776e20",
          9918 => x"6572726f",
          9919 => x"722e0000",
          9920 => x"0a256c75",
          9921 => x"20627974",
          9922 => x"65732025",
          9923 => x"73206174",
          9924 => x"20256c75",
          9925 => x"20627974",
          9926 => x"65732f73",
          9927 => x"65632e0a",
          9928 => x"00000000",
          9929 => x"72656164",
          9930 => x"00000000",
          9931 => x"303d2530",
          9932 => x"386c782c",
          9933 => x"20313d25",
          9934 => x"30386c78",
          9935 => x"2c20323d",
          9936 => x"2530386c",
          9937 => x"782c205f",
          9938 => x"494f423d",
          9939 => x"2530386c",
          9940 => x"78202530",
          9941 => x"386c7820",
          9942 => x"2530386c",
          9943 => x"780a0000",
          9944 => x"2530386c",
          9945 => x"58000000",
          9946 => x"3a202000",
          9947 => x"25303458",
          9948 => x"00000000",
          9949 => x"20202020",
          9950 => x"20202020",
          9951 => x"00000000",
          9952 => x"25303258",
          9953 => x"00000000",
          9954 => x"20200000",
          9955 => x"207c0000",
          9956 => x"7c000000",
          9957 => x"7a4f5300",
          9958 => x"0a2a2a20",
          9959 => x"25732028",
          9960 => x"00000000",
          9961 => x"30352f31",
          9962 => x"322f3230",
          9963 => x"32300000",
          9964 => x"76312e30",
          9965 => x"34660000",
          9966 => x"205a5055",
          9967 => x"2c207265",
          9968 => x"76202530",
          9969 => x"32782920",
          9970 => x"25732025",
          9971 => x"73202a2a",
          9972 => x"0a0a0000",
          9973 => x"5a505520",
          9974 => x"496e7465",
          9975 => x"72727570",
          9976 => x"74204861",
          9977 => x"6e646c65",
          9978 => x"72000000",
          9979 => x"54696d65",
          9980 => x"7220696e",
          9981 => x"74657272",
          9982 => x"75707400",
          9983 => x"50533220",
          9984 => x"696e7465",
          9985 => x"72727570",
          9986 => x"74000000",
          9987 => x"494f4354",
          9988 => x"4c205244",
          9989 => x"20696e74",
          9990 => x"65727275",
          9991 => x"70740000",
          9992 => x"494f4354",
          9993 => x"4c205752",
          9994 => x"20696e74",
          9995 => x"65727275",
          9996 => x"70740000",
          9997 => x"55415254",
          9998 => x"30205258",
          9999 => x"20696e74",
         10000 => x"65727275",
         10001 => x"70740000",
         10002 => x"55415254",
         10003 => x"30205458",
         10004 => x"20696e74",
         10005 => x"65727275",
         10006 => x"70740000",
         10007 => x"55415254",
         10008 => x"31205258",
         10009 => x"20696e74",
         10010 => x"65727275",
         10011 => x"70740000",
         10012 => x"55415254",
         10013 => x"31205458",
         10014 => x"20696e74",
         10015 => x"65727275",
         10016 => x"70740000",
         10017 => x"53657474",
         10018 => x"696e6720",
         10019 => x"75702074",
         10020 => x"696d6572",
         10021 => x"2e2e2e00",
         10022 => x"456e6162",
         10023 => x"6c696e67",
         10024 => x"2074696d",
         10025 => x"65722e2e",
         10026 => x"2e000000",
         10027 => x"6175746f",
         10028 => x"65786563",
         10029 => x"2e626174",
         10030 => x"00000000",
         10031 => x"7a4f532e",
         10032 => x"68737400",
         10033 => x"303a0000",
         10034 => x"4661696c",
         10035 => x"65642074",
         10036 => x"6f20696e",
         10037 => x"69746961",
         10038 => x"6c697365",
         10039 => x"20736420",
         10040 => x"63617264",
         10041 => x"20302c20",
         10042 => x"706c6561",
         10043 => x"73652069",
         10044 => x"6e697420",
         10045 => x"6d616e75",
         10046 => x"616c6c79",
         10047 => x"2e000000",
         10048 => x"2a200000",
         10049 => x"436c6561",
         10050 => x"72696e67",
         10051 => x"2e2e2e2e",
         10052 => x"00000000",
         10053 => x"436f7079",
         10054 => x"696e672e",
         10055 => x"2e2e0000",
         10056 => x"436f6d70",
         10057 => x"6172696e",
         10058 => x"672e2e2e",
         10059 => x"00000000",
         10060 => x"2530386c",
         10061 => x"78282530",
         10062 => x"3878292d",
         10063 => x"3e253038",
         10064 => x"6c782825",
         10065 => x"30387829",
         10066 => x"0a000000",
         10067 => x"44756d70",
         10068 => x"204d656d",
         10069 => x"6f727900",
         10070 => x"0a436f6d",
         10071 => x"706c6574",
         10072 => x"652e0000",
         10073 => x"2530386c",
         10074 => x"58202530",
         10075 => x"32582d00",
         10076 => x"3f3f3f00",
         10077 => x"2530386c",
         10078 => x"58202530",
         10079 => x"34582d00",
         10080 => x"2530386c",
         10081 => x"58202530",
         10082 => x"386c582d",
         10083 => x"00000000",
         10084 => x"45786563",
         10085 => x"7574696e",
         10086 => x"6720636f",
         10087 => x"64652040",
         10088 => x"20253038",
         10089 => x"6c78202e",
         10090 => x"2e2e0a00",
         10091 => x"43616c6c",
         10092 => x"696e6720",
         10093 => x"636f6465",
         10094 => x"20402025",
         10095 => x"30386c78",
         10096 => x"202e2e2e",
         10097 => x"0a000000",
         10098 => x"43616c6c",
         10099 => x"20726574",
         10100 => x"75726e65",
         10101 => x"6420636f",
         10102 => x"64652028",
         10103 => x"2564292e",
         10104 => x"0a000000",
         10105 => x"52657374",
         10106 => x"61727469",
         10107 => x"6e672061",
         10108 => x"70706c69",
         10109 => x"63617469",
         10110 => x"6f6e2e2e",
         10111 => x"2e000000",
         10112 => x"436f6c64",
         10113 => x"20726562",
         10114 => x"6f6f7469",
         10115 => x"6e672e2e",
         10116 => x"2e000000",
         10117 => x"5a505500",
         10118 => x"62696e00",
         10119 => x"25643a5c",
         10120 => x"25735c25",
         10121 => x"732e2573",
         10122 => x"00000000",
         10123 => x"25643a5c",
         10124 => x"25735c25",
         10125 => x"73000000",
         10126 => x"25643a5c",
         10127 => x"25730000",
         10128 => x"42616420",
         10129 => x"636f6d6d",
         10130 => x"616e642e",
         10131 => x"00000000",
         10132 => x"4d656d6f",
         10133 => x"72792065",
         10134 => x"78686175",
         10135 => x"73746564",
         10136 => x"2c206361",
         10137 => x"6e6e6f74",
         10138 => x"2070726f",
         10139 => x"63657373",
         10140 => x"20636f6d",
         10141 => x"6d616e64",
         10142 => x"2e000000",
         10143 => x"54657374",
         10144 => x"696e6720",
         10145 => x"7072696e",
         10146 => x"74660000",
         10147 => x"52756e6e",
         10148 => x"696e672e",
         10149 => x"2e2e0000",
         10150 => x"456e6162",
         10151 => x"6c696e67",
         10152 => x"20696e74",
         10153 => x"65727275",
         10154 => x"7074732e",
         10155 => x"2e2e0000",
         10156 => x"25642f25",
         10157 => x"642f2564",
         10158 => x"2025643a",
         10159 => x"25643a25",
         10160 => x"642e2564",
         10161 => x"25640a00",
         10162 => x"536f4320",
         10163 => x"436f6e66",
         10164 => x"69677572",
         10165 => x"6174696f",
         10166 => x"6e000000",
         10167 => x"20286672",
         10168 => x"6f6d2053",
         10169 => x"6f432063",
         10170 => x"6f6e6669",
         10171 => x"67290000",
         10172 => x"3a0a4465",
         10173 => x"76696365",
         10174 => x"7320696d",
         10175 => x"706c656d",
         10176 => x"656e7465",
         10177 => x"643a0000",
         10178 => x"20202020",
         10179 => x"57422053",
         10180 => x"4452414d",
         10181 => x"20202825",
         10182 => x"3038583a",
         10183 => x"25303858",
         10184 => x"292e0a00",
         10185 => x"20202020",
         10186 => x"53445241",
         10187 => x"4d202020",
         10188 => x"20202825",
         10189 => x"3038583a",
         10190 => x"25303858",
         10191 => x"292e0a00",
         10192 => x"20202020",
         10193 => x"494e534e",
         10194 => x"20425241",
         10195 => x"4d202825",
         10196 => x"3038583a",
         10197 => x"25303858",
         10198 => x"292e0a00",
         10199 => x"20202020",
         10200 => x"4252414d",
         10201 => x"20202020",
         10202 => x"20202825",
         10203 => x"3038583a",
         10204 => x"25303858",
         10205 => x"292e0a00",
         10206 => x"20202020",
         10207 => x"52414d20",
         10208 => x"20202020",
         10209 => x"20202825",
         10210 => x"3038583a",
         10211 => x"25303858",
         10212 => x"292e0a00",
         10213 => x"20202020",
         10214 => x"53442043",
         10215 => x"41524420",
         10216 => x"20202844",
         10217 => x"65766963",
         10218 => x"6573203d",
         10219 => x"25303264",
         10220 => x"292e0a00",
         10221 => x"20202020",
         10222 => x"54494d45",
         10223 => x"52312020",
         10224 => x"20202854",
         10225 => x"696d6572",
         10226 => x"7320203d",
         10227 => x"25303264",
         10228 => x"292e0a00",
         10229 => x"20202020",
         10230 => x"494e5452",
         10231 => x"20435452",
         10232 => x"4c202843",
         10233 => x"68616e6e",
         10234 => x"656c733d",
         10235 => x"25303264",
         10236 => x"292e0a00",
         10237 => x"20202020",
         10238 => x"57495348",
         10239 => x"424f4e45",
         10240 => x"20425553",
         10241 => x"00000000",
         10242 => x"20202020",
         10243 => x"57422049",
         10244 => x"32430000",
         10245 => x"20202020",
         10246 => x"494f4354",
         10247 => x"4c000000",
         10248 => x"20202020",
         10249 => x"50533200",
         10250 => x"20202020",
         10251 => x"53504900",
         10252 => x"41646472",
         10253 => x"65737365",
         10254 => x"733a0000",
         10255 => x"20202020",
         10256 => x"43505520",
         10257 => x"52657365",
         10258 => x"74205665",
         10259 => x"63746f72",
         10260 => x"20416464",
         10261 => x"72657373",
         10262 => x"203d2025",
         10263 => x"3038580a",
         10264 => x"00000000",
         10265 => x"20202020",
         10266 => x"43505520",
         10267 => x"4d656d6f",
         10268 => x"72792053",
         10269 => x"74617274",
         10270 => x"20416464",
         10271 => x"72657373",
         10272 => x"203d2025",
         10273 => x"3038580a",
         10274 => x"00000000",
         10275 => x"20202020",
         10276 => x"53746163",
         10277 => x"6b205374",
         10278 => x"61727420",
         10279 => x"41646472",
         10280 => x"65737320",
         10281 => x"20202020",
         10282 => x"203d2025",
         10283 => x"3038580a",
         10284 => x"00000000",
         10285 => x"4d697363",
         10286 => x"3a000000",
         10287 => x"20202020",
         10288 => x"5a505520",
         10289 => x"49642020",
         10290 => x"20202020",
         10291 => x"20202020",
         10292 => x"20202020",
         10293 => x"20202020",
         10294 => x"203d2025",
         10295 => x"3034580a",
         10296 => x"00000000",
         10297 => x"20202020",
         10298 => x"53797374",
         10299 => x"656d2043",
         10300 => x"6c6f636b",
         10301 => x"20467265",
         10302 => x"71202020",
         10303 => x"20202020",
         10304 => x"203d2025",
         10305 => x"642e2530",
         10306 => x"34644d48",
         10307 => x"7a0a0000",
         10308 => x"20202020",
         10309 => x"53445241",
         10310 => x"4d20436c",
         10311 => x"6f636b20",
         10312 => x"46726571",
         10313 => x"20202020",
         10314 => x"20202020",
         10315 => x"203d2025",
         10316 => x"642e2530",
         10317 => x"34644d48",
         10318 => x"7a0a0000",
         10319 => x"20202020",
         10320 => x"57697368",
         10321 => x"626f6e65",
         10322 => x"20534452",
         10323 => x"414d2043",
         10324 => x"6c6f636b",
         10325 => x"20467265",
         10326 => x"713d2025",
         10327 => x"642e2530",
         10328 => x"34644d48",
         10329 => x"7a0a0000",
         10330 => x"536d616c",
         10331 => x"6c000000",
         10332 => x"4d656469",
         10333 => x"756d0000",
         10334 => x"466c6578",
         10335 => x"00000000",
         10336 => x"45564f00",
         10337 => x"45564f6d",
         10338 => x"00000000",
         10339 => x"556e6b6e",
         10340 => x"6f776e00",
         10341 => x"0000a2f0",
         10342 => x"01000000",
         10343 => x"00000002",
         10344 => x"0000a2ec",
         10345 => x"01000000",
         10346 => x"00000003",
         10347 => x"0000a2e8",
         10348 => x"01000000",
         10349 => x"00000004",
         10350 => x"0000a2e4",
         10351 => x"01000000",
         10352 => x"00000005",
         10353 => x"0000a2e0",
         10354 => x"01000000",
         10355 => x"00000006",
         10356 => x"0000a2dc",
         10357 => x"01000000",
         10358 => x"00000007",
         10359 => x"0000a2d8",
         10360 => x"01000000",
         10361 => x"00000001",
         10362 => x"0000a2d4",
         10363 => x"01000000",
         10364 => x"00000008",
         10365 => x"0000a2d0",
         10366 => x"01000000",
         10367 => x"0000000b",
         10368 => x"0000a2cc",
         10369 => x"01000000",
         10370 => x"00000009",
         10371 => x"0000a2c8",
         10372 => x"01000000",
         10373 => x"0000000a",
         10374 => x"0000a2c4",
         10375 => x"04000000",
         10376 => x"0000000d",
         10377 => x"0000a2c0",
         10378 => x"04000000",
         10379 => x"0000000c",
         10380 => x"0000a2bc",
         10381 => x"04000000",
         10382 => x"0000000e",
         10383 => x"0000a2b8",
         10384 => x"03000000",
         10385 => x"0000000f",
         10386 => x"0000a2b4",
         10387 => x"04000000",
         10388 => x"0000000f",
         10389 => x"0000a2b0",
         10390 => x"04000000",
         10391 => x"00000010",
         10392 => x"0000a2ac",
         10393 => x"04000000",
         10394 => x"00000011",
         10395 => x"0000a2a8",
         10396 => x"03000000",
         10397 => x"00000012",
         10398 => x"0000a2a4",
         10399 => x"03000000",
         10400 => x"00000013",
         10401 => x"0000a2a0",
         10402 => x"03000000",
         10403 => x"00000014",
         10404 => x"0000a29c",
         10405 => x"03000000",
         10406 => x"00000015",
         10407 => x"1b5b4400",
         10408 => x"1b5b4300",
         10409 => x"1b5b4200",
         10410 => x"1b5b4100",
         10411 => x"1b5b367e",
         10412 => x"1b5b357e",
         10413 => x"1b5b347e",
         10414 => x"1b304600",
         10415 => x"1b5b337e",
         10416 => x"1b5b327e",
         10417 => x"1b5b317e",
         10418 => x"10000000",
         10419 => x"0e000000",
         10420 => x"0d000000",
         10421 => x"0b000000",
         10422 => x"08000000",
         10423 => x"06000000",
         10424 => x"05000000",
         10425 => x"04000000",
         10426 => x"03000000",
         10427 => x"02000000",
         10428 => x"01000000",
         10429 => x"68697374",
         10430 => x"6f727900",
         10431 => x"68697374",
         10432 => x"00000000",
         10433 => x"21000000",
         10434 => x"2530346c",
         10435 => x"75202025",
         10436 => x"730a0000",
         10437 => x"4661696c",
         10438 => x"65642074",
         10439 => x"6f207265",
         10440 => x"73657420",
         10441 => x"74686520",
         10442 => x"68697374",
         10443 => x"6f727920",
         10444 => x"66696c65",
         10445 => x"20746f20",
         10446 => x"454f462e",
         10447 => x"00000000",
         10448 => x"43616e6e",
         10449 => x"6f74206f",
         10450 => x"70656e2f",
         10451 => x"63726561",
         10452 => x"74652068",
         10453 => x"6973746f",
         10454 => x"72792066",
         10455 => x"696c652c",
         10456 => x"20646973",
         10457 => x"61626c69",
         10458 => x"6e672e00",
         10459 => x"53440000",
         10460 => x"222a3a3c",
         10461 => x"3e3f7c7f",
         10462 => x"00000000",
         10463 => x"2b2c3b3d",
         10464 => x"5b5d0000",
         10465 => x"46415400",
         10466 => x"46415433",
         10467 => x"32000000",
         10468 => x"ebfe904d",
         10469 => x"53444f53",
         10470 => x"352e3000",
         10471 => x"4e4f204e",
         10472 => x"414d4520",
         10473 => x"20202046",
         10474 => x"41543332",
         10475 => x"20202000",
         10476 => x"4e4f204e",
         10477 => x"414d4520",
         10478 => x"20202046",
         10479 => x"41542020",
         10480 => x"20202000",
         10481 => x"0000a36c",
         10482 => x"00000000",
         10483 => x"00000000",
         10484 => x"00000000",
         10485 => x"01030507",
         10486 => x"090e1012",
         10487 => x"1416181c",
         10488 => x"1e000000",
         10489 => x"809a4541",
         10490 => x"8e418f80",
         10491 => x"45454549",
         10492 => x"49498e8f",
         10493 => x"9092924f",
         10494 => x"994f5555",
         10495 => x"59999a9b",
         10496 => x"9c9d9e9f",
         10497 => x"41494f55",
         10498 => x"a5a5a6a7",
         10499 => x"a8a9aaab",
         10500 => x"acadaeaf",
         10501 => x"b0b1b2b3",
         10502 => x"b4b5b6b7",
         10503 => x"b8b9babb",
         10504 => x"bcbdbebf",
         10505 => x"c0c1c2c3",
         10506 => x"c4c5c6c7",
         10507 => x"c8c9cacb",
         10508 => x"cccdcecf",
         10509 => x"d0d1d2d3",
         10510 => x"d4d5d6d7",
         10511 => x"d8d9dadb",
         10512 => x"dcdddedf",
         10513 => x"e0e1e2e3",
         10514 => x"e4e5e6e7",
         10515 => x"e8e9eaeb",
         10516 => x"ecedeeef",
         10517 => x"f0f1f2f3",
         10518 => x"f4f5f6f7",
         10519 => x"f8f9fafb",
         10520 => x"fcfdfeff",
         10521 => x"2b2e2c3b",
         10522 => x"3d5b5d2f",
         10523 => x"5c222a3a",
         10524 => x"3c3e3f7c",
         10525 => x"7f000000",
         10526 => x"00010004",
         10527 => x"00100040",
         10528 => x"01000200",
         10529 => x"00000000",
         10530 => x"00010002",
         10531 => x"00040008",
         10532 => x"00100020",
         10533 => x"00000000",
         10534 => x"00c700fc",
         10535 => x"00e900e2",
         10536 => x"00e400e0",
         10537 => x"00e500e7",
         10538 => x"00ea00eb",
         10539 => x"00e800ef",
         10540 => x"00ee00ec",
         10541 => x"00c400c5",
         10542 => x"00c900e6",
         10543 => x"00c600f4",
         10544 => x"00f600f2",
         10545 => x"00fb00f9",
         10546 => x"00ff00d6",
         10547 => x"00dc00a2",
         10548 => x"00a300a5",
         10549 => x"20a70192",
         10550 => x"00e100ed",
         10551 => x"00f300fa",
         10552 => x"00f100d1",
         10553 => x"00aa00ba",
         10554 => x"00bf2310",
         10555 => x"00ac00bd",
         10556 => x"00bc00a1",
         10557 => x"00ab00bb",
         10558 => x"25912592",
         10559 => x"25932502",
         10560 => x"25242561",
         10561 => x"25622556",
         10562 => x"25552563",
         10563 => x"25512557",
         10564 => x"255d255c",
         10565 => x"255b2510",
         10566 => x"25142534",
         10567 => x"252c251c",
         10568 => x"2500253c",
         10569 => x"255e255f",
         10570 => x"255a2554",
         10571 => x"25692566",
         10572 => x"25602550",
         10573 => x"256c2567",
         10574 => x"25682564",
         10575 => x"25652559",
         10576 => x"25582552",
         10577 => x"2553256b",
         10578 => x"256a2518",
         10579 => x"250c2588",
         10580 => x"2584258c",
         10581 => x"25902580",
         10582 => x"03b100df",
         10583 => x"039303c0",
         10584 => x"03a303c3",
         10585 => x"00b503c4",
         10586 => x"03a60398",
         10587 => x"03a903b4",
         10588 => x"221e03c6",
         10589 => x"03b52229",
         10590 => x"226100b1",
         10591 => x"22652264",
         10592 => x"23202321",
         10593 => x"00f72248",
         10594 => x"00b02219",
         10595 => x"00b7221a",
         10596 => x"207f00b2",
         10597 => x"25a000a0",
         10598 => x"0061031a",
         10599 => x"00e00317",
         10600 => x"00f80307",
         10601 => x"00ff0001",
         10602 => x"01780100",
         10603 => x"01300132",
         10604 => x"01060139",
         10605 => x"0110014a",
         10606 => x"012e0179",
         10607 => x"01060180",
         10608 => x"004d0243",
         10609 => x"01810182",
         10610 => x"01820184",
         10611 => x"01840186",
         10612 => x"01870187",
         10613 => x"0189018a",
         10614 => x"018b018b",
         10615 => x"018d018e",
         10616 => x"018f0190",
         10617 => x"01910191",
         10618 => x"01930194",
         10619 => x"01f60196",
         10620 => x"01970198",
         10621 => x"0198023d",
         10622 => x"019b019c",
         10623 => x"019d0220",
         10624 => x"019f01a0",
         10625 => x"01a001a2",
         10626 => x"01a201a4",
         10627 => x"01a401a6",
         10628 => x"01a701a7",
         10629 => x"01a901aa",
         10630 => x"01ab01ac",
         10631 => x"01ac01ae",
         10632 => x"01af01af",
         10633 => x"01b101b2",
         10634 => x"01b301b3",
         10635 => x"01b501b5",
         10636 => x"01b701b8",
         10637 => x"01b801ba",
         10638 => x"01bb01bc",
         10639 => x"01bc01be",
         10640 => x"01f701c0",
         10641 => x"01c101c2",
         10642 => x"01c301c4",
         10643 => x"01c501c4",
         10644 => x"01c701c8",
         10645 => x"01c701ca",
         10646 => x"01cb01ca",
         10647 => x"01cd0110",
         10648 => x"01dd0001",
         10649 => x"018e01de",
         10650 => x"011201f3",
         10651 => x"000301f1",
         10652 => x"01f401f4",
         10653 => x"01f80128",
         10654 => x"02220112",
         10655 => x"023a0009",
         10656 => x"2c65023b",
         10657 => x"023b023d",
         10658 => x"2c66023f",
         10659 => x"02400241",
         10660 => x"02410246",
         10661 => x"010a0253",
         10662 => x"00400181",
         10663 => x"01860255",
         10664 => x"0189018a",
         10665 => x"0258018f",
         10666 => x"025a0190",
         10667 => x"025c025d",
         10668 => x"025e025f",
         10669 => x"01930261",
         10670 => x"02620194",
         10671 => x"02640265",
         10672 => x"02660267",
         10673 => x"01970196",
         10674 => x"026a2c62",
         10675 => x"026c026d",
         10676 => x"026e019c",
         10677 => x"02700271",
         10678 => x"019d0273",
         10679 => x"0274019f",
         10680 => x"02760277",
         10681 => x"02780279",
         10682 => x"027a027b",
         10683 => x"027c2c64",
         10684 => x"027e027f",
         10685 => x"01a60281",
         10686 => x"028201a9",
         10687 => x"02840285",
         10688 => x"02860287",
         10689 => x"01ae0244",
         10690 => x"01b101b2",
         10691 => x"0245028d",
         10692 => x"028e028f",
         10693 => x"02900291",
         10694 => x"01b7037b",
         10695 => x"000303fd",
         10696 => x"03fe03ff",
         10697 => x"03ac0004",
         10698 => x"03860388",
         10699 => x"0389038a",
         10700 => x"03b10311",
         10701 => x"03c20002",
         10702 => x"03a303a3",
         10703 => x"03c40308",
         10704 => x"03cc0003",
         10705 => x"038c038e",
         10706 => x"038f03d8",
         10707 => x"011803f2",
         10708 => x"000a03f9",
         10709 => x"03f303f4",
         10710 => x"03f503f6",
         10711 => x"03f703f7",
         10712 => x"03f903fa",
         10713 => x"03fa0430",
         10714 => x"03200450",
         10715 => x"07100460",
         10716 => x"0122048a",
         10717 => x"013604c1",
         10718 => x"010e04cf",
         10719 => x"000104c0",
         10720 => x"04d00144",
         10721 => x"05610426",
         10722 => x"00000000",
         10723 => x"1d7d0001",
         10724 => x"2c631e00",
         10725 => x"01961ea0",
         10726 => x"015a1f00",
         10727 => x"06081f10",
         10728 => x"06061f20",
         10729 => x"06081f30",
         10730 => x"06081f40",
         10731 => x"06061f51",
         10732 => x"00071f59",
         10733 => x"1f521f5b",
         10734 => x"1f541f5d",
         10735 => x"1f561f5f",
         10736 => x"1f600608",
         10737 => x"1f70000e",
         10738 => x"1fba1fbb",
         10739 => x"1fc81fc9",
         10740 => x"1fca1fcb",
         10741 => x"1fda1fdb",
         10742 => x"1ff81ff9",
         10743 => x"1fea1feb",
         10744 => x"1ffa1ffb",
         10745 => x"1f800608",
         10746 => x"1f900608",
         10747 => x"1fa00608",
         10748 => x"1fb00004",
         10749 => x"1fb81fb9",
         10750 => x"1fb21fbc",
         10751 => x"1fcc0001",
         10752 => x"1fc31fd0",
         10753 => x"06021fe0",
         10754 => x"06021fe5",
         10755 => x"00011fec",
         10756 => x"1ff30001",
         10757 => x"1ffc214e",
         10758 => x"00012132",
         10759 => x"21700210",
         10760 => x"21840001",
         10761 => x"218324d0",
         10762 => x"051a2c30",
         10763 => x"042f2c60",
         10764 => x"01022c67",
         10765 => x"01062c75",
         10766 => x"01022c80",
         10767 => x"01642d00",
         10768 => x"0826ff41",
         10769 => x"031a0000",
         10770 => x"00000000",
         10771 => x"000098a0",
         10772 => x"01020100",
         10773 => x"00000000",
         10774 => x"00000000",
         10775 => x"000098a8",
         10776 => x"01040100",
         10777 => x"00000000",
         10778 => x"00000000",
         10779 => x"000098b0",
         10780 => x"01140300",
         10781 => x"00000000",
         10782 => x"00000000",
         10783 => x"000098b8",
         10784 => x"012b0300",
         10785 => x"00000000",
         10786 => x"00000000",
         10787 => x"000098c0",
         10788 => x"01300300",
         10789 => x"00000000",
         10790 => x"00000000",
         10791 => x"000098c8",
         10792 => x"013c0400",
         10793 => x"00000000",
         10794 => x"00000000",
         10795 => x"000098d0",
         10796 => x"013d0400",
         10797 => x"00000000",
         10798 => x"00000000",
         10799 => x"000098d8",
         10800 => x"013f0400",
         10801 => x"00000000",
         10802 => x"00000000",
         10803 => x"000098e0",
         10804 => x"01400400",
         10805 => x"00000000",
         10806 => x"00000000",
         10807 => x"000098e8",
         10808 => x"01410400",
         10809 => x"00000000",
         10810 => x"00000000",
         10811 => x"000098ec",
         10812 => x"01420400",
         10813 => x"00000000",
         10814 => x"00000000",
         10815 => x"000098f0",
         10816 => x"01430400",
         10817 => x"00000000",
         10818 => x"00000000",
         10819 => x"000098f4",
         10820 => x"01500500",
         10821 => x"00000000",
         10822 => x"00000000",
         10823 => x"000098f8",
         10824 => x"01510500",
         10825 => x"00000000",
         10826 => x"00000000",
         10827 => x"000098fc",
         10828 => x"01540500",
         10829 => x"00000000",
         10830 => x"00000000",
         10831 => x"00009900",
         10832 => x"01550500",
         10833 => x"00000000",
         10834 => x"00000000",
         10835 => x"00009904",
         10836 => x"01790700",
         10837 => x"00000000",
         10838 => x"00000000",
         10839 => x"0000990c",
         10840 => x"01780700",
         10841 => x"00000000",
         10842 => x"00000000",
         10843 => x"00009910",
         10844 => x"01820800",
         10845 => x"00000000",
         10846 => x"00000000",
         10847 => x"00009918",
         10848 => x"01830800",
         10849 => x"00000000",
         10850 => x"00000000",
         10851 => x"00009920",
         10852 => x"01850800",
         10853 => x"00000000",
         10854 => x"00000000",
         10855 => x"00009928",
         10856 => x"01870800",
         10857 => x"00000000",
         10858 => x"00000000",
         10859 => x"00009930",
         10860 => x"018c0900",
         10861 => x"00000000",
         10862 => x"00000000",
         10863 => x"00009938",
         10864 => x"018d0900",
         10865 => x"00000000",
         10866 => x"00000000",
         10867 => x"00009940",
         10868 => x"018e0900",
         10869 => x"00000000",
         10870 => x"00000000",
         10871 => x"00009948",
         10872 => x"018f0900",
         10873 => x"00000000",
         10874 => x"00000000",
         10875 => x"00000000",
         10876 => x"00000000",
         10877 => x"00007fff",
         10878 => x"00000000",
         10879 => x"00007fff",
         10880 => x"00010000",
         10881 => x"00007fff",
         10882 => x"00010000",
         10883 => x"00810000",
         10884 => x"01000000",
         10885 => x"017fffff",
         10886 => x"00000000",
         10887 => x"00000000",
         10888 => x"00007800",
         10889 => x"00000000",
         10890 => x"05f5e100",
         10891 => x"05f5e100",
         10892 => x"05f5e100",
         10893 => x"00000000",
         10894 => x"01010101",
         10895 => x"01010101",
         10896 => x"01011001",
         10897 => x"01000000",
         10898 => x"00000000",
         10899 => x"00000000",
         10900 => x"00000000",
         10901 => x"00000000",
         10902 => x"00000000",
         10903 => x"00000000",
         10904 => x"00000000",
         10905 => x"00000000",
         10906 => x"00000000",
         10907 => x"00000000",
         10908 => x"00000000",
         10909 => x"00000000",
         10910 => x"00000000",
         10911 => x"00000000",
         10912 => x"00000000",
         10913 => x"00000000",
         10914 => x"00000000",
         10915 => x"00000000",
         10916 => x"00000000",
         10917 => x"00000000",
         10918 => x"00000000",
         10919 => x"00000000",
         10920 => x"00000000",
         10921 => x"00000000",
         10922 => x"0000a2f4",
         10923 => x"01000000",
         10924 => x"0000a2fc",
         10925 => x"01000000",
         10926 => x"0000a304",
         10927 => x"02000000",
         10928 => x"cce0f2f3",
         10929 => x"cecff6f7",
         10930 => x"f8f9fafb",
         10931 => x"fcfdfeff",
         10932 => x"e1c1c2c3",
         10933 => x"c4c5c6e2",
         10934 => x"e3e4e5e6",
         10935 => x"ebeeeff4",
         10936 => x"00616263",
         10937 => x"64656667",
         10938 => x"68696b6a",
         10939 => x"2f2a2e2d",
         10940 => x"20212223",
         10941 => x"24252627",
         10942 => x"28294f2c",
         10943 => x"512b5749",
         10944 => x"55010203",
         10945 => x"04050607",
         10946 => x"08090a0b",
         10947 => x"0c0d0e0f",
         10948 => x"10111213",
         10949 => x"14151617",
         10950 => x"18191a52",
         10951 => x"5954be3c",
         10952 => x"c7818283",
         10953 => x"84858687",
         10954 => x"88898a8b",
         10955 => x"8c8d8e8f",
         10956 => x"90919293",
         10957 => x"94959697",
         10958 => x"98999abc",
         10959 => x"8040a5c0",
         10960 => x"00e80000",
         10961 => x"00000000",
         10962 => x"00000000",
         10963 => x"00000000",
         10964 => x"00000000",
         10965 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

