-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b83ff",
             1 => x"f80d0b0b",
             2 => x"0b93b704",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"9b040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b92fe",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b8294",
           162 => x"b0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93830400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b80cf",
           171 => x"942d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b80d1",
           179 => x"802d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"95040b0b",
           269 => x"0b8ca404",
           270 => x"0b0b0b8c",
           271 => x"b3040b0b",
           272 => x"0b8cc204",
           273 => x"0b0b0b8c",
           274 => x"d1040b0b",
           275 => x"0b8ce004",
           276 => x"0b0b0b8c",
           277 => x"ef040b0b",
           278 => x"0b8cfe04",
           279 => x"0b0b0b8d",
           280 => x"8d040b0b",
           281 => x"0b8d9c04",
           282 => x"0b0b0b8d",
           283 => x"ab040b0b",
           284 => x"0b8dbb04",
           285 => x"0b0b0b8d",
           286 => x"cb040b0b",
           287 => x"0b8ddb04",
           288 => x"0b0b0b8d",
           289 => x"eb040b0b",
           290 => x"0b8dfb04",
           291 => x"0b0b0b8e",
           292 => x"8b040b0b",
           293 => x"0b8e9b04",
           294 => x"0b0b0b8e",
           295 => x"ab040b0b",
           296 => x"0b8ebb04",
           297 => x"0b0b0b8e",
           298 => x"cb040b0b",
           299 => x"0b8edb04",
           300 => x"0b0b0b8e",
           301 => x"eb040b0b",
           302 => x"0b8efb04",
           303 => x"0b0b0b8f",
           304 => x"8b040b0b",
           305 => x"0b8f9b04",
           306 => x"0b0b0b8f",
           307 => x"ab040b0b",
           308 => x"0b8fbb04",
           309 => x"0b0b0b8f",
           310 => x"cb040b0b",
           311 => x"0b8fdb04",
           312 => x"0b0b0b8f",
           313 => x"eb040b0b",
           314 => x"0b8ffb04",
           315 => x"0b0b0b90",
           316 => x"8b040b0b",
           317 => x"0b909b04",
           318 => x"0b0b0b90",
           319 => x"ab040b0b",
           320 => x"0b90bb04",
           321 => x"0b0b0b90",
           322 => x"cb040b0b",
           323 => x"0b90db04",
           324 => x"0b0b0b90",
           325 => x"eb040b0b",
           326 => x"0b90fb04",
           327 => x"0b0b0b91",
           328 => x"8b040b0b",
           329 => x"0b919b04",
           330 => x"0b0b0b91",
           331 => x"ab040b0b",
           332 => x"0b91bb04",
           333 => x"0b0b0b91",
           334 => x"cb040b0b",
           335 => x"0b91db04",
           336 => x"0b0b0b91",
           337 => x"eb040b0b",
           338 => x"0b91fb04",
           339 => x"0b0b0b92",
           340 => x"8b040b0b",
           341 => x"0b929b04",
           342 => x"0b0b0b92",
           343 => x"ab040b0b",
           344 => x"0b92bb04",
           345 => x"0b0b0b92",
           346 => x"cb04ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0482b5b4",
           386 => x"0c80f4c6",
           387 => x"2d82b5b4",
           388 => x"0882d090",
           389 => x"0482b5b4",
           390 => x"0cbed22d",
           391 => x"82b5b408",
           392 => x"82d09004",
           393 => x"82b5b40c",
           394 => x"bb832d82",
           395 => x"b5b40882",
           396 => x"d0900482",
           397 => x"b5b40cb4",
           398 => x"fc2d82b5",
           399 => x"b40882d0",
           400 => x"900482b5",
           401 => x"b40c94ab",
           402 => x"2d82b5b4",
           403 => x"0882d090",
           404 => x"0482b5b4",
           405 => x"0cbce22d",
           406 => x"82b5b408",
           407 => x"82d09004",
           408 => x"82b5b40c",
           409 => x"b5b22d82",
           410 => x"b5b40882",
           411 => x"d0900482",
           412 => x"b5b40caf",
           413 => x"ab2d82b5",
           414 => x"b40882d0",
           415 => x"900482b5",
           416 => x"b40c93d6",
           417 => x"2d82b5b4",
           418 => x"0882d090",
           419 => x"0482b5b4",
           420 => x"0c96be2d",
           421 => x"82b5b408",
           422 => x"82d09004",
           423 => x"82b5b40c",
           424 => x"97cb2d82",
           425 => x"b5b40882",
           426 => x"d0900482",
           427 => x"b5b40c80",
           428 => x"f7f02d82",
           429 => x"b5b40882",
           430 => x"d0900482",
           431 => x"b5b40c80",
           432 => x"f8ce2d82",
           433 => x"b5b40882",
           434 => x"d0900482",
           435 => x"b5b40c80",
           436 => x"f08a2d82",
           437 => x"b5b40882",
           438 => x"d0900482",
           439 => x"b5b40c80",
           440 => x"f2822d82",
           441 => x"b5b40882",
           442 => x"d0900482",
           443 => x"b5b40c80",
           444 => x"f3b52d82",
           445 => x"b5b40882",
           446 => x"d0900482",
           447 => x"b5b40c81",
           448 => x"d7912d82",
           449 => x"b5b40882",
           450 => x"d0900482",
           451 => x"b5b40c81",
           452 => x"e4822d82",
           453 => x"b5b40882",
           454 => x"d0900482",
           455 => x"b5b40c81",
           456 => x"dbf62d82",
           457 => x"b5b40882",
           458 => x"d0900482",
           459 => x"b5b40c81",
           460 => x"def32d82",
           461 => x"b5b40882",
           462 => x"d0900482",
           463 => x"b5b40c81",
           464 => x"e9912d82",
           465 => x"b5b40882",
           466 => x"d0900482",
           467 => x"b5b40c81",
           468 => x"f1f12d82",
           469 => x"b5b40882",
           470 => x"d0900482",
           471 => x"b5b40c81",
           472 => x"e2e42d82",
           473 => x"b5b40882",
           474 => x"d0900482",
           475 => x"b5b40c81",
           476 => x"ecb02d82",
           477 => x"b5b40882",
           478 => x"d0900482",
           479 => x"b5b40c81",
           480 => x"edcf2d82",
           481 => x"b5b40882",
           482 => x"d0900482",
           483 => x"b5b40c81",
           484 => x"edee2d82",
           485 => x"b5b40882",
           486 => x"d0900482",
           487 => x"b5b40c81",
           488 => x"f5d82d82",
           489 => x"b5b40882",
           490 => x"d0900482",
           491 => x"b5b40c81",
           492 => x"f3be2d82",
           493 => x"b5b40882",
           494 => x"d0900482",
           495 => x"b5b40c81",
           496 => x"f8ac2d82",
           497 => x"b5b40882",
           498 => x"d0900482",
           499 => x"b5b40c81",
           500 => x"eef22d82",
           501 => x"b5b40882",
           502 => x"d0900482",
           503 => x"b5b40c81",
           504 => x"fbac2d82",
           505 => x"b5b40882",
           506 => x"d0900482",
           507 => x"b5b40c81",
           508 => x"fcad2d82",
           509 => x"b5b40882",
           510 => x"d0900482",
           511 => x"b5b40c81",
           512 => x"e4e22d82",
           513 => x"b5b40882",
           514 => x"d0900482",
           515 => x"b5b40c81",
           516 => x"e4bb2d82",
           517 => x"b5b40882",
           518 => x"d0900482",
           519 => x"b5b40c81",
           520 => x"e5e62d82",
           521 => x"b5b40882",
           522 => x"d0900482",
           523 => x"b5b40c81",
           524 => x"efc92d82",
           525 => x"b5b40882",
           526 => x"d0900482",
           527 => x"b5b40c81",
           528 => x"fd9e2d82",
           529 => x"b5b40882",
           530 => x"d0900482",
           531 => x"b5b40c81",
           532 => x"ffa82d82",
           533 => x"b5b40882",
           534 => x"d0900482",
           535 => x"b5b40c82",
           536 => x"82ea2d82",
           537 => x"b5b40882",
           538 => x"d0900482",
           539 => x"b5b40c81",
           540 => x"d6b02d82",
           541 => x"b5b40882",
           542 => x"d0900482",
           543 => x"b5b40c82",
           544 => x"85d62d82",
           545 => x"b5b40882",
           546 => x"d0900482",
           547 => x"b5b40c82",
           548 => x"948b2d82",
           549 => x"b5b40882",
           550 => x"d0900482",
           551 => x"b5b40c82",
           552 => x"91f72d82",
           553 => x"b5b40882",
           554 => x"d0900482",
           555 => x"b5b40c81",
           556 => x"a7eb2d82",
           557 => x"b5b40882",
           558 => x"d0900482",
           559 => x"b5b40c81",
           560 => x"a9d52d82",
           561 => x"b5b40882",
           562 => x"d0900482",
           563 => x"b5b40c81",
           564 => x"abb92d82",
           565 => x"b5b40882",
           566 => x"d0900482",
           567 => x"b5b40c80",
           568 => x"f0b32d82",
           569 => x"b5b40882",
           570 => x"d0900482",
           571 => x"b5b40c80",
           572 => x"f1d72d82",
           573 => x"b5b40882",
           574 => x"d0900482",
           575 => x"b5b40c80",
           576 => x"f5bb2d82",
           577 => x"b5b40882",
           578 => x"d0900482",
           579 => x"b5b40c80",
           580 => x"d6962d82",
           581 => x"b5b40882",
           582 => x"d0900482",
           583 => x"b5b40c81",
           584 => x"a1ff2d82",
           585 => x"b5b40882",
           586 => x"d0900482",
           587 => x"b5b40c81",
           588 => x"a2a72d82",
           589 => x"b5b40882",
           590 => x"d0900482",
           591 => x"b5b40c81",
           592 => x"a69f2d82",
           593 => x"b5b40882",
           594 => x"d0900482",
           595 => x"b5b40c81",
           596 => x"9ee92d82",
           597 => x"b5b40882",
           598 => x"d090043c",
           599 => x"04000010",
           600 => x"10101010",
           601 => x"10101010",
           602 => x"10101010",
           603 => x"10101010",
           604 => x"10101010",
           605 => x"10101010",
           606 => x"10101010",
           607 => x"10105351",
           608 => x"04000073",
           609 => x"81ff0673",
           610 => x"83060981",
           611 => x"05830510",
           612 => x"10102b07",
           613 => x"72fc060c",
           614 => x"51510472",
           615 => x"72807281",
           616 => x"06ff0509",
           617 => x"72060571",
           618 => x"1052720a",
           619 => x"100a5372",
           620 => x"ed385151",
           621 => x"53510482",
           622 => x"b5a87082",
           623 => x"cd84278e",
           624 => x"38807170",
           625 => x"8405530c",
           626 => x"0b0b0b93",
           627 => x"ba048c81",
           628 => x"5180eecb",
           629 => x"040082b5",
           630 => x"b4080282",
           631 => x"b5b40cfb",
           632 => x"3d0d82b5",
           633 => x"b4088c05",
           634 => x"7082b5b4",
           635 => x"08fc050c",
           636 => x"82b5b408",
           637 => x"fc050854",
           638 => x"82b5b408",
           639 => x"88050853",
           640 => x"82ccfc08",
           641 => x"5254849a",
           642 => x"3f82b5a8",
           643 => x"087082b5",
           644 => x"b408f805",
           645 => x"0c82b5b4",
           646 => x"08f80508",
           647 => x"7082b5a8",
           648 => x"0c515487",
           649 => x"3d0d82b5",
           650 => x"b40c0482",
           651 => x"b5b40802",
           652 => x"82b5b40c",
           653 => x"fb3d0d82",
           654 => x"b5b40890",
           655 => x"05088511",
           656 => x"33708132",
           657 => x"70810651",
           658 => x"51515271",
           659 => x"8f38800b",
           660 => x"82b5b408",
           661 => x"8c050825",
           662 => x"83388d39",
           663 => x"800b82b5",
           664 => x"b408f405",
           665 => x"0c81c439",
           666 => x"82b5b408",
           667 => x"8c0508ff",
           668 => x"0582b5b4",
           669 => x"088c050c",
           670 => x"800b82b5",
           671 => x"b408f805",
           672 => x"0c82b5b4",
           673 => x"08880508",
           674 => x"82b5b408",
           675 => x"fc050c82",
           676 => x"b5b408f8",
           677 => x"05088a2e",
           678 => x"80f63880",
           679 => x"0b82b5b4",
           680 => x"088c0508",
           681 => x"2580e938",
           682 => x"82b5b408",
           683 => x"90050851",
           684 => x"abb23f82",
           685 => x"b5a80870",
           686 => x"82b5b408",
           687 => x"f8050c52",
           688 => x"82b5b408",
           689 => x"f80508ff",
           690 => x"2e098106",
           691 => x"8d38800b",
           692 => x"82b5b408",
           693 => x"f4050c80",
           694 => x"d23982b5",
           695 => x"b408fc05",
           696 => x"0882b5b4",
           697 => x"08f80508",
           698 => x"53537173",
           699 => x"3482b5b4",
           700 => x"088c0508",
           701 => x"ff0582b5",
           702 => x"b4088c05",
           703 => x"0c82b5b4",
           704 => x"08fc0508",
           705 => x"810582b5",
           706 => x"b408fc05",
           707 => x"0cff8039",
           708 => x"82b5b408",
           709 => x"fc050852",
           710 => x"80723482",
           711 => x"b5b40888",
           712 => x"05087082",
           713 => x"b5b408f4",
           714 => x"050c5282",
           715 => x"b5b408f4",
           716 => x"050882b5",
           717 => x"a80c873d",
           718 => x"0d82b5b4",
           719 => x"0c0482b5",
           720 => x"b4080282",
           721 => x"b5b40cf4",
           722 => x"3d0d860b",
           723 => x"82b5b408",
           724 => x"e5053482",
           725 => x"b5b40888",
           726 => x"050882b5",
           727 => x"b408e005",
           728 => x"0cfe0a0b",
           729 => x"82b5b408",
           730 => x"e8050c82",
           731 => x"b5b40890",
           732 => x"057082b5",
           733 => x"b408fc05",
           734 => x"0c82b5b4",
           735 => x"08fc0508",
           736 => x"5482b5b4",
           737 => x"088c0508",
           738 => x"5382b5b4",
           739 => x"08e00570",
           740 => x"53515481",
           741 => x"8d3f82b5",
           742 => x"a8087082",
           743 => x"b5b408dc",
           744 => x"050c82b5",
           745 => x"b408ec05",
           746 => x"0882b5b4",
           747 => x"08880508",
           748 => x"05515480",
           749 => x"743482b5",
           750 => x"b408dc05",
           751 => x"087082b5",
           752 => x"a80c548e",
           753 => x"3d0d82b5",
           754 => x"b40c0482",
           755 => x"b5b40802",
           756 => x"82b5b40c",
           757 => x"fb3d0d82",
           758 => x"b5b40890",
           759 => x"057082b5",
           760 => x"b408fc05",
           761 => x"0c82b5b4",
           762 => x"08fc0508",
           763 => x"5482b5b4",
           764 => x"088c0508",
           765 => x"5382b5b4",
           766 => x"08880508",
           767 => x"5254a33f",
           768 => x"82b5a808",
           769 => x"7082b5b4",
           770 => x"08f8050c",
           771 => x"82b5b408",
           772 => x"f8050870",
           773 => x"82b5a80c",
           774 => x"5154873d",
           775 => x"0d82b5b4",
           776 => x"0c0482b5",
           777 => x"b4080282",
           778 => x"b5b40ced",
           779 => x"3d0d800b",
           780 => x"82b5b408",
           781 => x"e4052382",
           782 => x"b5b40888",
           783 => x"05085380",
           784 => x"0b8c140c",
           785 => x"82b5b408",
           786 => x"88050885",
           787 => x"11337081",
           788 => x"2a708132",
           789 => x"70810651",
           790 => x"51515153",
           791 => x"72802e8d",
           792 => x"38ff0b82",
           793 => x"b5b408e0",
           794 => x"050c96ac",
           795 => x"3982b5b4",
           796 => x"088c0508",
           797 => x"53723353",
           798 => x"7282b5b4",
           799 => x"08f80534",
           800 => x"7281ff06",
           801 => x"5372802e",
           802 => x"95fa3882",
           803 => x"b5b4088c",
           804 => x"05088105",
           805 => x"82b5b408",
           806 => x"8c050c82",
           807 => x"b5b408e4",
           808 => x"05227081",
           809 => x"06515372",
           810 => x"802e958b",
           811 => x"3882b5b4",
           812 => x"08f80533",
           813 => x"53af7327",
           814 => x"81fc3882",
           815 => x"b5b408f8",
           816 => x"05335372",
           817 => x"b92681ee",
           818 => x"3882b5b4",
           819 => x"08f80533",
           820 => x"5372b02e",
           821 => x"09810680",
           822 => x"c53882b5",
           823 => x"b408e805",
           824 => x"3370982b",
           825 => x"70982c51",
           826 => x"515372b2",
           827 => x"3882b5b4",
           828 => x"08e40522",
           829 => x"70832a70",
           830 => x"81327081",
           831 => x"06515151",
           832 => x"5372802e",
           833 => x"993882b5",
           834 => x"b408e405",
           835 => x"22708280",
           836 => x"07515372",
           837 => x"82b5b408",
           838 => x"e40523fe",
           839 => x"d03982b5",
           840 => x"b408e805",
           841 => x"3370982b",
           842 => x"70982c70",
           843 => x"70832b72",
           844 => x"11731151",
           845 => x"51515351",
           846 => x"55537282",
           847 => x"b5b408e8",
           848 => x"053482b5",
           849 => x"b408e805",
           850 => x"335482b5",
           851 => x"b408f805",
           852 => x"337015d0",
           853 => x"11515153",
           854 => x"7282b5b4",
           855 => x"08e80534",
           856 => x"82b5b408",
           857 => x"e8053370",
           858 => x"982b7098",
           859 => x"2c515153",
           860 => x"7280258b",
           861 => x"3880ff0b",
           862 => x"82b5b408",
           863 => x"e8053482",
           864 => x"b5b408e4",
           865 => x"05227083",
           866 => x"2a708106",
           867 => x"51515372",
           868 => x"fddb3882",
           869 => x"b5b408e8",
           870 => x"05337088",
           871 => x"2b70902b",
           872 => x"70902c70",
           873 => x"882c5151",
           874 => x"51515372",
           875 => x"82b5b408",
           876 => x"ec0523fd",
           877 => x"b83982b5",
           878 => x"b408e405",
           879 => x"2270832a",
           880 => x"70810651",
           881 => x"51537280",
           882 => x"2e9d3882",
           883 => x"b5b408e8",
           884 => x"05337098",
           885 => x"2b70982c",
           886 => x"51515372",
           887 => x"8a38810b",
           888 => x"82b5b408",
           889 => x"e8053482",
           890 => x"b5b408f8",
           891 => x"0533e011",
           892 => x"82b5b408",
           893 => x"c4050c53",
           894 => x"82b5b408",
           895 => x"c4050880",
           896 => x"d8269294",
           897 => x"3882b5b4",
           898 => x"08c40508",
           899 => x"70822b82",
           900 => x"95fc1170",
           901 => x"08515151",
           902 => x"53720482",
           903 => x"b5b408e4",
           904 => x"05227090",
           905 => x"07515372",
           906 => x"82b5b408",
           907 => x"e4052382",
           908 => x"b5b408e4",
           909 => x"052270a0",
           910 => x"07515372",
           911 => x"82b5b408",
           912 => x"e40523fc",
           913 => x"a83982b5",
           914 => x"b408e405",
           915 => x"22708180",
           916 => x"07515372",
           917 => x"82b5b408",
           918 => x"e40523fc",
           919 => x"903982b5",
           920 => x"b408e405",
           921 => x"227080c0",
           922 => x"07515372",
           923 => x"82b5b408",
           924 => x"e40523fb",
           925 => x"f83982b5",
           926 => x"b408e405",
           927 => x"22708807",
           928 => x"51537282",
           929 => x"b5b408e4",
           930 => x"0523800b",
           931 => x"82b5b408",
           932 => x"e80534fb",
           933 => x"d83982b5",
           934 => x"b408e405",
           935 => x"22708407",
           936 => x"51537282",
           937 => x"b5b408e4",
           938 => x"0523fbc1",
           939 => x"39bf0b82",
           940 => x"b5b408fc",
           941 => x"053482b5",
           942 => x"b408ec05",
           943 => x"22ff1151",
           944 => x"537282b5",
           945 => x"b408ec05",
           946 => x"2380e30b",
           947 => x"82b5b408",
           948 => x"f805348d",
           949 => x"a83982b5",
           950 => x"b4089005",
           951 => x"0882b5b4",
           952 => x"08900508",
           953 => x"840582b5",
           954 => x"b4089005",
           955 => x"0c700851",
           956 => x"537282b5",
           957 => x"b408fc05",
           958 => x"3482b5b4",
           959 => x"08ec0522",
           960 => x"ff115153",
           961 => x"7282b5b4",
           962 => x"08ec0523",
           963 => x"8cef3982",
           964 => x"b5b40890",
           965 => x"050882b5",
           966 => x"b4089005",
           967 => x"08840582",
           968 => x"b5b40890",
           969 => x"050c7008",
           970 => x"82b5b408",
           971 => x"fc050c82",
           972 => x"b5b408e4",
           973 => x"05227083",
           974 => x"2a708106",
           975 => x"51515153",
           976 => x"72802eab",
           977 => x"3882b5b4",
           978 => x"08e80533",
           979 => x"70982b53",
           980 => x"72982c53",
           981 => x"82b5b408",
           982 => x"fc050852",
           983 => x"53adfa3f",
           984 => x"82b5a808",
           985 => x"537282b5",
           986 => x"b408f405",
           987 => x"23993982",
           988 => x"b5b408fc",
           989 => x"050851a8",
           990 => x"ac3f82b5",
           991 => x"a8085372",
           992 => x"82b5b408",
           993 => x"f4052382",
           994 => x"b5b408ec",
           995 => x"05225382",
           996 => x"b5b408f4",
           997 => x"05227371",
           998 => x"31545472",
           999 => x"82b5b408",
          1000 => x"ec05238b",
          1001 => x"d83982b5",
          1002 => x"b4089005",
          1003 => x"0882b5b4",
          1004 => x"08900508",
          1005 => x"840582b5",
          1006 => x"b4089005",
          1007 => x"0c700882",
          1008 => x"b5b408fc",
          1009 => x"050c82b5",
          1010 => x"b408e405",
          1011 => x"2270832a",
          1012 => x"70810651",
          1013 => x"51515372",
          1014 => x"802eab38",
          1015 => x"82b5b408",
          1016 => x"e8053370",
          1017 => x"982b5372",
          1018 => x"982c5382",
          1019 => x"b5b408fc",
          1020 => x"05085253",
          1021 => x"ace33f82",
          1022 => x"b5a80853",
          1023 => x"7282b5b4",
          1024 => x"08f40523",
          1025 => x"993982b5",
          1026 => x"b408fc05",
          1027 => x"0851a795",
          1028 => x"3f82b5a8",
          1029 => x"08537282",
          1030 => x"b5b408f4",
          1031 => x"052382b5",
          1032 => x"b408ec05",
          1033 => x"225382b5",
          1034 => x"b408f405",
          1035 => x"22737131",
          1036 => x"54547282",
          1037 => x"b5b408ec",
          1038 => x"05238ac1",
          1039 => x"3982b5b4",
          1040 => x"08e40522",
          1041 => x"70822a70",
          1042 => x"81065151",
          1043 => x"5372802e",
          1044 => x"a43882b5",
          1045 => x"b4089005",
          1046 => x"0882b5b4",
          1047 => x"08900508",
          1048 => x"840582b5",
          1049 => x"b4089005",
          1050 => x"0c700882",
          1051 => x"b5b408dc",
          1052 => x"050c53a2",
          1053 => x"3982b5b4",
          1054 => x"08900508",
          1055 => x"82b5b408",
          1056 => x"90050884",
          1057 => x"0582b5b4",
          1058 => x"0890050c",
          1059 => x"700882b5",
          1060 => x"b408dc05",
          1061 => x"0c5382b5",
          1062 => x"b408dc05",
          1063 => x"0882b5b4",
          1064 => x"08fc050c",
          1065 => x"82b5b408",
          1066 => x"fc050880",
          1067 => x"25a43882",
          1068 => x"b5b408e4",
          1069 => x"05227082",
          1070 => x"07515372",
          1071 => x"82b5b408",
          1072 => x"e4052382",
          1073 => x"b5b408fc",
          1074 => x"05083082",
          1075 => x"b5b408fc",
          1076 => x"050c82b5",
          1077 => x"b408e405",
          1078 => x"2270ffbf",
          1079 => x"06515372",
          1080 => x"82b5b408",
          1081 => x"e4052381",
          1082 => x"af39880b",
          1083 => x"82b5b408",
          1084 => x"f40523a9",
          1085 => x"3982b5b4",
          1086 => x"08e40522",
          1087 => x"7080c007",
          1088 => x"51537282",
          1089 => x"b5b408e4",
          1090 => x"052380f8",
          1091 => x"0b82b5b4",
          1092 => x"08f80534",
          1093 => x"900b82b5",
          1094 => x"b408f405",
          1095 => x"2382b5b4",
          1096 => x"08e40522",
          1097 => x"70822a70",
          1098 => x"81065151",
          1099 => x"5372802e",
          1100 => x"a43882b5",
          1101 => x"b4089005",
          1102 => x"0882b5b4",
          1103 => x"08900508",
          1104 => x"840582b5",
          1105 => x"b4089005",
          1106 => x"0c700882",
          1107 => x"b5b408d8",
          1108 => x"050c53a2",
          1109 => x"3982b5b4",
          1110 => x"08900508",
          1111 => x"82b5b408",
          1112 => x"90050884",
          1113 => x"0582b5b4",
          1114 => x"0890050c",
          1115 => x"700882b5",
          1116 => x"b408d805",
          1117 => x"0c5382b5",
          1118 => x"b408d805",
          1119 => x"0882b5b4",
          1120 => x"08fc050c",
          1121 => x"82b5b408",
          1122 => x"e4052270",
          1123 => x"cf065153",
          1124 => x"7282b5b4",
          1125 => x"08e40523",
          1126 => x"82b5b80b",
          1127 => x"82b5b408",
          1128 => x"f0050c82",
          1129 => x"b5b408f0",
          1130 => x"050882b5",
          1131 => x"b408f405",
          1132 => x"2282b5b4",
          1133 => x"08fc0508",
          1134 => x"71557054",
          1135 => x"565455af",
          1136 => x"953f82b5",
          1137 => x"a8085372",
          1138 => x"753482b5",
          1139 => x"b408f005",
          1140 => x"0882b5b4",
          1141 => x"08d4050c",
          1142 => x"82b5b408",
          1143 => x"f0050870",
          1144 => x"33515389",
          1145 => x"7327a438",
          1146 => x"82b5b408",
          1147 => x"f0050853",
          1148 => x"72335482",
          1149 => x"b5b408f8",
          1150 => x"05337015",
          1151 => x"df115151",
          1152 => x"537282b5",
          1153 => x"b408d005",
          1154 => x"34973982",
          1155 => x"b5b408f0",
          1156 => x"05085372",
          1157 => x"33b01151",
          1158 => x"537282b5",
          1159 => x"b408d005",
          1160 => x"3482b5b4",
          1161 => x"08d40508",
          1162 => x"5382b5b4",
          1163 => x"08d00533",
          1164 => x"733482b5",
          1165 => x"b408f005",
          1166 => x"08810582",
          1167 => x"b5b408f0",
          1168 => x"050c82b5",
          1169 => x"b408f405",
          1170 => x"22705382",
          1171 => x"b5b408fc",
          1172 => x"05085253",
          1173 => x"adcd3f82",
          1174 => x"b5a80870",
          1175 => x"82b5b408",
          1176 => x"fc050c53",
          1177 => x"82b5b408",
          1178 => x"fc050880",
          1179 => x"2e8438fe",
          1180 => x"b23982b5",
          1181 => x"b408f005",
          1182 => x"0882b5b8",
          1183 => x"54557254",
          1184 => x"74707531",
          1185 => x"51537282",
          1186 => x"b5b408fc",
          1187 => x"053482b5",
          1188 => x"b408e405",
          1189 => x"2270b206",
          1190 => x"51537280",
          1191 => x"2e943882",
          1192 => x"b5b408ec",
          1193 => x"0522ff11",
          1194 => x"51537282",
          1195 => x"b5b408ec",
          1196 => x"052382b5",
          1197 => x"b408e405",
          1198 => x"2270862a",
          1199 => x"70810651",
          1200 => x"51537280",
          1201 => x"2e80e738",
          1202 => x"82b5b408",
          1203 => x"ec052270",
          1204 => x"902b82b5",
          1205 => x"b408cc05",
          1206 => x"0c82b5b4",
          1207 => x"08cc0508",
          1208 => x"902c82b5",
          1209 => x"b408cc05",
          1210 => x"0c82b5b4",
          1211 => x"08f40522",
          1212 => x"51537290",
          1213 => x"2e098106",
          1214 => x"953882b5",
          1215 => x"b408cc05",
          1216 => x"08fe0553",
          1217 => x"7282b5b4",
          1218 => x"08c80523",
          1219 => x"933982b5",
          1220 => x"b408cc05",
          1221 => x"08ff0553",
          1222 => x"7282b5b4",
          1223 => x"08c80523",
          1224 => x"82b5b408",
          1225 => x"c8052282",
          1226 => x"b5b408ec",
          1227 => x"052382b5",
          1228 => x"b408e405",
          1229 => x"2270832a",
          1230 => x"70810651",
          1231 => x"51537280",
          1232 => x"2e80d038",
          1233 => x"82b5b408",
          1234 => x"e8053370",
          1235 => x"982b7098",
          1236 => x"2c82b5b4",
          1237 => x"08fc0533",
          1238 => x"57515153",
          1239 => x"72742497",
          1240 => x"3882b5b4",
          1241 => x"08e40522",
          1242 => x"70f70651",
          1243 => x"537282b5",
          1244 => x"b408e405",
          1245 => x"239d3982",
          1246 => x"b5b408e8",
          1247 => x"05335382",
          1248 => x"b5b408fc",
          1249 => x"05337371",
          1250 => x"31545472",
          1251 => x"82b5b408",
          1252 => x"e8053482",
          1253 => x"b5b408e4",
          1254 => x"05227083",
          1255 => x"2a708106",
          1256 => x"51515372",
          1257 => x"802eb138",
          1258 => x"82b5b408",
          1259 => x"e8053370",
          1260 => x"882b7090",
          1261 => x"2b70902c",
          1262 => x"70882c51",
          1263 => x"51515153",
          1264 => x"725482b5",
          1265 => x"b408ec05",
          1266 => x"22707531",
          1267 => x"51537282",
          1268 => x"b5b408ec",
          1269 => x"0523af39",
          1270 => x"82b5b408",
          1271 => x"fc053370",
          1272 => x"882b7090",
          1273 => x"2b70902c",
          1274 => x"70882c51",
          1275 => x"51515153",
          1276 => x"725482b5",
          1277 => x"b408ec05",
          1278 => x"22707531",
          1279 => x"51537282",
          1280 => x"b5b408ec",
          1281 => x"052382b5",
          1282 => x"b408e405",
          1283 => x"22708380",
          1284 => x"06515372",
          1285 => x"b03882b5",
          1286 => x"b408ec05",
          1287 => x"22ff1154",
          1288 => x"547282b5",
          1289 => x"b408ec05",
          1290 => x"2373902b",
          1291 => x"70902c51",
          1292 => x"53807325",
          1293 => x"903882b5",
          1294 => x"b4088805",
          1295 => x"0852a051",
          1296 => x"96903fd2",
          1297 => x"3982b5b4",
          1298 => x"08e40522",
          1299 => x"70812a70",
          1300 => x"81065151",
          1301 => x"5372802e",
          1302 => x"913882b5",
          1303 => x"b4088805",
          1304 => x"0852ad51",
          1305 => x"95ec3f80",
          1306 => x"c73982b5",
          1307 => x"b408e405",
          1308 => x"2270842a",
          1309 => x"70810651",
          1310 => x"51537280",
          1311 => x"2e903882",
          1312 => x"b5b40888",
          1313 => x"050852ab",
          1314 => x"5195c73f",
          1315 => x"a33982b5",
          1316 => x"b408e405",
          1317 => x"2270852a",
          1318 => x"70810651",
          1319 => x"51537280",
          1320 => x"2e8e3882",
          1321 => x"b5b40888",
          1322 => x"050852a0",
          1323 => x"5195a33f",
          1324 => x"82b5b408",
          1325 => x"e4052270",
          1326 => x"862a7081",
          1327 => x"06515153",
          1328 => x"72802eb1",
          1329 => x"3882b5b4",
          1330 => x"08880508",
          1331 => x"52b05195",
          1332 => x"813f82b5",
          1333 => x"b408f405",
          1334 => x"22537290",
          1335 => x"2e098106",
          1336 => x"943882b5",
          1337 => x"b4088805",
          1338 => x"085282b5",
          1339 => x"b408f805",
          1340 => x"335194de",
          1341 => x"3f82b5b4",
          1342 => x"08e40522",
          1343 => x"70882a70",
          1344 => x"81065151",
          1345 => x"5372802e",
          1346 => x"b03882b5",
          1347 => x"b408ec05",
          1348 => x"22ff1154",
          1349 => x"547282b5",
          1350 => x"b408ec05",
          1351 => x"2373902b",
          1352 => x"70902c51",
          1353 => x"53807325",
          1354 => x"903882b5",
          1355 => x"b4088805",
          1356 => x"0852b051",
          1357 => x"949c3fd2",
          1358 => x"3982b5b4",
          1359 => x"08e40522",
          1360 => x"70832a70",
          1361 => x"81065151",
          1362 => x"5372802e",
          1363 => x"b03882b5",
          1364 => x"b408e805",
          1365 => x"33ff1154",
          1366 => x"547282b5",
          1367 => x"b408e805",
          1368 => x"3473982b",
          1369 => x"70982c51",
          1370 => x"53807325",
          1371 => x"903882b5",
          1372 => x"b4088805",
          1373 => x"0852b051",
          1374 => x"93d83fd2",
          1375 => x"3982b5b4",
          1376 => x"08e40522",
          1377 => x"70872a70",
          1378 => x"81065151",
          1379 => x"5372b038",
          1380 => x"82b5b408",
          1381 => x"ec0522ff",
          1382 => x"11545472",
          1383 => x"82b5b408",
          1384 => x"ec052373",
          1385 => x"902b7090",
          1386 => x"2c515380",
          1387 => x"73259038",
          1388 => x"82b5b408",
          1389 => x"88050852",
          1390 => x"a0519396",
          1391 => x"3fd23982",
          1392 => x"b5b408f8",
          1393 => x"05335372",
          1394 => x"80e32e09",
          1395 => x"81069738",
          1396 => x"82b5b408",
          1397 => x"88050852",
          1398 => x"82b5b408",
          1399 => x"fc053351",
          1400 => x"92f03f81",
          1401 => x"ee3982b5",
          1402 => x"b408f805",
          1403 => x"33537280",
          1404 => x"f32e0981",
          1405 => x"0680cb38",
          1406 => x"82b5b408",
          1407 => x"f40522ff",
          1408 => x"11515372",
          1409 => x"82b5b408",
          1410 => x"f4052372",
          1411 => x"83ffff06",
          1412 => x"537283ff",
          1413 => x"ff2e81bb",
          1414 => x"3882b5b4",
          1415 => x"08880508",
          1416 => x"5282b5b4",
          1417 => x"08fc0508",
          1418 => x"70335282",
          1419 => x"b5b408fc",
          1420 => x"05088105",
          1421 => x"82b5b408",
          1422 => x"fc050c53",
          1423 => x"92943fff",
          1424 => x"b73982b5",
          1425 => x"b408f805",
          1426 => x"33537280",
          1427 => x"d32e0981",
          1428 => x"0680cb38",
          1429 => x"82b5b408",
          1430 => x"f40522ff",
          1431 => x"11515372",
          1432 => x"82b5b408",
          1433 => x"f4052372",
          1434 => x"83ffff06",
          1435 => x"537283ff",
          1436 => x"ff2e80df",
          1437 => x"3882b5b4",
          1438 => x"08880508",
          1439 => x"5282b5b4",
          1440 => x"08fc0508",
          1441 => x"70335253",
          1442 => x"91c83f82",
          1443 => x"b5b408fc",
          1444 => x"05088105",
          1445 => x"82b5b408",
          1446 => x"fc050cff",
          1447 => x"b73982b5",
          1448 => x"b408f005",
          1449 => x"0882b5b8",
          1450 => x"2ea93882",
          1451 => x"b5b40888",
          1452 => x"05085282",
          1453 => x"b5b408f0",
          1454 => x"0508ff05",
          1455 => x"82b5b408",
          1456 => x"f0050c82",
          1457 => x"b5b408f0",
          1458 => x"05087033",
          1459 => x"52539182",
          1460 => x"3fcc3982",
          1461 => x"b5b408e4",
          1462 => x"05227087",
          1463 => x"2a708106",
          1464 => x"51515372",
          1465 => x"802e80c3",
          1466 => x"3882b5b4",
          1467 => x"08ec0522",
          1468 => x"ff115454",
          1469 => x"7282b5b4",
          1470 => x"08ec0523",
          1471 => x"73902b70",
          1472 => x"902c5153",
          1473 => x"807325a3",
          1474 => x"3882b5b4",
          1475 => x"08880508",
          1476 => x"52a05190",
          1477 => x"bd3fd239",
          1478 => x"82b5b408",
          1479 => x"88050852",
          1480 => x"82b5b408",
          1481 => x"f8053351",
          1482 => x"90a83f80",
          1483 => x"0b82b5b4",
          1484 => x"08e40523",
          1485 => x"eab73982",
          1486 => x"b5b408f8",
          1487 => x"05335372",
          1488 => x"a52e0981",
          1489 => x"06a83881",
          1490 => x"0b82b5b4",
          1491 => x"08e40523",
          1492 => x"800b82b5",
          1493 => x"b408ec05",
          1494 => x"23800b82",
          1495 => x"b5b408e8",
          1496 => x"05348a0b",
          1497 => x"82b5b408",
          1498 => x"f40523ea",
          1499 => x"803982b5",
          1500 => x"b4088805",
          1501 => x"085282b5",
          1502 => x"b408f805",
          1503 => x"33518fd2",
          1504 => x"3fe9ea39",
          1505 => x"82b5b408",
          1506 => x"8805088c",
          1507 => x"11087082",
          1508 => x"b5b408e0",
          1509 => x"050c5153",
          1510 => x"82b5b408",
          1511 => x"e0050882",
          1512 => x"b5a80c95",
          1513 => x"3d0d82b5",
          1514 => x"b40c0482",
          1515 => x"b5b40802",
          1516 => x"82b5b40c",
          1517 => x"f73d0d80",
          1518 => x"0b82b5b4",
          1519 => x"08f00534",
          1520 => x"82b5b408",
          1521 => x"8c050853",
          1522 => x"80730c82",
          1523 => x"b5b40888",
          1524 => x"05087008",
          1525 => x"51537233",
          1526 => x"537282b5",
          1527 => x"b408f805",
          1528 => x"347281ff",
          1529 => x"065372a0",
          1530 => x"2e098106",
          1531 => x"913882b5",
          1532 => x"b4088805",
          1533 => x"08700881",
          1534 => x"05710c53",
          1535 => x"ce3982b5",
          1536 => x"b408f805",
          1537 => x"335372ad",
          1538 => x"2e098106",
          1539 => x"a438810b",
          1540 => x"82b5b408",
          1541 => x"f0053482",
          1542 => x"b5b40888",
          1543 => x"05087008",
          1544 => x"8105710c",
          1545 => x"70085153",
          1546 => x"723382b5",
          1547 => x"b408f805",
          1548 => x"3482b5b4",
          1549 => x"08f80533",
          1550 => x"5372b02e",
          1551 => x"09810681",
          1552 => x"dc3882b5",
          1553 => x"b4088805",
          1554 => x"08700881",
          1555 => x"05710c70",
          1556 => x"08515372",
          1557 => x"3382b5b4",
          1558 => x"08f80534",
          1559 => x"82b5b408",
          1560 => x"f8053382",
          1561 => x"b5b408e8",
          1562 => x"050c82b5",
          1563 => x"b408e805",
          1564 => x"0880e22e",
          1565 => x"b63882b5",
          1566 => x"b408e805",
          1567 => x"0880f82e",
          1568 => x"843880cd",
          1569 => x"39900b82",
          1570 => x"b5b408f4",
          1571 => x"053482b5",
          1572 => x"b4088805",
          1573 => x"08700881",
          1574 => x"05710c70",
          1575 => x"08515372",
          1576 => x"3382b5b4",
          1577 => x"08f80534",
          1578 => x"81a43982",
          1579 => x"0b82b5b4",
          1580 => x"08f40534",
          1581 => x"82b5b408",
          1582 => x"88050870",
          1583 => x"08810571",
          1584 => x"0c700851",
          1585 => x"53723382",
          1586 => x"b5b408f8",
          1587 => x"053480fe",
          1588 => x"3982b5b4",
          1589 => x"08f80533",
          1590 => x"5372a026",
          1591 => x"8d38810b",
          1592 => x"82b5b408",
          1593 => x"ec050c83",
          1594 => x"803982b5",
          1595 => x"b408f805",
          1596 => x"3353af73",
          1597 => x"27903882",
          1598 => x"b5b408f8",
          1599 => x"05335372",
          1600 => x"b9268338",
          1601 => x"8d39800b",
          1602 => x"82b5b408",
          1603 => x"ec050c82",
          1604 => x"d839880b",
          1605 => x"82b5b408",
          1606 => x"f40534b2",
          1607 => x"3982b5b4",
          1608 => x"08f80533",
          1609 => x"53af7327",
          1610 => x"903882b5",
          1611 => x"b408f805",
          1612 => x"335372b9",
          1613 => x"2683388d",
          1614 => x"39800b82",
          1615 => x"b5b408ec",
          1616 => x"050c82a5",
          1617 => x"398a0b82",
          1618 => x"b5b408f4",
          1619 => x"0534800b",
          1620 => x"82b5b408",
          1621 => x"fc050c82",
          1622 => x"b5b408f8",
          1623 => x"053353a0",
          1624 => x"732781cf",
          1625 => x"3882b5b4",
          1626 => x"08f80533",
          1627 => x"5380e073",
          1628 => x"27943882",
          1629 => x"b5b408f8",
          1630 => x"0533e011",
          1631 => x"51537282",
          1632 => x"b5b408f8",
          1633 => x"053482b5",
          1634 => x"b408f805",
          1635 => x"33d01151",
          1636 => x"537282b5",
          1637 => x"b408f805",
          1638 => x"3482b5b4",
          1639 => x"08f80533",
          1640 => x"53907327",
          1641 => x"ad3882b5",
          1642 => x"b408f805",
          1643 => x"33f91151",
          1644 => x"537282b5",
          1645 => x"b408f805",
          1646 => x"3482b5b4",
          1647 => x"08f80533",
          1648 => x"53728926",
          1649 => x"8d38800b",
          1650 => x"82b5b408",
          1651 => x"ec050c81",
          1652 => x"983982b5",
          1653 => x"b408f805",
          1654 => x"3382b5b4",
          1655 => x"08f40533",
          1656 => x"54547274",
          1657 => x"268d3880",
          1658 => x"0b82b5b4",
          1659 => x"08ec050c",
          1660 => x"80f73982",
          1661 => x"b5b408f4",
          1662 => x"05337082",
          1663 => x"b5b408fc",
          1664 => x"05082982",
          1665 => x"b5b408f8",
          1666 => x"05337012",
          1667 => x"82b5b408",
          1668 => x"fc050c82",
          1669 => x"b5b40888",
          1670 => x"05087008",
          1671 => x"8105710c",
          1672 => x"70085151",
          1673 => x"52555372",
          1674 => x"3382b5b4",
          1675 => x"08f80534",
          1676 => x"fea53982",
          1677 => x"b5b408f0",
          1678 => x"05335372",
          1679 => x"802e9038",
          1680 => x"82b5b408",
          1681 => x"fc050830",
          1682 => x"82b5b408",
          1683 => x"fc050c82",
          1684 => x"b5b4088c",
          1685 => x"050882b5",
          1686 => x"b408fc05",
          1687 => x"08710c53",
          1688 => x"810b82b5",
          1689 => x"b408ec05",
          1690 => x"0c82b5b4",
          1691 => x"08ec0508",
          1692 => x"82b5a80c",
          1693 => x"8b3d0d82",
          1694 => x"b5b40c04",
          1695 => x"82b5b408",
          1696 => x"0282b5b4",
          1697 => x"0cfd3d0d",
          1698 => x"82ccf808",
          1699 => x"5382b5b4",
          1700 => x"088c0508",
          1701 => x"5282b5b4",
          1702 => x"08880508",
          1703 => x"51df8c3f",
          1704 => x"82b5a808",
          1705 => x"7082b5a8",
          1706 => x"0c54853d",
          1707 => x"0d82b5b4",
          1708 => x"0c0482b5",
          1709 => x"b4080282",
          1710 => x"b5b40cf7",
          1711 => x"3d0d800b",
          1712 => x"82b5b408",
          1713 => x"f0053482",
          1714 => x"b5b4088c",
          1715 => x"05085380",
          1716 => x"730c82b5",
          1717 => x"b4088805",
          1718 => x"08700851",
          1719 => x"53723353",
          1720 => x"7282b5b4",
          1721 => x"08f80534",
          1722 => x"7281ff06",
          1723 => x"5372a02e",
          1724 => x"09810691",
          1725 => x"3882b5b4",
          1726 => x"08880508",
          1727 => x"70088105",
          1728 => x"710c53ce",
          1729 => x"3982b5b4",
          1730 => x"08f80533",
          1731 => x"5372ad2e",
          1732 => x"098106a4",
          1733 => x"38810b82",
          1734 => x"b5b408f0",
          1735 => x"053482b5",
          1736 => x"b4088805",
          1737 => x"08700881",
          1738 => x"05710c70",
          1739 => x"08515372",
          1740 => x"3382b5b4",
          1741 => x"08f80534",
          1742 => x"82b5b408",
          1743 => x"f8053353",
          1744 => x"72b02e09",
          1745 => x"810681dc",
          1746 => x"3882b5b4",
          1747 => x"08880508",
          1748 => x"70088105",
          1749 => x"710c7008",
          1750 => x"51537233",
          1751 => x"82b5b408",
          1752 => x"f8053482",
          1753 => x"b5b408f8",
          1754 => x"053382b5",
          1755 => x"b408e805",
          1756 => x"0c82b5b4",
          1757 => x"08e80508",
          1758 => x"80e22eb6",
          1759 => x"3882b5b4",
          1760 => x"08e80508",
          1761 => x"80f82e84",
          1762 => x"3880cd39",
          1763 => x"900b82b5",
          1764 => x"b408f405",
          1765 => x"3482b5b4",
          1766 => x"08880508",
          1767 => x"70088105",
          1768 => x"710c7008",
          1769 => x"51537233",
          1770 => x"82b5b408",
          1771 => x"f8053481",
          1772 => x"a439820b",
          1773 => x"82b5b408",
          1774 => x"f4053482",
          1775 => x"b5b40888",
          1776 => x"05087008",
          1777 => x"8105710c",
          1778 => x"70085153",
          1779 => x"723382b5",
          1780 => x"b408f805",
          1781 => x"3480fe39",
          1782 => x"82b5b408",
          1783 => x"f8053353",
          1784 => x"72a0268d",
          1785 => x"38810b82",
          1786 => x"b5b408ec",
          1787 => x"050c8380",
          1788 => x"3982b5b4",
          1789 => x"08f80533",
          1790 => x"53af7327",
          1791 => x"903882b5",
          1792 => x"b408f805",
          1793 => x"335372b9",
          1794 => x"2683388d",
          1795 => x"39800b82",
          1796 => x"b5b408ec",
          1797 => x"050c82d8",
          1798 => x"39880b82",
          1799 => x"b5b408f4",
          1800 => x"0534b239",
          1801 => x"82b5b408",
          1802 => x"f8053353",
          1803 => x"af732790",
          1804 => x"3882b5b4",
          1805 => x"08f80533",
          1806 => x"5372b926",
          1807 => x"83388d39",
          1808 => x"800b82b5",
          1809 => x"b408ec05",
          1810 => x"0c82a539",
          1811 => x"8a0b82b5",
          1812 => x"b408f405",
          1813 => x"34800b82",
          1814 => x"b5b408fc",
          1815 => x"050c82b5",
          1816 => x"b408f805",
          1817 => x"3353a073",
          1818 => x"2781cf38",
          1819 => x"82b5b408",
          1820 => x"f8053353",
          1821 => x"80e07327",
          1822 => x"943882b5",
          1823 => x"b408f805",
          1824 => x"33e01151",
          1825 => x"537282b5",
          1826 => x"b408f805",
          1827 => x"3482b5b4",
          1828 => x"08f80533",
          1829 => x"d0115153",
          1830 => x"7282b5b4",
          1831 => x"08f80534",
          1832 => x"82b5b408",
          1833 => x"f8053353",
          1834 => x"907327ad",
          1835 => x"3882b5b4",
          1836 => x"08f80533",
          1837 => x"f9115153",
          1838 => x"7282b5b4",
          1839 => x"08f80534",
          1840 => x"82b5b408",
          1841 => x"f8053353",
          1842 => x"7289268d",
          1843 => x"38800b82",
          1844 => x"b5b408ec",
          1845 => x"050c8198",
          1846 => x"3982b5b4",
          1847 => x"08f80533",
          1848 => x"82b5b408",
          1849 => x"f4053354",
          1850 => x"54727426",
          1851 => x"8d38800b",
          1852 => x"82b5b408",
          1853 => x"ec050c80",
          1854 => x"f73982b5",
          1855 => x"b408f405",
          1856 => x"337082b5",
          1857 => x"b408fc05",
          1858 => x"082982b5",
          1859 => x"b408f805",
          1860 => x"33701282",
          1861 => x"b5b408fc",
          1862 => x"050c82b5",
          1863 => x"b4088805",
          1864 => x"08700881",
          1865 => x"05710c70",
          1866 => x"08515152",
          1867 => x"55537233",
          1868 => x"82b5b408",
          1869 => x"f80534fe",
          1870 => x"a53982b5",
          1871 => x"b408f005",
          1872 => x"33537280",
          1873 => x"2e903882",
          1874 => x"b5b408fc",
          1875 => x"05083082",
          1876 => x"b5b408fc",
          1877 => x"050c82b5",
          1878 => x"b4088c05",
          1879 => x"0882b5b4",
          1880 => x"08fc0508",
          1881 => x"710c5381",
          1882 => x"0b82b5b4",
          1883 => x"08ec050c",
          1884 => x"82b5b408",
          1885 => x"ec050882",
          1886 => x"b5a80c8b",
          1887 => x"3d0d82b5",
          1888 => x"b40c0482",
          1889 => x"b5b40802",
          1890 => x"82b5b40c",
          1891 => x"fb3d0d80",
          1892 => x"0b82b5b4",
          1893 => x"08f8050c",
          1894 => x"82ccfc08",
          1895 => x"85113370",
          1896 => x"812a7081",
          1897 => x"32708106",
          1898 => x"51515151",
          1899 => x"5372802e",
          1900 => x"8d38ff0b",
          1901 => x"82b5b408",
          1902 => x"f4050c81",
          1903 => x"923982b5",
          1904 => x"b4088805",
          1905 => x"08537233",
          1906 => x"82b5b408",
          1907 => x"88050881",
          1908 => x"0582b5b4",
          1909 => x"0888050c",
          1910 => x"537282b5",
          1911 => x"b408fc05",
          1912 => x"347281ff",
          1913 => x"06537280",
          1914 => x"2eb03882",
          1915 => x"ccfc0882",
          1916 => x"ccfc0853",
          1917 => x"82b5b408",
          1918 => x"fc053352",
          1919 => x"90110851",
          1920 => x"53722d82",
          1921 => x"b5a80853",
          1922 => x"72802eff",
          1923 => x"b138ff0b",
          1924 => x"82b5b408",
          1925 => x"f8050cff",
          1926 => x"a53982cc",
          1927 => x"fc0882cc",
          1928 => x"fc085353",
          1929 => x"8a519013",
          1930 => x"0853722d",
          1931 => x"82b5a808",
          1932 => x"5372802e",
          1933 => x"8a38ff0b",
          1934 => x"82b5b408",
          1935 => x"f8050c82",
          1936 => x"b5b408f8",
          1937 => x"05087082",
          1938 => x"b5b408f4",
          1939 => x"050c5382",
          1940 => x"b5b408f4",
          1941 => x"050882b5",
          1942 => x"a80c873d",
          1943 => x"0d82b5b4",
          1944 => x"0c0482b5",
          1945 => x"b4080282",
          1946 => x"b5b40cfb",
          1947 => x"3d0d800b",
          1948 => x"82b5b408",
          1949 => x"f8050c82",
          1950 => x"b5b4088c",
          1951 => x"05088511",
          1952 => x"3370812a",
          1953 => x"70813270",
          1954 => x"81065151",
          1955 => x"51515372",
          1956 => x"802e8d38",
          1957 => x"ff0b82b5",
          1958 => x"b408f405",
          1959 => x"0c80f339",
          1960 => x"82b5b408",
          1961 => x"88050853",
          1962 => x"723382b5",
          1963 => x"b4088805",
          1964 => x"08810582",
          1965 => x"b5b40888",
          1966 => x"050c5372",
          1967 => x"82b5b408",
          1968 => x"fc053472",
          1969 => x"81ff0653",
          1970 => x"72802eb6",
          1971 => x"3882b5b4",
          1972 => x"088c0508",
          1973 => x"82b5b408",
          1974 => x"8c050853",
          1975 => x"82b5b408",
          1976 => x"fc053352",
          1977 => x"90110851",
          1978 => x"53722d82",
          1979 => x"b5a80853",
          1980 => x"72802eff",
          1981 => x"ab38ff0b",
          1982 => x"82b5b408",
          1983 => x"f8050cff",
          1984 => x"9f3982b5",
          1985 => x"b408f805",
          1986 => x"087082b5",
          1987 => x"b408f405",
          1988 => x"0c5382b5",
          1989 => x"b408f405",
          1990 => x"0882b5a8",
          1991 => x"0c873d0d",
          1992 => x"82b5b40c",
          1993 => x"0482b5b4",
          1994 => x"080282b5",
          1995 => x"b40cfe3d",
          1996 => x"0d82ccfc",
          1997 => x"085282b5",
          1998 => x"b4088805",
          1999 => x"0851933f",
          2000 => x"82b5a808",
          2001 => x"7082b5a8",
          2002 => x"0c53843d",
          2003 => x"0d82b5b4",
          2004 => x"0c0482b5",
          2005 => x"b4080282",
          2006 => x"b5b40cfb",
          2007 => x"3d0d82b5",
          2008 => x"b4088c05",
          2009 => x"08851133",
          2010 => x"70812a70",
          2011 => x"81327081",
          2012 => x"06515151",
          2013 => x"51537280",
          2014 => x"2e8d38ff",
          2015 => x"0b82b5b4",
          2016 => x"08fc050c",
          2017 => x"81cb3982",
          2018 => x"b5b4088c",
          2019 => x"05088511",
          2020 => x"3370822a",
          2021 => x"70810651",
          2022 => x"51515372",
          2023 => x"802e80db",
          2024 => x"3882b5b4",
          2025 => x"088c0508",
          2026 => x"82b5b408",
          2027 => x"8c050854",
          2028 => x"548c1408",
          2029 => x"88140825",
          2030 => x"9f3882b5",
          2031 => x"b4088c05",
          2032 => x"08700870",
          2033 => x"82b5b408",
          2034 => x"88050852",
          2035 => x"57545472",
          2036 => x"75347308",
          2037 => x"8105740c",
          2038 => x"82b5b408",
          2039 => x"8c05088c",
          2040 => x"11088105",
          2041 => x"8c120c82",
          2042 => x"b5b40888",
          2043 => x"05087082",
          2044 => x"b5b408fc",
          2045 => x"050c5153",
          2046 => x"80d73982",
          2047 => x"b5b4088c",
          2048 => x"050882b5",
          2049 => x"b4088c05",
          2050 => x"085382b5",
          2051 => x"b4088805",
          2052 => x"087081ff",
          2053 => x"06539012",
          2054 => x"08515454",
          2055 => x"722d82b5",
          2056 => x"a8085372",
          2057 => x"a33882b5",
          2058 => x"b4088c05",
          2059 => x"088c1108",
          2060 => x"81058c12",
          2061 => x"0c82b5b4",
          2062 => x"08880508",
          2063 => x"7082b5b4",
          2064 => x"08fc050c",
          2065 => x"51538a39",
          2066 => x"ff0b82b5",
          2067 => x"b408fc05",
          2068 => x"0c82b5b4",
          2069 => x"08fc0508",
          2070 => x"82b5a80c",
          2071 => x"873d0d82",
          2072 => x"b5b40c04",
          2073 => x"82b5b408",
          2074 => x"0282b5b4",
          2075 => x"0cf93d0d",
          2076 => x"82b5b408",
          2077 => x"88050885",
          2078 => x"11337081",
          2079 => x"32708106",
          2080 => x"51515152",
          2081 => x"71802e8d",
          2082 => x"38ff0b82",
          2083 => x"b5b408f8",
          2084 => x"050c8394",
          2085 => x"3982b5b4",
          2086 => x"08880508",
          2087 => x"85113370",
          2088 => x"862a7081",
          2089 => x"06515151",
          2090 => x"5271802e",
          2091 => x"80c53882",
          2092 => x"b5b40888",
          2093 => x"050882b5",
          2094 => x"b4088805",
          2095 => x"08535385",
          2096 => x"123370ff",
          2097 => x"bf065152",
          2098 => x"71851434",
          2099 => x"82b5b408",
          2100 => x"8805088c",
          2101 => x"11088105",
          2102 => x"8c120c82",
          2103 => x"b5b40888",
          2104 => x"05088411",
          2105 => x"337082b5",
          2106 => x"b408f805",
          2107 => x"0c515152",
          2108 => x"82b63982",
          2109 => x"b5b40888",
          2110 => x"05088511",
          2111 => x"3370822a",
          2112 => x"70810651",
          2113 => x"51515271",
          2114 => x"802e80d7",
          2115 => x"3882b5b4",
          2116 => x"08880508",
          2117 => x"70087033",
          2118 => x"82b5b408",
          2119 => x"fc050c51",
          2120 => x"5282b5b4",
          2121 => x"08fc0508",
          2122 => x"a93882b5",
          2123 => x"b4088805",
          2124 => x"0882b5b4",
          2125 => x"08880508",
          2126 => x"53538512",
          2127 => x"3370a007",
          2128 => x"51527185",
          2129 => x"1434ff0b",
          2130 => x"82b5b408",
          2131 => x"f8050c81",
          2132 => x"d73982b5",
          2133 => x"b4088805",
          2134 => x"08700881",
          2135 => x"05710c52",
          2136 => x"81a13982",
          2137 => x"b5b40888",
          2138 => x"050882b5",
          2139 => x"b4088805",
          2140 => x"08529411",
          2141 => x"08515271",
          2142 => x"2d82b5a8",
          2143 => x"087082b5",
          2144 => x"b408fc05",
          2145 => x"0c5282b5",
          2146 => x"b408fc05",
          2147 => x"08802580",
          2148 => x"f23882b5",
          2149 => x"b4088805",
          2150 => x"0882b5b4",
          2151 => x"08f4050c",
          2152 => x"82b5b408",
          2153 => x"88050885",
          2154 => x"113382b5",
          2155 => x"b408f005",
          2156 => x"0c5282b5",
          2157 => x"b408fc05",
          2158 => x"08ff2e09",
          2159 => x"81069538",
          2160 => x"82b5b408",
          2161 => x"f0050890",
          2162 => x"07527182",
          2163 => x"b5b408ec",
          2164 => x"05349339",
          2165 => x"82b5b408",
          2166 => x"f00508a0",
          2167 => x"07527182",
          2168 => x"b5b408ec",
          2169 => x"053482b5",
          2170 => x"b408f405",
          2171 => x"085282b5",
          2172 => x"b408ec05",
          2173 => x"33851334",
          2174 => x"ff0b82b5",
          2175 => x"b408f805",
          2176 => x"0ca63982",
          2177 => x"b5b40888",
          2178 => x"05088c11",
          2179 => x"0881058c",
          2180 => x"120c82b5",
          2181 => x"b408fc05",
          2182 => x"087081ff",
          2183 => x"067082b5",
          2184 => x"b408f805",
          2185 => x"0c515152",
          2186 => x"82b5b408",
          2187 => x"f8050882",
          2188 => x"b5a80c89",
          2189 => x"3d0d82b5",
          2190 => x"b40c0482",
          2191 => x"b5b40802",
          2192 => x"82b5b40c",
          2193 => x"fd3d0d82",
          2194 => x"b5b40888",
          2195 => x"050882b5",
          2196 => x"b408fc05",
          2197 => x"0c82b5b4",
          2198 => x"088c0508",
          2199 => x"82b5b408",
          2200 => x"f8050c82",
          2201 => x"b5b40890",
          2202 => x"0508802e",
          2203 => x"82a23882",
          2204 => x"b5b408f8",
          2205 => x"050882b5",
          2206 => x"b408fc05",
          2207 => x"082681ac",
          2208 => x"3882b5b4",
          2209 => x"08f80508",
          2210 => x"82b5b408",
          2211 => x"90050805",
          2212 => x"5182b5b4",
          2213 => x"08fc0508",
          2214 => x"71278190",
          2215 => x"3882b5b4",
          2216 => x"08fc0508",
          2217 => x"82b5b408",
          2218 => x"90050805",
          2219 => x"82b5b408",
          2220 => x"fc050c82",
          2221 => x"b5b408f8",
          2222 => x"050882b5",
          2223 => x"b4089005",
          2224 => x"080582b5",
          2225 => x"b408f805",
          2226 => x"0c82b5b4",
          2227 => x"08900508",
          2228 => x"810582b5",
          2229 => x"b4089005",
          2230 => x"0c82b5b4",
          2231 => x"08900508",
          2232 => x"ff0582b5",
          2233 => x"b4089005",
          2234 => x"0c82b5b4",
          2235 => x"08900508",
          2236 => x"802e819c",
          2237 => x"3882b5b4",
          2238 => x"08fc0508",
          2239 => x"ff0582b5",
          2240 => x"b408fc05",
          2241 => x"0c82b5b4",
          2242 => x"08f80508",
          2243 => x"ff0582b5",
          2244 => x"b408f805",
          2245 => x"0c82b5b4",
          2246 => x"08fc0508",
          2247 => x"82b5b408",
          2248 => x"f8050853",
          2249 => x"51713371",
          2250 => x"34ffae39",
          2251 => x"82b5b408",
          2252 => x"90050881",
          2253 => x"0582b5b4",
          2254 => x"0890050c",
          2255 => x"82b5b408",
          2256 => x"900508ff",
          2257 => x"0582b5b4",
          2258 => x"0890050c",
          2259 => x"82b5b408",
          2260 => x"90050880",
          2261 => x"2eba3882",
          2262 => x"b5b408f8",
          2263 => x"05085170",
          2264 => x"3382b5b4",
          2265 => x"08f80508",
          2266 => x"810582b5",
          2267 => x"b408f805",
          2268 => x"0c82b5b4",
          2269 => x"08fc0508",
          2270 => x"52527171",
          2271 => x"3482b5b4",
          2272 => x"08fc0508",
          2273 => x"810582b5",
          2274 => x"b408fc05",
          2275 => x"0cffad39",
          2276 => x"82b5b408",
          2277 => x"88050870",
          2278 => x"82b5a80c",
          2279 => x"51853d0d",
          2280 => x"82b5b40c",
          2281 => x"0482b5b4",
          2282 => x"080282b5",
          2283 => x"b40cfe3d",
          2284 => x"0d82b5b4",
          2285 => x"08880508",
          2286 => x"82b5b408",
          2287 => x"fc050c82",
          2288 => x"b5b408fc",
          2289 => x"05085271",
          2290 => x"3382b5b4",
          2291 => x"08fc0508",
          2292 => x"810582b5",
          2293 => x"b408fc05",
          2294 => x"0c7081ff",
          2295 => x"06515170",
          2296 => x"802e8338",
          2297 => x"da3982b5",
          2298 => x"b408fc05",
          2299 => x"08ff0582",
          2300 => x"b5b408fc",
          2301 => x"050c82b5",
          2302 => x"b408fc05",
          2303 => x"0882b5b4",
          2304 => x"08880508",
          2305 => x"317082b5",
          2306 => x"a80c5184",
          2307 => x"3d0d82b5",
          2308 => x"b40c0482",
          2309 => x"b5b40802",
          2310 => x"82b5b40c",
          2311 => x"fe3d0d82",
          2312 => x"b5b40888",
          2313 => x"050882b5",
          2314 => x"b408fc05",
          2315 => x"0c82b5b4",
          2316 => x"088c0508",
          2317 => x"52713382",
          2318 => x"b5b4088c",
          2319 => x"05088105",
          2320 => x"82b5b408",
          2321 => x"8c050c82",
          2322 => x"b5b408fc",
          2323 => x"05085351",
          2324 => x"70723482",
          2325 => x"b5b408fc",
          2326 => x"05088105",
          2327 => x"82b5b408",
          2328 => x"fc050c70",
          2329 => x"81ff0651",
          2330 => x"70802e84",
          2331 => x"38ffbe39",
          2332 => x"82b5b408",
          2333 => x"88050870",
          2334 => x"82b5a80c",
          2335 => x"51843d0d",
          2336 => x"82b5b40c",
          2337 => x"0482b5b4",
          2338 => x"080282b5",
          2339 => x"b40cfd3d",
          2340 => x"0d82b5b4",
          2341 => x"08880508",
          2342 => x"82b5b408",
          2343 => x"fc050c82",
          2344 => x"b5b4088c",
          2345 => x"050882b5",
          2346 => x"b408f805",
          2347 => x"0c82b5b4",
          2348 => x"08900508",
          2349 => x"802e80e5",
          2350 => x"3882b5b4",
          2351 => x"08900508",
          2352 => x"810582b5",
          2353 => x"b4089005",
          2354 => x"0c82b5b4",
          2355 => x"08900508",
          2356 => x"ff0582b5",
          2357 => x"b4089005",
          2358 => x"0c82b5b4",
          2359 => x"08900508",
          2360 => x"802eba38",
          2361 => x"82b5b408",
          2362 => x"f8050851",
          2363 => x"703382b5",
          2364 => x"b408f805",
          2365 => x"08810582",
          2366 => x"b5b408f8",
          2367 => x"050c82b5",
          2368 => x"b408fc05",
          2369 => x"08525271",
          2370 => x"713482b5",
          2371 => x"b408fc05",
          2372 => x"08810582",
          2373 => x"b5b408fc",
          2374 => x"050cffad",
          2375 => x"3982b5b4",
          2376 => x"08880508",
          2377 => x"7082b5a8",
          2378 => x"0c51853d",
          2379 => x"0d82b5b4",
          2380 => x"0c0482b5",
          2381 => x"b4080282",
          2382 => x"b5b40cfd",
          2383 => x"3d0d82b5",
          2384 => x"b4089005",
          2385 => x"08802e81",
          2386 => x"f43882b5",
          2387 => x"b4088c05",
          2388 => x"08527133",
          2389 => x"82b5b408",
          2390 => x"8c050881",
          2391 => x"0582b5b4",
          2392 => x"088c050c",
          2393 => x"82b5b408",
          2394 => x"88050870",
          2395 => x"337281ff",
          2396 => x"06535454",
          2397 => x"5171712e",
          2398 => x"843880ce",
          2399 => x"3982b5b4",
          2400 => x"08880508",
          2401 => x"52713382",
          2402 => x"b5b40888",
          2403 => x"05088105",
          2404 => x"82b5b408",
          2405 => x"88050c70",
          2406 => x"81ff0651",
          2407 => x"51708d38",
          2408 => x"800b82b5",
          2409 => x"b408fc05",
          2410 => x"0c819b39",
          2411 => x"82b5b408",
          2412 => x"900508ff",
          2413 => x"0582b5b4",
          2414 => x"0890050c",
          2415 => x"82b5b408",
          2416 => x"90050880",
          2417 => x"2e8438ff",
          2418 => x"813982b5",
          2419 => x"b4089005",
          2420 => x"08802e80",
          2421 => x"e83882b5",
          2422 => x"b4088805",
          2423 => x"08703352",
          2424 => x"53708d38",
          2425 => x"ff0b82b5",
          2426 => x"b408fc05",
          2427 => x"0c80d739",
          2428 => x"82b5b408",
          2429 => x"8c0508ff",
          2430 => x"0582b5b4",
          2431 => x"088c050c",
          2432 => x"82b5b408",
          2433 => x"8c050870",
          2434 => x"33525270",
          2435 => x"8c38810b",
          2436 => x"82b5b408",
          2437 => x"fc050cae",
          2438 => x"3982b5b4",
          2439 => x"08880508",
          2440 => x"703382b5",
          2441 => x"b4088c05",
          2442 => x"08703372",
          2443 => x"71317082",
          2444 => x"b5b408fc",
          2445 => x"050c5355",
          2446 => x"5252538a",
          2447 => x"39800b82",
          2448 => x"b5b408fc",
          2449 => x"050c82b5",
          2450 => x"b408fc05",
          2451 => x"0882b5a8",
          2452 => x"0c853d0d",
          2453 => x"82b5b40c",
          2454 => x"0482b5b4",
          2455 => x"080282b5",
          2456 => x"b40cfd3d",
          2457 => x"0d82b5b4",
          2458 => x"08880508",
          2459 => x"82b5b408",
          2460 => x"f8050c82",
          2461 => x"b5b4088c",
          2462 => x"05088d38",
          2463 => x"800b82b5",
          2464 => x"b408fc05",
          2465 => x"0c80ec39",
          2466 => x"82b5b408",
          2467 => x"f8050852",
          2468 => x"713382b5",
          2469 => x"b408f805",
          2470 => x"08810582",
          2471 => x"b5b408f8",
          2472 => x"050c7081",
          2473 => x"ff065151",
          2474 => x"70802e9f",
          2475 => x"3882b5b4",
          2476 => x"088c0508",
          2477 => x"ff0582b5",
          2478 => x"b4088c05",
          2479 => x"0c82b5b4",
          2480 => x"088c0508",
          2481 => x"ff2e8438",
          2482 => x"ffbe3982",
          2483 => x"b5b408f8",
          2484 => x"0508ff05",
          2485 => x"82b5b408",
          2486 => x"f8050c82",
          2487 => x"b5b408f8",
          2488 => x"050882b5",
          2489 => x"b4088805",
          2490 => x"08317082",
          2491 => x"b5b408fc",
          2492 => x"050c5182",
          2493 => x"b5b408fc",
          2494 => x"050882b5",
          2495 => x"a80c853d",
          2496 => x"0d82b5b4",
          2497 => x"0c0482b5",
          2498 => x"b4080282",
          2499 => x"b5b40cfe",
          2500 => x"3d0d82b5",
          2501 => x"b4088805",
          2502 => x"0882b5b4",
          2503 => x"08fc050c",
          2504 => x"82b5b408",
          2505 => x"90050880",
          2506 => x"2e80d438",
          2507 => x"82b5b408",
          2508 => x"90050881",
          2509 => x"0582b5b4",
          2510 => x"0890050c",
          2511 => x"82b5b408",
          2512 => x"900508ff",
          2513 => x"0582b5b4",
          2514 => x"0890050c",
          2515 => x"82b5b408",
          2516 => x"90050880",
          2517 => x"2ea93882",
          2518 => x"b5b4088c",
          2519 => x"05085170",
          2520 => x"82b5b408",
          2521 => x"fc050852",
          2522 => x"52717134",
          2523 => x"82b5b408",
          2524 => x"fc050881",
          2525 => x"0582b5b4",
          2526 => x"08fc050c",
          2527 => x"ffbe3982",
          2528 => x"b5b40888",
          2529 => x"05087082",
          2530 => x"b5a80c51",
          2531 => x"843d0d82",
          2532 => x"b5b40c04",
          2533 => x"82b5b408",
          2534 => x"0282b5b4",
          2535 => x"0cf93d0d",
          2536 => x"800b82b5",
          2537 => x"b408fc05",
          2538 => x"0c82b5b4",
          2539 => x"08880508",
          2540 => x"8025b938",
          2541 => x"82b5b408",
          2542 => x"88050830",
          2543 => x"82b5b408",
          2544 => x"88050c80",
          2545 => x"0b82b5b4",
          2546 => x"08f4050c",
          2547 => x"82b5b408",
          2548 => x"fc05088a",
          2549 => x"38810b82",
          2550 => x"b5b408f4",
          2551 => x"050c82b5",
          2552 => x"b408f405",
          2553 => x"0882b5b4",
          2554 => x"08fc050c",
          2555 => x"82b5b408",
          2556 => x"8c050880",
          2557 => x"25b93882",
          2558 => x"b5b4088c",
          2559 => x"05083082",
          2560 => x"b5b4088c",
          2561 => x"050c800b",
          2562 => x"82b5b408",
          2563 => x"f0050c82",
          2564 => x"b5b408fc",
          2565 => x"05088a38",
          2566 => x"810b82b5",
          2567 => x"b408f005",
          2568 => x"0c82b5b4",
          2569 => x"08f00508",
          2570 => x"82b5b408",
          2571 => x"fc050c80",
          2572 => x"5382b5b4",
          2573 => x"088c0508",
          2574 => x"5282b5b4",
          2575 => x"08880508",
          2576 => x"5182c53f",
          2577 => x"82b5a808",
          2578 => x"7082b5b4",
          2579 => x"08f8050c",
          2580 => x"5482b5b4",
          2581 => x"08fc0508",
          2582 => x"802e9038",
          2583 => x"82b5b408",
          2584 => x"f8050830",
          2585 => x"82b5b408",
          2586 => x"f8050c82",
          2587 => x"b5b408f8",
          2588 => x"05087082",
          2589 => x"b5a80c54",
          2590 => x"893d0d82",
          2591 => x"b5b40c04",
          2592 => x"82b5b408",
          2593 => x"0282b5b4",
          2594 => x"0cfb3d0d",
          2595 => x"800b82b5",
          2596 => x"b408fc05",
          2597 => x"0c82b5b4",
          2598 => x"08880508",
          2599 => x"80259938",
          2600 => x"82b5b408",
          2601 => x"88050830",
          2602 => x"82b5b408",
          2603 => x"88050c81",
          2604 => x"0b82b5b4",
          2605 => x"08fc050c",
          2606 => x"82b5b408",
          2607 => x"8c050880",
          2608 => x"25903882",
          2609 => x"b5b4088c",
          2610 => x"05083082",
          2611 => x"b5b4088c",
          2612 => x"050c8153",
          2613 => x"82b5b408",
          2614 => x"8c050852",
          2615 => x"82b5b408",
          2616 => x"88050851",
          2617 => x"81a23f82",
          2618 => x"b5a80870",
          2619 => x"82b5b408",
          2620 => x"f8050c54",
          2621 => x"82b5b408",
          2622 => x"fc050880",
          2623 => x"2e903882",
          2624 => x"b5b408f8",
          2625 => x"05083082",
          2626 => x"b5b408f8",
          2627 => x"050c82b5",
          2628 => x"b408f805",
          2629 => x"087082b5",
          2630 => x"a80c5487",
          2631 => x"3d0d82b5",
          2632 => x"b40c0482",
          2633 => x"b5b40802",
          2634 => x"82b5b40c",
          2635 => x"fd3d0d80",
          2636 => x"5382b5b4",
          2637 => x"088c0508",
          2638 => x"5282b5b4",
          2639 => x"08880508",
          2640 => x"5180c53f",
          2641 => x"82b5a808",
          2642 => x"7082b5a8",
          2643 => x"0c54853d",
          2644 => x"0d82b5b4",
          2645 => x"0c0482b5",
          2646 => x"b4080282",
          2647 => x"b5b40cfd",
          2648 => x"3d0d8153",
          2649 => x"82b5b408",
          2650 => x"8c050852",
          2651 => x"82b5b408",
          2652 => x"88050851",
          2653 => x"933f82b5",
          2654 => x"a8087082",
          2655 => x"b5a80c54",
          2656 => x"853d0d82",
          2657 => x"b5b40c04",
          2658 => x"82b5b408",
          2659 => x"0282b5b4",
          2660 => x"0cfd3d0d",
          2661 => x"810b82b5",
          2662 => x"b408fc05",
          2663 => x"0c800b82",
          2664 => x"b5b408f8",
          2665 => x"050c82b5",
          2666 => x"b4088c05",
          2667 => x"0882b5b4",
          2668 => x"08880508",
          2669 => x"27b93882",
          2670 => x"b5b408fc",
          2671 => x"0508802e",
          2672 => x"ae38800b",
          2673 => x"82b5b408",
          2674 => x"8c050824",
          2675 => x"a23882b5",
          2676 => x"b4088c05",
          2677 => x"081082b5",
          2678 => x"b4088c05",
          2679 => x"0c82b5b4",
          2680 => x"08fc0508",
          2681 => x"1082b5b4",
          2682 => x"08fc050c",
          2683 => x"ffb83982",
          2684 => x"b5b408fc",
          2685 => x"0508802e",
          2686 => x"80e13882",
          2687 => x"b5b4088c",
          2688 => x"050882b5",
          2689 => x"b4088805",
          2690 => x"0826ad38",
          2691 => x"82b5b408",
          2692 => x"88050882",
          2693 => x"b5b4088c",
          2694 => x"05083182",
          2695 => x"b5b40888",
          2696 => x"050c82b5",
          2697 => x"b408f805",
          2698 => x"0882b5b4",
          2699 => x"08fc0508",
          2700 => x"0782b5b4",
          2701 => x"08f8050c",
          2702 => x"82b5b408",
          2703 => x"fc050881",
          2704 => x"2a82b5b4",
          2705 => x"08fc050c",
          2706 => x"82b5b408",
          2707 => x"8c050881",
          2708 => x"2a82b5b4",
          2709 => x"088c050c",
          2710 => x"ff953982",
          2711 => x"b5b40890",
          2712 => x"0508802e",
          2713 => x"933882b5",
          2714 => x"b4088805",
          2715 => x"087082b5",
          2716 => x"b408f405",
          2717 => x"0c519139",
          2718 => x"82b5b408",
          2719 => x"f8050870",
          2720 => x"82b5b408",
          2721 => x"f4050c51",
          2722 => x"82b5b408",
          2723 => x"f4050882",
          2724 => x"b5a80c85",
          2725 => x"3d0d82b5",
          2726 => x"b40c04f9",
          2727 => x"3d0d7970",
          2728 => x"08705656",
          2729 => x"5874802e",
          2730 => x"80e33895",
          2731 => x"39750851",
          2732 => x"f1f33f82",
          2733 => x"b5a80815",
          2734 => x"780c8516",
          2735 => x"335480cd",
          2736 => x"39743354",
          2737 => x"73a02e09",
          2738 => x"81068638",
          2739 => x"811555f1",
          2740 => x"39805776",
          2741 => x"902982b0",
          2742 => x"a8057008",
          2743 => x"5256f1c5",
          2744 => x"3f82b5a8",
          2745 => x"08537452",
          2746 => x"750851f4",
          2747 => x"c53f82b5",
          2748 => x"a8088b38",
          2749 => x"84163354",
          2750 => x"73812eff",
          2751 => x"b0388117",
          2752 => x"7081ff06",
          2753 => x"58549977",
          2754 => x"27c938ff",
          2755 => x"547382b5",
          2756 => x"a80c893d",
          2757 => x"0d04ff3d",
          2758 => x"0d735271",
          2759 => x"9326818e",
          2760 => x"38718429",
          2761 => x"8294c005",
          2762 => x"52710804",
          2763 => x"829a8c51",
          2764 => x"81803982",
          2765 => x"9a985180",
          2766 => x"f939829a",
          2767 => x"ac5180f2",
          2768 => x"39829ac0",
          2769 => x"5180eb39",
          2770 => x"829ad051",
          2771 => x"80e43982",
          2772 => x"9ae05180",
          2773 => x"dd39829a",
          2774 => x"f45180d6",
          2775 => x"39829b84",
          2776 => x"5180cf39",
          2777 => x"829b9c51",
          2778 => x"80c83982",
          2779 => x"9bb45180",
          2780 => x"c139829b",
          2781 => x"cc51bb39",
          2782 => x"829be851",
          2783 => x"b539829b",
          2784 => x"fc51af39",
          2785 => x"829ca851",
          2786 => x"a939829c",
          2787 => x"bc51a339",
          2788 => x"829cdc51",
          2789 => x"9d39829c",
          2790 => x"f0519739",
          2791 => x"829d8851",
          2792 => x"9139829d",
          2793 => x"a0518b39",
          2794 => x"829db851",
          2795 => x"8539829d",
          2796 => x"c451e3cf",
          2797 => x"3f833d0d",
          2798 => x"04fb3d0d",
          2799 => x"77795656",
          2800 => x"7487e726",
          2801 => x"8a387452",
          2802 => x"7587e829",
          2803 => x"51903987",
          2804 => x"e8527451",
          2805 => x"facd3f82",
          2806 => x"b5a80852",
          2807 => x"7551fac3",
          2808 => x"3f82b5a8",
          2809 => x"08547953",
          2810 => x"7552829d",
          2811 => x"d451ffbb",
          2812 => x"e53f873d",
          2813 => x"0d04ec3d",
          2814 => x"0d660284",
          2815 => x"0580e305",
          2816 => x"335b5780",
          2817 => x"68783070",
          2818 => x"7a077325",
          2819 => x"51575959",
          2820 => x"78567787",
          2821 => x"ff268338",
          2822 => x"81567476",
          2823 => x"077081ff",
          2824 => x"06515593",
          2825 => x"56748182",
          2826 => x"38815376",
          2827 => x"528c3d70",
          2828 => x"525680fe",
          2829 => x"dc3f82b5",
          2830 => x"a8085782",
          2831 => x"b5a808b9",
          2832 => x"3882b5a8",
          2833 => x"0887c098",
          2834 => x"880c82b5",
          2835 => x"a8085996",
          2836 => x"3dd40554",
          2837 => x"84805377",
          2838 => x"52755181",
          2839 => x"83983f82",
          2840 => x"b5a80857",
          2841 => x"82b5a808",
          2842 => x"90387a55",
          2843 => x"74802e89",
          2844 => x"38741975",
          2845 => x"195959d7",
          2846 => x"39963dd8",
          2847 => x"0551818b",
          2848 => x"813f7630",
          2849 => x"70780780",
          2850 => x"257b3070",
          2851 => x"9f2a7206",
          2852 => x"51575156",
          2853 => x"74802e90",
          2854 => x"38829df8",
          2855 => x"5387c098",
          2856 => x"88085278",
          2857 => x"51fe923f",
          2858 => x"76567582",
          2859 => x"b5a80c96",
          2860 => x"3d0d04f8",
          2861 => x"3d0d7c02",
          2862 => x"8405b705",
          2863 => x"335859ff",
          2864 => x"5880537b",
          2865 => x"527a51fe",
          2866 => x"ad3f82b5",
          2867 => x"a808a638",
          2868 => x"76802e88",
          2869 => x"3876812e",
          2870 => x"9a389a39",
          2871 => x"62566155",
          2872 => x"605482b5",
          2873 => x"a8537f52",
          2874 => x"7e51782d",
          2875 => x"82b5a808",
          2876 => x"58833978",
          2877 => x"047782b5",
          2878 => x"a80c8a3d",
          2879 => x"0d04f33d",
          2880 => x"0d7f6163",
          2881 => x"028c0580",
          2882 => x"cf053373",
          2883 => x"73156841",
          2884 => x"5f5c5c5e",
          2885 => x"5e5e7a52",
          2886 => x"829e8051",
          2887 => x"ffb9b73f",
          2888 => x"829e8851",
          2889 => x"e0dd3f80",
          2890 => x"55747927",
          2891 => x"80fd387b",
          2892 => x"902e8938",
          2893 => x"7ba02ea6",
          2894 => x"3880c439",
          2895 => x"74185372",
          2896 => x"7a278e38",
          2897 => x"72225282",
          2898 => x"9e8c51ff",
          2899 => x"b9883f88",
          2900 => x"39829e98",
          2901 => x"51e0ac3f",
          2902 => x"82155580",
          2903 => x"c1397418",
          2904 => x"53727a27",
          2905 => x"8e387208",
          2906 => x"52829e80",
          2907 => x"51ffb8e6",
          2908 => x"3f883982",
          2909 => x"9e9451e0",
          2910 => x"8a3f8415",
          2911 => x"55a03974",
          2912 => x"1853727a",
          2913 => x"278e3872",
          2914 => x"3352829e",
          2915 => x"a051ffb8",
          2916 => x"c53f8839",
          2917 => x"829ea851",
          2918 => x"dfe93f81",
          2919 => x"155582cc",
          2920 => x"fc0852a0",
          2921 => x"51e3ab3f",
          2922 => x"feff3982",
          2923 => x"9eac51df",
          2924 => x"d23f8055",
          2925 => x"74792780",
          2926 => x"c6387418",
          2927 => x"70335553",
          2928 => x"8056727a",
          2929 => x"27833881",
          2930 => x"5680539f",
          2931 => x"74278338",
          2932 => x"81537573",
          2933 => x"067081ff",
          2934 => x"06515372",
          2935 => x"802e9038",
          2936 => x"7380fe26",
          2937 => x"8a3882cc",
          2938 => x"fc085273",
          2939 => x"51883982",
          2940 => x"ccfc0852",
          2941 => x"a051e2da",
          2942 => x"3f811555",
          2943 => x"ffb63982",
          2944 => x"9eb051de",
          2945 => x"fe3f7818",
          2946 => x"791c5c58",
          2947 => x"9cc03f82",
          2948 => x"b5a80898",
          2949 => x"2b70982c",
          2950 => x"515776a0",
          2951 => x"2e098106",
          2952 => x"aa389caa",
          2953 => x"3f82b5a8",
          2954 => x"08982b70",
          2955 => x"982c70a0",
          2956 => x"32703072",
          2957 => x"9b327030",
          2958 => x"70720773",
          2959 => x"75070651",
          2960 => x"58585957",
          2961 => x"51578073",
          2962 => x"24d83876",
          2963 => x"9b2e0981",
          2964 => x"06853880",
          2965 => x"538c397c",
          2966 => x"1e537278",
          2967 => x"26fdb738",
          2968 => x"ff537282",
          2969 => x"b5a80c8f",
          2970 => x"3d0d04fc",
          2971 => x"3d0d029b",
          2972 => x"0533829e",
          2973 => x"b453829e",
          2974 => x"b85255ff",
          2975 => x"b6d83f82",
          2976 => x"b4802251",
          2977 => x"a59b3f82",
          2978 => x"9ec45482",
          2979 => x"9ed05382",
          2980 => x"b4813352",
          2981 => x"829ed851",
          2982 => x"ffb6bb3f",
          2983 => x"74802e84",
          2984 => x"38a0cd3f",
          2985 => x"863d0d04",
          2986 => x"fe3d0d87",
          2987 => x"c0968008",
          2988 => x"53a5b73f",
          2989 => x"81519883",
          2990 => x"3f829ef4",
          2991 => x"5199983f",
          2992 => x"805197f7",
          2993 => x"3f72812a",
          2994 => x"70810651",
          2995 => x"5271802e",
          2996 => x"92388151",
          2997 => x"97e53f82",
          2998 => x"9f8c5198",
          2999 => x"fa3f8051",
          3000 => x"97d93f72",
          3001 => x"822a7081",
          3002 => x"06515271",
          3003 => x"802e9238",
          3004 => x"815197c7",
          3005 => x"3f829fa0",
          3006 => x"5198dc3f",
          3007 => x"805197bb",
          3008 => x"3f72832a",
          3009 => x"70810651",
          3010 => x"5271802e",
          3011 => x"92388151",
          3012 => x"97a93f82",
          3013 => x"9fb05198",
          3014 => x"be3f8051",
          3015 => x"979d3f72",
          3016 => x"842a7081",
          3017 => x"06515271",
          3018 => x"802e9238",
          3019 => x"8151978b",
          3020 => x"3f829fc4",
          3021 => x"5198a03f",
          3022 => x"805196ff",
          3023 => x"3f72852a",
          3024 => x"70810651",
          3025 => x"5271802e",
          3026 => x"92388151",
          3027 => x"96ed3f82",
          3028 => x"9fd85198",
          3029 => x"823f8051",
          3030 => x"96e13f72",
          3031 => x"862a7081",
          3032 => x"06515271",
          3033 => x"802e9238",
          3034 => x"815196cf",
          3035 => x"3f829fec",
          3036 => x"5197e43f",
          3037 => x"805196c3",
          3038 => x"3f72872a",
          3039 => x"70810651",
          3040 => x"5271802e",
          3041 => x"92388151",
          3042 => x"96b13f82",
          3043 => x"a0805197",
          3044 => x"c63f8051",
          3045 => x"96a53f72",
          3046 => x"882a7081",
          3047 => x"06515271",
          3048 => x"802e9238",
          3049 => x"81519693",
          3050 => x"3f82a094",
          3051 => x"5197a83f",
          3052 => x"80519687",
          3053 => x"3fa3bb3f",
          3054 => x"843d0d04",
          3055 => x"fb3d0d77",
          3056 => x"028405a3",
          3057 => x"05337055",
          3058 => x"56568052",
          3059 => x"7551eeb6",
          3060 => x"3f0b0b82",
          3061 => x"b0a43354",
          3062 => x"73a93881",
          3063 => x"5382a0d4",
          3064 => x"5282cca8",
          3065 => x"5180f7a9",
          3066 => x"3f82b5a8",
          3067 => x"08307082",
          3068 => x"b5a80807",
          3069 => x"80258271",
          3070 => x"31515154",
          3071 => x"730b0b82",
          3072 => x"b0a4340b",
          3073 => x"0b82b0a4",
          3074 => x"33547381",
          3075 => x"2e098106",
          3076 => x"af3882cc",
          3077 => x"a8537452",
          3078 => x"755181b1",
          3079 => x"da3f82b5",
          3080 => x"a808802e",
          3081 => x"8b3882b5",
          3082 => x"a80851da",
          3083 => x"d63f9139",
          3084 => x"82cca851",
          3085 => x"8183cb3f",
          3086 => x"820b0b0b",
          3087 => x"82b0a434",
          3088 => x"0b0b82b0",
          3089 => x"a4335473",
          3090 => x"822e0981",
          3091 => x"068c3882",
          3092 => x"a0e45374",
          3093 => x"527551a9",
          3094 => x"a23f800b",
          3095 => x"82b5a80c",
          3096 => x"873d0d04",
          3097 => x"cd3d0d80",
          3098 => x"707182cc",
          3099 => x"a40c405e",
          3100 => x"81527d51",
          3101 => x"80c5f53f",
          3102 => x"82b5a808",
          3103 => x"81ff065a",
          3104 => x"797e2e09",
          3105 => x"8106a338",
          3106 => x"973d5a83",
          3107 => x"5382a0ec",
          3108 => x"527951e7",
          3109 => x"f03f7d53",
          3110 => x"795282b6",
          3111 => x"d45180f5",
          3112 => x"8f3f82b5",
          3113 => x"a8087e2e",
          3114 => x"883882a0",
          3115 => x"f0518d95",
          3116 => x"39817040",
          3117 => x"5e82a1a8",
          3118 => x"51d9c83f",
          3119 => x"973d7047",
          3120 => x"5b80f852",
          3121 => x"7a51fdf4",
          3122 => x"3fb53dff",
          3123 => x"840551f3",
          3124 => x"ca3f82b5",
          3125 => x"a808902b",
          3126 => x"70902c51",
          3127 => x"5a7980c2",
          3128 => x"2e879938",
          3129 => x"7980c224",
          3130 => x"b23879bd",
          3131 => x"2e81d138",
          3132 => x"79bd2490",
          3133 => x"3879802e",
          3134 => x"ffbb3879",
          3135 => x"bc2e80da",
          3136 => x"388ac039",
          3137 => x"7980c02e",
          3138 => x"83953879",
          3139 => x"80c02485",
          3140 => x"c93879bf",
          3141 => x"2e828a38",
          3142 => x"8aa93979",
          3143 => x"80f92e89",
          3144 => x"c5387980",
          3145 => x"f9249238",
          3146 => x"7980c32e",
          3147 => x"87fa3879",
          3148 => x"80f82e89",
          3149 => x"8d388a8b",
          3150 => x"39798183",
          3151 => x"2e89f238",
          3152 => x"79818324",
          3153 => x"8b387981",
          3154 => x"822e89d7",
          3155 => x"3889f439",
          3156 => x"7981852e",
          3157 => x"89e73889",
          3158 => x"ea39b53d",
          3159 => x"ff801153",
          3160 => x"ff840551",
          3161 => x"d2cc3f82",
          3162 => x"b5a80880",
          3163 => x"2efec638",
          3164 => x"b53dfefc",
          3165 => x"1153ff84",
          3166 => x"0551d2b6",
          3167 => x"3f82b5a8",
          3168 => x"08802efe",
          3169 => x"b038b53d",
          3170 => x"fef81153",
          3171 => x"ff840551",
          3172 => x"d2a03f82",
          3173 => x"b5a80886",
          3174 => x"3882b5a8",
          3175 => x"084382a1",
          3176 => x"ac51d7df",
          3177 => x"3f64645d",
          3178 => x"5b7a7c27",
          3179 => x"81ea3862",
          3180 => x"5a797b70",
          3181 => x"84055d0c",
          3182 => x"7b7b26f5",
          3183 => x"3881d939",
          3184 => x"b53dff80",
          3185 => x"1153ff84",
          3186 => x"0551d1e6",
          3187 => x"3f82b5a8",
          3188 => x"08802efd",
          3189 => x"e038b53d",
          3190 => x"fefc1153",
          3191 => x"ff840551",
          3192 => x"d1d03f82",
          3193 => x"b5a80880",
          3194 => x"2efdca38",
          3195 => x"b53dfef8",
          3196 => x"1153ff84",
          3197 => x"0551d1ba",
          3198 => x"3f82b5a8",
          3199 => x"08802efd",
          3200 => x"b43882a1",
          3201 => x"bc51d6fb",
          3202 => x"3f645b7a",
          3203 => x"64278188",
          3204 => x"38625a7a",
          3205 => x"7081055c",
          3206 => x"337a3462",
          3207 => x"810543eb",
          3208 => x"39b53dff",
          3209 => x"801153ff",
          3210 => x"840551d1",
          3211 => x"853f82b5",
          3212 => x"a808802e",
          3213 => x"fcff38b5",
          3214 => x"3dfefc11",
          3215 => x"53ff8405",
          3216 => x"51d0ef3f",
          3217 => x"82b5a808",
          3218 => x"802efce9",
          3219 => x"38b53dfe",
          3220 => x"f81153ff",
          3221 => x"840551d0",
          3222 => x"d93f82b5",
          3223 => x"a808802e",
          3224 => x"fcd33882",
          3225 => x"a1c851d6",
          3226 => x"9a3f645b",
          3227 => x"7a6427a8",
          3228 => x"38627033",
          3229 => x"7c335f5b",
          3230 => x"5c797d2e",
          3231 => x"92387955",
          3232 => x"7b547a33",
          3233 => x"537a5282",
          3234 => x"a1d851ff",
          3235 => x"aec83f81",
          3236 => x"1b638105",
          3237 => x"445bd539",
          3238 => x"82a1f051",
          3239 => x"89a739b5",
          3240 => x"3dff8011",
          3241 => x"53ff8405",
          3242 => x"51d0873f",
          3243 => x"82b5a808",
          3244 => x"80df3882",
          3245 => x"b494335a",
          3246 => x"79802e89",
          3247 => x"3882b3cc",
          3248 => x"084580cd",
          3249 => x"3982b495",
          3250 => x"335a7980",
          3251 => x"2e883882",
          3252 => x"b3d40845",
          3253 => x"bc3982b4",
          3254 => x"96335a79",
          3255 => x"802e8838",
          3256 => x"82b3dc08",
          3257 => x"45ab3982",
          3258 => x"b497335a",
          3259 => x"79802e88",
          3260 => x"3882b3e4",
          3261 => x"08459a39",
          3262 => x"82b49233",
          3263 => x"5a79802e",
          3264 => x"883882b3",
          3265 => x"ec084589",
          3266 => x"3982b3fc",
          3267 => x"08fc8005",
          3268 => x"45b53dfe",
          3269 => x"fc1153ff",
          3270 => x"840551cf",
          3271 => x"953f82b5",
          3272 => x"a80880de",
          3273 => x"3882b494",
          3274 => x"335a7980",
          3275 => x"2e893882",
          3276 => x"b3d00844",
          3277 => x"80cc3982",
          3278 => x"b495335a",
          3279 => x"79802e88",
          3280 => x"3882b3d8",
          3281 => x"0844bb39",
          3282 => x"82b49633",
          3283 => x"5a79802e",
          3284 => x"883882b3",
          3285 => x"e00844aa",
          3286 => x"3982b497",
          3287 => x"335a7980",
          3288 => x"2e883882",
          3289 => x"b3e80844",
          3290 => x"993982b4",
          3291 => x"92335a79",
          3292 => x"802e8838",
          3293 => x"82b3f008",
          3294 => x"44883982",
          3295 => x"b3fc0888",
          3296 => x"0544b53d",
          3297 => x"fef81153",
          3298 => x"ff840551",
          3299 => x"cea43f82",
          3300 => x"b5a80880",
          3301 => x"2ea73880",
          3302 => x"635d5d7b",
          3303 => x"882e8338",
          3304 => x"815d7b90",
          3305 => x"32703070",
          3306 => x"72079f2a",
          3307 => x"70600651",
          3308 => x"515b5b79",
          3309 => x"802e8838",
          3310 => x"7ba02e83",
          3311 => x"38884382",
          3312 => x"a1f451d3",
          3313 => x"be3fa055",
          3314 => x"64546253",
          3315 => x"63526451",
          3316 => x"f2ac3f82",
          3317 => x"a2845186",
          3318 => x"ec39b53d",
          3319 => x"ff801153",
          3320 => x"ff840551",
          3321 => x"cdcc3f82",
          3322 => x"b5a80880",
          3323 => x"2ef9c638",
          3324 => x"b53dfefc",
          3325 => x"1153ff84",
          3326 => x"0551cdb6",
          3327 => x"3f82b5a8",
          3328 => x"08802ea4",
          3329 => x"38645a02",
          3330 => x"80cf0533",
          3331 => x"7a346481",
          3332 => x"0545b53d",
          3333 => x"fefc1153",
          3334 => x"ff840551",
          3335 => x"cd943f82",
          3336 => x"b5a808e1",
          3337 => x"38f98e39",
          3338 => x"64703354",
          3339 => x"5282a290",
          3340 => x"51ffaba2",
          3341 => x"3f80f852",
          3342 => x"7a51ccc0",
          3343 => x"3f7a467a",
          3344 => x"335a79ae",
          3345 => x"2ef8ee38",
          3346 => x"9f7a279f",
          3347 => x"38b53dfe",
          3348 => x"fc1153ff",
          3349 => x"840551cc",
          3350 => x"d93f82b5",
          3351 => x"a808802e",
          3352 => x"9138645a",
          3353 => x"0280cf05",
          3354 => x"337a3464",
          3355 => x"810545ff",
          3356 => x"b73982a2",
          3357 => x"9c51d28b",
          3358 => x"3fffad39",
          3359 => x"b53dfef4",
          3360 => x"1153ff84",
          3361 => x"0551c6a3",
          3362 => x"3f82b5a8",
          3363 => x"08802ef8",
          3364 => x"a438b53d",
          3365 => x"fef01153",
          3366 => x"ff840551",
          3367 => x"c68d3f82",
          3368 => x"b5a80880",
          3369 => x"2ea63861",
          3370 => x"5a0280c2",
          3371 => x"05227a70",
          3372 => x"82055c23",
          3373 => x"7942b53d",
          3374 => x"fef01153",
          3375 => x"ff840551",
          3376 => x"c5e93f82",
          3377 => x"b5a808df",
          3378 => x"38f7ea39",
          3379 => x"61702254",
          3380 => x"5282a2a4",
          3381 => x"51ffa9fe",
          3382 => x"3f80f852",
          3383 => x"7a51cb9c",
          3384 => x"3f7a467a",
          3385 => x"335a79ae",
          3386 => x"2ef7ca38",
          3387 => x"799f2687",
          3388 => x"38618205",
          3389 => x"42d639b5",
          3390 => x"3dfef011",
          3391 => x"53ff8405",
          3392 => x"51c5a83f",
          3393 => x"82b5a808",
          3394 => x"802e9338",
          3395 => x"615a0280",
          3396 => x"c205227a",
          3397 => x"7082055c",
          3398 => x"237942ff",
          3399 => x"af3982a2",
          3400 => x"9c51d0df",
          3401 => x"3fffa539",
          3402 => x"b53dfef4",
          3403 => x"1153ff84",
          3404 => x"0551c4f7",
          3405 => x"3f82b5a8",
          3406 => x"08802ef6",
          3407 => x"f838b53d",
          3408 => x"fef01153",
          3409 => x"ff840551",
          3410 => x"c4e13f82",
          3411 => x"b5a80880",
          3412 => x"2ea03861",
          3413 => x"61710c5a",
          3414 => x"61840542",
          3415 => x"b53dfef0",
          3416 => x"1153ff84",
          3417 => x"0551c4c3",
          3418 => x"3f82b5a8",
          3419 => x"08e538f6",
          3420 => x"c4396170",
          3421 => x"08545282",
          3422 => x"a2b051ff",
          3423 => x"a8d83f80",
          3424 => x"f8527a51",
          3425 => x"c9f63f7a",
          3426 => x"467a335a",
          3427 => x"79ae2ef6",
          3428 => x"a4389f7a",
          3429 => x"279b38b5",
          3430 => x"3dfef011",
          3431 => x"53ff8405",
          3432 => x"51c4883f",
          3433 => x"82b5a808",
          3434 => x"802e8d38",
          3435 => x"6161710c",
          3436 => x"5a618405",
          3437 => x"42ffbb39",
          3438 => x"82a29c51",
          3439 => x"cfc53fff",
          3440 => x"b139b53d",
          3441 => x"ff801153",
          3442 => x"ff840551",
          3443 => x"c9e43f82",
          3444 => x"b5a80880",
          3445 => x"2ef5de38",
          3446 => x"645282a2",
          3447 => x"bc51ffa7",
          3448 => x"f53f645a",
          3449 => x"7904b53d",
          3450 => x"ff801153",
          3451 => x"ff840551",
          3452 => x"c9c03f82",
          3453 => x"b5a80880",
          3454 => x"2ef5ba38",
          3455 => x"645282a2",
          3456 => x"d851ffa7",
          3457 => x"d13f645a",
          3458 => x"792d82b5",
          3459 => x"a808802e",
          3460 => x"f5a33882",
          3461 => x"b5a80852",
          3462 => x"82a2f451",
          3463 => x"ffa7b73f",
          3464 => x"f5933982",
          3465 => x"a39051ce",
          3466 => x"da3fffa7",
          3467 => x"8a3ff585",
          3468 => x"3982a3ac",
          3469 => x"51cecc3f",
          3470 => x"805affa8",
          3471 => x"3991b13f",
          3472 => x"f4f3397a",
          3473 => x"467a335a",
          3474 => x"79802ef4",
          3475 => x"e8387e7e",
          3476 => x"065a7980",
          3477 => x"2e81d638",
          3478 => x"b53dff84",
          3479 => x"055183d3",
          3480 => x"3f82b5a8",
          3481 => x"085d815c",
          3482 => x"7b822eb2",
          3483 => x"387b8224",
          3484 => x"89387b81",
          3485 => x"2e8c3880",
          3486 => x"cd397b83",
          3487 => x"2eb03880",
          3488 => x"c53982a3",
          3489 => x"c0567c55",
          3490 => x"82a3c454",
          3491 => x"805382a3",
          3492 => x"c852b53d",
          3493 => x"ffb00551",
          3494 => x"ffa9a33f",
          3495 => x"bb3982a3",
          3496 => x"e852b53d",
          3497 => x"ffb00551",
          3498 => x"ffa9933f",
          3499 => x"ab397c55",
          3500 => x"82a3c454",
          3501 => x"805382a3",
          3502 => x"d852b53d",
          3503 => x"ffb00551",
          3504 => x"ffa8fb3f",
          3505 => x"93397c54",
          3506 => x"805382a3",
          3507 => x"e452b53d",
          3508 => x"ffb00551",
          3509 => x"ffa8e73f",
          3510 => x"82ccf859",
          3511 => x"82b3cc58",
          3512 => x"82b5d857",
          3513 => x"80566555",
          3514 => x"805482d0",
          3515 => x"805382d0",
          3516 => x"8052b53d",
          3517 => x"ffb00551",
          3518 => x"ebb93f82",
          3519 => x"b5a80882",
          3520 => x"b5a80809",
          3521 => x"70307072",
          3522 => x"07802551",
          3523 => x"5c5c4080",
          3524 => x"5b7b8326",
          3525 => x"8338815b",
          3526 => x"797b065a",
          3527 => x"79802e8d",
          3528 => x"38811c70",
          3529 => x"81ff065d",
          3530 => x"5a7bfebc",
          3531 => x"387e8132",
          3532 => x"7e813207",
          3533 => x"5a798a38",
          3534 => x"7fff2e09",
          3535 => x"8106f2f5",
          3536 => x"3882a3ec",
          3537 => x"51ccbc3f",
          3538 => x"f2eb39f5",
          3539 => x"3d0d800b",
          3540 => x"82b5d834",
          3541 => x"87c0948c",
          3542 => x"70085455",
          3543 => x"87848052",
          3544 => x"7251e3bf",
          3545 => x"3f82b5a8",
          3546 => x"08902b75",
          3547 => x"08555387",
          3548 => x"84805273",
          3549 => x"51e3ac3f",
          3550 => x"7282b5a8",
          3551 => x"0807750c",
          3552 => x"87c0949c",
          3553 => x"70085455",
          3554 => x"87848052",
          3555 => x"7251e393",
          3556 => x"3f82b5a8",
          3557 => x"08902b75",
          3558 => x"08555387",
          3559 => x"84805273",
          3560 => x"51e3803f",
          3561 => x"7282b5a8",
          3562 => x"0807750c",
          3563 => x"8c80830b",
          3564 => x"87c09484",
          3565 => x"0c8c8083",
          3566 => x"0b87c094",
          3567 => x"940c82a3",
          3568 => x"fc51cbbf",
          3569 => x"3f80f5d3",
          3570 => x"5a80f8bf",
          3571 => x"5b830284",
          3572 => x"05990534",
          3573 => x"805c8d3d",
          3574 => x"e40582cc",
          3575 => x"fc0c89c4",
          3576 => x"3f93873f",
          3577 => x"82a49051",
          3578 => x"cb993f82",
          3579 => x"a4a451cb",
          3580 => x"923f82a4",
          3581 => x"b051cb8b",
          3582 => x"3f80dda8",
          3583 => x"5192e63f",
          3584 => x"8151ece7",
          3585 => x"3ff0dd3f",
          3586 => x"8004fe3d",
          3587 => x"0d805283",
          3588 => x"5371882b",
          3589 => x"5287d93f",
          3590 => x"82b5a808",
          3591 => x"81ff0672",
          3592 => x"07ff1454",
          3593 => x"52728025",
          3594 => x"e8387182",
          3595 => x"b5a80c84",
          3596 => x"3d0d04fc",
          3597 => x"3d0d7670",
          3598 => x"08545580",
          3599 => x"73525472",
          3600 => x"742e818a",
          3601 => x"38723351",
          3602 => x"70a02e09",
          3603 => x"81068638",
          3604 => x"811353f1",
          3605 => x"39723351",
          3606 => x"70a22e09",
          3607 => x"81068638",
          3608 => x"81135381",
          3609 => x"54725273",
          3610 => x"812e0981",
          3611 => x"069f3884",
          3612 => x"39811252",
          3613 => x"80723352",
          3614 => x"5470a22e",
          3615 => x"83388154",
          3616 => x"70802e9d",
          3617 => x"3873ea38",
          3618 => x"98398112",
          3619 => x"52807233",
          3620 => x"525470a0",
          3621 => x"2e833881",
          3622 => x"5470802e",
          3623 => x"843873ea",
          3624 => x"38807233",
          3625 => x"525470a0",
          3626 => x"2e098106",
          3627 => x"83388154",
          3628 => x"70a23270",
          3629 => x"30708025",
          3630 => x"76075151",
          3631 => x"5170802e",
          3632 => x"88388072",
          3633 => x"70810554",
          3634 => x"3471750c",
          3635 => x"72517082",
          3636 => x"b5a80c86",
          3637 => x"3d0d04fc",
          3638 => x"3d0d7653",
          3639 => x"7208802e",
          3640 => x"9238863d",
          3641 => x"fc055272",
          3642 => x"51ffbdbf",
          3643 => x"3f82b5a8",
          3644 => x"08853880",
          3645 => x"53833974",
          3646 => x"537282b5",
          3647 => x"a80c863d",
          3648 => x"0d04fc3d",
          3649 => x"0d768211",
          3650 => x"33ff0552",
          3651 => x"53815270",
          3652 => x"8b268198",
          3653 => x"38831333",
          3654 => x"ff055182",
          3655 => x"52709e26",
          3656 => x"818a3884",
          3657 => x"13335183",
          3658 => x"52709726",
          3659 => x"80fe3885",
          3660 => x"13335184",
          3661 => x"5270bb26",
          3662 => x"80f23886",
          3663 => x"13335185",
          3664 => x"5270bb26",
          3665 => x"80e63888",
          3666 => x"13225586",
          3667 => x"527487e7",
          3668 => x"2680d938",
          3669 => x"8a132254",
          3670 => x"87527387",
          3671 => x"e72680cc",
          3672 => x"38810b87",
          3673 => x"c0989c0c",
          3674 => x"722287c0",
          3675 => x"98bc0c82",
          3676 => x"133387c0",
          3677 => x"98b80c83",
          3678 => x"133387c0",
          3679 => x"98b40c84",
          3680 => x"133387c0",
          3681 => x"98b00c85",
          3682 => x"133387c0",
          3683 => x"98ac0c86",
          3684 => x"133387c0",
          3685 => x"98a80c74",
          3686 => x"87c098a4",
          3687 => x"0c7387c0",
          3688 => x"98a00c80",
          3689 => x"0b87c098",
          3690 => x"9c0c8052",
          3691 => x"7182b5a8",
          3692 => x"0c863d0d",
          3693 => x"04f33d0d",
          3694 => x"7f5b87c0",
          3695 => x"989c5d81",
          3696 => x"7d0c87c0",
          3697 => x"98bc085e",
          3698 => x"7d7b2387",
          3699 => x"c098b808",
          3700 => x"5a79821c",
          3701 => x"3487c098",
          3702 => x"b4085a79",
          3703 => x"831c3487",
          3704 => x"c098b008",
          3705 => x"5a79841c",
          3706 => x"3487c098",
          3707 => x"ac085a79",
          3708 => x"851c3487",
          3709 => x"c098a808",
          3710 => x"5a79861c",
          3711 => x"3487c098",
          3712 => x"a4085c7b",
          3713 => x"881c2387",
          3714 => x"c098a008",
          3715 => x"5a798a1c",
          3716 => x"23807d0c",
          3717 => x"7983ffff",
          3718 => x"06597b83",
          3719 => x"ffff0658",
          3720 => x"861b3357",
          3721 => x"851b3356",
          3722 => x"841b3355",
          3723 => x"831b3354",
          3724 => x"821b3353",
          3725 => x"7d83ffff",
          3726 => x"065282a4",
          3727 => x"c851ff9f",
          3728 => x"953f8f3d",
          3729 => x"0d04fb3d",
          3730 => x"0d029f05",
          3731 => x"3382b3c8",
          3732 => x"337081ff",
          3733 => x"06585555",
          3734 => x"87c09484",
          3735 => x"5175802e",
          3736 => x"863887c0",
          3737 => x"94945170",
          3738 => x"0870962a",
          3739 => x"70810653",
          3740 => x"54527080",
          3741 => x"2e8c3871",
          3742 => x"912a7081",
          3743 => x"06515170",
          3744 => x"d7387281",
          3745 => x"32708106",
          3746 => x"51517080",
          3747 => x"2e8d3871",
          3748 => x"932a7081",
          3749 => x"06515170",
          3750 => x"ffbe3873",
          3751 => x"81ff0651",
          3752 => x"87c09480",
          3753 => x"5270802e",
          3754 => x"863887c0",
          3755 => x"94905274",
          3756 => x"720c7482",
          3757 => x"b5a80c87",
          3758 => x"3d0d04ff",
          3759 => x"3d0d028f",
          3760 => x"05337030",
          3761 => x"709f2a51",
          3762 => x"52527082",
          3763 => x"b3c83483",
          3764 => x"3d0d04f9",
          3765 => x"3d0d02a7",
          3766 => x"05335877",
          3767 => x"8a2e0981",
          3768 => x"0687387a",
          3769 => x"528d51eb",
          3770 => x"3f82b3c8",
          3771 => x"337081ff",
          3772 => x"06585687",
          3773 => x"c0948453",
          3774 => x"76802e86",
          3775 => x"3887c094",
          3776 => x"94537208",
          3777 => x"70962a70",
          3778 => x"81065556",
          3779 => x"5472802e",
          3780 => x"8c387391",
          3781 => x"2a708106",
          3782 => x"515372d7",
          3783 => x"38748132",
          3784 => x"70810651",
          3785 => x"5372802e",
          3786 => x"8d387393",
          3787 => x"2a708106",
          3788 => x"515372ff",
          3789 => x"be387581",
          3790 => x"ff065387",
          3791 => x"c0948054",
          3792 => x"72802e86",
          3793 => x"3887c094",
          3794 => x"90547774",
          3795 => x"0c800b82",
          3796 => x"b5a80c89",
          3797 => x"3d0d04f9",
          3798 => x"3d0d7954",
          3799 => x"80743370",
          3800 => x"81ff0653",
          3801 => x"53577077",
          3802 => x"2e80fc38",
          3803 => x"7181ff06",
          3804 => x"811582b3",
          3805 => x"c8337081",
          3806 => x"ff065957",
          3807 => x"555887c0",
          3808 => x"94845175",
          3809 => x"802e8638",
          3810 => x"87c09494",
          3811 => x"51700870",
          3812 => x"962a7081",
          3813 => x"06535452",
          3814 => x"70802e8c",
          3815 => x"3871912a",
          3816 => x"70810651",
          3817 => x"5170d738",
          3818 => x"72813270",
          3819 => x"81065151",
          3820 => x"70802e8d",
          3821 => x"3871932a",
          3822 => x"70810651",
          3823 => x"5170ffbe",
          3824 => x"387481ff",
          3825 => x"065187c0",
          3826 => x"94805270",
          3827 => x"802e8638",
          3828 => x"87c09490",
          3829 => x"5277720c",
          3830 => x"81177433",
          3831 => x"7081ff06",
          3832 => x"53535770",
          3833 => x"ff863876",
          3834 => x"82b5a80c",
          3835 => x"893d0d04",
          3836 => x"fe3d0d82",
          3837 => x"b3c83370",
          3838 => x"81ff0654",
          3839 => x"5287c094",
          3840 => x"84517280",
          3841 => x"2e863887",
          3842 => x"c0949451",
          3843 => x"70087082",
          3844 => x"2a708106",
          3845 => x"51515170",
          3846 => x"802ee238",
          3847 => x"7181ff06",
          3848 => x"5187c094",
          3849 => x"80527080",
          3850 => x"2e863887",
          3851 => x"c0949052",
          3852 => x"71087081",
          3853 => x"ff0682b5",
          3854 => x"a80c5184",
          3855 => x"3d0d04ff",
          3856 => x"af3f82b5",
          3857 => x"a80881ff",
          3858 => x"0682b5a8",
          3859 => x"0c04fe3d",
          3860 => x"0d82b3c8",
          3861 => x"337081ff",
          3862 => x"06525387",
          3863 => x"c0948452",
          3864 => x"70802e86",
          3865 => x"3887c094",
          3866 => x"94527108",
          3867 => x"70822a70",
          3868 => x"81065151",
          3869 => x"51ff5270",
          3870 => x"802ea038",
          3871 => x"7281ff06",
          3872 => x"5187c094",
          3873 => x"80527080",
          3874 => x"2e863887",
          3875 => x"c0949052",
          3876 => x"71087098",
          3877 => x"2b70982c",
          3878 => x"51535171",
          3879 => x"82b5a80c",
          3880 => x"843d0d04",
          3881 => x"ff3d0d87",
          3882 => x"c09e8008",
          3883 => x"709c2a8a",
          3884 => x"06515170",
          3885 => x"802e84b4",
          3886 => x"3887c09e",
          3887 => x"a40882b3",
          3888 => x"cc0c87c0",
          3889 => x"9ea80882",
          3890 => x"b3d00c87",
          3891 => x"c09e9408",
          3892 => x"82b3d40c",
          3893 => x"87c09e98",
          3894 => x"0882b3d8",
          3895 => x"0c87c09e",
          3896 => x"9c0882b3",
          3897 => x"dc0c87c0",
          3898 => x"9ea00882",
          3899 => x"b3e00c87",
          3900 => x"c09eac08",
          3901 => x"82b3e40c",
          3902 => x"87c09eb0",
          3903 => x"0882b3e8",
          3904 => x"0c87c09e",
          3905 => x"b40882b3",
          3906 => x"ec0c87c0",
          3907 => x"9eb80882",
          3908 => x"b3f00c87",
          3909 => x"c09ebc08",
          3910 => x"82b3f40c",
          3911 => x"87c09ec0",
          3912 => x"0882b3f8",
          3913 => x"0c87c09e",
          3914 => x"c40882b3",
          3915 => x"fc0c87c0",
          3916 => x"9e800851",
          3917 => x"7082b480",
          3918 => x"2387c09e",
          3919 => x"840882b4",
          3920 => x"840c87c0",
          3921 => x"9e880882",
          3922 => x"b4880c87",
          3923 => x"c09e8c08",
          3924 => x"82b48c0c",
          3925 => x"810b82b4",
          3926 => x"9034800b",
          3927 => x"87c09e90",
          3928 => x"08708480",
          3929 => x"0a065152",
          3930 => x"5270802e",
          3931 => x"83388152",
          3932 => x"7182b491",
          3933 => x"34800b87",
          3934 => x"c09e9008",
          3935 => x"7088800a",
          3936 => x"06515252",
          3937 => x"70802e83",
          3938 => x"38815271",
          3939 => x"82b49234",
          3940 => x"800b87c0",
          3941 => x"9e900870",
          3942 => x"90800a06",
          3943 => x"51525270",
          3944 => x"802e8338",
          3945 => x"81527182",
          3946 => x"b4933480",
          3947 => x"0b87c09e",
          3948 => x"90087088",
          3949 => x"80800651",
          3950 => x"52527080",
          3951 => x"2e833881",
          3952 => x"527182b4",
          3953 => x"9434800b",
          3954 => x"87c09e90",
          3955 => x"0870a080",
          3956 => x"80065152",
          3957 => x"5270802e",
          3958 => x"83388152",
          3959 => x"7182b495",
          3960 => x"34800b87",
          3961 => x"c09e9008",
          3962 => x"70908080",
          3963 => x"06515252",
          3964 => x"70802e83",
          3965 => x"38815271",
          3966 => x"82b49634",
          3967 => x"800b87c0",
          3968 => x"9e900870",
          3969 => x"84808006",
          3970 => x"51525270",
          3971 => x"802e8338",
          3972 => x"81527182",
          3973 => x"b4973480",
          3974 => x"0b87c09e",
          3975 => x"90087082",
          3976 => x"80800651",
          3977 => x"52527080",
          3978 => x"2e833881",
          3979 => x"527182b4",
          3980 => x"9834800b",
          3981 => x"87c09e90",
          3982 => x"08708180",
          3983 => x"80065152",
          3984 => x"5270802e",
          3985 => x"83388152",
          3986 => x"7182b499",
          3987 => x"34800b87",
          3988 => x"c09e9008",
          3989 => x"7080c080",
          3990 => x"06515252",
          3991 => x"70802e83",
          3992 => x"38815271",
          3993 => x"82b49a34",
          3994 => x"800b87c0",
          3995 => x"9e900870",
          3996 => x"a0800651",
          3997 => x"52527080",
          3998 => x"2e833881",
          3999 => x"527182b4",
          4000 => x"9b3487c0",
          4001 => x"9e900870",
          4002 => x"98800670",
          4003 => x"8a2a5151",
          4004 => x"517082b4",
          4005 => x"9c34800b",
          4006 => x"87c09e90",
          4007 => x"08708480",
          4008 => x"06515252",
          4009 => x"70802e83",
          4010 => x"38815271",
          4011 => x"82b49d34",
          4012 => x"87c09e90",
          4013 => x"087083f0",
          4014 => x"0670842a",
          4015 => x"51515170",
          4016 => x"82b49e34",
          4017 => x"800b87c0",
          4018 => x"9e900870",
          4019 => x"88065152",
          4020 => x"5270802e",
          4021 => x"83388152",
          4022 => x"7182b49f",
          4023 => x"3487c09e",
          4024 => x"90087087",
          4025 => x"06515170",
          4026 => x"82b4a034",
          4027 => x"833d0d04",
          4028 => x"fb3d0d82",
          4029 => x"a4e051ff",
          4030 => x"bd893f82",
          4031 => x"b4903354",
          4032 => x"73802e89",
          4033 => x"3882a4f4",
          4034 => x"51ffbcf7",
          4035 => x"3f82a588",
          4036 => x"51ffbcef",
          4037 => x"3f82b492",
          4038 => x"33547380",
          4039 => x"2e943882",
          4040 => x"b3ec0882",
          4041 => x"b3f00811",
          4042 => x"545282a5",
          4043 => x"a051ff95",
          4044 => x"a53f82b4",
          4045 => x"97335473",
          4046 => x"802e9438",
          4047 => x"82b3e408",
          4048 => x"82b3e808",
          4049 => x"11545282",
          4050 => x"a5bc51ff",
          4051 => x"95883f82",
          4052 => x"b4943354",
          4053 => x"73802e94",
          4054 => x"3882b3cc",
          4055 => x"0882b3d0",
          4056 => x"08115452",
          4057 => x"82a5d851",
          4058 => x"ff94eb3f",
          4059 => x"82b49533",
          4060 => x"5473802e",
          4061 => x"943882b3",
          4062 => x"d40882b3",
          4063 => x"d8081154",
          4064 => x"5282a5f4",
          4065 => x"51ff94ce",
          4066 => x"3f82b496",
          4067 => x"33547380",
          4068 => x"2e943882",
          4069 => x"b3dc0882",
          4070 => x"b3e00811",
          4071 => x"545282a6",
          4072 => x"9051ff94",
          4073 => x"b13f82b4",
          4074 => x"9b335473",
          4075 => x"802e8e38",
          4076 => x"82b49c33",
          4077 => x"5282a6ac",
          4078 => x"51ff949a",
          4079 => x"3f82b49f",
          4080 => x"33547380",
          4081 => x"2e8e3882",
          4082 => x"b4a03352",
          4083 => x"82a6cc51",
          4084 => x"ff94833f",
          4085 => x"82b49d33",
          4086 => x"5473802e",
          4087 => x"8e3882b4",
          4088 => x"9e335282",
          4089 => x"a6ec51ff",
          4090 => x"93ec3f82",
          4091 => x"b4913354",
          4092 => x"73802e89",
          4093 => x"3882a78c",
          4094 => x"51ffbb87",
          4095 => x"3f82b493",
          4096 => x"33547380",
          4097 => x"2e893882",
          4098 => x"a7a051ff",
          4099 => x"baf53f82",
          4100 => x"b4983354",
          4101 => x"73802e89",
          4102 => x"3882a7ac",
          4103 => x"51ffbae3",
          4104 => x"3f82b499",
          4105 => x"33547380",
          4106 => x"2e893882",
          4107 => x"a7b851ff",
          4108 => x"bad13f82",
          4109 => x"b49a3354",
          4110 => x"73802e89",
          4111 => x"3882a7c4",
          4112 => x"51ffbabf",
          4113 => x"3f82a7d0",
          4114 => x"51ffbab7",
          4115 => x"3f82b3f4",
          4116 => x"085282a7",
          4117 => x"dc51ff92",
          4118 => x"fd3f82b3",
          4119 => x"f8085282",
          4120 => x"a88451ff",
          4121 => x"92f03f82",
          4122 => x"b3fc0852",
          4123 => x"82a8ac51",
          4124 => x"ff92e33f",
          4125 => x"82a8d451",
          4126 => x"ffba883f",
          4127 => x"82b48022",
          4128 => x"5282a8dc",
          4129 => x"51ff92ce",
          4130 => x"3f82b484",
          4131 => x"0856bd84",
          4132 => x"c0527551",
          4133 => x"d18d3f82",
          4134 => x"b5a808bd",
          4135 => x"84c02976",
          4136 => x"71315454",
          4137 => x"82b5a808",
          4138 => x"5282a984",
          4139 => x"51ff92a6",
          4140 => x"3f82b497",
          4141 => x"33547380",
          4142 => x"2ea93882",
          4143 => x"b4880856",
          4144 => x"bd84c052",
          4145 => x"7551d0db",
          4146 => x"3f82b5a8",
          4147 => x"08bd84c0",
          4148 => x"29767131",
          4149 => x"545482b5",
          4150 => x"a8085282",
          4151 => x"a9b051ff",
          4152 => x"91f43f82",
          4153 => x"b4923354",
          4154 => x"73802ea9",
          4155 => x"3882b48c",
          4156 => x"0856bd84",
          4157 => x"c0527551",
          4158 => x"d0a93f82",
          4159 => x"b5a808bd",
          4160 => x"84c02976",
          4161 => x"71315454",
          4162 => x"82b5a808",
          4163 => x"5282a9dc",
          4164 => x"51ff91c2",
          4165 => x"3f82a1f0",
          4166 => x"51ffb8e7",
          4167 => x"3f873d0d",
          4168 => x"04fe3d0d",
          4169 => x"02920533",
          4170 => x"ff055271",
          4171 => x"8426aa38",
          4172 => x"71842982",
          4173 => x"95900552",
          4174 => x"71080482",
          4175 => x"aa88519d",
          4176 => x"3982aa90",
          4177 => x"51973982",
          4178 => x"aa985191",
          4179 => x"3982aaa0",
          4180 => x"518b3982",
          4181 => x"aaa45185",
          4182 => x"3982aaac",
          4183 => x"51ffb8a3",
          4184 => x"3f843d0d",
          4185 => x"04718880",
          4186 => x"0c04800b",
          4187 => x"87c09684",
          4188 => x"0c0482b4",
          4189 => x"a40887c0",
          4190 => x"96840c04",
          4191 => x"fd3d0d76",
          4192 => x"982b7098",
          4193 => x"2c79982b",
          4194 => x"70982c72",
          4195 => x"10137082",
          4196 => x"2b515351",
          4197 => x"54515180",
          4198 => x"0b82aab8",
          4199 => x"12335553",
          4200 => x"7174259c",
          4201 => x"3882aab4",
          4202 => x"11081202",
          4203 => x"84059705",
          4204 => x"33713352",
          4205 => x"52527072",
          4206 => x"2e098106",
          4207 => x"83388153",
          4208 => x"7282b5a8",
          4209 => x"0c853d0d",
          4210 => x"04fc3d0d",
          4211 => x"78028405",
          4212 => x"9f053371",
          4213 => x"33545553",
          4214 => x"71802ea2",
          4215 => x"388851ff",
          4216 => x"bac33fa0",
          4217 => x"51ffbabd",
          4218 => x"3f8851ff",
          4219 => x"bab73f72",
          4220 => x"33ff0552",
          4221 => x"71733471",
          4222 => x"81ff0652",
          4223 => x"db397651",
          4224 => x"ffb7803f",
          4225 => x"73733486",
          4226 => x"3d0d04f6",
          4227 => x"3d0d7c02",
          4228 => x"8405b705",
          4229 => x"33028805",
          4230 => x"bb053382",
          4231 => x"b5803370",
          4232 => x"842982b4",
          4233 => x"a8057008",
          4234 => x"5159595a",
          4235 => x"58597480",
          4236 => x"2e863874",
          4237 => x"519ab23f",
          4238 => x"82b58033",
          4239 => x"70842982",
          4240 => x"b4a80581",
          4241 => x"19705458",
          4242 => x"565a9db3",
          4243 => x"3f82b5a8",
          4244 => x"08750c82",
          4245 => x"b5803370",
          4246 => x"842982b4",
          4247 => x"a8057008",
          4248 => x"51565a74",
          4249 => x"802ea638",
          4250 => x"75537852",
          4251 => x"7451c495",
          4252 => x"3f82b580",
          4253 => x"33810555",
          4254 => x"7482b580",
          4255 => x"347481ff",
          4256 => x"06559375",
          4257 => x"27873880",
          4258 => x"0b82b580",
          4259 => x"3477802e",
          4260 => x"b63882b4",
          4261 => x"fc085675",
          4262 => x"802eac38",
          4263 => x"82b4f833",
          4264 => x"5574a438",
          4265 => x"8c3dfc05",
          4266 => x"54765378",
          4267 => x"52755180",
          4268 => x"d9c13f82",
          4269 => x"b4fc0852",
          4270 => x"8a51818e",
          4271 => x"ce3f82b4",
          4272 => x"fc085180",
          4273 => x"dd9e3f8c",
          4274 => x"3d0d04fd",
          4275 => x"3d0d82b4",
          4276 => x"a8539354",
          4277 => x"72085271",
          4278 => x"802e8938",
          4279 => x"71519989",
          4280 => x"3f80730c",
          4281 => x"ff148414",
          4282 => x"54547380",
          4283 => x"25e63880",
          4284 => x"0b82b580",
          4285 => x"3482b4fc",
          4286 => x"08527180",
          4287 => x"2e953871",
          4288 => x"5180ddfe",
          4289 => x"3f82b4fc",
          4290 => x"085198dd",
          4291 => x"3f800b82",
          4292 => x"b4fc0c85",
          4293 => x"3d0d04dc",
          4294 => x"3d0d8157",
          4295 => x"805282b4",
          4296 => x"fc085180",
          4297 => x"e2eb3f82",
          4298 => x"b5a80880",
          4299 => x"d23882b4",
          4300 => x"fc085380",
          4301 => x"f852883d",
          4302 => x"70525681",
          4303 => x"8bb93f82",
          4304 => x"b5a80880",
          4305 => x"2eb93875",
          4306 => x"51c0da3f",
          4307 => x"82b5a808",
          4308 => x"55800b82",
          4309 => x"b5a80825",
          4310 => x"9d3882b5",
          4311 => x"a808ff05",
          4312 => x"70175555",
          4313 => x"80743475",
          4314 => x"53765281",
          4315 => x"1782ada8",
          4316 => x"5257ff8c",
          4317 => x"e13f74ff",
          4318 => x"2e098106",
          4319 => x"ffb038a6",
          4320 => x"3d0d04d9",
          4321 => x"3d0daa3d",
          4322 => x"08ad3d08",
          4323 => x"5a5a8170",
          4324 => x"58588052",
          4325 => x"82b4fc08",
          4326 => x"5180e1f5",
          4327 => x"3f82b5a8",
          4328 => x"08819538",
          4329 => x"ff0b82b4",
          4330 => x"fc085455",
          4331 => x"80f8528b",
          4332 => x"3d705256",
          4333 => x"818ac03f",
          4334 => x"82b5a808",
          4335 => x"802ea538",
          4336 => x"7551ffbf",
          4337 => x"e03f82b5",
          4338 => x"a8088118",
          4339 => x"5855800b",
          4340 => x"82b5a808",
          4341 => x"258e3882",
          4342 => x"b5a808ff",
          4343 => x"05701755",
          4344 => x"55807434",
          4345 => x"74097030",
          4346 => x"7072079f",
          4347 => x"2a515555",
          4348 => x"78772e85",
          4349 => x"3873ffac",
          4350 => x"3882b4fc",
          4351 => x"088c1108",
          4352 => x"535180e1",
          4353 => x"8c3f82b5",
          4354 => x"a808802e",
          4355 => x"893882ad",
          4356 => x"b451ffb2",
          4357 => x"ee3f7877",
          4358 => x"2e098106",
          4359 => x"9b387552",
          4360 => x"7951ffbf",
          4361 => x"ee3f7951",
          4362 => x"ffbefa3f",
          4363 => x"ab3d0854",
          4364 => x"82b5a808",
          4365 => x"74348058",
          4366 => x"7782b5a8",
          4367 => x"0ca93d0d",
          4368 => x"04f63d0d",
          4369 => x"7c7e715c",
          4370 => x"71723357",
          4371 => x"595a5873",
          4372 => x"a02e0981",
          4373 => x"06a23878",
          4374 => x"33780556",
          4375 => x"77762798",
          4376 => x"38811770",
          4377 => x"5b707133",
          4378 => x"56585573",
          4379 => x"a02e0981",
          4380 => x"06863875",
          4381 => x"7526ea38",
          4382 => x"80547388",
          4383 => x"2982b584",
          4384 => x"05700852",
          4385 => x"55ffbe9d",
          4386 => x"3f82b5a8",
          4387 => x"08537952",
          4388 => x"740851c1",
          4389 => x"9d3f82b5",
          4390 => x"a80880c6",
          4391 => x"38841533",
          4392 => x"5574812e",
          4393 => x"88387482",
          4394 => x"2e8838b6",
          4395 => x"39fce83f",
          4396 => x"ad39811a",
          4397 => x"5a8c3dfc",
          4398 => x"1153f805",
          4399 => x"51ffabf2",
          4400 => x"3f82b5a8",
          4401 => x"08802e9a",
          4402 => x"38ff1b53",
          4403 => x"78527751",
          4404 => x"fdb13f82",
          4405 => x"b5a80881",
          4406 => x"ff065574",
          4407 => x"85387454",
          4408 => x"91398114",
          4409 => x"7081ff06",
          4410 => x"51548274",
          4411 => x"27ff8b38",
          4412 => x"80547382",
          4413 => x"b5a80c8c",
          4414 => x"3d0d04d3",
          4415 => x"3d0db03d",
          4416 => x"08b23d08",
          4417 => x"b43d0859",
          4418 => x"5f5a800b",
          4419 => x"af3d3482",
          4420 => x"b5803382",
          4421 => x"b4fc0855",
          4422 => x"5b7381cb",
          4423 => x"387382b4",
          4424 => x"f8335555",
          4425 => x"73833881",
          4426 => x"5576802e",
          4427 => x"81bc3881",
          4428 => x"70760655",
          4429 => x"5673802e",
          4430 => x"81ad38a8",
          4431 => x"5197c03f",
          4432 => x"82b5a808",
          4433 => x"82b4fc0c",
          4434 => x"82b5a808",
          4435 => x"802e8192",
          4436 => x"38935376",
          4437 => x"5282b5a8",
          4438 => x"085180cc",
          4439 => x"b43f82b5",
          4440 => x"a808802e",
          4441 => x"8c3882ad",
          4442 => x"e051ffb0",
          4443 => x"963f80f7",
          4444 => x"3982b5a8",
          4445 => x"085b82b4",
          4446 => x"fc085380",
          4447 => x"f852903d",
          4448 => x"70525481",
          4449 => x"86f13f82",
          4450 => x"b5a80856",
          4451 => x"82b5a808",
          4452 => x"742e0981",
          4453 => x"0680d038",
          4454 => x"82b5a808",
          4455 => x"51ffbc85",
          4456 => x"3f82b5a8",
          4457 => x"0855800b",
          4458 => x"82b5a808",
          4459 => x"25a93882",
          4460 => x"b5a808ff",
          4461 => x"05701755",
          4462 => x"55807434",
          4463 => x"80537481",
          4464 => x"ff065275",
          4465 => x"51f8c43f",
          4466 => x"811b7081",
          4467 => x"ff065c54",
          4468 => x"937b2783",
          4469 => x"38805b74",
          4470 => x"ff2e0981",
          4471 => x"06ff9738",
          4472 => x"86397582",
          4473 => x"b4f83476",
          4474 => x"8c3882b4",
          4475 => x"fc08802e",
          4476 => x"8438f9d7",
          4477 => x"3f8f3d5d",
          4478 => x"ecd43f82",
          4479 => x"b5a80898",
          4480 => x"2b70982c",
          4481 => x"515978ff",
          4482 => x"2eee3878",
          4483 => x"81ff0682",
          4484 => x"ccd43370",
          4485 => x"982b7098",
          4486 => x"2c82ccd0",
          4487 => x"3370982b",
          4488 => x"70972c71",
          4489 => x"982c0570",
          4490 => x"842982aa",
          4491 => x"b4057008",
          4492 => x"15703351",
          4493 => x"51515159",
          4494 => x"5951595d",
          4495 => x"58815673",
          4496 => x"782e80e9",
          4497 => x"38777427",
          4498 => x"b4387481",
          4499 => x"800a2981",
          4500 => x"ff0a0570",
          4501 => x"982c5155",
          4502 => x"80752480",
          4503 => x"ce387653",
          4504 => x"74527751",
          4505 => x"f6963f82",
          4506 => x"b5a80881",
          4507 => x"ff065473",
          4508 => x"802ed738",
          4509 => x"7482ccd0",
          4510 => x"348156b1",
          4511 => x"39748180",
          4512 => x"0a298180",
          4513 => x"0a057098",
          4514 => x"2c7081ff",
          4515 => x"06565155",
          4516 => x"73952697",
          4517 => x"38765374",
          4518 => x"527751f5",
          4519 => x"df3f82b5",
          4520 => x"a80881ff",
          4521 => x"065473cc",
          4522 => x"38d33980",
          4523 => x"5675802e",
          4524 => x"80ca3881",
          4525 => x"1c557482",
          4526 => x"ccd43474",
          4527 => x"982b7098",
          4528 => x"2c82ccd0",
          4529 => x"3370982b",
          4530 => x"70982c70",
          4531 => x"10117082",
          4532 => x"2b82aab8",
          4533 => x"11335e51",
          4534 => x"51515758",
          4535 => x"51557477",
          4536 => x"2e098106",
          4537 => x"fe923882",
          4538 => x"aabc1408",
          4539 => x"7d0c800b",
          4540 => x"82ccd434",
          4541 => x"800b82cc",
          4542 => x"d0349239",
          4543 => x"7582ccd4",
          4544 => x"347582cc",
          4545 => x"d03478af",
          4546 => x"3d34757d",
          4547 => x"0c7e5473",
          4548 => x"9526fde1",
          4549 => x"38738429",
          4550 => x"8295a405",
          4551 => x"54730804",
          4552 => x"82ccdc33",
          4553 => x"54737e2e",
          4554 => x"fdcb3882",
          4555 => x"ccd83355",
          4556 => x"737527ab",
          4557 => x"3874982b",
          4558 => x"70982c51",
          4559 => x"55737524",
          4560 => x"9e38741a",
          4561 => x"54733381",
          4562 => x"15347481",
          4563 => x"800a2981",
          4564 => x"ff0a0570",
          4565 => x"982c82cc",
          4566 => x"dc335651",
          4567 => x"55df3982",
          4568 => x"ccdc3381",
          4569 => x"11565474",
          4570 => x"82ccdc34",
          4571 => x"731a54ae",
          4572 => x"3d337434",
          4573 => x"82ccd833",
          4574 => x"54737e25",
          4575 => x"89388114",
          4576 => x"547382cc",
          4577 => x"d83482cc",
          4578 => x"dc337081",
          4579 => x"800a2981",
          4580 => x"ff0a0570",
          4581 => x"982c82cc",
          4582 => x"d8335a51",
          4583 => x"56567477",
          4584 => x"25a33874",
          4585 => x"1a703352",
          4586 => x"54ffaef9",
          4587 => x"3f748180",
          4588 => x"0a298180",
          4589 => x"0a057098",
          4590 => x"2c82ccd8",
          4591 => x"33565155",
          4592 => x"737524df",
          4593 => x"3882ccdc",
          4594 => x"3370982b",
          4595 => x"70982c82",
          4596 => x"ccd8335a",
          4597 => x"51565674",
          4598 => x"7725fc99",
          4599 => x"388851ff",
          4600 => x"aec33f74",
          4601 => x"81800a29",
          4602 => x"81800a05",
          4603 => x"70982c82",
          4604 => x"ccd83356",
          4605 => x"51557375",
          4606 => x"24e338fb",
          4607 => x"f839837a",
          4608 => x"34800b81",
          4609 => x"1b3482cc",
          4610 => x"dc538052",
          4611 => x"82a2f051",
          4612 => x"f3b73f81",
          4613 => x"e43982cc",
          4614 => x"dc337081",
          4615 => x"ff065555",
          4616 => x"73802efb",
          4617 => x"d03882cc",
          4618 => x"d833ff05",
          4619 => x"547382cc",
          4620 => x"d834ff15",
          4621 => x"547382cc",
          4622 => x"dc348851",
          4623 => x"ffade63f",
          4624 => x"82ccdc33",
          4625 => x"70982b70",
          4626 => x"982c82cc",
          4627 => x"d8335751",
          4628 => x"56577474",
          4629 => x"25a83874",
          4630 => x"1a548114",
          4631 => x"33743473",
          4632 => x"3351ffad",
          4633 => x"c03f7481",
          4634 => x"800a2981",
          4635 => x"800a0570",
          4636 => x"982c82cc",
          4637 => x"d8335851",
          4638 => x"55757524",
          4639 => x"da38a051",
          4640 => x"ffada23f",
          4641 => x"82ccdc33",
          4642 => x"70982b70",
          4643 => x"982c82cc",
          4644 => x"d8335751",
          4645 => x"56577474",
          4646 => x"24fada38",
          4647 => x"8851ffad",
          4648 => x"843f7481",
          4649 => x"800a2981",
          4650 => x"800a0570",
          4651 => x"982c82cc",
          4652 => x"d8335851",
          4653 => x"55757525",
          4654 => x"e338fab9",
          4655 => x"3982ccd8",
          4656 => x"337a0554",
          4657 => x"8074348a",
          4658 => x"51ffacd9",
          4659 => x"3f82ccd8",
          4660 => x"527951f6",
          4661 => x"ec3f82b5",
          4662 => x"a80881ff",
          4663 => x"06547396",
          4664 => x"3882ccd8",
          4665 => x"33547380",
          4666 => x"2e8f3881",
          4667 => x"53735279",
          4668 => x"51f2983f",
          4669 => x"8439807a",
          4670 => x"34800b82",
          4671 => x"ccdc3480",
          4672 => x"0b82ccd8",
          4673 => x"347982b5",
          4674 => x"a80caf3d",
          4675 => x"0d0482cc",
          4676 => x"dc335473",
          4677 => x"802ef9dd",
          4678 => x"388851ff",
          4679 => x"ac873f82",
          4680 => x"ccdc33ff",
          4681 => x"05547382",
          4682 => x"ccdc3473",
          4683 => x"81ff0654",
          4684 => x"e23982cc",
          4685 => x"dc3382cc",
          4686 => x"d8335555",
          4687 => x"73752ef9",
          4688 => x"b438ff14",
          4689 => x"547382cc",
          4690 => x"d8347498",
          4691 => x"2b70982c",
          4692 => x"7581ff06",
          4693 => x"56515574",
          4694 => x"7425a838",
          4695 => x"741a5481",
          4696 => x"14337434",
          4697 => x"733351ff",
          4698 => x"abbb3f74",
          4699 => x"81800a29",
          4700 => x"81800a05",
          4701 => x"70982c82",
          4702 => x"ccd83358",
          4703 => x"51557575",
          4704 => x"24da38a0",
          4705 => x"51ffab9d",
          4706 => x"3f82ccdc",
          4707 => x"3370982b",
          4708 => x"70982c82",
          4709 => x"ccd83357",
          4710 => x"51565774",
          4711 => x"7424f8d5",
          4712 => x"388851ff",
          4713 => x"aaff3f74",
          4714 => x"81800a29",
          4715 => x"81800a05",
          4716 => x"70982c82",
          4717 => x"ccd83358",
          4718 => x"51557575",
          4719 => x"25e338f8",
          4720 => x"b43982cc",
          4721 => x"dc337081",
          4722 => x"ff0682cc",
          4723 => x"d8335956",
          4724 => x"54747727",
          4725 => x"f89f3881",
          4726 => x"14547382",
          4727 => x"ccdc3474",
          4728 => x"1a703352",
          4729 => x"54ffaabd",
          4730 => x"3f82ccdc",
          4731 => x"337081ff",
          4732 => x"0682ccd8",
          4733 => x"33585654",
          4734 => x"757526db",
          4735 => x"38f7f639",
          4736 => x"82ccdc53",
          4737 => x"805282a2",
          4738 => x"f051efbd",
          4739 => x"3f800b82",
          4740 => x"ccdc3480",
          4741 => x"0b82ccd8",
          4742 => x"34f7da39",
          4743 => x"7ab03882",
          4744 => x"b4f40855",
          4745 => x"74802ea6",
          4746 => x"387451ff",
          4747 => x"b2f73f82",
          4748 => x"b5a80882",
          4749 => x"ccd83482",
          4750 => x"b5a80881",
          4751 => x"ff068105",
          4752 => x"53745279",
          4753 => x"51ffb4bd",
          4754 => x"3f935b81",
          4755 => x"c0397a84",
          4756 => x"2982b4a8",
          4757 => x"05fc1108",
          4758 => x"56547480",
          4759 => x"2ea73874",
          4760 => x"51ffb2c1",
          4761 => x"3f82b5a8",
          4762 => x"0882ccd8",
          4763 => x"3482b5a8",
          4764 => x"0881ff06",
          4765 => x"81055374",
          4766 => x"527951ff",
          4767 => x"b4873fff",
          4768 => x"1b5480fa",
          4769 => x"39730855",
          4770 => x"74802ef6",
          4771 => x"e8387451",
          4772 => x"ffb2923f",
          4773 => x"99397a93",
          4774 => x"2e098106",
          4775 => x"ae3882b4",
          4776 => x"a8085574",
          4777 => x"802ea438",
          4778 => x"7451ffb1",
          4779 => x"f83f82b5",
          4780 => x"a80882cc",
          4781 => x"d83482b5",
          4782 => x"a80881ff",
          4783 => x"06810553",
          4784 => x"74527951",
          4785 => x"ffb3be3f",
          4786 => x"80c3397a",
          4787 => x"842982b4",
          4788 => x"ac057008",
          4789 => x"56547480",
          4790 => x"2eab3874",
          4791 => x"51ffb1c5",
          4792 => x"3f82b5a8",
          4793 => x"0882ccd8",
          4794 => x"3482b5a8",
          4795 => x"0881ff06",
          4796 => x"81055374",
          4797 => x"527951ff",
          4798 => x"b38b3f81",
          4799 => x"1b547381",
          4800 => x"ff065b89",
          4801 => x"397482cc",
          4802 => x"d834747a",
          4803 => x"3482ccdc",
          4804 => x"5382ccd8",
          4805 => x"33527951",
          4806 => x"edaf3ff5",
          4807 => x"d83982cc",
          4808 => x"dc337081",
          4809 => x"ff0682cc",
          4810 => x"d8335956",
          4811 => x"54747727",
          4812 => x"f5c33881",
          4813 => x"14547382",
          4814 => x"ccdc3474",
          4815 => x"1a703352",
          4816 => x"54ffa7e1",
          4817 => x"3ff5ae39",
          4818 => x"82ccdc33",
          4819 => x"5473802e",
          4820 => x"f5a33888",
          4821 => x"51ffa7cd",
          4822 => x"3f82ccdc",
          4823 => x"33ff0554",
          4824 => x"7382ccdc",
          4825 => x"34f58e39",
          4826 => x"f93d0d83",
          4827 => x"dff40b82",
          4828 => x"b5a00c82",
          4829 => x"800b82b5",
          4830 => x"9c239080",
          4831 => x"53805283",
          4832 => x"dff451ff",
          4833 => x"b7803f82",
          4834 => x"b5a00854",
          4835 => x"80587774",
          4836 => x"34815776",
          4837 => x"81153482",
          4838 => x"b5a00854",
          4839 => x"77841534",
          4840 => x"76851534",
          4841 => x"82b5a008",
          4842 => x"54778615",
          4843 => x"34768715",
          4844 => x"3482b5a0",
          4845 => x"0882b59c",
          4846 => x"22ff05fe",
          4847 => x"80800770",
          4848 => x"83ffff06",
          4849 => x"70882a58",
          4850 => x"51555674",
          4851 => x"88173473",
          4852 => x"89173482",
          4853 => x"b59c2270",
          4854 => x"882982b5",
          4855 => x"a00805f8",
          4856 => x"11515555",
          4857 => x"77821534",
          4858 => x"76831534",
          4859 => x"893d0d04",
          4860 => x"ff3d0d73",
          4861 => x"52815184",
          4862 => x"72278f38",
          4863 => x"fb12832a",
          4864 => x"82117083",
          4865 => x"ffff0651",
          4866 => x"51517082",
          4867 => x"b5a80c83",
          4868 => x"3d0d04f9",
          4869 => x"3d0d02a6",
          4870 => x"05220284",
          4871 => x"05aa0522",
          4872 => x"710582b5",
          4873 => x"a0087183",
          4874 => x"2b711174",
          4875 => x"832b7311",
          4876 => x"70338112",
          4877 => x"3371882b",
          4878 => x"0702a405",
          4879 => x"ae052271",
          4880 => x"81ffff06",
          4881 => x"0770882a",
          4882 => x"53515259",
          4883 => x"545b5b57",
          4884 => x"53545571",
          4885 => x"77347081",
          4886 => x"183482b5",
          4887 => x"a0081475",
          4888 => x"882a5254",
          4889 => x"70821534",
          4890 => x"74831534",
          4891 => x"82b5a008",
          4892 => x"70177033",
          4893 => x"81123371",
          4894 => x"882b0770",
          4895 => x"832b8fff",
          4896 => x"f8065152",
          4897 => x"56527105",
          4898 => x"7383ffff",
          4899 => x"0670882a",
          4900 => x"54545171",
          4901 => x"82123472",
          4902 => x"81ff0653",
          4903 => x"72831234",
          4904 => x"82b5a008",
          4905 => x"16567176",
          4906 => x"34728117",
          4907 => x"34893d0d",
          4908 => x"04fb3d0d",
          4909 => x"82b5a008",
          4910 => x"0284059e",
          4911 => x"05227083",
          4912 => x"2b721186",
          4913 => x"11338712",
          4914 => x"33718b2b",
          4915 => x"71832b07",
          4916 => x"585b5952",
          4917 => x"55527205",
          4918 => x"84123385",
          4919 => x"13337188",
          4920 => x"2b077088",
          4921 => x"2a545656",
          4922 => x"52708413",
          4923 => x"34738513",
          4924 => x"3482b5a0",
          4925 => x"08701484",
          4926 => x"11338512",
          4927 => x"33718b2b",
          4928 => x"71832b07",
          4929 => x"56595752",
          4930 => x"72058612",
          4931 => x"33871333",
          4932 => x"71882b07",
          4933 => x"70882a54",
          4934 => x"56565270",
          4935 => x"86133473",
          4936 => x"87133482",
          4937 => x"b5a00813",
          4938 => x"70338112",
          4939 => x"3371882b",
          4940 => x"077081ff",
          4941 => x"ff067088",
          4942 => x"2a535153",
          4943 => x"53537173",
          4944 => x"34708114",
          4945 => x"34873d0d",
          4946 => x"04fa3d0d",
          4947 => x"02a20522",
          4948 => x"82b5a008",
          4949 => x"71832b71",
          4950 => x"11703381",
          4951 => x"12337188",
          4952 => x"2b077088",
          4953 => x"29157033",
          4954 => x"81123371",
          4955 => x"982b7190",
          4956 => x"2b07535f",
          4957 => x"5355525a",
          4958 => x"56575354",
          4959 => x"71802580",
          4960 => x"f6387251",
          4961 => x"feab3f82",
          4962 => x"b5a00870",
          4963 => x"16703381",
          4964 => x"1233718b",
          4965 => x"2b71832b",
          4966 => x"07741170",
          4967 => x"33811233",
          4968 => x"71882b07",
          4969 => x"70832b8f",
          4970 => x"fff80651",
          4971 => x"52545153",
          4972 => x"5a585372",
          4973 => x"0574882a",
          4974 => x"54527282",
          4975 => x"13347383",
          4976 => x"133482b5",
          4977 => x"a0087016",
          4978 => x"70338112",
          4979 => x"33718b2b",
          4980 => x"71832b07",
          4981 => x"56595755",
          4982 => x"72057033",
          4983 => x"81123371",
          4984 => x"882b0770",
          4985 => x"81ffff06",
          4986 => x"70882a57",
          4987 => x"51525852",
          4988 => x"72743471",
          4989 => x"81153488",
          4990 => x"3d0d04fb",
          4991 => x"3d0d82b5",
          4992 => x"a0080284",
          4993 => x"059e0522",
          4994 => x"70832b72",
          4995 => x"11821133",
          4996 => x"83123371",
          4997 => x"8b2b7183",
          4998 => x"2b07595b",
          4999 => x"59525652",
          5000 => x"73057133",
          5001 => x"81133371",
          5002 => x"882b0702",
          5003 => x"8c05a205",
          5004 => x"22710770",
          5005 => x"882a5351",
          5006 => x"53535371",
          5007 => x"73347081",
          5008 => x"143482b5",
          5009 => x"a0087015",
          5010 => x"70338112",
          5011 => x"33718b2b",
          5012 => x"71832b07",
          5013 => x"56595752",
          5014 => x"72058212",
          5015 => x"33831333",
          5016 => x"71882b07",
          5017 => x"70882a54",
          5018 => x"55565270",
          5019 => x"82133472",
          5020 => x"83133482",
          5021 => x"b5a00814",
          5022 => x"82113383",
          5023 => x"12337188",
          5024 => x"2b0782b5",
          5025 => x"a80c5254",
          5026 => x"873d0d04",
          5027 => x"f73d0d7b",
          5028 => x"82b5a008",
          5029 => x"31832a70",
          5030 => x"83ffff06",
          5031 => x"70535753",
          5032 => x"fda73f82",
          5033 => x"b5a00876",
          5034 => x"832b7111",
          5035 => x"82113383",
          5036 => x"1233718b",
          5037 => x"2b71832b",
          5038 => x"07751170",
          5039 => x"33811233",
          5040 => x"71982b71",
          5041 => x"902b0753",
          5042 => x"42405153",
          5043 => x"5b585559",
          5044 => x"54728025",
          5045 => x"8d388280",
          5046 => x"80527551",
          5047 => x"fe9d3f81",
          5048 => x"84398414",
          5049 => x"33851533",
          5050 => x"718b2b71",
          5051 => x"832b0776",
          5052 => x"1179882a",
          5053 => x"53515558",
          5054 => x"55768614",
          5055 => x"347581ff",
          5056 => x"06567587",
          5057 => x"143482b5",
          5058 => x"a0087019",
          5059 => x"84123385",
          5060 => x"13337188",
          5061 => x"2b077088",
          5062 => x"2a54575b",
          5063 => x"56537284",
          5064 => x"16347385",
          5065 => x"163482b5",
          5066 => x"a0081853",
          5067 => x"800b8614",
          5068 => x"34800b87",
          5069 => x"143482b5",
          5070 => x"a0085376",
          5071 => x"84143475",
          5072 => x"85143482",
          5073 => x"b5a00818",
          5074 => x"70338112",
          5075 => x"3371882b",
          5076 => x"07708280",
          5077 => x"80077088",
          5078 => x"2a535155",
          5079 => x"56547474",
          5080 => x"34728115",
          5081 => x"348b3d0d",
          5082 => x"04ff3d0d",
          5083 => x"735282b5",
          5084 => x"a0088438",
          5085 => x"f7f23f71",
          5086 => x"802e8638",
          5087 => x"7151fe8c",
          5088 => x"3f833d0d",
          5089 => x"04f53d0d",
          5090 => x"807e5258",
          5091 => x"f8e23f82",
          5092 => x"b5a80883",
          5093 => x"ffff0682",
          5094 => x"b5a00884",
          5095 => x"11338512",
          5096 => x"3371882b",
          5097 => x"07705f59",
          5098 => x"56585a81",
          5099 => x"ffff5975",
          5100 => x"782e80cb",
          5101 => x"38758829",
          5102 => x"17703381",
          5103 => x"12337188",
          5104 => x"2b077081",
          5105 => x"ffff0679",
          5106 => x"317083ff",
          5107 => x"ff06707f",
          5108 => x"27525351",
          5109 => x"56595577",
          5110 => x"79278a38",
          5111 => x"73802e85",
          5112 => x"3875785a",
          5113 => x"5b841533",
          5114 => x"85163371",
          5115 => x"882b0757",
          5116 => x"5475c238",
          5117 => x"7881ffff",
          5118 => x"2e85387a",
          5119 => x"79595680",
          5120 => x"76832b82",
          5121 => x"b5a00811",
          5122 => x"70338112",
          5123 => x"3371882b",
          5124 => x"077081ff",
          5125 => x"ff065152",
          5126 => x"5a565c55",
          5127 => x"73752e83",
          5128 => x"38815580",
          5129 => x"54797826",
          5130 => x"81cc3874",
          5131 => x"5474802e",
          5132 => x"81c43877",
          5133 => x"7a2e0981",
          5134 => x"06893875",
          5135 => x"51f8f23f",
          5136 => x"81ac3982",
          5137 => x"80805379",
          5138 => x"527551f7",
          5139 => x"c63f82b5",
          5140 => x"a008701c",
          5141 => x"86113387",
          5142 => x"1233718b",
          5143 => x"2b71832b",
          5144 => x"07535a5e",
          5145 => x"5574057a",
          5146 => x"177083ff",
          5147 => x"ff067088",
          5148 => x"2a5c5956",
          5149 => x"54788415",
          5150 => x"347681ff",
          5151 => x"06577685",
          5152 => x"153482b5",
          5153 => x"a0087583",
          5154 => x"2b711172",
          5155 => x"1e861133",
          5156 => x"87123371",
          5157 => x"882b0770",
          5158 => x"882a535b",
          5159 => x"5e535a56",
          5160 => x"54738619",
          5161 => x"34758719",
          5162 => x"3482b5a0",
          5163 => x"08701c84",
          5164 => x"11338512",
          5165 => x"33718b2b",
          5166 => x"71832b07",
          5167 => x"535d5a55",
          5168 => x"74055478",
          5169 => x"86153476",
          5170 => x"87153482",
          5171 => x"b5a00870",
          5172 => x"16711d84",
          5173 => x"11338512",
          5174 => x"3371882b",
          5175 => x"0770882a",
          5176 => x"535a5f52",
          5177 => x"56547384",
          5178 => x"16347585",
          5179 => x"163482b5",
          5180 => x"a0081b84",
          5181 => x"05547382",
          5182 => x"b5a80c8d",
          5183 => x"3d0d04fe",
          5184 => x"3d0d7452",
          5185 => x"82b5a008",
          5186 => x"8438f4dc",
          5187 => x"3f715371",
          5188 => x"802e8b38",
          5189 => x"7151fced",
          5190 => x"3f82b5a8",
          5191 => x"08537282",
          5192 => x"b5a80c84",
          5193 => x"3d0d04ee",
          5194 => x"3d0d6466",
          5195 => x"405c8070",
          5196 => x"424082b5",
          5197 => x"a008602e",
          5198 => x"09810684",
          5199 => x"38f4a93f",
          5200 => x"7b8e387e",
          5201 => x"51ffb83f",
          5202 => x"82b5a808",
          5203 => x"5483c739",
          5204 => x"7e8b387b",
          5205 => x"51fc923f",
          5206 => x"7e5483ba",
          5207 => x"397e51f5",
          5208 => x"8f3f82b5",
          5209 => x"a80883ff",
          5210 => x"ff0682b5",
          5211 => x"a0087d71",
          5212 => x"31832a70",
          5213 => x"83ffff06",
          5214 => x"70832b73",
          5215 => x"11703381",
          5216 => x"12337188",
          5217 => x"2b077075",
          5218 => x"317083ff",
          5219 => x"ff067088",
          5220 => x"29fc0573",
          5221 => x"88291a70",
          5222 => x"33811233",
          5223 => x"71882b07",
          5224 => x"70902b53",
          5225 => x"444e5348",
          5226 => x"41525c54",
          5227 => x"5b415c56",
          5228 => x"5b5b7380",
          5229 => x"258f3876",
          5230 => x"81ffff06",
          5231 => x"75317083",
          5232 => x"ffff0642",
          5233 => x"54821633",
          5234 => x"83173371",
          5235 => x"882b0770",
          5236 => x"88291c70",
          5237 => x"33811233",
          5238 => x"71982b71",
          5239 => x"902b0753",
          5240 => x"47455256",
          5241 => x"54738025",
          5242 => x"8b387875",
          5243 => x"317083ff",
          5244 => x"ff064154",
          5245 => x"777b2781",
          5246 => x"fe386018",
          5247 => x"54737b2e",
          5248 => x"0981068f",
          5249 => x"387851f6",
          5250 => x"c03f7a83",
          5251 => x"ffff0658",
          5252 => x"81e5397f",
          5253 => x"8e387a74",
          5254 => x"24893878",
          5255 => x"51f6aa3f",
          5256 => x"81a5397f",
          5257 => x"18557a75",
          5258 => x"2480c838",
          5259 => x"791d8211",
          5260 => x"33831233",
          5261 => x"71882b07",
          5262 => x"535754f4",
          5263 => x"f43f8052",
          5264 => x"7851f7b7",
          5265 => x"3f82b5a8",
          5266 => x"0883ffff",
          5267 => x"067e547c",
          5268 => x"5370832b",
          5269 => x"82b5a008",
          5270 => x"11840553",
          5271 => x"5559ff9f",
          5272 => x"da3f82b5",
          5273 => x"a0081484",
          5274 => x"057583ff",
          5275 => x"ff06595c",
          5276 => x"81853960",
          5277 => x"15547a74",
          5278 => x"2480d438",
          5279 => x"7851f5c9",
          5280 => x"3f82b5a0",
          5281 => x"081d8211",
          5282 => x"33831233",
          5283 => x"71882b07",
          5284 => x"534354f4",
          5285 => x"9c3f8052",
          5286 => x"7851f6df",
          5287 => x"3f82b5a8",
          5288 => x"0883ffff",
          5289 => x"067e547c",
          5290 => x"5370832b",
          5291 => x"82b5a008",
          5292 => x"11840553",
          5293 => x"5559ff9f",
          5294 => x"823f82b5",
          5295 => x"a0081484",
          5296 => x"05606205",
          5297 => x"19555c73",
          5298 => x"83ffff06",
          5299 => x"58a9397b",
          5300 => x"7f5254f9",
          5301 => x"b03f82b5",
          5302 => x"a8085c82",
          5303 => x"b5a80880",
          5304 => x"2e93387d",
          5305 => x"53735282",
          5306 => x"b5a80851",
          5307 => x"ffa3963f",
          5308 => x"7351f798",
          5309 => x"3f7a587a",
          5310 => x"78279938",
          5311 => x"80537a52",
          5312 => x"7851f28f",
          5313 => x"3f7a1983",
          5314 => x"2b82b5a0",
          5315 => x"08058405",
          5316 => x"51f6f93f",
          5317 => x"7b547382",
          5318 => x"b5a80c94",
          5319 => x"3d0d04fc",
          5320 => x"3d0d7777",
          5321 => x"29705254",
          5322 => x"fbd53f82",
          5323 => x"b5a80855",
          5324 => x"82b5a808",
          5325 => x"802e8e38",
          5326 => x"73538052",
          5327 => x"82b5a808",
          5328 => x"51ffa7c2",
          5329 => x"3f7482b5",
          5330 => x"a80c863d",
          5331 => x"0d04ff3d",
          5332 => x"0d028f05",
          5333 => x"33518152",
          5334 => x"70722687",
          5335 => x"3882b5a4",
          5336 => x"11335271",
          5337 => x"82b5a80c",
          5338 => x"833d0d04",
          5339 => x"fc3d0d02",
          5340 => x"9b053302",
          5341 => x"84059f05",
          5342 => x"33565383",
          5343 => x"51728126",
          5344 => x"80e03872",
          5345 => x"842b87c0",
          5346 => x"928c1153",
          5347 => x"51885474",
          5348 => x"802e8438",
          5349 => x"81885473",
          5350 => x"720c87c0",
          5351 => x"928c1151",
          5352 => x"81710c85",
          5353 => x"0b87c098",
          5354 => x"8c0c7052",
          5355 => x"71087082",
          5356 => x"06515170",
          5357 => x"802e8a38",
          5358 => x"87c0988c",
          5359 => x"085170ec",
          5360 => x"387108fc",
          5361 => x"80800652",
          5362 => x"71923887",
          5363 => x"c0988c08",
          5364 => x"5170802e",
          5365 => x"87387182",
          5366 => x"b5a41434",
          5367 => x"82b5a413",
          5368 => x"33517082",
          5369 => x"b5a80c86",
          5370 => x"3d0d04f3",
          5371 => x"3d0d6062",
          5372 => x"64028c05",
          5373 => x"bf053357",
          5374 => x"40585b83",
          5375 => x"74525afe",
          5376 => x"cd3f82b5",
          5377 => x"a8088106",
          5378 => x"7a545271",
          5379 => x"81be3871",
          5380 => x"7275842b",
          5381 => x"87c09280",
          5382 => x"1187c092",
          5383 => x"8c1287c0",
          5384 => x"92841341",
          5385 => x"5a40575a",
          5386 => x"58850b87",
          5387 => x"c0988c0c",
          5388 => x"767d0c84",
          5389 => x"760c7508",
          5390 => x"70852a70",
          5391 => x"81065153",
          5392 => x"5471802e",
          5393 => x"8e387b08",
          5394 => x"52717b70",
          5395 => x"81055d34",
          5396 => x"81195980",
          5397 => x"74a20653",
          5398 => x"5371732e",
          5399 => x"83388153",
          5400 => x"7883ff26",
          5401 => x"8f387280",
          5402 => x"2e8a3887",
          5403 => x"c0988c08",
          5404 => x"5271c338",
          5405 => x"87c0988c",
          5406 => x"08527180",
          5407 => x"2e873878",
          5408 => x"84802e99",
          5409 => x"3881760c",
          5410 => x"87c0928c",
          5411 => x"15537208",
          5412 => x"70820651",
          5413 => x"5271f738",
          5414 => x"ff1a5a8d",
          5415 => x"39848017",
          5416 => x"81197081",
          5417 => x"ff065a53",
          5418 => x"5779802e",
          5419 => x"903873fc",
          5420 => x"80800652",
          5421 => x"7187387d",
          5422 => x"7826feed",
          5423 => x"3873fc80",
          5424 => x"80065271",
          5425 => x"802e8338",
          5426 => x"81527153",
          5427 => x"7282b5a8",
          5428 => x"0c8f3d0d",
          5429 => x"04f33d0d",
          5430 => x"60626402",
          5431 => x"8c05bf05",
          5432 => x"33574058",
          5433 => x"5b835980",
          5434 => x"745258fc",
          5435 => x"e13f82b5",
          5436 => x"a8088106",
          5437 => x"79545271",
          5438 => x"782e0981",
          5439 => x"0681b138",
          5440 => x"7774842b",
          5441 => x"87c09280",
          5442 => x"1187c092",
          5443 => x"8c1287c0",
          5444 => x"92841340",
          5445 => x"595f565a",
          5446 => x"850b87c0",
          5447 => x"988c0c76",
          5448 => x"7d0c8276",
          5449 => x"0c805875",
          5450 => x"0870842a",
          5451 => x"70810651",
          5452 => x"53547180",
          5453 => x"2e8c387a",
          5454 => x"7081055c",
          5455 => x"337c0c81",
          5456 => x"18587381",
          5457 => x"2a708106",
          5458 => x"51527180",
          5459 => x"2e8a3887",
          5460 => x"c0988c08",
          5461 => x"5271d038",
          5462 => x"87c0988c",
          5463 => x"08527180",
          5464 => x"2e873877",
          5465 => x"84802e99",
          5466 => x"3881760c",
          5467 => x"87c0928c",
          5468 => x"15537208",
          5469 => x"70820651",
          5470 => x"5271f738",
          5471 => x"ff19598d",
          5472 => x"39811a70",
          5473 => x"81ff0684",
          5474 => x"8019595b",
          5475 => x"5278802e",
          5476 => x"903873fc",
          5477 => x"80800652",
          5478 => x"7187387d",
          5479 => x"7a26fef8",
          5480 => x"3873fc80",
          5481 => x"80065271",
          5482 => x"802e8338",
          5483 => x"81527153",
          5484 => x"7282b5a8",
          5485 => x"0c8f3d0d",
          5486 => x"04fa3d0d",
          5487 => x"7a028405",
          5488 => x"a3053302",
          5489 => x"8805a705",
          5490 => x"33715454",
          5491 => x"5657fafe",
          5492 => x"3f82b5a8",
          5493 => x"08810653",
          5494 => x"83547280",
          5495 => x"fe38850b",
          5496 => x"87c0988c",
          5497 => x"0c815671",
          5498 => x"762e80dc",
          5499 => x"38717624",
          5500 => x"93387484",
          5501 => x"2b87c092",
          5502 => x"8c115454",
          5503 => x"71802e8d",
          5504 => x"3880d439",
          5505 => x"71832e80",
          5506 => x"c63880cb",
          5507 => x"39720870",
          5508 => x"812a7081",
          5509 => x"06515152",
          5510 => x"71802e8a",
          5511 => x"3887c098",
          5512 => x"8c085271",
          5513 => x"e83887c0",
          5514 => x"988c0852",
          5515 => x"71963881",
          5516 => x"730c87c0",
          5517 => x"928c1453",
          5518 => x"72087082",
          5519 => x"06515271",
          5520 => x"f7389639",
          5521 => x"80569239",
          5522 => x"88800a77",
          5523 => x"0c853981",
          5524 => x"80770c72",
          5525 => x"56833984",
          5526 => x"56755473",
          5527 => x"82b5a80c",
          5528 => x"883d0d04",
          5529 => x"fe3d0d74",
          5530 => x"81113371",
          5531 => x"3371882b",
          5532 => x"0782b5a8",
          5533 => x"0c535184",
          5534 => x"3d0d04fd",
          5535 => x"3d0d7583",
          5536 => x"11338212",
          5537 => x"3371902b",
          5538 => x"71882b07",
          5539 => x"81143370",
          5540 => x"7207882b",
          5541 => x"75337107",
          5542 => x"82b5a80c",
          5543 => x"52535456",
          5544 => x"5452853d",
          5545 => x"0d04ff3d",
          5546 => x"0d730284",
          5547 => x"05920522",
          5548 => x"52527072",
          5549 => x"70810554",
          5550 => x"3470882a",
          5551 => x"51707234",
          5552 => x"833d0d04",
          5553 => x"ff3d0d73",
          5554 => x"75525270",
          5555 => x"72708105",
          5556 => x"54347088",
          5557 => x"2a517072",
          5558 => x"70810554",
          5559 => x"3470882a",
          5560 => x"51707270",
          5561 => x"81055434",
          5562 => x"70882a51",
          5563 => x"70723483",
          5564 => x"3d0d04fe",
          5565 => x"3d0d7675",
          5566 => x"77545451",
          5567 => x"70802e92",
          5568 => x"38717081",
          5569 => x"05533373",
          5570 => x"70810555",
          5571 => x"34ff1151",
          5572 => x"eb39843d",
          5573 => x"0d04fe3d",
          5574 => x"0d757776",
          5575 => x"54525372",
          5576 => x"72708105",
          5577 => x"5434ff11",
          5578 => x"5170f438",
          5579 => x"843d0d04",
          5580 => x"fc3d0d78",
          5581 => x"77795656",
          5582 => x"53747081",
          5583 => x"05563374",
          5584 => x"70810556",
          5585 => x"33717131",
          5586 => x"ff165652",
          5587 => x"52527280",
          5588 => x"2e863871",
          5589 => x"802ee238",
          5590 => x"7182b5a8",
          5591 => x"0c863d0d",
          5592 => x"04fe3d0d",
          5593 => x"74765451",
          5594 => x"89397173",
          5595 => x"2e8a3881",
          5596 => x"11517033",
          5597 => x"5271f338",
          5598 => x"703382b5",
          5599 => x"a80c843d",
          5600 => x"0d04800b",
          5601 => x"82b5a80c",
          5602 => x"04800b82",
          5603 => x"b5a80c04",
          5604 => x"f73d0d7b",
          5605 => x"56800b83",
          5606 => x"1733565a",
          5607 => x"747a2e80",
          5608 => x"d6388154",
          5609 => x"b0160853",
          5610 => x"b4167053",
          5611 => x"81173352",
          5612 => x"59faa23f",
          5613 => x"82b5a808",
          5614 => x"7a2e0981",
          5615 => x"06b73882",
          5616 => x"b5a80883",
          5617 => x"1734b016",
          5618 => x"0870a418",
          5619 => x"08319c18",
          5620 => x"08595658",
          5621 => x"7477279f",
          5622 => x"38821633",
          5623 => x"5574822e",
          5624 => x"09810693",
          5625 => x"38815476",
          5626 => x"18537852",
          5627 => x"81163351",
          5628 => x"f9e33f83",
          5629 => x"39815a79",
          5630 => x"82b5a80c",
          5631 => x"8b3d0d04",
          5632 => x"fa3d0d78",
          5633 => x"7a565680",
          5634 => x"5774b017",
          5635 => x"082eaf38",
          5636 => x"7551fefc",
          5637 => x"3f82b5a8",
          5638 => x"085782b5",
          5639 => x"a8089f38",
          5640 => x"81547453",
          5641 => x"b4165281",
          5642 => x"163351f7",
          5643 => x"be3f82b5",
          5644 => x"a808802e",
          5645 => x"8538ff55",
          5646 => x"815774b0",
          5647 => x"170c7682",
          5648 => x"b5a80c88",
          5649 => x"3d0d04f8",
          5650 => x"3d0d7a70",
          5651 => x"5257fec0",
          5652 => x"3f82b5a8",
          5653 => x"085882b5",
          5654 => x"a8088191",
          5655 => x"38763355",
          5656 => x"74832e09",
          5657 => x"810680f0",
          5658 => x"38841733",
          5659 => x"5978812e",
          5660 => x"09810680",
          5661 => x"e3388480",
          5662 => x"5382b5a8",
          5663 => x"0852b417",
          5664 => x"705256fd",
          5665 => x"913f82d4",
          5666 => x"d55284b2",
          5667 => x"1751fc96",
          5668 => x"3f848b85",
          5669 => x"a4d25275",
          5670 => x"51fca93f",
          5671 => x"868a85e4",
          5672 => x"f2528498",
          5673 => x"1751fc9c",
          5674 => x"3f901708",
          5675 => x"52849c17",
          5676 => x"51fc913f",
          5677 => x"8c170852",
          5678 => x"84a01751",
          5679 => x"fc863fa0",
          5680 => x"17088105",
          5681 => x"70b0190c",
          5682 => x"79555375",
          5683 => x"52811733",
          5684 => x"51f8823f",
          5685 => x"77841834",
          5686 => x"80538052",
          5687 => x"81173351",
          5688 => x"f9d73f82",
          5689 => x"b5a80880",
          5690 => x"2e833881",
          5691 => x"587782b5",
          5692 => x"a80c8a3d",
          5693 => x"0d04fb3d",
          5694 => x"0d77fe1a",
          5695 => x"981208fe",
          5696 => x"05555654",
          5697 => x"80567473",
          5698 => x"278d388a",
          5699 => x"14227571",
          5700 => x"29ac1608",
          5701 => x"05575375",
          5702 => x"82b5a80c",
          5703 => x"873d0d04",
          5704 => x"f93d0d7a",
          5705 => x"7a700856",
          5706 => x"54578177",
          5707 => x"2781df38",
          5708 => x"76981508",
          5709 => x"2781d738",
          5710 => x"ff743354",
          5711 => x"5872822e",
          5712 => x"80f53872",
          5713 => x"82248938",
          5714 => x"72812e8d",
          5715 => x"3881bf39",
          5716 => x"72832e81",
          5717 => x"8e3881b6",
          5718 => x"3976812a",
          5719 => x"1770892a",
          5720 => x"a4160805",
          5721 => x"53745255",
          5722 => x"fd963f82",
          5723 => x"b5a80881",
          5724 => x"9f387483",
          5725 => x"ff0614b4",
          5726 => x"11338117",
          5727 => x"70892aa4",
          5728 => x"18080555",
          5729 => x"76545757",
          5730 => x"53fcf53f",
          5731 => x"82b5a808",
          5732 => x"80fe3874",
          5733 => x"83ff0614",
          5734 => x"b4113370",
          5735 => x"882b7807",
          5736 => x"79810671",
          5737 => x"842a5c52",
          5738 => x"58515372",
          5739 => x"80e23875",
          5740 => x"9fff0658",
          5741 => x"80da3976",
          5742 => x"882aa415",
          5743 => x"08055273",
          5744 => x"51fcbd3f",
          5745 => x"82b5a808",
          5746 => x"80c63876",
          5747 => x"1083fe06",
          5748 => x"7405b405",
          5749 => x"51f98d3f",
          5750 => x"82b5a808",
          5751 => x"83ffff06",
          5752 => x"58ae3976",
          5753 => x"872aa415",
          5754 => x"08055273",
          5755 => x"51fc913f",
          5756 => x"82b5a808",
          5757 => x"9b387682",
          5758 => x"2b83fc06",
          5759 => x"7405b405",
          5760 => x"51f8f83f",
          5761 => x"82b5a808",
          5762 => x"f00a0658",
          5763 => x"83398158",
          5764 => x"7782b5a8",
          5765 => x"0c893d0d",
          5766 => x"04f83d0d",
          5767 => x"7a7c7e5a",
          5768 => x"58568259",
          5769 => x"81772782",
          5770 => x"9e387698",
          5771 => x"17082782",
          5772 => x"96387533",
          5773 => x"5372792e",
          5774 => x"819d3872",
          5775 => x"79248938",
          5776 => x"72812e8d",
          5777 => x"38828039",
          5778 => x"72832e81",
          5779 => x"b83881f7",
          5780 => x"3976812a",
          5781 => x"1770892a",
          5782 => x"a4180805",
          5783 => x"53765255",
          5784 => x"fb9e3f82",
          5785 => x"b5a80859",
          5786 => x"82b5a808",
          5787 => x"81d93874",
          5788 => x"83ff0616",
          5789 => x"b4058116",
          5790 => x"78810659",
          5791 => x"56547753",
          5792 => x"76802e8f",
          5793 => x"3877842b",
          5794 => x"9ff00674",
          5795 => x"338f0671",
          5796 => x"07515372",
          5797 => x"7434810b",
          5798 => x"83173474",
          5799 => x"892aa417",
          5800 => x"08055275",
          5801 => x"51fad93f",
          5802 => x"82b5a808",
          5803 => x"5982b5a8",
          5804 => x"08819438",
          5805 => x"7483ff06",
          5806 => x"16b40578",
          5807 => x"842a5454",
          5808 => x"768f3877",
          5809 => x"882a7433",
          5810 => x"81f00671",
          5811 => x"8f060751",
          5812 => x"53727434",
          5813 => x"80ec3976",
          5814 => x"882aa417",
          5815 => x"08055275",
          5816 => x"51fa9d3f",
          5817 => x"82b5a808",
          5818 => x"5982b5a8",
          5819 => x"0880d838",
          5820 => x"7783ffff",
          5821 => x"06527610",
          5822 => x"83fe0676",
          5823 => x"05b40551",
          5824 => x"f7a43fbe",
          5825 => x"3976872a",
          5826 => x"a4170805",
          5827 => x"527551f9",
          5828 => x"ef3f82b5",
          5829 => x"a8085982",
          5830 => x"b5a808ab",
          5831 => x"3877f00a",
          5832 => x"0677822b",
          5833 => x"83fc0670",
          5834 => x"18b40570",
          5835 => x"54515454",
          5836 => x"f6c93f82",
          5837 => x"b5a8088f",
          5838 => x"0a067407",
          5839 => x"527251f7",
          5840 => x"833f810b",
          5841 => x"83173478",
          5842 => x"82b5a80c",
          5843 => x"8a3d0d04",
          5844 => x"f83d0d7a",
          5845 => x"7c7e7208",
          5846 => x"59565659",
          5847 => x"817527a4",
          5848 => x"38749817",
          5849 => x"08279d38",
          5850 => x"73802eaa",
          5851 => x"38ff5373",
          5852 => x"527551fd",
          5853 => x"a43f82b5",
          5854 => x"a8085482",
          5855 => x"b5a80880",
          5856 => x"f2389339",
          5857 => x"825480eb",
          5858 => x"39815480",
          5859 => x"e63982b5",
          5860 => x"a8085480",
          5861 => x"de397452",
          5862 => x"7851fb84",
          5863 => x"3f82b5a8",
          5864 => x"085882b5",
          5865 => x"a808802e",
          5866 => x"80c73882",
          5867 => x"b5a80881",
          5868 => x"2ed23882",
          5869 => x"b5a808ff",
          5870 => x"2ecf3880",
          5871 => x"53745275",
          5872 => x"51fcd63f",
          5873 => x"82b5a808",
          5874 => x"c5389816",
          5875 => x"08fe1190",
          5876 => x"18085755",
          5877 => x"57747427",
          5878 => x"90388115",
          5879 => x"90170c84",
          5880 => x"16338107",
          5881 => x"54738417",
          5882 => x"34775576",
          5883 => x"7826ffa6",
          5884 => x"38805473",
          5885 => x"82b5a80c",
          5886 => x"8a3d0d04",
          5887 => x"f63d0d7c",
          5888 => x"7e710859",
          5889 => x"5b5b7995",
          5890 => x"388c1708",
          5891 => x"5877802e",
          5892 => x"88389817",
          5893 => x"087826b2",
          5894 => x"388158ae",
          5895 => x"3979527a",
          5896 => x"51f9fd3f",
          5897 => x"81557482",
          5898 => x"b5a80827",
          5899 => x"82e03882",
          5900 => x"b5a80855",
          5901 => x"82b5a808",
          5902 => x"ff2e82d2",
          5903 => x"38981708",
          5904 => x"82b5a808",
          5905 => x"2682c738",
          5906 => x"79589017",
          5907 => x"08705654",
          5908 => x"73802e82",
          5909 => x"b938777a",
          5910 => x"2e098106",
          5911 => x"80e23881",
          5912 => x"1a569817",
          5913 => x"08762683",
          5914 => x"38825675",
          5915 => x"527a51f9",
          5916 => x"af3f8059",
          5917 => x"82b5a808",
          5918 => x"812e0981",
          5919 => x"06863882",
          5920 => x"b5a80859",
          5921 => x"82b5a808",
          5922 => x"09703070",
          5923 => x"72078025",
          5924 => x"707c0782",
          5925 => x"b5a80854",
          5926 => x"51515555",
          5927 => x"7381ef38",
          5928 => x"82b5a808",
          5929 => x"802e9538",
          5930 => x"8c170854",
          5931 => x"81742790",
          5932 => x"38739818",
          5933 => x"08278938",
          5934 => x"73588539",
          5935 => x"7580db38",
          5936 => x"77568116",
          5937 => x"56981708",
          5938 => x"76268938",
          5939 => x"82567578",
          5940 => x"2681ac38",
          5941 => x"75527a51",
          5942 => x"f8c63f82",
          5943 => x"b5a80880",
          5944 => x"2eb83880",
          5945 => x"5982b5a8",
          5946 => x"08812e09",
          5947 => x"81068638",
          5948 => x"82b5a808",
          5949 => x"5982b5a8",
          5950 => x"08097030",
          5951 => x"70720780",
          5952 => x"25707c07",
          5953 => x"51515555",
          5954 => x"7380f838",
          5955 => x"75782e09",
          5956 => x"8106ffae",
          5957 => x"38735580",
          5958 => x"f539ff53",
          5959 => x"75527651",
          5960 => x"f9f73f82",
          5961 => x"b5a80882",
          5962 => x"b5a80830",
          5963 => x"7082b5a8",
          5964 => x"08078025",
          5965 => x"51555579",
          5966 => x"802e9438",
          5967 => x"73802e8f",
          5968 => x"38755379",
          5969 => x"527651f9",
          5970 => x"d03f82b5",
          5971 => x"a8085574",
          5972 => x"a538758c",
          5973 => x"180c9817",
          5974 => x"08fe0590",
          5975 => x"18085654",
          5976 => x"74742686",
          5977 => x"38ff1590",
          5978 => x"180c8417",
          5979 => x"33810754",
          5980 => x"73841834",
          5981 => x"9739ff56",
          5982 => x"74812e90",
          5983 => x"388c3980",
          5984 => x"558c3982",
          5985 => x"b5a80855",
          5986 => x"85398156",
          5987 => x"75557482",
          5988 => x"b5a80c8c",
          5989 => x"3d0d04f8",
          5990 => x"3d0d7a70",
          5991 => x"5255f3f0",
          5992 => x"3f82b5a8",
          5993 => x"08588156",
          5994 => x"82b5a808",
          5995 => x"80d8387b",
          5996 => x"527451f6",
          5997 => x"c13f82b5",
          5998 => x"a80882b5",
          5999 => x"a808b017",
          6000 => x"0c598480",
          6001 => x"537752b4",
          6002 => x"15705257",
          6003 => x"f2c83f77",
          6004 => x"56843981",
          6005 => x"16568a15",
          6006 => x"22587578",
          6007 => x"27973881",
          6008 => x"54751953",
          6009 => x"76528115",
          6010 => x"3351ede9",
          6011 => x"3f82b5a8",
          6012 => x"08802edf",
          6013 => x"388a1522",
          6014 => x"76327030",
          6015 => x"70720770",
          6016 => x"9f2a5351",
          6017 => x"56567582",
          6018 => x"b5a80c8a",
          6019 => x"3d0d04f8",
          6020 => x"3d0d7a7c",
          6021 => x"71085856",
          6022 => x"5774f080",
          6023 => x"0a2680f1",
          6024 => x"38749f06",
          6025 => x"537280e9",
          6026 => x"38749018",
          6027 => x"0c881708",
          6028 => x"5473aa38",
          6029 => x"75335382",
          6030 => x"73278838",
          6031 => x"a8160854",
          6032 => x"739b3874",
          6033 => x"852a5382",
          6034 => x"0b881722",
          6035 => x"5a587279",
          6036 => x"2780fe38",
          6037 => x"a8160898",
          6038 => x"180c80cd",
          6039 => x"398a1622",
          6040 => x"70892b54",
          6041 => x"58727526",
          6042 => x"b2387352",
          6043 => x"7651f5b0",
          6044 => x"3f82b5a8",
          6045 => x"085482b5",
          6046 => x"a808ff2e",
          6047 => x"bd38810b",
          6048 => x"82b5a808",
          6049 => x"278b3898",
          6050 => x"160882b5",
          6051 => x"a8082685",
          6052 => x"388258bd",
          6053 => x"39747331",
          6054 => x"55cb3973",
          6055 => x"527551f4",
          6056 => x"d53f82b5",
          6057 => x"a8089818",
          6058 => x"0c739418",
          6059 => x"0c981708",
          6060 => x"53825872",
          6061 => x"802e9a38",
          6062 => x"85398158",
          6063 => x"94397489",
          6064 => x"2a139818",
          6065 => x"0c7483ff",
          6066 => x"0616b405",
          6067 => x"9c180c80",
          6068 => x"587782b5",
          6069 => x"a80c8a3d",
          6070 => x"0d04f83d",
          6071 => x"0d7a7008",
          6072 => x"901208a0",
          6073 => x"05595754",
          6074 => x"f0800a77",
          6075 => x"27863880",
          6076 => x"0b98150c",
          6077 => x"98140853",
          6078 => x"84557280",
          6079 => x"2e81cb38",
          6080 => x"7683ff06",
          6081 => x"587781b5",
          6082 => x"38811398",
          6083 => x"150c9414",
          6084 => x"08557492",
          6085 => x"3876852a",
          6086 => x"88172256",
          6087 => x"53747326",
          6088 => x"819b3880",
          6089 => x"c0398a16",
          6090 => x"22ff0577",
          6091 => x"892a0653",
          6092 => x"72818a38",
          6093 => x"74527351",
          6094 => x"f3e63f82",
          6095 => x"b5a80853",
          6096 => x"8255810b",
          6097 => x"82b5a808",
          6098 => x"2780ff38",
          6099 => x"815582b5",
          6100 => x"a808ff2e",
          6101 => x"80f43898",
          6102 => x"160882b5",
          6103 => x"a8082680",
          6104 => x"ca387b8a",
          6105 => x"38779815",
          6106 => x"0c845580",
          6107 => x"dd399414",
          6108 => x"08527351",
          6109 => x"f9863f82",
          6110 => x"b5a80853",
          6111 => x"875582b5",
          6112 => x"a808802e",
          6113 => x"80c43882",
          6114 => x"5582b5a8",
          6115 => x"08812eba",
          6116 => x"38815582",
          6117 => x"b5a808ff",
          6118 => x"2eb03882",
          6119 => x"b5a80852",
          6120 => x"7551fbf3",
          6121 => x"3f82b5a8",
          6122 => x"08a03872",
          6123 => x"94150c72",
          6124 => x"527551f2",
          6125 => x"c13f82b5",
          6126 => x"a8089815",
          6127 => x"0c769015",
          6128 => x"0c7716b4",
          6129 => x"059c150c",
          6130 => x"80557482",
          6131 => x"b5a80c8a",
          6132 => x"3d0d04f7",
          6133 => x"3d0d7b7d",
          6134 => x"71085b5b",
          6135 => x"57805276",
          6136 => x"51fcac3f",
          6137 => x"82b5a808",
          6138 => x"5482b5a8",
          6139 => x"0880ec38",
          6140 => x"82b5a808",
          6141 => x"56981708",
          6142 => x"527851f0",
          6143 => x"833f82b5",
          6144 => x"a8085482",
          6145 => x"b5a80880",
          6146 => x"d23882b5",
          6147 => x"a8089c18",
          6148 => x"08703351",
          6149 => x"54587281",
          6150 => x"e52e0981",
          6151 => x"06833881",
          6152 => x"5882b5a8",
          6153 => x"08557283",
          6154 => x"38815577",
          6155 => x"75075372",
          6156 => x"802e8e38",
          6157 => x"81165675",
          6158 => x"7a2e0981",
          6159 => x"068838a5",
          6160 => x"3982b5a8",
          6161 => x"08568152",
          6162 => x"7651fd8e",
          6163 => x"3f82b5a8",
          6164 => x"085482b5",
          6165 => x"a808802e",
          6166 => x"ff9b3873",
          6167 => x"842e0981",
          6168 => x"06833887",
          6169 => x"547382b5",
          6170 => x"a80c8b3d",
          6171 => x"0d04fd3d",
          6172 => x"0d769a11",
          6173 => x"5254ebec",
          6174 => x"3f82b5a8",
          6175 => x"0883ffff",
          6176 => x"06767033",
          6177 => x"51535371",
          6178 => x"832e0981",
          6179 => x"06903894",
          6180 => x"1451ebd0",
          6181 => x"3f82b5a8",
          6182 => x"08902b73",
          6183 => x"07537282",
          6184 => x"b5a80c85",
          6185 => x"3d0d04fc",
          6186 => x"3d0d7779",
          6187 => x"7083ffff",
          6188 => x"06549a12",
          6189 => x"535555eb",
          6190 => x"ed3f7670",
          6191 => x"33515372",
          6192 => x"832e0981",
          6193 => x"068b3873",
          6194 => x"902a5294",
          6195 => x"1551ebd6",
          6196 => x"3f863d0d",
          6197 => x"04f73d0d",
          6198 => x"7b7d5b55",
          6199 => x"8475085a",
          6200 => x"58981508",
          6201 => x"802e818a",
          6202 => x"38981508",
          6203 => x"527851ee",
          6204 => x"8f3f82b5",
          6205 => x"a8085882",
          6206 => x"b5a80880",
          6207 => x"f5389c15",
          6208 => x"08703355",
          6209 => x"53738638",
          6210 => x"845880e6",
          6211 => x"398b1333",
          6212 => x"70bf0670",
          6213 => x"81ff0658",
          6214 => x"51537286",
          6215 => x"163482b5",
          6216 => x"a8085373",
          6217 => x"81e52e83",
          6218 => x"38815373",
          6219 => x"ae2ea938",
          6220 => x"81707406",
          6221 => x"54577280",
          6222 => x"2e9e3875",
          6223 => x"8f2e9938",
          6224 => x"82b5a808",
          6225 => x"76df0654",
          6226 => x"5472882e",
          6227 => x"09810683",
          6228 => x"38765473",
          6229 => x"7a2ea038",
          6230 => x"80527451",
          6231 => x"fafc3f82",
          6232 => x"b5a80858",
          6233 => x"82b5a808",
          6234 => x"89389815",
          6235 => x"08fefa38",
          6236 => x"8639800b",
          6237 => x"98160c77",
          6238 => x"82b5a80c",
          6239 => x"8b3d0d04",
          6240 => x"fb3d0d77",
          6241 => x"70085754",
          6242 => x"81527351",
          6243 => x"fcc53f82",
          6244 => x"b5a80855",
          6245 => x"82b5a808",
          6246 => x"b4389814",
          6247 => x"08527551",
          6248 => x"ecde3f82",
          6249 => x"b5a80855",
          6250 => x"82b5a808",
          6251 => x"a038a053",
          6252 => x"82b5a808",
          6253 => x"529c1408",
          6254 => x"51eadb3f",
          6255 => x"8b53a014",
          6256 => x"529c1408",
          6257 => x"51eaac3f",
          6258 => x"810b8317",
          6259 => x"347482b5",
          6260 => x"a80c873d",
          6261 => x"0d04fd3d",
          6262 => x"0d757008",
          6263 => x"98120854",
          6264 => x"70535553",
          6265 => x"ec9a3f82",
          6266 => x"b5a8088d",
          6267 => x"389c1308",
          6268 => x"53e57334",
          6269 => x"810b8315",
          6270 => x"34853d0d",
          6271 => x"04fa3d0d",
          6272 => x"787a5757",
          6273 => x"800b8917",
          6274 => x"34981708",
          6275 => x"802e8182",
          6276 => x"38807089",
          6277 => x"18555555",
          6278 => x"9c170814",
          6279 => x"70338116",
          6280 => x"56515271",
          6281 => x"a02ea838",
          6282 => x"71852e09",
          6283 => x"81068438",
          6284 => x"81e55273",
          6285 => x"892e0981",
          6286 => x"068b38ae",
          6287 => x"73708105",
          6288 => x"55348115",
          6289 => x"55717370",
          6290 => x"81055534",
          6291 => x"8115558a",
          6292 => x"7427c538",
          6293 => x"75158805",
          6294 => x"52800b81",
          6295 => x"13349c17",
          6296 => x"08528b12",
          6297 => x"33881734",
          6298 => x"9c17089c",
          6299 => x"115252e8",
          6300 => x"8a3f82b5",
          6301 => x"a808760c",
          6302 => x"961251e7",
          6303 => x"e73f82b5",
          6304 => x"a8088617",
          6305 => x"23981251",
          6306 => x"e7da3f82",
          6307 => x"b5a80884",
          6308 => x"1723883d",
          6309 => x"0d04f33d",
          6310 => x"0d7f7008",
          6311 => x"5e5b8061",
          6312 => x"70335155",
          6313 => x"5573af2e",
          6314 => x"83388155",
          6315 => x"7380dc2e",
          6316 => x"91387480",
          6317 => x"2e8c3894",
          6318 => x"1d08881c",
          6319 => x"0caa3981",
          6320 => x"15418061",
          6321 => x"70335656",
          6322 => x"5673af2e",
          6323 => x"09810683",
          6324 => x"38815673",
          6325 => x"80dc3270",
          6326 => x"30708025",
          6327 => x"78075151",
          6328 => x"5473dc38",
          6329 => x"73881c0c",
          6330 => x"60703351",
          6331 => x"54739f26",
          6332 => x"9638ff80",
          6333 => x"0bab1c34",
          6334 => x"80527a51",
          6335 => x"f6913f82",
          6336 => x"b5a80855",
          6337 => x"85983991",
          6338 => x"3d61a01d",
          6339 => x"5c5a5e8b",
          6340 => x"53a05279",
          6341 => x"51e7ff3f",
          6342 => x"80705957",
          6343 => x"88793355",
          6344 => x"5c73ae2e",
          6345 => x"09810680",
          6346 => x"d4387818",
          6347 => x"7033811a",
          6348 => x"71ae3270",
          6349 => x"30709f2a",
          6350 => x"73822607",
          6351 => x"5151535a",
          6352 => x"5754738c",
          6353 => x"38791754",
          6354 => x"75743481",
          6355 => x"1757db39",
          6356 => x"75af3270",
          6357 => x"30709f2a",
          6358 => x"51515475",
          6359 => x"80dc2e8c",
          6360 => x"3873802e",
          6361 => x"873875a0",
          6362 => x"2682bd38",
          6363 => x"77197e0c",
          6364 => x"a454a076",
          6365 => x"2782bd38",
          6366 => x"a05482b8",
          6367 => x"39781870",
          6368 => x"33811a5a",
          6369 => x"5754a076",
          6370 => x"2781fc38",
          6371 => x"75af3270",
          6372 => x"307780dc",
          6373 => x"32703072",
          6374 => x"80257180",
          6375 => x"25075151",
          6376 => x"56515573",
          6377 => x"802eac38",
          6378 => x"84398118",
          6379 => x"5880781a",
          6380 => x"70335155",
          6381 => x"5573af2e",
          6382 => x"09810683",
          6383 => x"38815573",
          6384 => x"80dc3270",
          6385 => x"30708025",
          6386 => x"77075151",
          6387 => x"5473db38",
          6388 => x"81b53975",
          6389 => x"ae2e0981",
          6390 => x"06833881",
          6391 => x"54767c27",
          6392 => x"74075473",
          6393 => x"802ea238",
          6394 => x"7b8b3270",
          6395 => x"3077ae32",
          6396 => x"70307280",
          6397 => x"25719f2a",
          6398 => x"07535156",
          6399 => x"51557481",
          6400 => x"a7388857",
          6401 => x"8b5cfef5",
          6402 => x"3975982b",
          6403 => x"54738025",
          6404 => x"8c387580",
          6405 => x"ff0682ae",
          6406 => x"f0113357",
          6407 => x"547551e6",
          6408 => x"e13f82b5",
          6409 => x"a808802e",
          6410 => x"b2387818",
          6411 => x"7033811a",
          6412 => x"71545a56",
          6413 => x"54e6d23f",
          6414 => x"82b5a808",
          6415 => x"802e80e8",
          6416 => x"38ff1c54",
          6417 => x"76742780",
          6418 => x"df387917",
          6419 => x"54757434",
          6420 => x"81177a11",
          6421 => x"55577474",
          6422 => x"34a73975",
          6423 => x"5282ae90",
          6424 => x"51e5fe3f",
          6425 => x"82b5a808",
          6426 => x"bf38ff9f",
          6427 => x"16547399",
          6428 => x"268938e0",
          6429 => x"167081ff",
          6430 => x"06575479",
          6431 => x"17547574",
          6432 => x"34811757",
          6433 => x"fdf73977",
          6434 => x"197e0c76",
          6435 => x"802e9938",
          6436 => x"79335473",
          6437 => x"81e52e09",
          6438 => x"81068438",
          6439 => x"857a3484",
          6440 => x"54a07627",
          6441 => x"8f388b39",
          6442 => x"865581f2",
          6443 => x"39845680",
          6444 => x"f3398054",
          6445 => x"738b1b34",
          6446 => x"807b0858",
          6447 => x"527a51f2",
          6448 => x"ce3f82b5",
          6449 => x"a8085682",
          6450 => x"b5a80880",
          6451 => x"d738981b",
          6452 => x"08527651",
          6453 => x"e6aa3f82",
          6454 => x"b5a80856",
          6455 => x"82b5a808",
          6456 => x"80c2389c",
          6457 => x"1b087033",
          6458 => x"55557380",
          6459 => x"2effbe38",
          6460 => x"8b1533bf",
          6461 => x"06547386",
          6462 => x"1c348b15",
          6463 => x"3370832a",
          6464 => x"70810651",
          6465 => x"55587392",
          6466 => x"388b5379",
          6467 => x"527451e4",
          6468 => x"9f3f82b5",
          6469 => x"a808802e",
          6470 => x"8b387552",
          6471 => x"7a51f3ba",
          6472 => x"3fff9f39",
          6473 => x"75ab1c33",
          6474 => x"57557480",
          6475 => x"2ebb3874",
          6476 => x"842e0981",
          6477 => x"0680e738",
          6478 => x"75852a70",
          6479 => x"81067782",
          6480 => x"2a585154",
          6481 => x"73802e96",
          6482 => x"38758106",
          6483 => x"5473802e",
          6484 => x"fbb538ff",
          6485 => x"800bab1c",
          6486 => x"34805580",
          6487 => x"c1397581",
          6488 => x"065473ba",
          6489 => x"388555b6",
          6490 => x"3975822a",
          6491 => x"70810651",
          6492 => x"5473ab38",
          6493 => x"861b3370",
          6494 => x"842a7081",
          6495 => x"06515555",
          6496 => x"73802ee1",
          6497 => x"38901b08",
          6498 => x"83ff061d",
          6499 => x"b405527c",
          6500 => x"51f5db3f",
          6501 => x"82b5a808",
          6502 => x"881c0cfa",
          6503 => x"ea397482",
          6504 => x"b5a80c8f",
          6505 => x"3d0d04f6",
          6506 => x"3d0d7c5b",
          6507 => x"ff7b0870",
          6508 => x"71735559",
          6509 => x"5c555973",
          6510 => x"802e81c6",
          6511 => x"38757081",
          6512 => x"05573370",
          6513 => x"a0265252",
          6514 => x"71ba2e8d",
          6515 => x"3870ee38",
          6516 => x"71ba2e09",
          6517 => x"810681a5",
          6518 => x"387333d0",
          6519 => x"117081ff",
          6520 => x"06515253",
          6521 => x"70892691",
          6522 => x"38821473",
          6523 => x"81ff06d0",
          6524 => x"05565271",
          6525 => x"762e80f7",
          6526 => x"38800b82",
          6527 => x"aee05955",
          6528 => x"77087a55",
          6529 => x"57767081",
          6530 => x"05583374",
          6531 => x"70810556",
          6532 => x"33ff9f12",
          6533 => x"53535370",
          6534 => x"99268938",
          6535 => x"e0137081",
          6536 => x"ff065451",
          6537 => x"ff9f1251",
          6538 => x"70992689",
          6539 => x"38e01270",
          6540 => x"81ff0653",
          6541 => x"51723070",
          6542 => x"9f2a5151",
          6543 => x"72722e09",
          6544 => x"81068538",
          6545 => x"70ffbe38",
          6546 => x"72307477",
          6547 => x"32703070",
          6548 => x"72079f2a",
          6549 => x"739f2a07",
          6550 => x"53545451",
          6551 => x"70802e8f",
          6552 => x"38811584",
          6553 => x"19595583",
          6554 => x"7525ff94",
          6555 => x"388b3974",
          6556 => x"83248638",
          6557 => x"74767c0c",
          6558 => x"59785186",
          6559 => x"3982ccf4",
          6560 => x"33517082",
          6561 => x"b5a80c8c",
          6562 => x"3d0d04fa",
          6563 => x"3d0d7856",
          6564 => x"800b8317",
          6565 => x"34ff0bb0",
          6566 => x"170c7952",
          6567 => x"7551e2e0",
          6568 => x"3f845582",
          6569 => x"b5a80881",
          6570 => x"803884b2",
          6571 => x"1651dfb4",
          6572 => x"3f82b5a8",
          6573 => x"0883ffff",
          6574 => x"06548355",
          6575 => x"7382d4d5",
          6576 => x"2e098106",
          6577 => x"80e33880",
          6578 => x"0bb41733",
          6579 => x"56577481",
          6580 => x"e92e0981",
          6581 => x"06833881",
          6582 => x"577481eb",
          6583 => x"32703070",
          6584 => x"80257907",
          6585 => x"51515473",
          6586 => x"8a387481",
          6587 => x"e82e0981",
          6588 => x"06b53883",
          6589 => x"5382aea0",
          6590 => x"5280ea16",
          6591 => x"51e0b13f",
          6592 => x"82b5a808",
          6593 => x"5582b5a8",
          6594 => x"08802e9d",
          6595 => x"38855382",
          6596 => x"aea45281",
          6597 => x"861651e0",
          6598 => x"973f82b5",
          6599 => x"a8085582",
          6600 => x"b5a80880",
          6601 => x"2e833882",
          6602 => x"557482b5",
          6603 => x"a80c883d",
          6604 => x"0d04f23d",
          6605 => x"0d610284",
          6606 => x"0580cb05",
          6607 => x"33585580",
          6608 => x"750c6051",
          6609 => x"fce13f82",
          6610 => x"b5a80858",
          6611 => x"8b56800b",
          6612 => x"82b5a808",
          6613 => x"2486fc38",
          6614 => x"82b5a808",
          6615 => x"842982cc",
          6616 => x"e0057008",
          6617 => x"55538c56",
          6618 => x"73802e86",
          6619 => x"e6387375",
          6620 => x"0c7681fe",
          6621 => x"06743354",
          6622 => x"5772802e",
          6623 => x"ae388114",
          6624 => x"3351d7ca",
          6625 => x"3f82b5a8",
          6626 => x"0881ff06",
          6627 => x"70810654",
          6628 => x"55729838",
          6629 => x"76802e86",
          6630 => x"b8387482",
          6631 => x"2a708106",
          6632 => x"51538a56",
          6633 => x"7286ac38",
          6634 => x"86a73980",
          6635 => x"74347781",
          6636 => x"15348152",
          6637 => x"81143351",
          6638 => x"d7b23f82",
          6639 => x"b5a80881",
          6640 => x"ff067081",
          6641 => x"06545583",
          6642 => x"56728687",
          6643 => x"3876802e",
          6644 => x"8f387482",
          6645 => x"2a708106",
          6646 => x"51538a56",
          6647 => x"7285f438",
          6648 => x"80705374",
          6649 => x"525bfda3",
          6650 => x"3f82b5a8",
          6651 => x"0881ff06",
          6652 => x"5776822e",
          6653 => x"09810680",
          6654 => x"e2388c3d",
          6655 => x"74565883",
          6656 => x"5683f615",
          6657 => x"33705853",
          6658 => x"72802e8d",
          6659 => x"3883fa15",
          6660 => x"51dce83f",
          6661 => x"82b5a808",
          6662 => x"57767870",
          6663 => x"84055a0c",
          6664 => x"ff169016",
          6665 => x"56567580",
          6666 => x"25d73880",
          6667 => x"0b8d3d54",
          6668 => x"56727084",
          6669 => x"0554085b",
          6670 => x"83577a80",
          6671 => x"2e95387a",
          6672 => x"527351fc",
          6673 => x"c63f82b5",
          6674 => x"a80881ff",
          6675 => x"06578177",
          6676 => x"27893881",
          6677 => x"16568376",
          6678 => x"27d73881",
          6679 => x"5676842e",
          6680 => x"84f1388d",
          6681 => x"56768126",
          6682 => x"84e938bf",
          6683 => x"1451dbf4",
          6684 => x"3f82b5a8",
          6685 => x"0883ffff",
          6686 => x"06537284",
          6687 => x"802e0981",
          6688 => x"0684d038",
          6689 => x"80ca1451",
          6690 => x"dbda3f82",
          6691 => x"b5a80883",
          6692 => x"ffff0658",
          6693 => x"778d3880",
          6694 => x"d81451db",
          6695 => x"de3f82b5",
          6696 => x"a8085877",
          6697 => x"9c150c80",
          6698 => x"c4143382",
          6699 => x"153480c4",
          6700 => x"1433ff11",
          6701 => x"7081ff06",
          6702 => x"5154558d",
          6703 => x"56728126",
          6704 => x"84913874",
          6705 => x"81ff0678",
          6706 => x"712980c1",
          6707 => x"16335259",
          6708 => x"53728a15",
          6709 => x"2372802e",
          6710 => x"8b38ff13",
          6711 => x"73065372",
          6712 => x"802e8638",
          6713 => x"8d5683eb",
          6714 => x"3980c514",
          6715 => x"51daf53f",
          6716 => x"82b5a808",
          6717 => x"5382b5a8",
          6718 => x"08881523",
          6719 => x"728f0657",
          6720 => x"8d567683",
          6721 => x"ce3880c7",
          6722 => x"1451dad8",
          6723 => x"3f82b5a8",
          6724 => x"0883ffff",
          6725 => x"0655748d",
          6726 => x"3880d414",
          6727 => x"51dadc3f",
          6728 => x"82b5a808",
          6729 => x"5580c214",
          6730 => x"51dab93f",
          6731 => x"82b5a808",
          6732 => x"83ffff06",
          6733 => x"538d5672",
          6734 => x"802e8397",
          6735 => x"38881422",
          6736 => x"78147184",
          6737 => x"2a055a5a",
          6738 => x"78752683",
          6739 => x"86388a14",
          6740 => x"22527479",
          6741 => x"3151feff",
          6742 => x"ca3f82b5",
          6743 => x"a8085582",
          6744 => x"b5a80880",
          6745 => x"2e82ec38",
          6746 => x"82b5a808",
          6747 => x"80ffffff",
          6748 => x"f5268338",
          6749 => x"83577483",
          6750 => x"fff52683",
          6751 => x"38825774",
          6752 => x"9ff52685",
          6753 => x"38815789",
          6754 => x"398d5676",
          6755 => x"802e82c3",
          6756 => x"38821570",
          6757 => x"98160c7b",
          6758 => x"a0160c73",
          6759 => x"1c70a417",
          6760 => x"0c7a1dac",
          6761 => x"170c5455",
          6762 => x"76832e09",
          6763 => x"8106af38",
          6764 => x"80de1451",
          6765 => x"d9ae3f82",
          6766 => x"b5a80883",
          6767 => x"ffff0653",
          6768 => x"8d567282",
          6769 => x"8e387982",
          6770 => x"8a3880e0",
          6771 => x"1451d9ab",
          6772 => x"3f82b5a8",
          6773 => x"08a8150c",
          6774 => x"74822b53",
          6775 => x"a2398d56",
          6776 => x"79802e81",
          6777 => x"ee387713",
          6778 => x"a8150c74",
          6779 => x"15537682",
          6780 => x"2e8d3874",
          6781 => x"10157081",
          6782 => x"2a768106",
          6783 => x"05515383",
          6784 => x"ff13892a",
          6785 => x"538d5672",
          6786 => x"9c150826",
          6787 => x"81c538ff",
          6788 => x"0b90150c",
          6789 => x"ff0b8c15",
          6790 => x"0cff800b",
          6791 => x"84153476",
          6792 => x"832e0981",
          6793 => x"06819238",
          6794 => x"80e41451",
          6795 => x"d8b63f82",
          6796 => x"b5a80883",
          6797 => x"ffff0653",
          6798 => x"72812e09",
          6799 => x"810680f9",
          6800 => x"38811b52",
          6801 => x"7351dbb8",
          6802 => x"3f82b5a8",
          6803 => x"0880ea38",
          6804 => x"82b5a808",
          6805 => x"84153484",
          6806 => x"b21451d8",
          6807 => x"873f82b5",
          6808 => x"a80883ff",
          6809 => x"ff065372",
          6810 => x"82d4d52e",
          6811 => x"09810680",
          6812 => x"c838b414",
          6813 => x"51d8843f",
          6814 => x"82b5a808",
          6815 => x"848b85a4",
          6816 => x"d22e0981",
          6817 => x"06b33884",
          6818 => x"981451d7",
          6819 => x"ee3f82b5",
          6820 => x"a808868a",
          6821 => x"85e4f22e",
          6822 => x"0981069d",
          6823 => x"38849c14",
          6824 => x"51d7d83f",
          6825 => x"82b5a808",
          6826 => x"90150c84",
          6827 => x"a01451d7",
          6828 => x"ca3f82b5",
          6829 => x"a8088c15",
          6830 => x"0c767434",
          6831 => x"82ccf022",
          6832 => x"81055372",
          6833 => x"82ccf023",
          6834 => x"72861523",
          6835 => x"800b9415",
          6836 => x"0c805675",
          6837 => x"82b5a80c",
          6838 => x"903d0d04",
          6839 => x"fb3d0d77",
          6840 => x"54895573",
          6841 => x"802eb938",
          6842 => x"73085372",
          6843 => x"802eb138",
          6844 => x"72335271",
          6845 => x"802ea938",
          6846 => x"86132284",
          6847 => x"15225752",
          6848 => x"71762e09",
          6849 => x"81069938",
          6850 => x"81133351",
          6851 => x"d0c03f82",
          6852 => x"b5a80881",
          6853 => x"06527188",
          6854 => x"38717408",
          6855 => x"54558339",
          6856 => x"80537873",
          6857 => x"710c5274",
          6858 => x"82b5a80c",
          6859 => x"873d0d04",
          6860 => x"fa3d0d02",
          6861 => x"ab05337a",
          6862 => x"58893dfc",
          6863 => x"055256f4",
          6864 => x"e63f8b54",
          6865 => x"800b82b5",
          6866 => x"a80824bc",
          6867 => x"3882b5a8",
          6868 => x"08842982",
          6869 => x"cce00570",
          6870 => x"08555573",
          6871 => x"802e8438",
          6872 => x"80743478",
          6873 => x"5473802e",
          6874 => x"84388074",
          6875 => x"3478750c",
          6876 => x"75547580",
          6877 => x"2e923880",
          6878 => x"53893d70",
          6879 => x"53840551",
          6880 => x"f7b03f82",
          6881 => x"b5a80854",
          6882 => x"7382b5a8",
          6883 => x"0c883d0d",
          6884 => x"04eb3d0d",
          6885 => x"67028405",
          6886 => x"80e70533",
          6887 => x"59598954",
          6888 => x"78802e84",
          6889 => x"c83877bf",
          6890 => x"06705498",
          6891 => x"3dd00553",
          6892 => x"993d8405",
          6893 => x"5258f6fa",
          6894 => x"3f82b5a8",
          6895 => x"085582b5",
          6896 => x"a80884a4",
          6897 => x"387a5c68",
          6898 => x"528c3d70",
          6899 => x"5256edc6",
          6900 => x"3f82b5a8",
          6901 => x"085582b5",
          6902 => x"a8089238",
          6903 => x"0280d705",
          6904 => x"3370982b",
          6905 => x"55577380",
          6906 => x"25833886",
          6907 => x"55779c06",
          6908 => x"5473802e",
          6909 => x"81ab3874",
          6910 => x"802e9538",
          6911 => x"74842e09",
          6912 => x"8106aa38",
          6913 => x"7551eaf8",
          6914 => x"3f82b5a8",
          6915 => x"08559e39",
          6916 => x"02b20533",
          6917 => x"91065473",
          6918 => x"81b83877",
          6919 => x"822a7081",
          6920 => x"06515473",
          6921 => x"802e8e38",
          6922 => x"885583bc",
          6923 => x"39778807",
          6924 => x"587483b4",
          6925 => x"3877832a",
          6926 => x"70810651",
          6927 => x"5473802e",
          6928 => x"81af3862",
          6929 => x"527a51e8",
          6930 => x"a53f82b5",
          6931 => x"a8085682",
          6932 => x"88b20a52",
          6933 => x"628e0551",
          6934 => x"d4ea3f62",
          6935 => x"54a00b8b",
          6936 => x"15348053",
          6937 => x"62527a51",
          6938 => x"e8bd3f80",
          6939 => x"52629c05",
          6940 => x"51d4d13f",
          6941 => x"7a54810b",
          6942 => x"83153475",
          6943 => x"802e80f1",
          6944 => x"387ab011",
          6945 => x"08515480",
          6946 => x"53755297",
          6947 => x"3dd40551",
          6948 => x"ddbe3f82",
          6949 => x"b5a80855",
          6950 => x"82b5a808",
          6951 => x"82ca38b7",
          6952 => x"397482c4",
          6953 => x"3802b205",
          6954 => x"3370842a",
          6955 => x"70810651",
          6956 => x"55567380",
          6957 => x"2e863884",
          6958 => x"5582ad39",
          6959 => x"77812a70",
          6960 => x"81065154",
          6961 => x"73802ea9",
          6962 => x"38758106",
          6963 => x"5473802e",
          6964 => x"a0388755",
          6965 => x"82923973",
          6966 => x"527a51d6",
          6967 => x"a33f82b5",
          6968 => x"a8087bff",
          6969 => x"188c120c",
          6970 => x"555582b5",
          6971 => x"a80881f8",
          6972 => x"3877832a",
          6973 => x"70810651",
          6974 => x"5473802e",
          6975 => x"86387780",
          6976 => x"c007587a",
          6977 => x"b01108a0",
          6978 => x"1b0c63a4",
          6979 => x"1b0c6353",
          6980 => x"705257e6",
          6981 => x"d93f82b5",
          6982 => x"a80882b5",
          6983 => x"a808881b",
          6984 => x"0c639c05",
          6985 => x"525ad2d3",
          6986 => x"3f82b5a8",
          6987 => x"0882b5a8",
          6988 => x"088c1b0c",
          6989 => x"777a0c56",
          6990 => x"86172284",
          6991 => x"1a237790",
          6992 => x"1a34800b",
          6993 => x"911a3480",
          6994 => x"0b9c1a0c",
          6995 => x"800b941a",
          6996 => x"0c77852a",
          6997 => x"70810651",
          6998 => x"5473802e",
          6999 => x"818d3882",
          7000 => x"b5a80880",
          7001 => x"2e818438",
          7002 => x"82b5a808",
          7003 => x"941a0c8a",
          7004 => x"17227089",
          7005 => x"2b7b5259",
          7006 => x"57a83976",
          7007 => x"527851d7",
          7008 => x"9f3f82b5",
          7009 => x"a8085782",
          7010 => x"b5a80881",
          7011 => x"26833882",
          7012 => x"5582b5a8",
          7013 => x"08ff2e09",
          7014 => x"81068338",
          7015 => x"79557578",
          7016 => x"31567430",
          7017 => x"70760780",
          7018 => x"25515477",
          7019 => x"76278a38",
          7020 => x"81707506",
          7021 => x"555a73c3",
          7022 => x"3876981a",
          7023 => x"0c74a938",
          7024 => x"7583ff06",
          7025 => x"5473802e",
          7026 => x"a2387652",
          7027 => x"7a51d6a6",
          7028 => x"3f82b5a8",
          7029 => x"08853882",
          7030 => x"558e3975",
          7031 => x"892a82b5",
          7032 => x"a808059c",
          7033 => x"1a0c8439",
          7034 => x"80790c74",
          7035 => x"547382b5",
          7036 => x"a80c973d",
          7037 => x"0d04f23d",
          7038 => x"0d606365",
          7039 => x"6440405d",
          7040 => x"59807e0c",
          7041 => x"903dfc05",
          7042 => x"527851f9",
          7043 => x"cf3f82b5",
          7044 => x"a8085582",
          7045 => x"b5a8088a",
          7046 => x"38911933",
          7047 => x"5574802e",
          7048 => x"86387456",
          7049 => x"82c43990",
          7050 => x"19338106",
          7051 => x"55875674",
          7052 => x"802e82b6",
          7053 => x"38953982",
          7054 => x"0b911a34",
          7055 => x"825682aa",
          7056 => x"39810b91",
          7057 => x"1a348156",
          7058 => x"82a0398c",
          7059 => x"1908941a",
          7060 => x"08315574",
          7061 => x"7c278338",
          7062 => x"745c7b80",
          7063 => x"2e828938",
          7064 => x"94190870",
          7065 => x"83ff0656",
          7066 => x"567481b2",
          7067 => x"387e8a11",
          7068 => x"22ff0577",
          7069 => x"892a065b",
          7070 => x"5579a838",
          7071 => x"75873888",
          7072 => x"1908558f",
          7073 => x"39981908",
          7074 => x"527851d5",
          7075 => x"933f82b5",
          7076 => x"a8085581",
          7077 => x"7527ff9f",
          7078 => x"3874ff2e",
          7079 => x"ffa33874",
          7080 => x"981a0c98",
          7081 => x"1908527e",
          7082 => x"51d4cb3f",
          7083 => x"82b5a808",
          7084 => x"802eff83",
          7085 => x"3882b5a8",
          7086 => x"081a7c89",
          7087 => x"2a595777",
          7088 => x"802e80d6",
          7089 => x"38771a7f",
          7090 => x"8a112258",
          7091 => x"5c557575",
          7092 => x"27853875",
          7093 => x"7a315877",
          7094 => x"5476537c",
          7095 => x"52811b33",
          7096 => x"51ca883f",
          7097 => x"82b5a808",
          7098 => x"fed7387e",
          7099 => x"83113356",
          7100 => x"5674802e",
          7101 => x"9f38b016",
          7102 => x"08773155",
          7103 => x"74782794",
          7104 => x"38848053",
          7105 => x"b41652b0",
          7106 => x"16087731",
          7107 => x"892b7d05",
          7108 => x"51cfe03f",
          7109 => x"77892b56",
          7110 => x"b939769c",
          7111 => x"1a0c9419",
          7112 => x"0883ff06",
          7113 => x"84807131",
          7114 => x"57557b76",
          7115 => x"2783387b",
          7116 => x"569c1908",
          7117 => x"527e51d1",
          7118 => x"c73f82b5",
          7119 => x"a808fe81",
          7120 => x"38755394",
          7121 => x"190883ff",
          7122 => x"061fb405",
          7123 => x"527c51cf",
          7124 => x"a23f7b76",
          7125 => x"317e0817",
          7126 => x"7f0c761e",
          7127 => x"941b0818",
          7128 => x"941c0c5e",
          7129 => x"5cfdf339",
          7130 => x"80567582",
          7131 => x"b5a80c90",
          7132 => x"3d0d04f2",
          7133 => x"3d0d6063",
          7134 => x"65644040",
          7135 => x"5d58807e",
          7136 => x"0c903dfc",
          7137 => x"05527751",
          7138 => x"f6d23f82",
          7139 => x"b5a80855",
          7140 => x"82b5a808",
          7141 => x"8a389118",
          7142 => x"33557480",
          7143 => x"2e863874",
          7144 => x"5683b839",
          7145 => x"90183370",
          7146 => x"812a7081",
          7147 => x"06515656",
          7148 => x"87567480",
          7149 => x"2e83a438",
          7150 => x"9539820b",
          7151 => x"91193482",
          7152 => x"56839839",
          7153 => x"810b9119",
          7154 => x"34815683",
          7155 => x"8e399418",
          7156 => x"087c1156",
          7157 => x"56747627",
          7158 => x"84387509",
          7159 => x"5c7b802e",
          7160 => x"82ec3894",
          7161 => x"18087083",
          7162 => x"ff065656",
          7163 => x"7481fd38",
          7164 => x"7e8a1122",
          7165 => x"ff057789",
          7166 => x"2a065c55",
          7167 => x"7abf3875",
          7168 => x"8c388818",
          7169 => x"0855749c",
          7170 => x"387a5285",
          7171 => x"39981808",
          7172 => x"527751d7",
          7173 => x"e73f82b5",
          7174 => x"a8085582",
          7175 => x"b5a80880",
          7176 => x"2e82ab38",
          7177 => x"74812eff",
          7178 => x"913874ff",
          7179 => x"2eff9538",
          7180 => x"7498190c",
          7181 => x"88180885",
          7182 => x"38748819",
          7183 => x"0c7e55b0",
          7184 => x"15089c19",
          7185 => x"082e0981",
          7186 => x"068d3874",
          7187 => x"51cec13f",
          7188 => x"82b5a808",
          7189 => x"feee3898",
          7190 => x"1808527e",
          7191 => x"51d1973f",
          7192 => x"82b5a808",
          7193 => x"802efed2",
          7194 => x"3882b5a8",
          7195 => x"081b7c89",
          7196 => x"2a5a5778",
          7197 => x"802e80d5",
          7198 => x"38781b7f",
          7199 => x"8a112258",
          7200 => x"5b557575",
          7201 => x"27853875",
          7202 => x"7b315978",
          7203 => x"5476537c",
          7204 => x"52811a33",
          7205 => x"51c8be3f",
          7206 => x"82b5a808",
          7207 => x"fea6387e",
          7208 => x"b0110878",
          7209 => x"31565674",
          7210 => x"79279b38",
          7211 => x"848053b0",
          7212 => x"16087731",
          7213 => x"892b7d05",
          7214 => x"52b41651",
          7215 => x"ccb53f7e",
          7216 => x"55800b83",
          7217 => x"16347889",
          7218 => x"2b5680db",
          7219 => x"398c1808",
          7220 => x"94190826",
          7221 => x"93387e51",
          7222 => x"cdb63f82",
          7223 => x"b5a808fd",
          7224 => x"e3387e77",
          7225 => x"b0120c55",
          7226 => x"769c190c",
          7227 => x"94180883",
          7228 => x"ff068480",
          7229 => x"71315755",
          7230 => x"7b762783",
          7231 => x"387b569c",
          7232 => x"1808527e",
          7233 => x"51cdf93f",
          7234 => x"82b5a808",
          7235 => x"fdb63875",
          7236 => x"537c5294",
          7237 => x"180883ff",
          7238 => x"061fb405",
          7239 => x"51cbd43f",
          7240 => x"7e55810b",
          7241 => x"8316347b",
          7242 => x"76317e08",
          7243 => x"177f0c76",
          7244 => x"1e941a08",
          7245 => x"1870941c",
          7246 => x"0c8c1b08",
          7247 => x"58585e5c",
          7248 => x"74762783",
          7249 => x"38755574",
          7250 => x"8c190cfd",
          7251 => x"90399018",
          7252 => x"3380c007",
          7253 => x"55749019",
          7254 => x"34805675",
          7255 => x"82b5a80c",
          7256 => x"903d0d04",
          7257 => x"f83d0d7a",
          7258 => x"8b3dfc05",
          7259 => x"53705256",
          7260 => x"f2ea3f82",
          7261 => x"b5a80857",
          7262 => x"82b5a808",
          7263 => x"80fb3890",
          7264 => x"16337086",
          7265 => x"2a708106",
          7266 => x"51555573",
          7267 => x"802e80e9",
          7268 => x"38a01608",
          7269 => x"527851cc",
          7270 => x"e73f82b5",
          7271 => x"a8085782",
          7272 => x"b5a80880",
          7273 => x"d438a416",
          7274 => x"088b1133",
          7275 => x"a0075555",
          7276 => x"738b1634",
          7277 => x"88160853",
          7278 => x"74527508",
          7279 => x"51dde83f",
          7280 => x"8c160852",
          7281 => x"9c1551c9",
          7282 => x"fb3f8288",
          7283 => x"b20a5296",
          7284 => x"1551c9f0",
          7285 => x"3f765292",
          7286 => x"1551c9ca",
          7287 => x"3f785481",
          7288 => x"0b831534",
          7289 => x"7851ccdf",
          7290 => x"3f82b5a8",
          7291 => x"08901733",
          7292 => x"81bf0655",
          7293 => x"57739017",
          7294 => x"347682b5",
          7295 => x"a80c8a3d",
          7296 => x"0d04fc3d",
          7297 => x"0d767052",
          7298 => x"54fed93f",
          7299 => x"82b5a808",
          7300 => x"5382b5a8",
          7301 => x"089c3886",
          7302 => x"3dfc0552",
          7303 => x"7351f1bc",
          7304 => x"3f82b5a8",
          7305 => x"085382b5",
          7306 => x"a8088738",
          7307 => x"82b5a808",
          7308 => x"740c7282",
          7309 => x"b5a80c86",
          7310 => x"3d0d04ff",
          7311 => x"3d0d843d",
          7312 => x"51e6e43f",
          7313 => x"8b52800b",
          7314 => x"82b5a808",
          7315 => x"248b3882",
          7316 => x"b5a80882",
          7317 => x"ccf43480",
          7318 => x"527182b5",
          7319 => x"a80c833d",
          7320 => x"0d04ef3d",
          7321 => x"0d805393",
          7322 => x"3dd00552",
          7323 => x"943d51e9",
          7324 => x"c13f82b5",
          7325 => x"a8085582",
          7326 => x"b5a80880",
          7327 => x"e0387658",
          7328 => x"6352933d",
          7329 => x"d40551e0",
          7330 => x"8d3f82b5",
          7331 => x"a8085582",
          7332 => x"b5a808bc",
          7333 => x"380280c7",
          7334 => x"05337098",
          7335 => x"2b555673",
          7336 => x"80258938",
          7337 => x"767a9412",
          7338 => x"0c54b239",
          7339 => x"02a20533",
          7340 => x"70842a70",
          7341 => x"81065155",
          7342 => x"5673802e",
          7343 => x"9e38767f",
          7344 => x"53705254",
          7345 => x"dba83f82",
          7346 => x"b5a80894",
          7347 => x"150c8e39",
          7348 => x"82b5a808",
          7349 => x"842e0981",
          7350 => x"06833885",
          7351 => x"557482b5",
          7352 => x"a80c933d",
          7353 => x"0d04e43d",
          7354 => x"0d6f6f5b",
          7355 => x"5b807a34",
          7356 => x"80539e3d",
          7357 => x"ffb80552",
          7358 => x"9f3d51e8",
          7359 => x"b53f82b5",
          7360 => x"a8085782",
          7361 => x"b5a80882",
          7362 => x"fc387b43",
          7363 => x"7a7c9411",
          7364 => x"08475558",
          7365 => x"64547380",
          7366 => x"2e81ed38",
          7367 => x"a052933d",
          7368 => x"705255d5",
          7369 => x"ea3f82b5",
          7370 => x"a8085782",
          7371 => x"b5a80882",
          7372 => x"d4386852",
          7373 => x"7b51c9c8",
          7374 => x"3f82b5a8",
          7375 => x"085782b5",
          7376 => x"a80882c1",
          7377 => x"3869527b",
          7378 => x"51daa33f",
          7379 => x"82b5a808",
          7380 => x"45765274",
          7381 => x"51d5b83f",
          7382 => x"82b5a808",
          7383 => x"5782b5a8",
          7384 => x"0882a238",
          7385 => x"80527451",
          7386 => x"daeb3f82",
          7387 => x"b5a80857",
          7388 => x"82b5a808",
          7389 => x"a4386952",
          7390 => x"7b51d9f2",
          7391 => x"3f7382b5",
          7392 => x"a8082ea6",
          7393 => x"38765274",
          7394 => x"51d6cf3f",
          7395 => x"82b5a808",
          7396 => x"5782b5a8",
          7397 => x"08802ecc",
          7398 => x"3876842e",
          7399 => x"09810686",
          7400 => x"38825781",
          7401 => x"e0397681",
          7402 => x"dc389e3d",
          7403 => x"ffbc0552",
          7404 => x"7451dcc9",
          7405 => x"3f76903d",
          7406 => x"78118111",
          7407 => x"3351565a",
          7408 => x"5673802e",
          7409 => x"913802b9",
          7410 => x"05558116",
          7411 => x"81167033",
          7412 => x"56565673",
          7413 => x"f5388116",
          7414 => x"54737826",
          7415 => x"81903875",
          7416 => x"802e9938",
          7417 => x"78168105",
          7418 => x"55ff186f",
          7419 => x"11ff18ff",
          7420 => x"18585855",
          7421 => x"58743374",
          7422 => x"3475ee38",
          7423 => x"ff186f11",
          7424 => x"5558af74",
          7425 => x"34fe8d39",
          7426 => x"777b2e09",
          7427 => x"81068a38",
          7428 => x"ff186f11",
          7429 => x"5558af74",
          7430 => x"34800b82",
          7431 => x"ccf43370",
          7432 => x"842982ae",
          7433 => x"e0057008",
          7434 => x"7033525c",
          7435 => x"56565673",
          7436 => x"762e8d38",
          7437 => x"8116701a",
          7438 => x"70335155",
          7439 => x"5673f538",
          7440 => x"82165473",
          7441 => x"7826a738",
          7442 => x"80557476",
          7443 => x"27913874",
          7444 => x"19547333",
          7445 => x"7a708105",
          7446 => x"5c348115",
          7447 => x"55ec39ba",
          7448 => x"7a708105",
          7449 => x"5c3474ff",
          7450 => x"2e098106",
          7451 => x"85389157",
          7452 => x"94396e18",
          7453 => x"81195954",
          7454 => x"73337a70",
          7455 => x"81055c34",
          7456 => x"7a7826ee",
          7457 => x"38807a34",
          7458 => x"7682b5a8",
          7459 => x"0c9e3d0d",
          7460 => x"04f73d0d",
          7461 => x"7b7d8d3d",
          7462 => x"fc055471",
          7463 => x"535755ec",
          7464 => x"bb3f82b5",
          7465 => x"a8085382",
          7466 => x"b5a80882",
          7467 => x"fa389115",
          7468 => x"33537282",
          7469 => x"f2388c15",
          7470 => x"08547376",
          7471 => x"27923890",
          7472 => x"15337081",
          7473 => x"2a708106",
          7474 => x"51545772",
          7475 => x"83387356",
          7476 => x"94150854",
          7477 => x"80709417",
          7478 => x"0c587578",
          7479 => x"2e829738",
          7480 => x"798a1122",
          7481 => x"70892b59",
          7482 => x"51537378",
          7483 => x"2eb73876",
          7484 => x"52ff1651",
          7485 => x"fee8ac3f",
          7486 => x"82b5a808",
          7487 => x"ff157854",
          7488 => x"70535553",
          7489 => x"fee89c3f",
          7490 => x"82b5a808",
          7491 => x"73269638",
          7492 => x"76307075",
          7493 => x"06709418",
          7494 => x"0c777131",
          7495 => x"98180857",
          7496 => x"585153b1",
          7497 => x"39881508",
          7498 => x"5473a638",
          7499 => x"73527451",
          7500 => x"cdca3f82",
          7501 => x"b5a80854",
          7502 => x"82b5a808",
          7503 => x"812e819a",
          7504 => x"3882b5a8",
          7505 => x"08ff2e81",
          7506 => x"9b3882b5",
          7507 => x"a8088816",
          7508 => x"0c739816",
          7509 => x"0c73802e",
          7510 => x"819c3876",
          7511 => x"762780dc",
          7512 => x"38757731",
          7513 => x"94160818",
          7514 => x"94170c90",
          7515 => x"16337081",
          7516 => x"2a708106",
          7517 => x"51555a56",
          7518 => x"72802e9a",
          7519 => x"38735274",
          7520 => x"51ccf93f",
          7521 => x"82b5a808",
          7522 => x"5482b5a8",
          7523 => x"08943882",
          7524 => x"b5a80856",
          7525 => x"a7397352",
          7526 => x"7451c784",
          7527 => x"3f82b5a8",
          7528 => x"085473ff",
          7529 => x"2ebe3881",
          7530 => x"7427af38",
          7531 => x"79537398",
          7532 => x"140827a6",
          7533 => x"38739816",
          7534 => x"0cffa039",
          7535 => x"94150816",
          7536 => x"94160c75",
          7537 => x"83ff0653",
          7538 => x"72802eaa",
          7539 => x"38735279",
          7540 => x"51c6a33f",
          7541 => x"82b5a808",
          7542 => x"9438820b",
          7543 => x"91163482",
          7544 => x"5380c439",
          7545 => x"810b9116",
          7546 => x"348153bb",
          7547 => x"3975892a",
          7548 => x"82b5a808",
          7549 => x"05589415",
          7550 => x"08548c15",
          7551 => x"08742790",
          7552 => x"38738c16",
          7553 => x"0c901533",
          7554 => x"80c00753",
          7555 => x"72901634",
          7556 => x"7383ff06",
          7557 => x"5372802e",
          7558 => x"8c38779c",
          7559 => x"16082e85",
          7560 => x"38779c16",
          7561 => x"0c805372",
          7562 => x"82b5a80c",
          7563 => x"8b3d0d04",
          7564 => x"f93d0d79",
          7565 => x"56895475",
          7566 => x"802e818a",
          7567 => x"38805389",
          7568 => x"3dfc0552",
          7569 => x"8a3d8405",
          7570 => x"51e1e73f",
          7571 => x"82b5a808",
          7572 => x"5582b5a8",
          7573 => x"0880ea38",
          7574 => x"77760c7a",
          7575 => x"527551d8",
          7576 => x"b53f82b5",
          7577 => x"a8085582",
          7578 => x"b5a80880",
          7579 => x"c338ab16",
          7580 => x"3370982b",
          7581 => x"55578074",
          7582 => x"24a23886",
          7583 => x"16337084",
          7584 => x"2a708106",
          7585 => x"51555773",
          7586 => x"802ead38",
          7587 => x"9c160852",
          7588 => x"7751d3da",
          7589 => x"3f82b5a8",
          7590 => x"0888170c",
          7591 => x"77548614",
          7592 => x"22841723",
          7593 => x"74527551",
          7594 => x"cee53f82",
          7595 => x"b5a80855",
          7596 => x"74842e09",
          7597 => x"81068538",
          7598 => x"85558639",
          7599 => x"74802e84",
          7600 => x"3880760c",
          7601 => x"74547382",
          7602 => x"b5a80c89",
          7603 => x"3d0d04fc",
          7604 => x"3d0d7687",
          7605 => x"3dfc0553",
          7606 => x"705253e7",
          7607 => x"ff3f82b5",
          7608 => x"a8088738",
          7609 => x"82b5a808",
          7610 => x"730c863d",
          7611 => x"0d04fb3d",
          7612 => x"0d777989",
          7613 => x"3dfc0554",
          7614 => x"71535654",
          7615 => x"e7de3f82",
          7616 => x"b5a80853",
          7617 => x"82b5a808",
          7618 => x"80df3874",
          7619 => x"933882b5",
          7620 => x"a8085273",
          7621 => x"51cdf83f",
          7622 => x"82b5a808",
          7623 => x"5380ca39",
          7624 => x"82b5a808",
          7625 => x"527351d3",
          7626 => x"ac3f82b5",
          7627 => x"a8085382",
          7628 => x"b5a80884",
          7629 => x"2e098106",
          7630 => x"85388053",
          7631 => x"873982b5",
          7632 => x"a808a638",
          7633 => x"74527351",
          7634 => x"d5b33f72",
          7635 => x"527351cf",
          7636 => x"893f82b5",
          7637 => x"a8088432",
          7638 => x"70307072",
          7639 => x"079f2c70",
          7640 => x"82b5a808",
          7641 => x"06515154",
          7642 => x"547282b5",
          7643 => x"a80c873d",
          7644 => x"0d04ee3d",
          7645 => x"0d655780",
          7646 => x"53893d70",
          7647 => x"53963d52",
          7648 => x"56dfaf3f",
          7649 => x"82b5a808",
          7650 => x"5582b5a8",
          7651 => x"08b23864",
          7652 => x"527551d6",
          7653 => x"813f82b5",
          7654 => x"a8085582",
          7655 => x"b5a808a0",
          7656 => x"380280cb",
          7657 => x"05337098",
          7658 => x"2b555873",
          7659 => x"80258538",
          7660 => x"86558d39",
          7661 => x"76802e88",
          7662 => x"38765275",
          7663 => x"51d4be3f",
          7664 => x"7482b5a8",
          7665 => x"0c943d0d",
          7666 => x"04f03d0d",
          7667 => x"6365555c",
          7668 => x"8053923d",
          7669 => x"ec055293",
          7670 => x"3d51ded6",
          7671 => x"3f82b5a8",
          7672 => x"085b82b5",
          7673 => x"a8088280",
          7674 => x"387c740c",
          7675 => x"73089811",
          7676 => x"08fe1190",
          7677 => x"13085956",
          7678 => x"58557574",
          7679 => x"26913875",
          7680 => x"7c0c81e4",
          7681 => x"39815b81",
          7682 => x"cc39825b",
          7683 => x"81c73982",
          7684 => x"b5a80875",
          7685 => x"33555973",
          7686 => x"812e0981",
          7687 => x"06bf3882",
          7688 => x"755f5776",
          7689 => x"52923df0",
          7690 => x"0551c1f4",
          7691 => x"3f82b5a8",
          7692 => x"08ff2ed1",
          7693 => x"3882b5a8",
          7694 => x"08812ece",
          7695 => x"3882b5a8",
          7696 => x"08307082",
          7697 => x"b5a80807",
          7698 => x"80257a05",
          7699 => x"81197f53",
          7700 => x"595a5498",
          7701 => x"14087726",
          7702 => x"ca3880f9",
          7703 => x"39a41508",
          7704 => x"82b5a808",
          7705 => x"57587598",
          7706 => x"38775281",
          7707 => x"187d5258",
          7708 => x"ffbf8d3f",
          7709 => x"82b5a808",
          7710 => x"5b82b5a8",
          7711 => x"0880d638",
          7712 => x"7c703377",
          7713 => x"12ff1a5d",
          7714 => x"52565474",
          7715 => x"822e0981",
          7716 => x"069e38b4",
          7717 => x"1451ffbb",
          7718 => x"cb3f82b5",
          7719 => x"a80883ff",
          7720 => x"ff067030",
          7721 => x"7080251b",
          7722 => x"8219595b",
          7723 => x"51549b39",
          7724 => x"b41451ff",
          7725 => x"bbc53f82",
          7726 => x"b5a808f0",
          7727 => x"0a067030",
          7728 => x"7080251b",
          7729 => x"8419595b",
          7730 => x"51547583",
          7731 => x"ff067a58",
          7732 => x"5679ff92",
          7733 => x"38787c0c",
          7734 => x"7c799012",
          7735 => x"0c841133",
          7736 => x"81075654",
          7737 => x"74841534",
          7738 => x"7a82b5a8",
          7739 => x"0c923d0d",
          7740 => x"04f93d0d",
          7741 => x"798a3dfc",
          7742 => x"05537052",
          7743 => x"57e3dd3f",
          7744 => x"82b5a808",
          7745 => x"5682b5a8",
          7746 => x"0881a838",
          7747 => x"91173356",
          7748 => x"7581a038",
          7749 => x"90173370",
          7750 => x"812a7081",
          7751 => x"06515555",
          7752 => x"87557380",
          7753 => x"2e818e38",
          7754 => x"94170854",
          7755 => x"738c1808",
          7756 => x"27818038",
          7757 => x"739b3882",
          7758 => x"b5a80853",
          7759 => x"88170852",
          7760 => x"7651c48c",
          7761 => x"3f82b5a8",
          7762 => x"08748819",
          7763 => x"0c5680c9",
          7764 => x"39981708",
          7765 => x"527651ff",
          7766 => x"bfc63f82",
          7767 => x"b5a808ff",
          7768 => x"2e098106",
          7769 => x"83388156",
          7770 => x"82b5a808",
          7771 => x"812e0981",
          7772 => x"06853882",
          7773 => x"56a33975",
          7774 => x"a0387754",
          7775 => x"82b5a808",
          7776 => x"98150827",
          7777 => x"94389817",
          7778 => x"085382b5",
          7779 => x"a8085276",
          7780 => x"51c3bd3f",
          7781 => x"82b5a808",
          7782 => x"56941708",
          7783 => x"8c180c90",
          7784 => x"173380c0",
          7785 => x"07547390",
          7786 => x"18347580",
          7787 => x"2e853875",
          7788 => x"91183475",
          7789 => x"557482b5",
          7790 => x"a80c893d",
          7791 => x"0d04e23d",
          7792 => x"0d8253a0",
          7793 => x"3dffa405",
          7794 => x"52a13d51",
          7795 => x"dae43f82",
          7796 => x"b5a80855",
          7797 => x"82b5a808",
          7798 => x"81f53878",
          7799 => x"45a13d08",
          7800 => x"52953d70",
          7801 => x"5258d1ae",
          7802 => x"3f82b5a8",
          7803 => x"085582b5",
          7804 => x"a80881db",
          7805 => x"380280fb",
          7806 => x"05337085",
          7807 => x"2a708106",
          7808 => x"51555686",
          7809 => x"557381c7",
          7810 => x"3875982b",
          7811 => x"54807424",
          7812 => x"81bd3802",
          7813 => x"80d60533",
          7814 => x"70810658",
          7815 => x"54875576",
          7816 => x"81ad386b",
          7817 => x"527851cc",
          7818 => x"c53f82b5",
          7819 => x"a8087484",
          7820 => x"2a708106",
          7821 => x"51555673",
          7822 => x"802e80d4",
          7823 => x"38785482",
          7824 => x"b5a80894",
          7825 => x"15082e81",
          7826 => x"8638735a",
          7827 => x"82b5a808",
          7828 => x"5c76528a",
          7829 => x"3d705254",
          7830 => x"c7b53f82",
          7831 => x"b5a80855",
          7832 => x"82b5a808",
          7833 => x"80e93882",
          7834 => x"b5a80852",
          7835 => x"7351cce5",
          7836 => x"3f82b5a8",
          7837 => x"085582b5",
          7838 => x"a8088638",
          7839 => x"875580cf",
          7840 => x"3982b5a8",
          7841 => x"08842e88",
          7842 => x"3882b5a8",
          7843 => x"0880c038",
          7844 => x"7751cec2",
          7845 => x"3f82b5a8",
          7846 => x"0882b5a8",
          7847 => x"08307082",
          7848 => x"b5a80807",
          7849 => x"80255155",
          7850 => x"5575802e",
          7851 => x"94387380",
          7852 => x"2e8f3880",
          7853 => x"53755277",
          7854 => x"51c1953f",
          7855 => x"82b5a808",
          7856 => x"55748c38",
          7857 => x"7851ffba",
          7858 => x"fe3f82b5",
          7859 => x"a8085574",
          7860 => x"82b5a80c",
          7861 => x"a03d0d04",
          7862 => x"e93d0d82",
          7863 => x"53993dc0",
          7864 => x"05529a3d",
          7865 => x"51d8cb3f",
          7866 => x"82b5a808",
          7867 => x"5482b5a8",
          7868 => x"0882b038",
          7869 => x"785e6952",
          7870 => x"8e3d7052",
          7871 => x"58cf973f",
          7872 => x"82b5a808",
          7873 => x"5482b5a8",
          7874 => x"08863888",
          7875 => x"54829439",
          7876 => x"82b5a808",
          7877 => x"842e0981",
          7878 => x"06828838",
          7879 => x"0280df05",
          7880 => x"3370852a",
          7881 => x"81065155",
          7882 => x"86547481",
          7883 => x"f638785a",
          7884 => x"74528a3d",
          7885 => x"705257c1",
          7886 => x"c33f82b5",
          7887 => x"a8087555",
          7888 => x"5682b5a8",
          7889 => x"08833887",
          7890 => x"5482b5a8",
          7891 => x"08812e09",
          7892 => x"81068338",
          7893 => x"825482b5",
          7894 => x"a808ff2e",
          7895 => x"09810686",
          7896 => x"38815481",
          7897 => x"b4397381",
          7898 => x"b03882b5",
          7899 => x"a8085278",
          7900 => x"51c4a43f",
          7901 => x"82b5a808",
          7902 => x"5482b5a8",
          7903 => x"08819a38",
          7904 => x"8b53a052",
          7905 => x"b41951ff",
          7906 => x"b78c3f78",
          7907 => x"54ae0bb4",
          7908 => x"15347854",
          7909 => x"900bbf15",
          7910 => x"348288b2",
          7911 => x"0a5280ca",
          7912 => x"1951ffb6",
          7913 => x"9f3f7553",
          7914 => x"78b41153",
          7915 => x"51c9f83f",
          7916 => x"a05378b4",
          7917 => x"115380d4",
          7918 => x"0551ffb6",
          7919 => x"b63f7854",
          7920 => x"ae0b80d5",
          7921 => x"15347f53",
          7922 => x"7880d411",
          7923 => x"5351c9d7",
          7924 => x"3f785481",
          7925 => x"0b831534",
          7926 => x"7751cba4",
          7927 => x"3f82b5a8",
          7928 => x"085482b5",
          7929 => x"a808b238",
          7930 => x"8288b20a",
          7931 => x"52649605",
          7932 => x"51ffb5d0",
          7933 => x"3f755364",
          7934 => x"527851c9",
          7935 => x"aa3f6454",
          7936 => x"900b8b15",
          7937 => x"34785481",
          7938 => x"0b831534",
          7939 => x"7851ffb8",
          7940 => x"b63f82b5",
          7941 => x"a808548b",
          7942 => x"39805375",
          7943 => x"527651ff",
          7944 => x"beae3f73",
          7945 => x"82b5a80c",
          7946 => x"993d0d04",
          7947 => x"da3d0da9",
          7948 => x"3d840551",
          7949 => x"d2f13f82",
          7950 => x"53a83dff",
          7951 => x"840552a9",
          7952 => x"3d51d5ee",
          7953 => x"3f82b5a8",
          7954 => x"085582b5",
          7955 => x"a80882d3",
          7956 => x"38784da9",
          7957 => x"3d08529d",
          7958 => x"3d705258",
          7959 => x"ccb83f82",
          7960 => x"b5a80855",
          7961 => x"82b5a808",
          7962 => x"82b93802",
          7963 => x"819b0533",
          7964 => x"81a00654",
          7965 => x"86557382",
          7966 => x"aa38a053",
          7967 => x"a43d0852",
          7968 => x"a83dff88",
          7969 => x"0551ffb4",
          7970 => x"ea3fac53",
          7971 => x"7752923d",
          7972 => x"705254ff",
          7973 => x"b4dd3faa",
          7974 => x"3d085273",
          7975 => x"51cbf73f",
          7976 => x"82b5a808",
          7977 => x"5582b5a8",
          7978 => x"08953863",
          7979 => x"6f2e0981",
          7980 => x"06883865",
          7981 => x"a23d082e",
          7982 => x"92388855",
          7983 => x"81e53982",
          7984 => x"b5a80884",
          7985 => x"2e098106",
          7986 => x"81b83873",
          7987 => x"51c9b13f",
          7988 => x"82b5a808",
          7989 => x"5582b5a8",
          7990 => x"0881c838",
          7991 => x"68569353",
          7992 => x"a83dff95",
          7993 => x"05528d16",
          7994 => x"51ffb487",
          7995 => x"3f02af05",
          7996 => x"338b1734",
          7997 => x"8b163370",
          7998 => x"842a7081",
          7999 => x"06515555",
          8000 => x"73893874",
          8001 => x"a0075473",
          8002 => x"8b173478",
          8003 => x"54810b83",
          8004 => x"15348b16",
          8005 => x"3370842a",
          8006 => x"70810651",
          8007 => x"55557380",
          8008 => x"2e80e538",
          8009 => x"6e642e80",
          8010 => x"df387552",
          8011 => x"7851c6be",
          8012 => x"3f82b5a8",
          8013 => x"08527851",
          8014 => x"ffb7bb3f",
          8015 => x"825582b5",
          8016 => x"a808802e",
          8017 => x"80dd3882",
          8018 => x"b5a80852",
          8019 => x"7851ffb5",
          8020 => x"af3f82b5",
          8021 => x"a8087980",
          8022 => x"d4115858",
          8023 => x"5582b5a8",
          8024 => x"0880c038",
          8025 => x"81163354",
          8026 => x"73ae2e09",
          8027 => x"81069938",
          8028 => x"63537552",
          8029 => x"7651c6af",
          8030 => x"3f785481",
          8031 => x"0b831534",
          8032 => x"873982b5",
          8033 => x"a8089c38",
          8034 => x"7751c8ca",
          8035 => x"3f82b5a8",
          8036 => x"085582b5",
          8037 => x"a8088c38",
          8038 => x"7851ffb5",
          8039 => x"aa3f82b5",
          8040 => x"a8085574",
          8041 => x"82b5a80c",
          8042 => x"a83d0d04",
          8043 => x"ed3d0d02",
          8044 => x"80db0533",
          8045 => x"02840580",
          8046 => x"df053357",
          8047 => x"57825395",
          8048 => x"3dd00552",
          8049 => x"963d51d2",
          8050 => x"e93f82b5",
          8051 => x"a8085582",
          8052 => x"b5a80880",
          8053 => x"cf38785a",
          8054 => x"6552953d",
          8055 => x"d40551c9",
          8056 => x"b53f82b5",
          8057 => x"a8085582",
          8058 => x"b5a808b8",
          8059 => x"380280cf",
          8060 => x"053381a0",
          8061 => x"06548655",
          8062 => x"73aa3875",
          8063 => x"a7066171",
          8064 => x"098b1233",
          8065 => x"71067a74",
          8066 => x"06075157",
          8067 => x"5556748b",
          8068 => x"15347854",
          8069 => x"810b8315",
          8070 => x"347851ff",
          8071 => x"b4a93f82",
          8072 => x"b5a80855",
          8073 => x"7482b5a8",
          8074 => x"0c953d0d",
          8075 => x"04ef3d0d",
          8076 => x"64568253",
          8077 => x"933dd005",
          8078 => x"52943d51",
          8079 => x"d1f43f82",
          8080 => x"b5a80855",
          8081 => x"82b5a808",
          8082 => x"80cb3876",
          8083 => x"58635293",
          8084 => x"3dd40551",
          8085 => x"c8c03f82",
          8086 => x"b5a80855",
          8087 => x"82b5a808",
          8088 => x"b4380280",
          8089 => x"c7053381",
          8090 => x"a0065486",
          8091 => x"5573a638",
          8092 => x"84162286",
          8093 => x"17227190",
          8094 => x"2b075354",
          8095 => x"961f51ff",
          8096 => x"b0c23f76",
          8097 => x"54810b83",
          8098 => x"15347651",
          8099 => x"ffb3b83f",
          8100 => x"82b5a808",
          8101 => x"557482b5",
          8102 => x"a80c933d",
          8103 => x"0d04ea3d",
          8104 => x"0d696b5c",
          8105 => x"5a805398",
          8106 => x"3dd00552",
          8107 => x"993d51d1",
          8108 => x"813f82b5",
          8109 => x"a80882b5",
          8110 => x"a8083070",
          8111 => x"82b5a808",
          8112 => x"07802551",
          8113 => x"55577980",
          8114 => x"2e818538",
          8115 => x"81707506",
          8116 => x"55557380",
          8117 => x"2e80f938",
          8118 => x"7b5d805f",
          8119 => x"80528d3d",
          8120 => x"705254ff",
          8121 => x"bea93f82",
          8122 => x"b5a80857",
          8123 => x"82b5a808",
          8124 => x"80d13874",
          8125 => x"527351c3",
          8126 => x"dc3f82b5",
          8127 => x"a8085782",
          8128 => x"b5a808bf",
          8129 => x"3882b5a8",
          8130 => x"0882b5a8",
          8131 => x"08655b59",
          8132 => x"56781881",
          8133 => x"197b1856",
          8134 => x"59557433",
          8135 => x"74348116",
          8136 => x"568a7827",
          8137 => x"ec388b56",
          8138 => x"751a5480",
          8139 => x"74347580",
          8140 => x"2e9e38ff",
          8141 => x"16701b70",
          8142 => x"33515556",
          8143 => x"73a02ee8",
          8144 => x"388e3976",
          8145 => x"842e0981",
          8146 => x"06863880",
          8147 => x"7a348057",
          8148 => x"76307078",
          8149 => x"07802551",
          8150 => x"547a802e",
          8151 => x"80c13873",
          8152 => x"802ebc38",
          8153 => x"7ba01108",
          8154 => x"5351ffb1",
          8155 => x"933f82b5",
          8156 => x"a8085782",
          8157 => x"b5a808a7",
          8158 => x"387b7033",
          8159 => x"555580c3",
          8160 => x"5673832e",
          8161 => x"8b3880e4",
          8162 => x"5673842e",
          8163 => x"8338a756",
          8164 => x"7515b405",
          8165 => x"51ffade3",
          8166 => x"3f82b5a8",
          8167 => x"087b0c76",
          8168 => x"82b5a80c",
          8169 => x"983d0d04",
          8170 => x"e63d0d82",
          8171 => x"539c3dff",
          8172 => x"b805529d",
          8173 => x"3d51cefa",
          8174 => x"3f82b5a8",
          8175 => x"0882b5a8",
          8176 => x"08565482",
          8177 => x"b5a80883",
          8178 => x"98388b53",
          8179 => x"a0528b3d",
          8180 => x"705259ff",
          8181 => x"aec03f73",
          8182 => x"6d703370",
          8183 => x"81ff0652",
          8184 => x"5755579f",
          8185 => x"742781bc",
          8186 => x"38785874",
          8187 => x"81ff066d",
          8188 => x"81054e70",
          8189 => x"5255ffaf",
          8190 => x"893f82b5",
          8191 => x"a808802e",
          8192 => x"a5386c70",
          8193 => x"33705357",
          8194 => x"54ffaefd",
          8195 => x"3f82b5a8",
          8196 => x"08802e8d",
          8197 => x"3874882b",
          8198 => x"76076d81",
          8199 => x"054e5586",
          8200 => x"3982b5a8",
          8201 => x"0855ff9f",
          8202 => x"157083ff",
          8203 => x"ff065154",
          8204 => x"7399268a",
          8205 => x"38e01570",
          8206 => x"83ffff06",
          8207 => x"565480ff",
          8208 => x"75278738",
          8209 => x"82adf015",
          8210 => x"33557480",
          8211 => x"2ea33874",
          8212 => x"5282aff0",
          8213 => x"51ffae89",
          8214 => x"3f82b5a8",
          8215 => x"08933881",
          8216 => x"ff752788",
          8217 => x"38768926",
          8218 => x"88388b39",
          8219 => x"8a772786",
          8220 => x"38865581",
          8221 => x"ec3981ff",
          8222 => x"75278f38",
          8223 => x"74882a54",
          8224 => x"73787081",
          8225 => x"055a3481",
          8226 => x"17577478",
          8227 => x"7081055a",
          8228 => x"3481176d",
          8229 => x"70337081",
          8230 => x"ff065257",
          8231 => x"5557739f",
          8232 => x"26fec838",
          8233 => x"8b3d3354",
          8234 => x"86557381",
          8235 => x"e52e81b1",
          8236 => x"3876802e",
          8237 => x"993802a7",
          8238 => x"05557615",
          8239 => x"70335154",
          8240 => x"73a02e09",
          8241 => x"81068738",
          8242 => x"ff175776",
          8243 => x"ed387941",
          8244 => x"80438052",
          8245 => x"913d7052",
          8246 => x"55ffbab3",
          8247 => x"3f82b5a8",
          8248 => x"085482b5",
          8249 => x"a80880f7",
          8250 => x"38815274",
          8251 => x"51ffbfe5",
          8252 => x"3f82b5a8",
          8253 => x"085482b5",
          8254 => x"a8088d38",
          8255 => x"7680c438",
          8256 => x"6754e574",
          8257 => x"3480c639",
          8258 => x"82b5a808",
          8259 => x"842e0981",
          8260 => x"0680cc38",
          8261 => x"80547674",
          8262 => x"2e80c438",
          8263 => x"81527451",
          8264 => x"ffbdb03f",
          8265 => x"82b5a808",
          8266 => x"5482b5a8",
          8267 => x"08b138a0",
          8268 => x"5382b5a8",
          8269 => x"08526751",
          8270 => x"ffabdb3f",
          8271 => x"6754880b",
          8272 => x"8b15348b",
          8273 => x"53785267",
          8274 => x"51ffaba7",
          8275 => x"3f795481",
          8276 => x"0b831534",
          8277 => x"7951ffad",
          8278 => x"ee3f82b5",
          8279 => x"a8085473",
          8280 => x"557482b5",
          8281 => x"a80c9c3d",
          8282 => x"0d04f23d",
          8283 => x"0d606202",
          8284 => x"880580cb",
          8285 => x"0533933d",
          8286 => x"fc055572",
          8287 => x"54405e5a",
          8288 => x"d2da3f82",
          8289 => x"b5a80858",
          8290 => x"82b5a808",
          8291 => x"82bd3891",
          8292 => x"1a335877",
          8293 => x"82b5387c",
          8294 => x"802e9738",
          8295 => x"8c1a0859",
          8296 => x"78903890",
          8297 => x"1a337081",
          8298 => x"2a708106",
          8299 => x"51555573",
          8300 => x"90388754",
          8301 => x"82973982",
          8302 => x"58829039",
          8303 => x"8158828b",
          8304 => x"397e8a11",
          8305 => x"2270892b",
          8306 => x"70557f54",
          8307 => x"565656fe",
          8308 => x"ced13fff",
          8309 => x"147d0670",
          8310 => x"30707207",
          8311 => x"9f2a82b5",
          8312 => x"a808058c",
          8313 => x"19087c40",
          8314 => x"5a5d5555",
          8315 => x"81772788",
          8316 => x"38981608",
          8317 => x"77268338",
          8318 => x"82577677",
          8319 => x"56598056",
          8320 => x"74527951",
          8321 => x"ffae993f",
          8322 => x"81157f55",
          8323 => x"55981408",
          8324 => x"75268338",
          8325 => x"825582b5",
          8326 => x"a808812e",
          8327 => x"ff993882",
          8328 => x"b5a808ff",
          8329 => x"2eff9538",
          8330 => x"82b5a808",
          8331 => x"8e388116",
          8332 => x"56757b2e",
          8333 => x"09810687",
          8334 => x"38933974",
          8335 => x"59805674",
          8336 => x"772e0981",
          8337 => x"06ffb938",
          8338 => x"875880ff",
          8339 => x"397d802e",
          8340 => x"ba38787b",
          8341 => x"55557a80",
          8342 => x"2eb43881",
          8343 => x"15567381",
          8344 => x"2e098106",
          8345 => x"8338ff56",
          8346 => x"75537452",
          8347 => x"7e51ffaf",
          8348 => x"a83f82b5",
          8349 => x"a8085882",
          8350 => x"b5a80880",
          8351 => x"ce387481",
          8352 => x"16ff1656",
          8353 => x"565c73d3",
          8354 => x"388439ff",
          8355 => x"195c7e7c",
          8356 => x"8c120c55",
          8357 => x"7d802eb3",
          8358 => x"3878881b",
          8359 => x"0c7c8c1b",
          8360 => x"0c901a33",
          8361 => x"80c00754",
          8362 => x"73901b34",
          8363 => x"981508fe",
          8364 => x"05901608",
          8365 => x"57547574",
          8366 => x"26913875",
          8367 => x"7b319016",
          8368 => x"0c841533",
          8369 => x"81075473",
          8370 => x"84163477",
          8371 => x"547382b5",
          8372 => x"a80c903d",
          8373 => x"0d04e93d",
          8374 => x"0d6b6d02",
          8375 => x"880580eb",
          8376 => x"05339d3d",
          8377 => x"545a5c59",
          8378 => x"c5bd3f8b",
          8379 => x"56800b82",
          8380 => x"b5a80824",
          8381 => x"8bf83882",
          8382 => x"b5a80884",
          8383 => x"2982cce0",
          8384 => x"05700851",
          8385 => x"5574802e",
          8386 => x"84388075",
          8387 => x"3482b5a8",
          8388 => x"0881ff06",
          8389 => x"5f81527e",
          8390 => x"51ffa0d0",
          8391 => x"3f82b5a8",
          8392 => x"0881ff06",
          8393 => x"70810656",
          8394 => x"57835674",
          8395 => x"8bc03876",
          8396 => x"822a7081",
          8397 => x"0651558a",
          8398 => x"56748bb2",
          8399 => x"38993dfc",
          8400 => x"05538352",
          8401 => x"7e51ffa4",
          8402 => x"f03f82b5",
          8403 => x"a8089938",
          8404 => x"67557480",
          8405 => x"2e923874",
          8406 => x"82808026",
          8407 => x"8b38ff15",
          8408 => x"75065574",
          8409 => x"802e8338",
          8410 => x"81487880",
          8411 => x"2e873884",
          8412 => x"80792692",
          8413 => x"38788180",
          8414 => x"0a268b38",
          8415 => x"ff197906",
          8416 => x"5574802e",
          8417 => x"86389356",
          8418 => x"8ae43978",
          8419 => x"892a6e89",
          8420 => x"2a70892b",
          8421 => x"77594843",
          8422 => x"597a8338",
          8423 => x"81566130",
          8424 => x"70802577",
          8425 => x"07515591",
          8426 => x"56748ac2",
          8427 => x"38993df8",
          8428 => x"05538152",
          8429 => x"7e51ffa4",
          8430 => x"803f8156",
          8431 => x"82b5a808",
          8432 => x"8aac3877",
          8433 => x"832a7077",
          8434 => x"0682b5a8",
          8435 => x"08435645",
          8436 => x"748338bf",
          8437 => x"4166558e",
          8438 => x"56607526",
          8439 => x"8a903874",
          8440 => x"61317048",
          8441 => x"5580ff75",
          8442 => x"278a8338",
          8443 => x"93567881",
          8444 => x"802689fa",
          8445 => x"3877812a",
          8446 => x"70810656",
          8447 => x"4374802e",
          8448 => x"95387787",
          8449 => x"06557482",
          8450 => x"2e838d38",
          8451 => x"77810655",
          8452 => x"74802e83",
          8453 => x"83387781",
          8454 => x"06559356",
          8455 => x"825e7480",
          8456 => x"2e89cb38",
          8457 => x"785a7d83",
          8458 => x"2e098106",
          8459 => x"80e13878",
          8460 => x"ae386691",
          8461 => x"2a57810b",
          8462 => x"82b09422",
          8463 => x"565a7480",
          8464 => x"2e9d3874",
          8465 => x"77269838",
          8466 => x"82b09456",
          8467 => x"79108217",
          8468 => x"70225757",
          8469 => x"5a74802e",
          8470 => x"86387675",
          8471 => x"27ee3879",
          8472 => x"526651fe",
          8473 => x"c9bd3f82",
          8474 => x"b5a80884",
          8475 => x"29848705",
          8476 => x"70892a5e",
          8477 => x"55a05c80",
          8478 => x"0b82b5a8",
          8479 => x"08fc808a",
          8480 => x"055644fd",
          8481 => x"fff00a75",
          8482 => x"2780ec38",
          8483 => x"88d33978",
          8484 => x"ae38668c",
          8485 => x"2a57810b",
          8486 => x"82b08422",
          8487 => x"565a7480",
          8488 => x"2e9d3874",
          8489 => x"77269838",
          8490 => x"82b08456",
          8491 => x"79108217",
          8492 => x"70225757",
          8493 => x"5a74802e",
          8494 => x"86387675",
          8495 => x"27ee3879",
          8496 => x"526651fe",
          8497 => x"c8dd3f82",
          8498 => x"b5a80810",
          8499 => x"84055782",
          8500 => x"b5a8089f",
          8501 => x"f5269638",
          8502 => x"810b82b5",
          8503 => x"a8081082",
          8504 => x"b5a80805",
          8505 => x"7111722a",
          8506 => x"83055956",
          8507 => x"5e83ff17",
          8508 => x"892a5d81",
          8509 => x"5ca04460",
          8510 => x"1c7d1165",
          8511 => x"05697012",
          8512 => x"ff057130",
          8513 => x"70720674",
          8514 => x"315c5259",
          8515 => x"5759407d",
          8516 => x"832e0981",
          8517 => x"06893876",
          8518 => x"1c601841",
          8519 => x"5c843976",
          8520 => x"1d5d7990",
          8521 => x"29187062",
          8522 => x"31685851",
          8523 => x"55747626",
          8524 => x"87af3875",
          8525 => x"7c317d31",
          8526 => x"7a537065",
          8527 => x"315255fe",
          8528 => x"c7e13f82",
          8529 => x"b5a80858",
          8530 => x"7d832e09",
          8531 => x"81069b38",
          8532 => x"82b5a808",
          8533 => x"83fff526",
          8534 => x"80dd3878",
          8535 => x"87833879",
          8536 => x"812a5978",
          8537 => x"fdbe3886",
          8538 => x"f8397d82",
          8539 => x"2e098106",
          8540 => x"80c53883",
          8541 => x"fff50b82",
          8542 => x"b5a80827",
          8543 => x"a038788f",
          8544 => x"38791a55",
          8545 => x"7480c026",
          8546 => x"86387459",
          8547 => x"fd963962",
          8548 => x"81065574",
          8549 => x"802e8f38",
          8550 => x"835efd88",
          8551 => x"3982b5a8",
          8552 => x"089ff526",
          8553 => x"92387886",
          8554 => x"b838791a",
          8555 => x"59818079",
          8556 => x"27fcf138",
          8557 => x"86ab3980",
          8558 => x"557d812e",
          8559 => x"09810683",
          8560 => x"387d559f",
          8561 => x"f578278b",
          8562 => x"38748106",
          8563 => x"558e5674",
          8564 => x"869c3884",
          8565 => x"80538052",
          8566 => x"7a51ffa2",
          8567 => x"b93f8b53",
          8568 => x"82aeac52",
          8569 => x"7a51ffa2",
          8570 => x"8a3f8480",
          8571 => x"528b1b51",
          8572 => x"ffa1b33f",
          8573 => x"798d1c34",
          8574 => x"7b83ffff",
          8575 => x"06528e1b",
          8576 => x"51ffa1a2",
          8577 => x"3f810b90",
          8578 => x"1c347d83",
          8579 => x"32703070",
          8580 => x"962a8480",
          8581 => x"06545155",
          8582 => x"911b51ff",
          8583 => x"a1883f66",
          8584 => x"557483ff",
          8585 => x"ff269038",
          8586 => x"7483ffff",
          8587 => x"0652931b",
          8588 => x"51ffa0f2",
          8589 => x"3f8a3974",
          8590 => x"52a01b51",
          8591 => x"ffa1853f",
          8592 => x"f80b951c",
          8593 => x"34bf5298",
          8594 => x"1b51ffa0",
          8595 => x"d93f81ff",
          8596 => x"529a1b51",
          8597 => x"ffa0cf3f",
          8598 => x"60529c1b",
          8599 => x"51ffa0e4",
          8600 => x"3f7d832e",
          8601 => x"09810680",
          8602 => x"cb388288",
          8603 => x"b20a5280",
          8604 => x"c31b51ff",
          8605 => x"a0ce3f7c",
          8606 => x"52a41b51",
          8607 => x"ffa0c53f",
          8608 => x"8252ac1b",
          8609 => x"51ffa0bc",
          8610 => x"3f8152b0",
          8611 => x"1b51ffa0",
          8612 => x"953f8652",
          8613 => x"b21b51ff",
          8614 => x"a08c3fff",
          8615 => x"800b80c0",
          8616 => x"1c34a90b",
          8617 => x"80c21c34",
          8618 => x"935382ae",
          8619 => x"b85280c7",
          8620 => x"1b51ae39",
          8621 => x"8288b20a",
          8622 => x"52a71b51",
          8623 => x"ffa0853f",
          8624 => x"7c83ffff",
          8625 => x"0652961b",
          8626 => x"51ff9fda",
          8627 => x"3fff800b",
          8628 => x"a41c34a9",
          8629 => x"0ba61c34",
          8630 => x"935382ae",
          8631 => x"cc52ab1b",
          8632 => x"51ffa08f",
          8633 => x"3f82d4d5",
          8634 => x"5283fe1b",
          8635 => x"705259ff",
          8636 => x"9fb43f81",
          8637 => x"5460537a",
          8638 => x"527e51ff",
          8639 => x"9bd73f81",
          8640 => x"5682b5a8",
          8641 => x"0883e738",
          8642 => x"7d832e09",
          8643 => x"810680ee",
          8644 => x"38755460",
          8645 => x"8605537a",
          8646 => x"527e51ff",
          8647 => x"9bb73f84",
          8648 => x"80538052",
          8649 => x"7a51ff9f",
          8650 => x"ed3f848b",
          8651 => x"85a4d252",
          8652 => x"7a51ff9f",
          8653 => x"8f3f868a",
          8654 => x"85e4f252",
          8655 => x"83e41b51",
          8656 => x"ff9f813f",
          8657 => x"ff185283",
          8658 => x"e81b51ff",
          8659 => x"9ef63f82",
          8660 => x"5283ec1b",
          8661 => x"51ff9eec",
          8662 => x"3f82d4d5",
          8663 => x"527851ff",
          8664 => x"9ec43f75",
          8665 => x"54608705",
          8666 => x"537a527e",
          8667 => x"51ff9ae5",
          8668 => x"3f755460",
          8669 => x"16537a52",
          8670 => x"7e51ff9a",
          8671 => x"d83f6553",
          8672 => x"80527a51",
          8673 => x"ff9f8f3f",
          8674 => x"7f568058",
          8675 => x"7d832e09",
          8676 => x"81069a38",
          8677 => x"f8527a51",
          8678 => x"ff9ea93f",
          8679 => x"ff52841b",
          8680 => x"51ff9ea0",
          8681 => x"3ff00a52",
          8682 => x"881b5191",
          8683 => x"3987ffff",
          8684 => x"f8557d81",
          8685 => x"2e8338f8",
          8686 => x"5574527a",
          8687 => x"51ff9e84",
          8688 => x"3f7c5561",
          8689 => x"57746226",
          8690 => x"83387457",
          8691 => x"76547553",
          8692 => x"7a527e51",
          8693 => x"ff99fe3f",
          8694 => x"82b5a808",
          8695 => x"82873884",
          8696 => x"805382b5",
          8697 => x"a808527a",
          8698 => x"51ff9eaa",
          8699 => x"3f761675",
          8700 => x"78315656",
          8701 => x"74cd3881",
          8702 => x"18587780",
          8703 => x"2eff8d38",
          8704 => x"79557d83",
          8705 => x"2e833863",
          8706 => x"55615774",
          8707 => x"62268338",
          8708 => x"74577654",
          8709 => x"75537a52",
          8710 => x"7e51ff99",
          8711 => x"b83f82b5",
          8712 => x"a80881c1",
          8713 => x"38761675",
          8714 => x"78315656",
          8715 => x"74db388c",
          8716 => x"567d832e",
          8717 => x"93388656",
          8718 => x"6683ffff",
          8719 => x"268a3884",
          8720 => x"567d822e",
          8721 => x"83388156",
          8722 => x"64810658",
          8723 => x"7780fe38",
          8724 => x"84805377",
          8725 => x"527a51ff",
          8726 => x"9dbc3f82",
          8727 => x"d4d55278",
          8728 => x"51ff9cc2",
          8729 => x"3f83be1b",
          8730 => x"55777534",
          8731 => x"810b8116",
          8732 => x"34810b82",
          8733 => x"16347783",
          8734 => x"16347584",
          8735 => x"16346067",
          8736 => x"055680fd",
          8737 => x"c1527551",
          8738 => x"fec1983f",
          8739 => x"fe0b8516",
          8740 => x"3482b5a8",
          8741 => x"08822abf",
          8742 => x"07567586",
          8743 => x"163482b5",
          8744 => x"a8088716",
          8745 => x"34605283",
          8746 => x"c61b51ff",
          8747 => x"9c963f66",
          8748 => x"5283ca1b",
          8749 => x"51ff9c8c",
          8750 => x"3f815477",
          8751 => x"537a527e",
          8752 => x"51ff9891",
          8753 => x"3f815682",
          8754 => x"b5a808a2",
          8755 => x"38805380",
          8756 => x"527e51ff",
          8757 => x"99e33f81",
          8758 => x"5682b5a8",
          8759 => x"08903889",
          8760 => x"398e568a",
          8761 => x"39815686",
          8762 => x"3982b5a8",
          8763 => x"08567582",
          8764 => x"b5a80c99",
          8765 => x"3d0d04f5",
          8766 => x"3d0d7d60",
          8767 => x"5b598079",
          8768 => x"60ff055a",
          8769 => x"57577678",
          8770 => x"25b4388d",
          8771 => x"3df81155",
          8772 => x"558153fc",
          8773 => x"15527951",
          8774 => x"c9dc3f7a",
          8775 => x"812e0981",
          8776 => x"069c388c",
          8777 => x"3d335574",
          8778 => x"8d2edb38",
          8779 => x"74767081",
          8780 => x"05583481",
          8781 => x"1757748a",
          8782 => x"2e098106",
          8783 => x"c9388076",
          8784 => x"34785576",
          8785 => x"83387655",
          8786 => x"7482b5a8",
          8787 => x"0c8d3d0d",
          8788 => x"04f73d0d",
          8789 => x"7b028405",
          8790 => x"b3053359",
          8791 => x"57778a2e",
          8792 => x"09810687",
          8793 => x"388d5276",
          8794 => x"51e73f84",
          8795 => x"17085680",
          8796 => x"7624be38",
          8797 => x"88170877",
          8798 => x"178c0556",
          8799 => x"59777534",
          8800 => x"811656bb",
          8801 => x"7625a138",
          8802 => x"8b3dfc05",
          8803 => x"5475538c",
          8804 => x"17527608",
          8805 => x"51cbdc3f",
          8806 => x"79763270",
          8807 => x"30707207",
          8808 => x"9f2a7030",
          8809 => x"53515656",
          8810 => x"7584180c",
          8811 => x"81198818",
          8812 => x"0c8b3d0d",
          8813 => x"04f93d0d",
          8814 => x"79841108",
          8815 => x"56568075",
          8816 => x"24a73889",
          8817 => x"3dfc0554",
          8818 => x"74538c16",
          8819 => x"52750851",
          8820 => x"cba13f82",
          8821 => x"b5a80891",
          8822 => x"38841608",
          8823 => x"782e0981",
          8824 => x"06873888",
          8825 => x"16085583",
          8826 => x"39ff5574",
          8827 => x"82b5a80c",
          8828 => x"893d0d04",
          8829 => x"fd3d0d75",
          8830 => x"5480cc53",
          8831 => x"80527351",
          8832 => x"ff9a933f",
          8833 => x"76740c85",
          8834 => x"3d0d04ea",
          8835 => x"3d0d0280",
          8836 => x"e305336a",
          8837 => x"53863d70",
          8838 => x"535454d8",
          8839 => x"3f735272",
          8840 => x"51feae3f",
          8841 => x"7251ff8d",
          8842 => x"3f983d0d",
          8843 => x"04000000",
          8844 => x"00ffffff",
          8845 => x"ff00ffff",
          8846 => x"ffff00ff",
          8847 => x"ffffff00",
          8848 => x"00002ba8",
          8849 => x"00002b2c",
          8850 => x"00002b33",
          8851 => x"00002b3a",
          8852 => x"00002b41",
          8853 => x"00002b48",
          8854 => x"00002b4f",
          8855 => x"00002b56",
          8856 => x"00002b5d",
          8857 => x"00002b64",
          8858 => x"00002b6b",
          8859 => x"00002b72",
          8860 => x"00002b78",
          8861 => x"00002b7e",
          8862 => x"00002b84",
          8863 => x"00002b8a",
          8864 => x"00002b90",
          8865 => x"00002b96",
          8866 => x"00002b9c",
          8867 => x"00002ba2",
          8868 => x"0000413b",
          8869 => x"00004141",
          8870 => x"00004147",
          8871 => x"0000414d",
          8872 => x"00004153",
          8873 => x"00004720",
          8874 => x"00004816",
          8875 => x"0000490e",
          8876 => x"00004b48",
          8877 => x"000047fe",
          8878 => x"000045f5",
          8879 => x"000049c2",
          8880 => x"00004b1e",
          8881 => x"00004a00",
          8882 => x"00004a96",
          8883 => x"00004a1c",
          8884 => x"000048bd",
          8885 => x"000045f5",
          8886 => x"0000490e",
          8887 => x"00004932",
          8888 => x"000049c2",
          8889 => x"000045f5",
          8890 => x"000045f5",
          8891 => x"00004a1c",
          8892 => x"00004a96",
          8893 => x"00004b1e",
          8894 => x"00004b48",
          8895 => x"00000e2f",
          8896 => x"00001718",
          8897 => x"00001718",
          8898 => x"00000e5e",
          8899 => x"00001718",
          8900 => x"00001718",
          8901 => x"00001718",
          8902 => x"00001718",
          8903 => x"00001718",
          8904 => x"00001718",
          8905 => x"00001718",
          8906 => x"00000e1b",
          8907 => x"00001718",
          8908 => x"00000e46",
          8909 => x"00000e76",
          8910 => x"00001718",
          8911 => x"00001718",
          8912 => x"00001718",
          8913 => x"00001718",
          8914 => x"00001718",
          8915 => x"00001718",
          8916 => x"00001718",
          8917 => x"00001718",
          8918 => x"00001718",
          8919 => x"00001718",
          8920 => x"00001718",
          8921 => x"00001718",
          8922 => x"00001718",
          8923 => x"00001718",
          8924 => x"00001718",
          8925 => x"00001718",
          8926 => x"00001718",
          8927 => x"00001718",
          8928 => x"00001718",
          8929 => x"00001718",
          8930 => x"00001718",
          8931 => x"00001718",
          8932 => x"00001718",
          8933 => x"00001718",
          8934 => x"00001718",
          8935 => x"00001718",
          8936 => x"00001718",
          8937 => x"00001718",
          8938 => x"00001718",
          8939 => x"00001718",
          8940 => x"00001718",
          8941 => x"00001718",
          8942 => x"00001718",
          8943 => x"00001718",
          8944 => x"00001718",
          8945 => x"00001718",
          8946 => x"00000fa6",
          8947 => x"00001718",
          8948 => x"00001718",
          8949 => x"00001718",
          8950 => x"00001718",
          8951 => x"00001114",
          8952 => x"00001718",
          8953 => x"00001718",
          8954 => x"00001718",
          8955 => x"00001718",
          8956 => x"00001718",
          8957 => x"00001718",
          8958 => x"00001718",
          8959 => x"00001718",
          8960 => x"00001718",
          8961 => x"00001718",
          8962 => x"00000ed6",
          8963 => x"0000103d",
          8964 => x"00000ead",
          8965 => x"00000ead",
          8966 => x"00000ead",
          8967 => x"00001718",
          8968 => x"0000103d",
          8969 => x"00001718",
          8970 => x"00001718",
          8971 => x"00000e96",
          8972 => x"00001718",
          8973 => x"00001718",
          8974 => x"000010ea",
          8975 => x"000010f5",
          8976 => x"00001718",
          8977 => x"00001718",
          8978 => x"00000f0f",
          8979 => x"00001718",
          8980 => x"0000111d",
          8981 => x"00001718",
          8982 => x"00001718",
          8983 => x"00001114",
          8984 => x"64696e69",
          8985 => x"74000000",
          8986 => x"64696f63",
          8987 => x"746c0000",
          8988 => x"66696e69",
          8989 => x"74000000",
          8990 => x"666c6f61",
          8991 => x"64000000",
          8992 => x"66657865",
          8993 => x"63000000",
          8994 => x"6d636c65",
          8995 => x"61720000",
          8996 => x"6d636f70",
          8997 => x"79000000",
          8998 => x"6d646966",
          8999 => x"66000000",
          9000 => x"6d64756d",
          9001 => x"70000000",
          9002 => x"6d656200",
          9003 => x"6d656800",
          9004 => x"6d657700",
          9005 => x"68696400",
          9006 => x"68696500",
          9007 => x"68666400",
          9008 => x"68666500",
          9009 => x"63616c6c",
          9010 => x"00000000",
          9011 => x"6a6d7000",
          9012 => x"72657374",
          9013 => x"61727400",
          9014 => x"72657365",
          9015 => x"74000000",
          9016 => x"696e666f",
          9017 => x"00000000",
          9018 => x"74657374",
          9019 => x"00000000",
          9020 => x"74626173",
          9021 => x"69630000",
          9022 => x"6d626173",
          9023 => x"69630000",
          9024 => x"6b696c6f",
          9025 => x"00000000",
          9026 => x"65640000",
          9027 => x"4469736b",
          9028 => x"20457272",
          9029 => x"6f720a00",
          9030 => x"496e7465",
          9031 => x"726e616c",
          9032 => x"20657272",
          9033 => x"6f722e0a",
          9034 => x"00000000",
          9035 => x"4469736b",
          9036 => x"206e6f74",
          9037 => x"20726561",
          9038 => x"64792e0a",
          9039 => x"00000000",
          9040 => x"4e6f2066",
          9041 => x"696c6520",
          9042 => x"666f756e",
          9043 => x"642e0a00",
          9044 => x"4e6f2070",
          9045 => x"61746820",
          9046 => x"666f756e",
          9047 => x"642e0a00",
          9048 => x"496e7661",
          9049 => x"6c696420",
          9050 => x"66696c65",
          9051 => x"6e616d65",
          9052 => x"2e0a0000",
          9053 => x"41636365",
          9054 => x"73732064",
          9055 => x"656e6965",
          9056 => x"642e0a00",
          9057 => x"46696c65",
          9058 => x"20616c72",
          9059 => x"65616479",
          9060 => x"20657869",
          9061 => x"7374732e",
          9062 => x"0a000000",
          9063 => x"46696c65",
          9064 => x"2068616e",
          9065 => x"646c6520",
          9066 => x"696e7661",
          9067 => x"6c69642e",
          9068 => x"0a000000",
          9069 => x"53442069",
          9070 => x"73207772",
          9071 => x"69746520",
          9072 => x"70726f74",
          9073 => x"65637465",
          9074 => x"642e0a00",
          9075 => x"44726976",
          9076 => x"65206e75",
          9077 => x"6d626572",
          9078 => x"20697320",
          9079 => x"696e7661",
          9080 => x"6c69642e",
          9081 => x"0a000000",
          9082 => x"4469736b",
          9083 => x"206e6f74",
          9084 => x"20656e61",
          9085 => x"626c6564",
          9086 => x"2e0a0000",
          9087 => x"4e6f2063",
          9088 => x"6f6d7061",
          9089 => x"7469626c",
          9090 => x"65206669",
          9091 => x"6c657379",
          9092 => x"7374656d",
          9093 => x"20666f75",
          9094 => x"6e64206f",
          9095 => x"6e206469",
          9096 => x"736b2e0a",
          9097 => x"00000000",
          9098 => x"466f726d",
          9099 => x"61742061",
          9100 => x"626f7274",
          9101 => x"65642e0a",
          9102 => x"00000000",
          9103 => x"54696d65",
          9104 => x"6f75742c",
          9105 => x"206f7065",
          9106 => x"72617469",
          9107 => x"6f6e2063",
          9108 => x"616e6365",
          9109 => x"6c6c6564",
          9110 => x"2e0a0000",
          9111 => x"46696c65",
          9112 => x"20697320",
          9113 => x"6c6f636b",
          9114 => x"65642e0a",
          9115 => x"00000000",
          9116 => x"496e7375",
          9117 => x"66666963",
          9118 => x"69656e74",
          9119 => x"206d656d",
          9120 => x"6f72792e",
          9121 => x"0a000000",
          9122 => x"546f6f20",
          9123 => x"6d616e79",
          9124 => x"206f7065",
          9125 => x"6e206669",
          9126 => x"6c65732e",
          9127 => x"0a000000",
          9128 => x"50617261",
          9129 => x"6d657465",
          9130 => x"72732069",
          9131 => x"6e636f72",
          9132 => x"72656374",
          9133 => x"2e0a0000",
          9134 => x"53756363",
          9135 => x"6573732e",
          9136 => x"0a000000",
          9137 => x"556e6b6e",
          9138 => x"6f776e20",
          9139 => x"6572726f",
          9140 => x"722e0a00",
          9141 => x"0a256c75",
          9142 => x"20627974",
          9143 => x"65732025",
          9144 => x"73206174",
          9145 => x"20256c75",
          9146 => x"20627974",
          9147 => x"65732f73",
          9148 => x"65632e0a",
          9149 => x"00000000",
          9150 => x"72656164",
          9151 => x"00000000",
          9152 => x"25303858",
          9153 => x"00000000",
          9154 => x"3a202000",
          9155 => x"25303458",
          9156 => x"00000000",
          9157 => x"20202020",
          9158 => x"20202020",
          9159 => x"00000000",
          9160 => x"25303258",
          9161 => x"00000000",
          9162 => x"20200000",
          9163 => x"207c0000",
          9164 => x"7c0d0a00",
          9165 => x"7a4f5300",
          9166 => x"0a2a2a20",
          9167 => x"25732028",
          9168 => x"00000000",
          9169 => x"30322f30",
          9170 => x"352f3230",
          9171 => x"32300000",
          9172 => x"76312e30",
          9173 => x"32000000",
          9174 => x"205a5055",
          9175 => x"2c207265",
          9176 => x"76202530",
          9177 => x"32782920",
          9178 => x"25732025",
          9179 => x"73202a2a",
          9180 => x"0a0a0000",
          9181 => x"5a505520",
          9182 => x"496e7465",
          9183 => x"72727570",
          9184 => x"74204861",
          9185 => x"6e646c65",
          9186 => x"720a0000",
          9187 => x"54696d65",
          9188 => x"7220696e",
          9189 => x"74657272",
          9190 => x"7570740a",
          9191 => x"00000000",
          9192 => x"50533220",
          9193 => x"696e7465",
          9194 => x"72727570",
          9195 => x"740a0000",
          9196 => x"494f4354",
          9197 => x"4c205244",
          9198 => x"20696e74",
          9199 => x"65727275",
          9200 => x"70740a00",
          9201 => x"494f4354",
          9202 => x"4c205752",
          9203 => x"20696e74",
          9204 => x"65727275",
          9205 => x"70740a00",
          9206 => x"55415254",
          9207 => x"30205258",
          9208 => x"20696e74",
          9209 => x"65727275",
          9210 => x"70740a00",
          9211 => x"55415254",
          9212 => x"30205458",
          9213 => x"20696e74",
          9214 => x"65727275",
          9215 => x"70740a00",
          9216 => x"55415254",
          9217 => x"31205258",
          9218 => x"20696e74",
          9219 => x"65727275",
          9220 => x"70740a00",
          9221 => x"55415254",
          9222 => x"31205458",
          9223 => x"20696e74",
          9224 => x"65727275",
          9225 => x"70740a00",
          9226 => x"53657474",
          9227 => x"696e6720",
          9228 => x"75702074",
          9229 => x"696d6572",
          9230 => x"2e2e2e0a",
          9231 => x"00000000",
          9232 => x"456e6162",
          9233 => x"6c696e67",
          9234 => x"2074696d",
          9235 => x"65722e2e",
          9236 => x"2e0a0000",
          9237 => x"6175746f",
          9238 => x"65786563",
          9239 => x"2e626174",
          9240 => x"00000000",
          9241 => x"7a4f532e",
          9242 => x"68737400",
          9243 => x"303a0000",
          9244 => x"4661696c",
          9245 => x"65642074",
          9246 => x"6f20696e",
          9247 => x"69746961",
          9248 => x"6c697365",
          9249 => x"20736420",
          9250 => x"63617264",
          9251 => x"20302c20",
          9252 => x"706c6561",
          9253 => x"73652069",
          9254 => x"6e697420",
          9255 => x"6d616e75",
          9256 => x"616c6c79",
          9257 => x"2e000000",
          9258 => x"2a200000",
          9259 => x"436c6561",
          9260 => x"72696e67",
          9261 => x"2e2e2e2e",
          9262 => x"00000000",
          9263 => x"436f7079",
          9264 => x"696e672e",
          9265 => x"2e2e0000",
          9266 => x"436f6d70",
          9267 => x"6172696e",
          9268 => x"672e2e2e",
          9269 => x"00000000",
          9270 => x"2530386c",
          9271 => x"78282530",
          9272 => x"3878292d",
          9273 => x"3e253038",
          9274 => x"6c782825",
          9275 => x"30387829",
          9276 => x"0a000000",
          9277 => x"44756d70",
          9278 => x"204d656d",
          9279 => x"6f72790a",
          9280 => x"00000000",
          9281 => x"0a436f6d",
          9282 => x"706c6574",
          9283 => x"652e0a00",
          9284 => x"25303858",
          9285 => x"20253032",
          9286 => x"582d0000",
          9287 => x"3f3f3f0a",
          9288 => x"00000000",
          9289 => x"25303858",
          9290 => x"20253034",
          9291 => x"582d0000",
          9292 => x"25303858",
          9293 => x"20253038",
          9294 => x"582d0000",
          9295 => x"45786563",
          9296 => x"7574696e",
          9297 => x"6720636f",
          9298 => x"64652040",
          9299 => x"20253038",
          9300 => x"78202e2e",
          9301 => x"2e0a0000",
          9302 => x"43616c6c",
          9303 => x"696e6720",
          9304 => x"636f6465",
          9305 => x"20402025",
          9306 => x"30387820",
          9307 => x"2e2e2e0a",
          9308 => x"00000000",
          9309 => x"43616c6c",
          9310 => x"20726574",
          9311 => x"75726e65",
          9312 => x"6420636f",
          9313 => x"64652028",
          9314 => x"2564292e",
          9315 => x"0a000000",
          9316 => x"52657374",
          9317 => x"61727469",
          9318 => x"6e672061",
          9319 => x"70706c69",
          9320 => x"63617469",
          9321 => x"6f6e2e2e",
          9322 => x"2e0a0000",
          9323 => x"436f6c64",
          9324 => x"20726562",
          9325 => x"6f6f7469",
          9326 => x"6e672e2e",
          9327 => x"2e0a0000",
          9328 => x"5a505500",
          9329 => x"62696e00",
          9330 => x"25643a5c",
          9331 => x"25735c25",
          9332 => x"732e2573",
          9333 => x"00000000",
          9334 => x"25643a5c",
          9335 => x"25735c25",
          9336 => x"73000000",
          9337 => x"25643a5c",
          9338 => x"25730000",
          9339 => x"42616420",
          9340 => x"636f6d6d",
          9341 => x"616e642e",
          9342 => x"00000000",
          9343 => x"48454c4c",
          9344 => x"4f203120",
          9345 => x"46524f4d",
          9346 => x"20505249",
          9347 => x"4e544600",
          9348 => x"48454c4c",
          9349 => x"4f203220",
          9350 => x"46524f4d",
          9351 => x"20505249",
          9352 => x"4e544600",
          9353 => x"52756e6e",
          9354 => x"696e672e",
          9355 => x"2e2e0a00",
          9356 => x"456e6162",
          9357 => x"6c696e67",
          9358 => x"20696e74",
          9359 => x"65727275",
          9360 => x"7074732e",
          9361 => x"2e2e0a00",
          9362 => x"25642f25",
          9363 => x"642f2564",
          9364 => x"2025643a",
          9365 => x"25643a25",
          9366 => x"642e2564",
          9367 => x"25640a00",
          9368 => x"536f4320",
          9369 => x"436f6e66",
          9370 => x"69677572",
          9371 => x"6174696f",
          9372 => x"6e000000",
          9373 => x"20286672",
          9374 => x"6f6d2053",
          9375 => x"6f432063",
          9376 => x"6f6e6669",
          9377 => x"67290000",
          9378 => x"3a0a4465",
          9379 => x"76696365",
          9380 => x"7320696d",
          9381 => x"706c656d",
          9382 => x"656e7465",
          9383 => x"643a0a00",
          9384 => x"20202020",
          9385 => x"57422053",
          9386 => x"4452414d",
          9387 => x"20202825",
          9388 => x"3038583a",
          9389 => x"25303858",
          9390 => x"292e0a00",
          9391 => x"20202020",
          9392 => x"53445241",
          9393 => x"4d202020",
          9394 => x"20202825",
          9395 => x"3038583a",
          9396 => x"25303858",
          9397 => x"292e0a00",
          9398 => x"20202020",
          9399 => x"494e534e",
          9400 => x"20425241",
          9401 => x"4d202825",
          9402 => x"3038583a",
          9403 => x"25303858",
          9404 => x"292e0a00",
          9405 => x"20202020",
          9406 => x"4252414d",
          9407 => x"20202020",
          9408 => x"20202825",
          9409 => x"3038583a",
          9410 => x"25303858",
          9411 => x"292e0a00",
          9412 => x"20202020",
          9413 => x"52414d20",
          9414 => x"20202020",
          9415 => x"20202825",
          9416 => x"3038583a",
          9417 => x"25303858",
          9418 => x"292e0a00",
          9419 => x"20202020",
          9420 => x"53442043",
          9421 => x"41524420",
          9422 => x"20202844",
          9423 => x"65766963",
          9424 => x"6573203d",
          9425 => x"25303264",
          9426 => x"292e0a00",
          9427 => x"20202020",
          9428 => x"54494d45",
          9429 => x"52312020",
          9430 => x"20202854",
          9431 => x"696d6572",
          9432 => x"7320203d",
          9433 => x"25303264",
          9434 => x"292e0a00",
          9435 => x"20202020",
          9436 => x"494e5452",
          9437 => x"20435452",
          9438 => x"4c202843",
          9439 => x"68616e6e",
          9440 => x"656c733d",
          9441 => x"25303264",
          9442 => x"292e0a00",
          9443 => x"20202020",
          9444 => x"57495348",
          9445 => x"424f4e45",
          9446 => x"20425553",
          9447 => x"0a000000",
          9448 => x"20202020",
          9449 => x"57422049",
          9450 => x"32430a00",
          9451 => x"20202020",
          9452 => x"494f4354",
          9453 => x"4c0a0000",
          9454 => x"20202020",
          9455 => x"5053320a",
          9456 => x"00000000",
          9457 => x"20202020",
          9458 => x"5350490a",
          9459 => x"00000000",
          9460 => x"41646472",
          9461 => x"65737365",
          9462 => x"733a0a00",
          9463 => x"20202020",
          9464 => x"43505520",
          9465 => x"52657365",
          9466 => x"74205665",
          9467 => x"63746f72",
          9468 => x"20416464",
          9469 => x"72657373",
          9470 => x"203d2025",
          9471 => x"3038580a",
          9472 => x"00000000",
          9473 => x"20202020",
          9474 => x"43505520",
          9475 => x"4d656d6f",
          9476 => x"72792053",
          9477 => x"74617274",
          9478 => x"20416464",
          9479 => x"72657373",
          9480 => x"203d2025",
          9481 => x"3038580a",
          9482 => x"00000000",
          9483 => x"20202020",
          9484 => x"53746163",
          9485 => x"6b205374",
          9486 => x"61727420",
          9487 => x"41646472",
          9488 => x"65737320",
          9489 => x"20202020",
          9490 => x"203d2025",
          9491 => x"3038580a",
          9492 => x"00000000",
          9493 => x"4d697363",
          9494 => x"3a0a0000",
          9495 => x"20202020",
          9496 => x"5a505520",
          9497 => x"49642020",
          9498 => x"20202020",
          9499 => x"20202020",
          9500 => x"20202020",
          9501 => x"20202020",
          9502 => x"203d2025",
          9503 => x"3034580a",
          9504 => x"00000000",
          9505 => x"20202020",
          9506 => x"53797374",
          9507 => x"656d2043",
          9508 => x"6c6f636b",
          9509 => x"20467265",
          9510 => x"71202020",
          9511 => x"20202020",
          9512 => x"203d2025",
          9513 => x"642e2530",
          9514 => x"34644d48",
          9515 => x"7a0a0000",
          9516 => x"20202020",
          9517 => x"53445241",
          9518 => x"4d20436c",
          9519 => x"6f636b20",
          9520 => x"46726571",
          9521 => x"20202020",
          9522 => x"20202020",
          9523 => x"203d2025",
          9524 => x"642e2530",
          9525 => x"34644d48",
          9526 => x"7a0a0000",
          9527 => x"20202020",
          9528 => x"57697368",
          9529 => x"626f6e65",
          9530 => x"20534452",
          9531 => x"414d2043",
          9532 => x"6c6f636b",
          9533 => x"20467265",
          9534 => x"713d2025",
          9535 => x"642e2530",
          9536 => x"34644d48",
          9537 => x"7a0a0000",
          9538 => x"536d616c",
          9539 => x"6c000000",
          9540 => x"4d656469",
          9541 => x"756d0000",
          9542 => x"466c6578",
          9543 => x"00000000",
          9544 => x"45564f00",
          9545 => x"45564f6d",
          9546 => x"696e0000",
          9547 => x"556e6b6e",
          9548 => x"6f776e00",
          9549 => x"00009690",
          9550 => x"01000000",
          9551 => x"00000002",
          9552 => x"0000968c",
          9553 => x"01000000",
          9554 => x"00000003",
          9555 => x"00009688",
          9556 => x"01000000",
          9557 => x"00000004",
          9558 => x"00009684",
          9559 => x"01000000",
          9560 => x"00000005",
          9561 => x"00009680",
          9562 => x"01000000",
          9563 => x"00000006",
          9564 => x"0000967c",
          9565 => x"01000000",
          9566 => x"00000007",
          9567 => x"00009678",
          9568 => x"01000000",
          9569 => x"00000001",
          9570 => x"00009674",
          9571 => x"01000000",
          9572 => x"00000008",
          9573 => x"00009670",
          9574 => x"01000000",
          9575 => x"0000000b",
          9576 => x"0000966c",
          9577 => x"01000000",
          9578 => x"00000009",
          9579 => x"00009668",
          9580 => x"01000000",
          9581 => x"0000000a",
          9582 => x"00009664",
          9583 => x"04000000",
          9584 => x"0000000d",
          9585 => x"00009660",
          9586 => x"04000000",
          9587 => x"0000000c",
          9588 => x"0000965c",
          9589 => x"04000000",
          9590 => x"0000000e",
          9591 => x"00009658",
          9592 => x"03000000",
          9593 => x"0000000f",
          9594 => x"00009654",
          9595 => x"04000000",
          9596 => x"0000000f",
          9597 => x"00009650",
          9598 => x"04000000",
          9599 => x"00000010",
          9600 => x"0000964c",
          9601 => x"04000000",
          9602 => x"00000011",
          9603 => x"00009648",
          9604 => x"03000000",
          9605 => x"00000012",
          9606 => x"00009644",
          9607 => x"03000000",
          9608 => x"00000013",
          9609 => x"00009640",
          9610 => x"03000000",
          9611 => x"00000014",
          9612 => x"0000963c",
          9613 => x"03000000",
          9614 => x"00000015",
          9615 => x"1b5b4400",
          9616 => x"1b5b4300",
          9617 => x"1b5b4200",
          9618 => x"1b5b4100",
          9619 => x"1b5b367e",
          9620 => x"1b5b357e",
          9621 => x"1b5b347e",
          9622 => x"1b304600",
          9623 => x"1b5b337e",
          9624 => x"1b5b327e",
          9625 => x"1b5b317e",
          9626 => x"10000000",
          9627 => x"0e000000",
          9628 => x"0d000000",
          9629 => x"0b000000",
          9630 => x"08000000",
          9631 => x"06000000",
          9632 => x"05000000",
          9633 => x"04000000",
          9634 => x"03000000",
          9635 => x"02000000",
          9636 => x"01000000",
          9637 => x"68697374",
          9638 => x"6f727900",
          9639 => x"68697374",
          9640 => x"00000000",
          9641 => x"21000000",
          9642 => x"25303464",
          9643 => x"20202573",
          9644 => x"0a000000",
          9645 => x"4661696c",
          9646 => x"65642074",
          9647 => x"6f207265",
          9648 => x"73657420",
          9649 => x"74686520",
          9650 => x"68697374",
          9651 => x"6f727920",
          9652 => x"66696c65",
          9653 => x"20746f20",
          9654 => x"454f462e",
          9655 => x"0a000000",
          9656 => x"43616e6e",
          9657 => x"6f74206f",
          9658 => x"70656e2f",
          9659 => x"63726561",
          9660 => x"74652068",
          9661 => x"6973746f",
          9662 => x"72792066",
          9663 => x"696c652c",
          9664 => x"20646973",
          9665 => x"61626c69",
          9666 => x"6e672e00",
          9667 => x"53440000",
          9668 => x"222a2b2c",
          9669 => x"3a3b3c3d",
          9670 => x"3e3f5b5d",
          9671 => x"7c7f0000",
          9672 => x"46415400",
          9673 => x"46415433",
          9674 => x"32000000",
          9675 => x"ebfe904d",
          9676 => x"53444f53",
          9677 => x"352e3000",
          9678 => x"4e4f204e",
          9679 => x"414d4520",
          9680 => x"20202046",
          9681 => x"41543332",
          9682 => x"20202000",
          9683 => x"4e4f204e",
          9684 => x"414d4520",
          9685 => x"20202046",
          9686 => x"41542020",
          9687 => x"20202000",
          9688 => x"0000970c",
          9689 => x"00000000",
          9690 => x"00000000",
          9691 => x"00000000",
          9692 => x"809a4541",
          9693 => x"8e418f80",
          9694 => x"45454549",
          9695 => x"49498e8f",
          9696 => x"9092924f",
          9697 => x"994f5555",
          9698 => x"59999a9b",
          9699 => x"9c9d9e9f",
          9700 => x"41494f55",
          9701 => x"a5a5a6a7",
          9702 => x"a8a9aaab",
          9703 => x"acadaeaf",
          9704 => x"b0b1b2b3",
          9705 => x"b4b5b6b7",
          9706 => x"b8b9babb",
          9707 => x"bcbdbebf",
          9708 => x"c0c1c2c3",
          9709 => x"c4c5c6c7",
          9710 => x"c8c9cacb",
          9711 => x"cccdcecf",
          9712 => x"d0d1d2d3",
          9713 => x"d4d5d6d7",
          9714 => x"d8d9dadb",
          9715 => x"dcdddedf",
          9716 => x"e0e1e2e3",
          9717 => x"e4e5e6e7",
          9718 => x"e8e9eaeb",
          9719 => x"ecedeeef",
          9720 => x"f0f1f2f3",
          9721 => x"f4f5f6f7",
          9722 => x"f8f9fafb",
          9723 => x"fcfdfeff",
          9724 => x"2b2e2c3b",
          9725 => x"3d5b5d2f",
          9726 => x"5c222a3a",
          9727 => x"3c3e3f7c",
          9728 => x"7f000000",
          9729 => x"00010004",
          9730 => x"00100040",
          9731 => x"01000200",
          9732 => x"00000000",
          9733 => x"00010002",
          9734 => x"00040008",
          9735 => x"00100020",
          9736 => x"00000000",
          9737 => x"00000000",
          9738 => x"00008c60",
          9739 => x"01020100",
          9740 => x"00000000",
          9741 => x"00000000",
          9742 => x"00008c68",
          9743 => x"01040100",
          9744 => x"00000000",
          9745 => x"00000000",
          9746 => x"00008c70",
          9747 => x"01140300",
          9748 => x"00000000",
          9749 => x"00000000",
          9750 => x"00008c78",
          9751 => x"012b0300",
          9752 => x"00000000",
          9753 => x"00000000",
          9754 => x"00008c80",
          9755 => x"01300300",
          9756 => x"00000000",
          9757 => x"00000000",
          9758 => x"00008c88",
          9759 => x"013c0400",
          9760 => x"00000000",
          9761 => x"00000000",
          9762 => x"00008c90",
          9763 => x"013d0400",
          9764 => x"00000000",
          9765 => x"00000000",
          9766 => x"00008c98",
          9767 => x"013f0400",
          9768 => x"00000000",
          9769 => x"00000000",
          9770 => x"00008ca0",
          9771 => x"01400400",
          9772 => x"00000000",
          9773 => x"00000000",
          9774 => x"00008ca8",
          9775 => x"01410400",
          9776 => x"00000000",
          9777 => x"00000000",
          9778 => x"00008cac",
          9779 => x"01420400",
          9780 => x"00000000",
          9781 => x"00000000",
          9782 => x"00008cb0",
          9783 => x"01430400",
          9784 => x"00000000",
          9785 => x"00000000",
          9786 => x"00008cb4",
          9787 => x"01500500",
          9788 => x"00000000",
          9789 => x"00000000",
          9790 => x"00008cb8",
          9791 => x"01510500",
          9792 => x"00000000",
          9793 => x"00000000",
          9794 => x"00008cbc",
          9795 => x"01540500",
          9796 => x"00000000",
          9797 => x"00000000",
          9798 => x"00008cc0",
          9799 => x"01550500",
          9800 => x"00000000",
          9801 => x"00000000",
          9802 => x"00008cc4",
          9803 => x"01790700",
          9804 => x"00000000",
          9805 => x"00000000",
          9806 => x"00008ccc",
          9807 => x"01780700",
          9808 => x"00000000",
          9809 => x"00000000",
          9810 => x"00008cd0",
          9811 => x"01820800",
          9812 => x"00000000",
          9813 => x"00000000",
          9814 => x"00008cd8",
          9815 => x"01830800",
          9816 => x"00000000",
          9817 => x"00000000",
          9818 => x"00008ce0",
          9819 => x"01850800",
          9820 => x"00000000",
          9821 => x"00000000",
          9822 => x"00008ce8",
          9823 => x"01870800",
          9824 => x"00000000",
          9825 => x"00000000",
          9826 => x"00008cf0",
          9827 => x"018c0900",
          9828 => x"00000000",
          9829 => x"00000000",
          9830 => x"00008cf8",
          9831 => x"018d0900",
          9832 => x"00000000",
          9833 => x"00000000",
          9834 => x"00008d00",
          9835 => x"018e0900",
          9836 => x"00000000",
          9837 => x"00000000",
          9838 => x"00008d08",
          9839 => x"018f0900",
          9840 => x"00000000",
          9841 => x"00000000",
          9842 => x"00000000",
          9843 => x"00000000",
          9844 => x"00007fff",
          9845 => x"00000000",
          9846 => x"00007fff",
          9847 => x"00010000",
          9848 => x"00007fff",
          9849 => x"00010000",
          9850 => x"00810000",
          9851 => x"01000000",
          9852 => x"017fffff",
          9853 => x"00000000",
          9854 => x"00000000",
          9855 => x"00007800",
          9856 => x"00000000",
          9857 => x"05f5e100",
          9858 => x"05f5e100",
          9859 => x"05f5e100",
          9860 => x"00000000",
          9861 => x"01010101",
          9862 => x"01010101",
          9863 => x"01011001",
          9864 => x"01000000",
          9865 => x"00000000",
          9866 => x"00000000",
          9867 => x"00000000",
          9868 => x"00000000",
          9869 => x"00000000",
          9870 => x"00000000",
          9871 => x"00000000",
          9872 => x"00000000",
          9873 => x"00000000",
          9874 => x"00000000",
          9875 => x"00000000",
          9876 => x"00000000",
          9877 => x"00000000",
          9878 => x"00000000",
          9879 => x"00000000",
          9880 => x"00000000",
          9881 => x"00000000",
          9882 => x"00000000",
          9883 => x"00000000",
          9884 => x"00000000",
          9885 => x"00000000",
          9886 => x"00000000",
          9887 => x"00000000",
          9888 => x"00000000",
          9889 => x"00009694",
          9890 => x"01000000",
          9891 => x"0000969c",
          9892 => x"01000000",
          9893 => x"000096a4",
          9894 => x"02000000",
          9895 => x"00000000",
          9896 => x"00000000",
          9897 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

