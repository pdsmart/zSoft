-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"ff",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"80",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"9a",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"c3",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"c5",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"e8",
           386 => x"8d",
           387 => x"e8",
           388 => x"90",
           389 => x"e8",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"82",
           395 => x"82",
           396 => x"82",
           397 => x"af",
           398 => x"bb",
           399 => x"d8",
           400 => x"bb",
           401 => x"ad",
           402 => x"e8",
           403 => x"90",
           404 => x"e8",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"82",
           418 => x"82",
           419 => x"82",
           420 => x"96",
           421 => x"bb",
           422 => x"d8",
           423 => x"bb",
           424 => x"cd",
           425 => x"e8",
           426 => x"90",
           427 => x"e8",
           428 => x"b7",
           429 => x"e8",
           430 => x"90",
           431 => x"e8",
           432 => x"95",
           433 => x"e8",
           434 => x"90",
           435 => x"e8",
           436 => x"d2",
           437 => x"e8",
           438 => x"90",
           439 => x"e8",
           440 => x"c9",
           441 => x"e8",
           442 => x"90",
           443 => x"e8",
           444 => x"fc",
           445 => x"e8",
           446 => x"90",
           447 => x"e8",
           448 => x"f0",
           449 => x"e8",
           450 => x"90",
           451 => x"e8",
           452 => x"e1",
           453 => x"e8",
           454 => x"90",
           455 => x"e8",
           456 => x"d5",
           457 => x"e8",
           458 => x"90",
           459 => x"e8",
           460 => x"d2",
           461 => x"e8",
           462 => x"90",
           463 => x"e8",
           464 => x"f0",
           465 => x"e8",
           466 => x"90",
           467 => x"e8",
           468 => x"d0",
           469 => x"e8",
           470 => x"90",
           471 => x"e8",
           472 => x"c3",
           473 => x"e8",
           474 => x"90",
           475 => x"e8",
           476 => x"8f",
           477 => x"e8",
           478 => x"90",
           479 => x"e8",
           480 => x"ae",
           481 => x"e8",
           482 => x"90",
           483 => x"e8",
           484 => x"cd",
           485 => x"e8",
           486 => x"90",
           487 => x"e8",
           488 => x"b7",
           489 => x"e8",
           490 => x"90",
           491 => x"e8",
           492 => x"9d",
           493 => x"e8",
           494 => x"90",
           495 => x"e8",
           496 => x"8b",
           497 => x"e8",
           498 => x"90",
           499 => x"e8",
           500 => x"d1",
           501 => x"e8",
           502 => x"90",
           503 => x"e8",
           504 => x"8b",
           505 => x"e8",
           506 => x"90",
           507 => x"e8",
           508 => x"8c",
           509 => x"e8",
           510 => x"90",
           511 => x"e8",
           512 => x"c1",
           513 => x"e8",
           514 => x"90",
           515 => x"e8",
           516 => x"9a",
           517 => x"e8",
           518 => x"90",
           519 => x"e8",
           520 => x"c5",
           521 => x"e8",
           522 => x"90",
           523 => x"e8",
           524 => x"a8",
           525 => x"e8",
           526 => x"90",
           527 => x"e8",
           528 => x"fd",
           529 => x"e8",
           530 => x"90",
           531 => x"e8",
           532 => x"87",
           533 => x"e8",
           534 => x"90",
           535 => x"e8",
           536 => x"c9",
           537 => x"e8",
           538 => x"90",
           539 => x"e8",
           540 => x"8f",
           541 => x"e8",
           542 => x"90",
           543 => x"e8",
           544 => x"b5",
           545 => x"e8",
           546 => x"90",
           547 => x"e8",
           548 => x"ea",
           549 => x"e8",
           550 => x"90",
           551 => x"e8",
           552 => x"d6",
           553 => x"e8",
           554 => x"90",
           555 => x"e8",
           556 => x"ca",
           557 => x"e8",
           558 => x"90",
           559 => x"e8",
           560 => x"b4",
           561 => x"e8",
           562 => x"90",
           563 => x"e8",
           564 => x"98",
           565 => x"e8",
           566 => x"90",
           567 => x"e8",
           568 => x"fb",
           569 => x"e8",
           570 => x"90",
           571 => x"e8",
           572 => x"9f",
           573 => x"e8",
           574 => x"90",
           575 => x"e8",
           576 => x"82",
           577 => x"e8",
           578 => x"90",
           579 => x"e8",
           580 => x"98",
           581 => x"e8",
           582 => x"90",
           583 => x"e8",
           584 => x"de",
           585 => x"e8",
           586 => x"90",
           587 => x"e8",
           588 => x"86",
           589 => x"e8",
           590 => x"90",
           591 => x"e8",
           592 => x"fe",
           593 => x"e8",
           594 => x"90",
           595 => x"e8",
           596 => x"c8",
           597 => x"e8",
           598 => x"90",
           599 => x"00",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"00",
           609 => x"ff",
           610 => x"06",
           611 => x"83",
           612 => x"10",
           613 => x"fc",
           614 => x"51",
           615 => x"80",
           616 => x"ff",
           617 => x"06",
           618 => x"52",
           619 => x"0a",
           620 => x"38",
           621 => x"51",
           622 => x"dc",
           623 => x"b8",
           624 => x"80",
           625 => x"05",
           626 => x"0b",
           627 => x"04",
           628 => x"80",
           629 => x"00",
           630 => x"08",
           631 => x"e8",
           632 => x"0d",
           633 => x"08",
           634 => x"82",
           635 => x"fc",
           636 => x"bb",
           637 => x"05",
           638 => x"bb",
           639 => x"05",
           640 => x"d3",
           641 => x"54",
           642 => x"82",
           643 => x"70",
           644 => x"08",
           645 => x"82",
           646 => x"f8",
           647 => x"82",
           648 => x"51",
           649 => x"0d",
           650 => x"0c",
           651 => x"e8",
           652 => x"bb",
           653 => x"3d",
           654 => x"e8",
           655 => x"08",
           656 => x"70",
           657 => x"81",
           658 => x"51",
           659 => x"38",
           660 => x"bb",
           661 => x"05",
           662 => x"38",
           663 => x"0b",
           664 => x"08",
           665 => x"81",
           666 => x"bb",
           667 => x"05",
           668 => x"82",
           669 => x"8c",
           670 => x"0b",
           671 => x"08",
           672 => x"82",
           673 => x"88",
           674 => x"bb",
           675 => x"05",
           676 => x"e8",
           677 => x"08",
           678 => x"f6",
           679 => x"82",
           680 => x"8c",
           681 => x"80",
           682 => x"bb",
           683 => x"05",
           684 => x"90",
           685 => x"dc",
           686 => x"bb",
           687 => x"05",
           688 => x"bb",
           689 => x"05",
           690 => x"09",
           691 => x"38",
           692 => x"bb",
           693 => x"05",
           694 => x"39",
           695 => x"08",
           696 => x"82",
           697 => x"f8",
           698 => x"53",
           699 => x"82",
           700 => x"8c",
           701 => x"05",
           702 => x"08",
           703 => x"82",
           704 => x"fc",
           705 => x"05",
           706 => x"08",
           707 => x"ff",
           708 => x"bb",
           709 => x"05",
           710 => x"72",
           711 => x"e8",
           712 => x"08",
           713 => x"e8",
           714 => x"0c",
           715 => x"e8",
           716 => x"08",
           717 => x"0c",
           718 => x"82",
           719 => x"04",
           720 => x"08",
           721 => x"e8",
           722 => x"0d",
           723 => x"bb",
           724 => x"05",
           725 => x"e8",
           726 => x"08",
           727 => x"08",
           728 => x"fe",
           729 => x"bb",
           730 => x"05",
           731 => x"e8",
           732 => x"70",
           733 => x"08",
           734 => x"82",
           735 => x"fc",
           736 => x"82",
           737 => x"8c",
           738 => x"82",
           739 => x"e0",
           740 => x"51",
           741 => x"3f",
           742 => x"08",
           743 => x"e8",
           744 => x"0c",
           745 => x"08",
           746 => x"82",
           747 => x"88",
           748 => x"51",
           749 => x"34",
           750 => x"08",
           751 => x"70",
           752 => x"0c",
           753 => x"0d",
           754 => x"0c",
           755 => x"e8",
           756 => x"bb",
           757 => x"3d",
           758 => x"e8",
           759 => x"70",
           760 => x"08",
           761 => x"82",
           762 => x"fc",
           763 => x"82",
           764 => x"8c",
           765 => x"82",
           766 => x"88",
           767 => x"54",
           768 => x"bb",
           769 => x"82",
           770 => x"f8",
           771 => x"bb",
           772 => x"05",
           773 => x"bb",
           774 => x"54",
           775 => x"82",
           776 => x"04",
           777 => x"08",
           778 => x"e8",
           779 => x"0d",
           780 => x"bb",
           781 => x"05",
           782 => x"e8",
           783 => x"08",
           784 => x"8c",
           785 => x"bb",
           786 => x"05",
           787 => x"33",
           788 => x"70",
           789 => x"81",
           790 => x"51",
           791 => x"80",
           792 => x"ff",
           793 => x"e8",
           794 => x"0c",
           795 => x"82",
           796 => x"8c",
           797 => x"72",
           798 => x"82",
           799 => x"f8",
           800 => x"81",
           801 => x"72",
           802 => x"fa",
           803 => x"e8",
           804 => x"08",
           805 => x"bb",
           806 => x"05",
           807 => x"e8",
           808 => x"22",
           809 => x"51",
           810 => x"2e",
           811 => x"82",
           812 => x"f8",
           813 => x"af",
           814 => x"fc",
           815 => x"e8",
           816 => x"33",
           817 => x"26",
           818 => x"82",
           819 => x"f8",
           820 => x"72",
           821 => x"81",
           822 => x"38",
           823 => x"08",
           824 => x"70",
           825 => x"98",
           826 => x"53",
           827 => x"82",
           828 => x"e4",
           829 => x"83",
           830 => x"32",
           831 => x"51",
           832 => x"72",
           833 => x"38",
           834 => x"08",
           835 => x"70",
           836 => x"51",
           837 => x"bb",
           838 => x"05",
           839 => x"39",
           840 => x"08",
           841 => x"70",
           842 => x"98",
           843 => x"83",
           844 => x"73",
           845 => x"51",
           846 => x"53",
           847 => x"e8",
           848 => x"34",
           849 => x"08",
           850 => x"54",
           851 => x"08",
           852 => x"70",
           853 => x"51",
           854 => x"82",
           855 => x"e8",
           856 => x"bb",
           857 => x"05",
           858 => x"2b",
           859 => x"51",
           860 => x"80",
           861 => x"80",
           862 => x"bb",
           863 => x"05",
           864 => x"e8",
           865 => x"22",
           866 => x"70",
           867 => x"51",
           868 => x"db",
           869 => x"e8",
           870 => x"33",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"bb",
           876 => x"05",
           877 => x"39",
           878 => x"08",
           879 => x"70",
           880 => x"81",
           881 => x"53",
           882 => x"9d",
           883 => x"e8",
           884 => x"33",
           885 => x"70",
           886 => x"51",
           887 => x"38",
           888 => x"bb",
           889 => x"05",
           890 => x"e8",
           891 => x"33",
           892 => x"bb",
           893 => x"05",
           894 => x"bb",
           895 => x"05",
           896 => x"26",
           897 => x"82",
           898 => x"c4",
           899 => x"82",
           900 => x"d8",
           901 => x"51",
           902 => x"72",
           903 => x"e8",
           904 => x"22",
           905 => x"51",
           906 => x"bb",
           907 => x"05",
           908 => x"e8",
           909 => x"22",
           910 => x"51",
           911 => x"bb",
           912 => x"05",
           913 => x"39",
           914 => x"08",
           915 => x"70",
           916 => x"51",
           917 => x"bb",
           918 => x"05",
           919 => x"39",
           920 => x"08",
           921 => x"70",
           922 => x"51",
           923 => x"bb",
           924 => x"05",
           925 => x"39",
           926 => x"08",
           927 => x"70",
           928 => x"53",
           929 => x"e8",
           930 => x"23",
           931 => x"bb",
           932 => x"05",
           933 => x"39",
           934 => x"08",
           935 => x"70",
           936 => x"53",
           937 => x"e8",
           938 => x"23",
           939 => x"bf",
           940 => x"e8",
           941 => x"34",
           942 => x"08",
           943 => x"ff",
           944 => x"72",
           945 => x"08",
           946 => x"80",
           947 => x"bb",
           948 => x"05",
           949 => x"39",
           950 => x"08",
           951 => x"82",
           952 => x"90",
           953 => x"05",
           954 => x"08",
           955 => x"70",
           956 => x"72",
           957 => x"08",
           958 => x"82",
           959 => x"ec",
           960 => x"11",
           961 => x"82",
           962 => x"ec",
           963 => x"ef",
           964 => x"e8",
           965 => x"08",
           966 => x"08",
           967 => x"84",
           968 => x"e8",
           969 => x"0c",
           970 => x"bb",
           971 => x"05",
           972 => x"e8",
           973 => x"22",
           974 => x"70",
           975 => x"51",
           976 => x"80",
           977 => x"82",
           978 => x"e8",
           979 => x"98",
           980 => x"98",
           981 => x"bb",
           982 => x"05",
           983 => x"a2",
           984 => x"bb",
           985 => x"72",
           986 => x"08",
           987 => x"99",
           988 => x"e8",
           989 => x"08",
           990 => x"3f",
           991 => x"08",
           992 => x"bb",
           993 => x"05",
           994 => x"e8",
           995 => x"22",
           996 => x"e8",
           997 => x"22",
           998 => x"54",
           999 => x"bb",
          1000 => x"05",
          1001 => x"39",
          1002 => x"08",
          1003 => x"82",
          1004 => x"90",
          1005 => x"05",
          1006 => x"08",
          1007 => x"70",
          1008 => x"e8",
          1009 => x"0c",
          1010 => x"08",
          1011 => x"70",
          1012 => x"81",
          1013 => x"51",
          1014 => x"2e",
          1015 => x"bb",
          1016 => x"05",
          1017 => x"2b",
          1018 => x"2c",
          1019 => x"e8",
          1020 => x"08",
          1021 => x"c1",
          1022 => x"dc",
          1023 => x"82",
          1024 => x"f4",
          1025 => x"39",
          1026 => x"08",
          1027 => x"51",
          1028 => x"82",
          1029 => x"53",
          1030 => x"e8",
          1031 => x"23",
          1032 => x"08",
          1033 => x"53",
          1034 => x"08",
          1035 => x"73",
          1036 => x"54",
          1037 => x"e8",
          1038 => x"23",
          1039 => x"82",
          1040 => x"e4",
          1041 => x"82",
          1042 => x"06",
          1043 => x"72",
          1044 => x"38",
          1045 => x"08",
          1046 => x"82",
          1047 => x"90",
          1048 => x"05",
          1049 => x"08",
          1050 => x"70",
          1051 => x"e8",
          1052 => x"0c",
          1053 => x"82",
          1054 => x"90",
          1055 => x"bb",
          1056 => x"05",
          1057 => x"82",
          1058 => x"90",
          1059 => x"08",
          1060 => x"08",
          1061 => x"53",
          1062 => x"08",
          1063 => x"82",
          1064 => x"fc",
          1065 => x"bb",
          1066 => x"05",
          1067 => x"a4",
          1068 => x"e8",
          1069 => x"22",
          1070 => x"51",
          1071 => x"bb",
          1072 => x"05",
          1073 => x"e8",
          1074 => x"08",
          1075 => x"e8",
          1076 => x"0c",
          1077 => x"08",
          1078 => x"70",
          1079 => x"51",
          1080 => x"bb",
          1081 => x"05",
          1082 => x"39",
          1083 => x"bb",
          1084 => x"05",
          1085 => x"82",
          1086 => x"e4",
          1087 => x"80",
          1088 => x"53",
          1089 => x"e8",
          1090 => x"23",
          1091 => x"82",
          1092 => x"f8",
          1093 => x"0b",
          1094 => x"08",
          1095 => x"82",
          1096 => x"e4",
          1097 => x"82",
          1098 => x"06",
          1099 => x"72",
          1100 => x"38",
          1101 => x"08",
          1102 => x"82",
          1103 => x"90",
          1104 => x"05",
          1105 => x"08",
          1106 => x"70",
          1107 => x"e8",
          1108 => x"0c",
          1109 => x"82",
          1110 => x"90",
          1111 => x"bb",
          1112 => x"05",
          1113 => x"82",
          1114 => x"90",
          1115 => x"08",
          1116 => x"08",
          1117 => x"53",
          1118 => x"08",
          1119 => x"82",
          1120 => x"fc",
          1121 => x"bb",
          1122 => x"05",
          1123 => x"06",
          1124 => x"82",
          1125 => x"e4",
          1126 => x"bb",
          1127 => x"bb",
          1128 => x"05",
          1129 => x"e8",
          1130 => x"08",
          1131 => x"08",
          1132 => x"82",
          1133 => x"fc",
          1134 => x"55",
          1135 => x"54",
          1136 => x"3f",
          1137 => x"08",
          1138 => x"34",
          1139 => x"08",
          1140 => x"82",
          1141 => x"d4",
          1142 => x"bb",
          1143 => x"05",
          1144 => x"51",
          1145 => x"27",
          1146 => x"bb",
          1147 => x"05",
          1148 => x"33",
          1149 => x"e8",
          1150 => x"33",
          1151 => x"11",
          1152 => x"72",
          1153 => x"08",
          1154 => x"97",
          1155 => x"e8",
          1156 => x"08",
          1157 => x"b0",
          1158 => x"72",
          1159 => x"08",
          1160 => x"82",
          1161 => x"d4",
          1162 => x"82",
          1163 => x"d0",
          1164 => x"34",
          1165 => x"08",
          1166 => x"81",
          1167 => x"e8",
          1168 => x"0c",
          1169 => x"08",
          1170 => x"70",
          1171 => x"e8",
          1172 => x"08",
          1173 => x"ab",
          1174 => x"dc",
          1175 => x"bb",
          1176 => x"05",
          1177 => x"bb",
          1178 => x"05",
          1179 => x"84",
          1180 => x"39",
          1181 => x"08",
          1182 => x"82",
          1183 => x"55",
          1184 => x"70",
          1185 => x"53",
          1186 => x"e8",
          1187 => x"34",
          1188 => x"08",
          1189 => x"70",
          1190 => x"53",
          1191 => x"94",
          1192 => x"e8",
          1193 => x"22",
          1194 => x"53",
          1195 => x"e8",
          1196 => x"23",
          1197 => x"08",
          1198 => x"70",
          1199 => x"81",
          1200 => x"53",
          1201 => x"80",
          1202 => x"bb",
          1203 => x"05",
          1204 => x"2b",
          1205 => x"08",
          1206 => x"82",
          1207 => x"cc",
          1208 => x"2c",
          1209 => x"08",
          1210 => x"82",
          1211 => x"f4",
          1212 => x"53",
          1213 => x"09",
          1214 => x"38",
          1215 => x"08",
          1216 => x"fe",
          1217 => x"82",
          1218 => x"c8",
          1219 => x"39",
          1220 => x"08",
          1221 => x"ff",
          1222 => x"82",
          1223 => x"c8",
          1224 => x"bb",
          1225 => x"05",
          1226 => x"e8",
          1227 => x"23",
          1228 => x"08",
          1229 => x"70",
          1230 => x"81",
          1231 => x"53",
          1232 => x"80",
          1233 => x"bb",
          1234 => x"05",
          1235 => x"2b",
          1236 => x"82",
          1237 => x"fc",
          1238 => x"51",
          1239 => x"74",
          1240 => x"82",
          1241 => x"e4",
          1242 => x"f7",
          1243 => x"72",
          1244 => x"08",
          1245 => x"9d",
          1246 => x"e8",
          1247 => x"33",
          1248 => x"e8",
          1249 => x"33",
          1250 => x"54",
          1251 => x"bb",
          1252 => x"05",
          1253 => x"e8",
          1254 => x"22",
          1255 => x"70",
          1256 => x"51",
          1257 => x"2e",
          1258 => x"bb",
          1259 => x"05",
          1260 => x"2b",
          1261 => x"70",
          1262 => x"88",
          1263 => x"51",
          1264 => x"54",
          1265 => x"08",
          1266 => x"70",
          1267 => x"53",
          1268 => x"e8",
          1269 => x"23",
          1270 => x"bb",
          1271 => x"05",
          1272 => x"2b",
          1273 => x"70",
          1274 => x"88",
          1275 => x"51",
          1276 => x"54",
          1277 => x"08",
          1278 => x"70",
          1279 => x"53",
          1280 => x"e8",
          1281 => x"23",
          1282 => x"08",
          1283 => x"70",
          1284 => x"51",
          1285 => x"38",
          1286 => x"08",
          1287 => x"ff",
          1288 => x"72",
          1289 => x"08",
          1290 => x"73",
          1291 => x"90",
          1292 => x"80",
          1293 => x"38",
          1294 => x"08",
          1295 => x"52",
          1296 => x"ee",
          1297 => x"82",
          1298 => x"e4",
          1299 => x"81",
          1300 => x"06",
          1301 => x"72",
          1302 => x"38",
          1303 => x"08",
          1304 => x"52",
          1305 => x"ca",
          1306 => x"39",
          1307 => x"08",
          1308 => x"70",
          1309 => x"81",
          1310 => x"53",
          1311 => x"90",
          1312 => x"e8",
          1313 => x"08",
          1314 => x"8a",
          1315 => x"39",
          1316 => x"08",
          1317 => x"70",
          1318 => x"81",
          1319 => x"53",
          1320 => x"8e",
          1321 => x"e8",
          1322 => x"08",
          1323 => x"8a",
          1324 => x"bb",
          1325 => x"05",
          1326 => x"2a",
          1327 => x"51",
          1328 => x"80",
          1329 => x"82",
          1330 => x"88",
          1331 => x"b0",
          1332 => x"3f",
          1333 => x"08",
          1334 => x"53",
          1335 => x"09",
          1336 => x"38",
          1337 => x"08",
          1338 => x"52",
          1339 => x"08",
          1340 => x"51",
          1341 => x"82",
          1342 => x"e4",
          1343 => x"88",
          1344 => x"06",
          1345 => x"72",
          1346 => x"38",
          1347 => x"08",
          1348 => x"ff",
          1349 => x"72",
          1350 => x"08",
          1351 => x"73",
          1352 => x"90",
          1353 => x"80",
          1354 => x"38",
          1355 => x"08",
          1356 => x"52",
          1357 => x"fa",
          1358 => x"82",
          1359 => x"e4",
          1360 => x"83",
          1361 => x"06",
          1362 => x"72",
          1363 => x"38",
          1364 => x"08",
          1365 => x"ff",
          1366 => x"72",
          1367 => x"08",
          1368 => x"73",
          1369 => x"98",
          1370 => x"80",
          1371 => x"38",
          1372 => x"08",
          1373 => x"52",
          1374 => x"b6",
          1375 => x"82",
          1376 => x"e4",
          1377 => x"87",
          1378 => x"06",
          1379 => x"72",
          1380 => x"bb",
          1381 => x"05",
          1382 => x"54",
          1383 => x"bb",
          1384 => x"05",
          1385 => x"2b",
          1386 => x"51",
          1387 => x"25",
          1388 => x"bb",
          1389 => x"05",
          1390 => x"51",
          1391 => x"d2",
          1392 => x"e8",
          1393 => x"33",
          1394 => x"e3",
          1395 => x"06",
          1396 => x"bb",
          1397 => x"05",
          1398 => x"bb",
          1399 => x"05",
          1400 => x"ce",
          1401 => x"39",
          1402 => x"08",
          1403 => x"53",
          1404 => x"2e",
          1405 => x"80",
          1406 => x"bb",
          1407 => x"05",
          1408 => x"51",
          1409 => x"bb",
          1410 => x"05",
          1411 => x"ff",
          1412 => x"72",
          1413 => x"2e",
          1414 => x"82",
          1415 => x"88",
          1416 => x"82",
          1417 => x"fc",
          1418 => x"33",
          1419 => x"e8",
          1420 => x"08",
          1421 => x"bb",
          1422 => x"05",
          1423 => x"f2",
          1424 => x"39",
          1425 => x"08",
          1426 => x"53",
          1427 => x"2e",
          1428 => x"80",
          1429 => x"bb",
          1430 => x"05",
          1431 => x"51",
          1432 => x"bb",
          1433 => x"05",
          1434 => x"ff",
          1435 => x"72",
          1436 => x"2e",
          1437 => x"82",
          1438 => x"88",
          1439 => x"82",
          1440 => x"fc",
          1441 => x"33",
          1442 => x"a6",
          1443 => x"e8",
          1444 => x"08",
          1445 => x"bb",
          1446 => x"05",
          1447 => x"39",
          1448 => x"08",
          1449 => x"82",
          1450 => x"a9",
          1451 => x"e8",
          1452 => x"08",
          1453 => x"e8",
          1454 => x"08",
          1455 => x"bb",
          1456 => x"05",
          1457 => x"e8",
          1458 => x"08",
          1459 => x"53",
          1460 => x"cc",
          1461 => x"e8",
          1462 => x"22",
          1463 => x"70",
          1464 => x"51",
          1465 => x"2e",
          1466 => x"82",
          1467 => x"ec",
          1468 => x"11",
          1469 => x"82",
          1470 => x"ec",
          1471 => x"90",
          1472 => x"2c",
          1473 => x"73",
          1474 => x"82",
          1475 => x"88",
          1476 => x"a0",
          1477 => x"3f",
          1478 => x"bb",
          1479 => x"05",
          1480 => x"bb",
          1481 => x"05",
          1482 => x"86",
          1483 => x"82",
          1484 => x"e4",
          1485 => x"b7",
          1486 => x"e8",
          1487 => x"33",
          1488 => x"2e",
          1489 => x"a8",
          1490 => x"82",
          1491 => x"e4",
          1492 => x"0b",
          1493 => x"08",
          1494 => x"80",
          1495 => x"e8",
          1496 => x"34",
          1497 => x"bb",
          1498 => x"05",
          1499 => x"39",
          1500 => x"08",
          1501 => x"52",
          1502 => x"08",
          1503 => x"51",
          1504 => x"e9",
          1505 => x"bb",
          1506 => x"05",
          1507 => x"08",
          1508 => x"e8",
          1509 => x"0c",
          1510 => x"bb",
          1511 => x"05",
          1512 => x"dc",
          1513 => x"0d",
          1514 => x"0c",
          1515 => x"e8",
          1516 => x"bb",
          1517 => x"3d",
          1518 => x"ac",
          1519 => x"bb",
          1520 => x"05",
          1521 => x"bb",
          1522 => x"05",
          1523 => x"dd",
          1524 => x"dc",
          1525 => x"bb",
          1526 => x"85",
          1527 => x"bb",
          1528 => x"82",
          1529 => x"02",
          1530 => x"0c",
          1531 => x"80",
          1532 => x"e8",
          1533 => x"0c",
          1534 => x"08",
          1535 => x"70",
          1536 => x"81",
          1537 => x"06",
          1538 => x"51",
          1539 => x"2e",
          1540 => x"0b",
          1541 => x"08",
          1542 => x"81",
          1543 => x"bb",
          1544 => x"05",
          1545 => x"33",
          1546 => x"08",
          1547 => x"81",
          1548 => x"e8",
          1549 => x"0c",
          1550 => x"bb",
          1551 => x"05",
          1552 => x"ff",
          1553 => x"80",
          1554 => x"82",
          1555 => x"82",
          1556 => x"53",
          1557 => x"08",
          1558 => x"52",
          1559 => x"51",
          1560 => x"82",
          1561 => x"53",
          1562 => x"ff",
          1563 => x"0b",
          1564 => x"08",
          1565 => x"ff",
          1566 => x"d3",
          1567 => x"d3",
          1568 => x"53",
          1569 => x"13",
          1570 => x"2d",
          1571 => x"08",
          1572 => x"2e",
          1573 => x"0b",
          1574 => x"08",
          1575 => x"82",
          1576 => x"f8",
          1577 => x"82",
          1578 => x"f4",
          1579 => x"82",
          1580 => x"f4",
          1581 => x"bb",
          1582 => x"3d",
          1583 => x"e8",
          1584 => x"bb",
          1585 => x"82",
          1586 => x"fb",
          1587 => x"0b",
          1588 => x"08",
          1589 => x"82",
          1590 => x"8c",
          1591 => x"11",
          1592 => x"2a",
          1593 => x"70",
          1594 => x"51",
          1595 => x"72",
          1596 => x"38",
          1597 => x"bb",
          1598 => x"05",
          1599 => x"39",
          1600 => x"08",
          1601 => x"53",
          1602 => x"bb",
          1603 => x"05",
          1604 => x"82",
          1605 => x"88",
          1606 => x"72",
          1607 => x"08",
          1608 => x"72",
          1609 => x"53",
          1610 => x"b6",
          1611 => x"e8",
          1612 => x"08",
          1613 => x"08",
          1614 => x"53",
          1615 => x"08",
          1616 => x"52",
          1617 => x"51",
          1618 => x"82",
          1619 => x"53",
          1620 => x"ff",
          1621 => x"0b",
          1622 => x"08",
          1623 => x"ff",
          1624 => x"bb",
          1625 => x"05",
          1626 => x"bb",
          1627 => x"05",
          1628 => x"bb",
          1629 => x"05",
          1630 => x"dc",
          1631 => x"0d",
          1632 => x"0c",
          1633 => x"e8",
          1634 => x"bb",
          1635 => x"3d",
          1636 => x"b0",
          1637 => x"bb",
          1638 => x"05",
          1639 => x"3f",
          1640 => x"08",
          1641 => x"dc",
          1642 => x"3d",
          1643 => x"e8",
          1644 => x"bb",
          1645 => x"82",
          1646 => x"fb",
          1647 => x"bb",
          1648 => x"05",
          1649 => x"33",
          1650 => x"70",
          1651 => x"81",
          1652 => x"51",
          1653 => x"80",
          1654 => x"ff",
          1655 => x"e8",
          1656 => x"0c",
          1657 => x"82",
          1658 => x"8c",
          1659 => x"11",
          1660 => x"2a",
          1661 => x"51",
          1662 => x"72",
          1663 => x"db",
          1664 => x"e8",
          1665 => x"08",
          1666 => x"08",
          1667 => x"54",
          1668 => x"08",
          1669 => x"25",
          1670 => x"bb",
          1671 => x"05",
          1672 => x"70",
          1673 => x"08",
          1674 => x"52",
          1675 => x"72",
          1676 => x"08",
          1677 => x"0c",
          1678 => x"08",
          1679 => x"8c",
          1680 => x"05",
          1681 => x"82",
          1682 => x"88",
          1683 => x"82",
          1684 => x"fc",
          1685 => x"53",
          1686 => x"82",
          1687 => x"8c",
          1688 => x"bb",
          1689 => x"05",
          1690 => x"bb",
          1691 => x"05",
          1692 => x"ff",
          1693 => x"12",
          1694 => x"54",
          1695 => x"bb",
          1696 => x"72",
          1697 => x"bb",
          1698 => x"05",
          1699 => x"08",
          1700 => x"12",
          1701 => x"e8",
          1702 => x"08",
          1703 => x"e8",
          1704 => x"0c",
          1705 => x"39",
          1706 => x"bb",
          1707 => x"05",
          1708 => x"e8",
          1709 => x"08",
          1710 => x"0c",
          1711 => x"82",
          1712 => x"04",
          1713 => x"08",
          1714 => x"e8",
          1715 => x"0d",
          1716 => x"08",
          1717 => x"85",
          1718 => x"81",
          1719 => x"06",
          1720 => x"52",
          1721 => x"8d",
          1722 => x"82",
          1723 => x"f8",
          1724 => x"94",
          1725 => x"e8",
          1726 => x"08",
          1727 => x"70",
          1728 => x"81",
          1729 => x"51",
          1730 => x"2e",
          1731 => x"82",
          1732 => x"88",
          1733 => x"bb",
          1734 => x"05",
          1735 => x"85",
          1736 => x"ff",
          1737 => x"52",
          1738 => x"34",
          1739 => x"08",
          1740 => x"8c",
          1741 => x"05",
          1742 => x"82",
          1743 => x"88",
          1744 => x"11",
          1745 => x"bb",
          1746 => x"05",
          1747 => x"52",
          1748 => x"82",
          1749 => x"88",
          1750 => x"11",
          1751 => x"2a",
          1752 => x"51",
          1753 => x"71",
          1754 => x"d7",
          1755 => x"e8",
          1756 => x"08",
          1757 => x"33",
          1758 => x"08",
          1759 => x"51",
          1760 => x"e8",
          1761 => x"08",
          1762 => x"bb",
          1763 => x"05",
          1764 => x"e8",
          1765 => x"08",
          1766 => x"12",
          1767 => x"07",
          1768 => x"85",
          1769 => x"0b",
          1770 => x"08",
          1771 => x"81",
          1772 => x"bb",
          1773 => x"05",
          1774 => x"81",
          1775 => x"52",
          1776 => x"82",
          1777 => x"88",
          1778 => x"bb",
          1779 => x"05",
          1780 => x"11",
          1781 => x"71",
          1782 => x"dc",
          1783 => x"bb",
          1784 => x"05",
          1785 => x"bb",
          1786 => x"05",
          1787 => x"80",
          1788 => x"bb",
          1789 => x"05",
          1790 => x"e8",
          1791 => x"0c",
          1792 => x"08",
          1793 => x"85",
          1794 => x"bb",
          1795 => x"05",
          1796 => x"bb",
          1797 => x"05",
          1798 => x"09",
          1799 => x"38",
          1800 => x"08",
          1801 => x"90",
          1802 => x"82",
          1803 => x"ec",
          1804 => x"39",
          1805 => x"08",
          1806 => x"a0",
          1807 => x"82",
          1808 => x"ec",
          1809 => x"bb",
          1810 => x"05",
          1811 => x"bb",
          1812 => x"05",
          1813 => x"34",
          1814 => x"bb",
          1815 => x"05",
          1816 => x"82",
          1817 => x"88",
          1818 => x"11",
          1819 => x"8c",
          1820 => x"bb",
          1821 => x"05",
          1822 => x"ff",
          1823 => x"bb",
          1824 => x"05",
          1825 => x"52",
          1826 => x"08",
          1827 => x"82",
          1828 => x"89",
          1829 => x"bb",
          1830 => x"82",
          1831 => x"02",
          1832 => x"0c",
          1833 => x"82",
          1834 => x"88",
          1835 => x"bb",
          1836 => x"05",
          1837 => x"e8",
          1838 => x"08",
          1839 => x"08",
          1840 => x"82",
          1841 => x"90",
          1842 => x"2e",
          1843 => x"82",
          1844 => x"f8",
          1845 => x"bb",
          1846 => x"05",
          1847 => x"ac",
          1848 => x"e8",
          1849 => x"08",
          1850 => x"08",
          1851 => x"05",
          1852 => x"e8",
          1853 => x"08",
          1854 => x"90",
          1855 => x"e8",
          1856 => x"08",
          1857 => x"08",
          1858 => x"05",
          1859 => x"08",
          1860 => x"82",
          1861 => x"f8",
          1862 => x"bb",
          1863 => x"05",
          1864 => x"bb",
          1865 => x"05",
          1866 => x"e8",
          1867 => x"08",
          1868 => x"bb",
          1869 => x"05",
          1870 => x"e8",
          1871 => x"08",
          1872 => x"bb",
          1873 => x"05",
          1874 => x"e8",
          1875 => x"08",
          1876 => x"9c",
          1877 => x"e8",
          1878 => x"08",
          1879 => x"bb",
          1880 => x"05",
          1881 => x"e8",
          1882 => x"08",
          1883 => x"bb",
          1884 => x"05",
          1885 => x"e8",
          1886 => x"08",
          1887 => x"08",
          1888 => x"53",
          1889 => x"71",
          1890 => x"39",
          1891 => x"08",
          1892 => x"81",
          1893 => x"e8",
          1894 => x"0c",
          1895 => x"08",
          1896 => x"ff",
          1897 => x"e8",
          1898 => x"0c",
          1899 => x"08",
          1900 => x"80",
          1901 => x"82",
          1902 => x"f8",
          1903 => x"70",
          1904 => x"e8",
          1905 => x"08",
          1906 => x"bb",
          1907 => x"05",
          1908 => x"e8",
          1909 => x"08",
          1910 => x"71",
          1911 => x"e8",
          1912 => x"08",
          1913 => x"bb",
          1914 => x"05",
          1915 => x"39",
          1916 => x"08",
          1917 => x"70",
          1918 => x"0c",
          1919 => x"0d",
          1920 => x"0c",
          1921 => x"e8",
          1922 => x"bb",
          1923 => x"3d",
          1924 => x"e8",
          1925 => x"08",
          1926 => x"08",
          1927 => x"82",
          1928 => x"fc",
          1929 => x"71",
          1930 => x"e8",
          1931 => x"08",
          1932 => x"bb",
          1933 => x"05",
          1934 => x"ff",
          1935 => x"70",
          1936 => x"38",
          1937 => x"bb",
          1938 => x"05",
          1939 => x"82",
          1940 => x"fc",
          1941 => x"bb",
          1942 => x"05",
          1943 => x"e8",
          1944 => x"08",
          1945 => x"bb",
          1946 => x"84",
          1947 => x"bb",
          1948 => x"82",
          1949 => x"02",
          1950 => x"0c",
          1951 => x"82",
          1952 => x"88",
          1953 => x"bb",
          1954 => x"05",
          1955 => x"e8",
          1956 => x"08",
          1957 => x"82",
          1958 => x"8c",
          1959 => x"05",
          1960 => x"08",
          1961 => x"82",
          1962 => x"fc",
          1963 => x"51",
          1964 => x"82",
          1965 => x"fc",
          1966 => x"05",
          1967 => x"08",
          1968 => x"70",
          1969 => x"51",
          1970 => x"84",
          1971 => x"39",
          1972 => x"08",
          1973 => x"70",
          1974 => x"0c",
          1975 => x"0d",
          1976 => x"0c",
          1977 => x"e8",
          1978 => x"bb",
          1979 => x"3d",
          1980 => x"e8",
          1981 => x"08",
          1982 => x"08",
          1983 => x"82",
          1984 => x"8c",
          1985 => x"bb",
          1986 => x"05",
          1987 => x"e8",
          1988 => x"08",
          1989 => x"e5",
          1990 => x"e8",
          1991 => x"08",
          1992 => x"bb",
          1993 => x"05",
          1994 => x"e8",
          1995 => x"08",
          1996 => x"bb",
          1997 => x"05",
          1998 => x"e8",
          1999 => x"08",
          2000 => x"38",
          2001 => x"08",
          2002 => x"51",
          2003 => x"bb",
          2004 => x"05",
          2005 => x"82",
          2006 => x"f8",
          2007 => x"bb",
          2008 => x"05",
          2009 => x"71",
          2010 => x"bb",
          2011 => x"05",
          2012 => x"82",
          2013 => x"fc",
          2014 => x"ad",
          2015 => x"e8",
          2016 => x"08",
          2017 => x"dc",
          2018 => x"3d",
          2019 => x"e8",
          2020 => x"bb",
          2021 => x"82",
          2022 => x"fd",
          2023 => x"bb",
          2024 => x"05",
          2025 => x"81",
          2026 => x"bb",
          2027 => x"05",
          2028 => x"33",
          2029 => x"08",
          2030 => x"81",
          2031 => x"e8",
          2032 => x"0c",
          2033 => x"08",
          2034 => x"70",
          2035 => x"ff",
          2036 => x"54",
          2037 => x"2e",
          2038 => x"ce",
          2039 => x"e8",
          2040 => x"08",
          2041 => x"82",
          2042 => x"88",
          2043 => x"05",
          2044 => x"08",
          2045 => x"70",
          2046 => x"51",
          2047 => x"38",
          2048 => x"bb",
          2049 => x"05",
          2050 => x"39",
          2051 => x"08",
          2052 => x"ff",
          2053 => x"e8",
          2054 => x"0c",
          2055 => x"08",
          2056 => x"80",
          2057 => x"ff",
          2058 => x"bb",
          2059 => x"05",
          2060 => x"80",
          2061 => x"bb",
          2062 => x"05",
          2063 => x"52",
          2064 => x"38",
          2065 => x"bb",
          2066 => x"05",
          2067 => x"39",
          2068 => x"08",
          2069 => x"ff",
          2070 => x"e8",
          2071 => x"0c",
          2072 => x"08",
          2073 => x"70",
          2074 => x"70",
          2075 => x"0b",
          2076 => x"08",
          2077 => x"ae",
          2078 => x"e8",
          2079 => x"08",
          2080 => x"bb",
          2081 => x"05",
          2082 => x"72",
          2083 => x"82",
          2084 => x"fc",
          2085 => x"55",
          2086 => x"8a",
          2087 => x"82",
          2088 => x"fc",
          2089 => x"bb",
          2090 => x"05",
          2091 => x"dc",
          2092 => x"0d",
          2093 => x"0c",
          2094 => x"e8",
          2095 => x"bb",
          2096 => x"3d",
          2097 => x"e8",
          2098 => x"08",
          2099 => x"08",
          2100 => x"82",
          2101 => x"8c",
          2102 => x"38",
          2103 => x"bb",
          2104 => x"05",
          2105 => x"39",
          2106 => x"08",
          2107 => x"52",
          2108 => x"bb",
          2109 => x"05",
          2110 => x"82",
          2111 => x"f8",
          2112 => x"81",
          2113 => x"51",
          2114 => x"9f",
          2115 => x"e8",
          2116 => x"08",
          2117 => x"bb",
          2118 => x"05",
          2119 => x"e8",
          2120 => x"08",
          2121 => x"38",
          2122 => x"82",
          2123 => x"f8",
          2124 => x"05",
          2125 => x"08",
          2126 => x"82",
          2127 => x"f8",
          2128 => x"bb",
          2129 => x"05",
          2130 => x"82",
          2131 => x"fc",
          2132 => x"82",
          2133 => x"fc",
          2134 => x"bb",
          2135 => x"3d",
          2136 => x"e8",
          2137 => x"bb",
          2138 => x"82",
          2139 => x"fe",
          2140 => x"bb",
          2141 => x"05",
          2142 => x"e8",
          2143 => x"0c",
          2144 => x"08",
          2145 => x"80",
          2146 => x"38",
          2147 => x"08",
          2148 => x"81",
          2149 => x"e8",
          2150 => x"0c",
          2151 => x"08",
          2152 => x"ff",
          2153 => x"e8",
          2154 => x"0c",
          2155 => x"08",
          2156 => x"80",
          2157 => x"82",
          2158 => x"8c",
          2159 => x"70",
          2160 => x"08",
          2161 => x"52",
          2162 => x"34",
          2163 => x"08",
          2164 => x"81",
          2165 => x"e8",
          2166 => x"0c",
          2167 => x"82",
          2168 => x"88",
          2169 => x"82",
          2170 => x"51",
          2171 => x"82",
          2172 => x"04",
          2173 => x"08",
          2174 => x"e8",
          2175 => x"0d",
          2176 => x"bb",
          2177 => x"05",
          2178 => x"e8",
          2179 => x"08",
          2180 => x"38",
          2181 => x"08",
          2182 => x"30",
          2183 => x"08",
          2184 => x"80",
          2185 => x"e8",
          2186 => x"0c",
          2187 => x"08",
          2188 => x"8a",
          2189 => x"82",
          2190 => x"f4",
          2191 => x"bb",
          2192 => x"05",
          2193 => x"e8",
          2194 => x"0c",
          2195 => x"08",
          2196 => x"80",
          2197 => x"82",
          2198 => x"8c",
          2199 => x"82",
          2200 => x"8c",
          2201 => x"0b",
          2202 => x"08",
          2203 => x"82",
          2204 => x"fc",
          2205 => x"38",
          2206 => x"bb",
          2207 => x"05",
          2208 => x"e8",
          2209 => x"08",
          2210 => x"08",
          2211 => x"80",
          2212 => x"e8",
          2213 => x"08",
          2214 => x"e8",
          2215 => x"08",
          2216 => x"3f",
          2217 => x"08",
          2218 => x"e8",
          2219 => x"0c",
          2220 => x"e8",
          2221 => x"08",
          2222 => x"38",
          2223 => x"08",
          2224 => x"30",
          2225 => x"08",
          2226 => x"82",
          2227 => x"f8",
          2228 => x"82",
          2229 => x"54",
          2230 => x"82",
          2231 => x"04",
          2232 => x"08",
          2233 => x"e8",
          2234 => x"0d",
          2235 => x"bb",
          2236 => x"05",
          2237 => x"e8",
          2238 => x"08",
          2239 => x"38",
          2240 => x"08",
          2241 => x"30",
          2242 => x"08",
          2243 => x"81",
          2244 => x"e8",
          2245 => x"0c",
          2246 => x"08",
          2247 => x"80",
          2248 => x"82",
          2249 => x"8c",
          2250 => x"82",
          2251 => x"8c",
          2252 => x"53",
          2253 => x"08",
          2254 => x"52",
          2255 => x"08",
          2256 => x"51",
          2257 => x"82",
          2258 => x"70",
          2259 => x"08",
          2260 => x"54",
          2261 => x"08",
          2262 => x"80",
          2263 => x"82",
          2264 => x"f8",
          2265 => x"82",
          2266 => x"f8",
          2267 => x"bb",
          2268 => x"05",
          2269 => x"bb",
          2270 => x"87",
          2271 => x"bb",
          2272 => x"82",
          2273 => x"02",
          2274 => x"0c",
          2275 => x"80",
          2276 => x"e8",
          2277 => x"08",
          2278 => x"e8",
          2279 => x"08",
          2280 => x"3f",
          2281 => x"08",
          2282 => x"dc",
          2283 => x"3d",
          2284 => x"e8",
          2285 => x"bb",
          2286 => x"82",
          2287 => x"fd",
          2288 => x"53",
          2289 => x"08",
          2290 => x"52",
          2291 => x"08",
          2292 => x"51",
          2293 => x"bb",
          2294 => x"82",
          2295 => x"54",
          2296 => x"82",
          2297 => x"04",
          2298 => x"08",
          2299 => x"e8",
          2300 => x"0d",
          2301 => x"bb",
          2302 => x"05",
          2303 => x"82",
          2304 => x"f8",
          2305 => x"bb",
          2306 => x"05",
          2307 => x"e8",
          2308 => x"08",
          2309 => x"82",
          2310 => x"fc",
          2311 => x"2e",
          2312 => x"0b",
          2313 => x"08",
          2314 => x"24",
          2315 => x"bb",
          2316 => x"05",
          2317 => x"bb",
          2318 => x"05",
          2319 => x"e8",
          2320 => x"08",
          2321 => x"e8",
          2322 => x"0c",
          2323 => x"82",
          2324 => x"fc",
          2325 => x"2e",
          2326 => x"82",
          2327 => x"8c",
          2328 => x"bb",
          2329 => x"05",
          2330 => x"38",
          2331 => x"08",
          2332 => x"82",
          2333 => x"8c",
          2334 => x"82",
          2335 => x"88",
          2336 => x"bb",
          2337 => x"05",
          2338 => x"e8",
          2339 => x"08",
          2340 => x"e8",
          2341 => x"0c",
          2342 => x"08",
          2343 => x"81",
          2344 => x"e8",
          2345 => x"0c",
          2346 => x"08",
          2347 => x"81",
          2348 => x"e8",
          2349 => x"0c",
          2350 => x"82",
          2351 => x"90",
          2352 => x"2e",
          2353 => x"bb",
          2354 => x"05",
          2355 => x"bb",
          2356 => x"05",
          2357 => x"39",
          2358 => x"08",
          2359 => x"70",
          2360 => x"08",
          2361 => x"51",
          2362 => x"08",
          2363 => x"82",
          2364 => x"85",
          2365 => x"bb",
          2366 => x"82",
          2367 => x"02",
          2368 => x"0c",
          2369 => x"80",
          2370 => x"e8",
          2371 => x"34",
          2372 => x"08",
          2373 => x"53",
          2374 => x"82",
          2375 => x"88",
          2376 => x"08",
          2377 => x"33",
          2378 => x"bb",
          2379 => x"05",
          2380 => x"ff",
          2381 => x"a0",
          2382 => x"06",
          2383 => x"bb",
          2384 => x"05",
          2385 => x"81",
          2386 => x"53",
          2387 => x"bb",
          2388 => x"05",
          2389 => x"ad",
          2390 => x"06",
          2391 => x"0b",
          2392 => x"08",
          2393 => x"82",
          2394 => x"88",
          2395 => x"08",
          2396 => x"0c",
          2397 => x"53",
          2398 => x"bb",
          2399 => x"05",
          2400 => x"e8",
          2401 => x"33",
          2402 => x"2e",
          2403 => x"81",
          2404 => x"bb",
          2405 => x"05",
          2406 => x"81",
          2407 => x"70",
          2408 => x"72",
          2409 => x"e8",
          2410 => x"34",
          2411 => x"08",
          2412 => x"82",
          2413 => x"e8",
          2414 => x"bb",
          2415 => x"05",
          2416 => x"2e",
          2417 => x"bb",
          2418 => x"05",
          2419 => x"2e",
          2420 => x"cd",
          2421 => x"82",
          2422 => x"f4",
          2423 => x"bb",
          2424 => x"05",
          2425 => x"81",
          2426 => x"70",
          2427 => x"72",
          2428 => x"e8",
          2429 => x"34",
          2430 => x"82",
          2431 => x"e8",
          2432 => x"34",
          2433 => x"08",
          2434 => x"70",
          2435 => x"71",
          2436 => x"51",
          2437 => x"82",
          2438 => x"f8",
          2439 => x"fe",
          2440 => x"e8",
          2441 => x"33",
          2442 => x"26",
          2443 => x"0b",
          2444 => x"08",
          2445 => x"83",
          2446 => x"bb",
          2447 => x"05",
          2448 => x"73",
          2449 => x"82",
          2450 => x"f8",
          2451 => x"72",
          2452 => x"38",
          2453 => x"0b",
          2454 => x"08",
          2455 => x"82",
          2456 => x"0b",
          2457 => x"08",
          2458 => x"b2",
          2459 => x"e8",
          2460 => x"33",
          2461 => x"27",
          2462 => x"bb",
          2463 => x"05",
          2464 => x"b9",
          2465 => x"8d",
          2466 => x"82",
          2467 => x"ec",
          2468 => x"a5",
          2469 => x"82",
          2470 => x"f4",
          2471 => x"0b",
          2472 => x"08",
          2473 => x"82",
          2474 => x"f8",
          2475 => x"a0",
          2476 => x"cf",
          2477 => x"e8",
          2478 => x"33",
          2479 => x"73",
          2480 => x"82",
          2481 => x"f8",
          2482 => x"11",
          2483 => x"82",
          2484 => x"f8",
          2485 => x"bb",
          2486 => x"05",
          2487 => x"51",
          2488 => x"bb",
          2489 => x"05",
          2490 => x"e8",
          2491 => x"33",
          2492 => x"27",
          2493 => x"bb",
          2494 => x"05",
          2495 => x"51",
          2496 => x"bb",
          2497 => x"05",
          2498 => x"e8",
          2499 => x"33",
          2500 => x"26",
          2501 => x"0b",
          2502 => x"08",
          2503 => x"81",
          2504 => x"bb",
          2505 => x"05",
          2506 => x"e8",
          2507 => x"33",
          2508 => x"74",
          2509 => x"80",
          2510 => x"e8",
          2511 => x"0c",
          2512 => x"82",
          2513 => x"f4",
          2514 => x"82",
          2515 => x"fc",
          2516 => x"82",
          2517 => x"f8",
          2518 => x"12",
          2519 => x"08",
          2520 => x"82",
          2521 => x"88",
          2522 => x"08",
          2523 => x"0c",
          2524 => x"51",
          2525 => x"72",
          2526 => x"e8",
          2527 => x"34",
          2528 => x"82",
          2529 => x"f0",
          2530 => x"72",
          2531 => x"38",
          2532 => x"08",
          2533 => x"30",
          2534 => x"08",
          2535 => x"82",
          2536 => x"8c",
          2537 => x"bb",
          2538 => x"05",
          2539 => x"53",
          2540 => x"bb",
          2541 => x"05",
          2542 => x"e8",
          2543 => x"08",
          2544 => x"0c",
          2545 => x"82",
          2546 => x"04",
          2547 => x"08",
          2548 => x"e8",
          2549 => x"0d",
          2550 => x"bb",
          2551 => x"05",
          2552 => x"e8",
          2553 => x"08",
          2554 => x"0c",
          2555 => x"08",
          2556 => x"70",
          2557 => x"72",
          2558 => x"82",
          2559 => x"f8",
          2560 => x"81",
          2561 => x"72",
          2562 => x"81",
          2563 => x"82",
          2564 => x"88",
          2565 => x"08",
          2566 => x"0c",
          2567 => x"82",
          2568 => x"f8",
          2569 => x"72",
          2570 => x"81",
          2571 => x"81",
          2572 => x"e8",
          2573 => x"34",
          2574 => x"08",
          2575 => x"70",
          2576 => x"71",
          2577 => x"51",
          2578 => x"82",
          2579 => x"f8",
          2580 => x"bb",
          2581 => x"05",
          2582 => x"b0",
          2583 => x"06",
          2584 => x"82",
          2585 => x"88",
          2586 => x"08",
          2587 => x"0c",
          2588 => x"53",
          2589 => x"bb",
          2590 => x"05",
          2591 => x"e8",
          2592 => x"33",
          2593 => x"08",
          2594 => x"82",
          2595 => x"e8",
          2596 => x"e2",
          2597 => x"82",
          2598 => x"e8",
          2599 => x"f8",
          2600 => x"80",
          2601 => x"0b",
          2602 => x"08",
          2603 => x"82",
          2604 => x"88",
          2605 => x"08",
          2606 => x"0c",
          2607 => x"53",
          2608 => x"bb",
          2609 => x"05",
          2610 => x"39",
          2611 => x"bb",
          2612 => x"05",
          2613 => x"e8",
          2614 => x"08",
          2615 => x"05",
          2616 => x"08",
          2617 => x"33",
          2618 => x"08",
          2619 => x"80",
          2620 => x"bb",
          2621 => x"05",
          2622 => x"a0",
          2623 => x"81",
          2624 => x"e8",
          2625 => x"0c",
          2626 => x"82",
          2627 => x"f8",
          2628 => x"af",
          2629 => x"38",
          2630 => x"08",
          2631 => x"53",
          2632 => x"83",
          2633 => x"80",
          2634 => x"e8",
          2635 => x"0c",
          2636 => x"88",
          2637 => x"e8",
          2638 => x"34",
          2639 => x"bb",
          2640 => x"05",
          2641 => x"73",
          2642 => x"82",
          2643 => x"f8",
          2644 => x"72",
          2645 => x"38",
          2646 => x"0b",
          2647 => x"08",
          2648 => x"82",
          2649 => x"0b",
          2650 => x"08",
          2651 => x"80",
          2652 => x"e8",
          2653 => x"0c",
          2654 => x"08",
          2655 => x"53",
          2656 => x"81",
          2657 => x"bb",
          2658 => x"05",
          2659 => x"e0",
          2660 => x"38",
          2661 => x"08",
          2662 => x"e0",
          2663 => x"72",
          2664 => x"08",
          2665 => x"82",
          2666 => x"f8",
          2667 => x"11",
          2668 => x"82",
          2669 => x"f8",
          2670 => x"bb",
          2671 => x"05",
          2672 => x"73",
          2673 => x"82",
          2674 => x"f8",
          2675 => x"11",
          2676 => x"82",
          2677 => x"f8",
          2678 => x"bb",
          2679 => x"05",
          2680 => x"89",
          2681 => x"80",
          2682 => x"e8",
          2683 => x"0c",
          2684 => x"82",
          2685 => x"f8",
          2686 => x"bb",
          2687 => x"05",
          2688 => x"72",
          2689 => x"38",
          2690 => x"bb",
          2691 => x"05",
          2692 => x"39",
          2693 => x"08",
          2694 => x"70",
          2695 => x"08",
          2696 => x"29",
          2697 => x"08",
          2698 => x"70",
          2699 => x"e8",
          2700 => x"0c",
          2701 => x"08",
          2702 => x"70",
          2703 => x"71",
          2704 => x"51",
          2705 => x"53",
          2706 => x"bb",
          2707 => x"05",
          2708 => x"39",
          2709 => x"08",
          2710 => x"53",
          2711 => x"90",
          2712 => x"e8",
          2713 => x"08",
          2714 => x"e8",
          2715 => x"0c",
          2716 => x"08",
          2717 => x"82",
          2718 => x"fc",
          2719 => x"0c",
          2720 => x"82",
          2721 => x"ec",
          2722 => x"bb",
          2723 => x"05",
          2724 => x"dc",
          2725 => x"0d",
          2726 => x"0c",
          2727 => x"0d",
          2728 => x"70",
          2729 => x"74",
          2730 => x"e3",
          2731 => x"75",
          2732 => x"d1",
          2733 => x"dc",
          2734 => x"0c",
          2735 => x"54",
          2736 => x"74",
          2737 => x"a0",
          2738 => x"06",
          2739 => x"15",
          2740 => x"80",
          2741 => x"29",
          2742 => x"05",
          2743 => x"56",
          2744 => x"82",
          2745 => x"53",
          2746 => x"08",
          2747 => x"3f",
          2748 => x"08",
          2749 => x"16",
          2750 => x"81",
          2751 => x"38",
          2752 => x"81",
          2753 => x"54",
          2754 => x"c9",
          2755 => x"73",
          2756 => x"0c",
          2757 => x"04",
          2758 => x"73",
          2759 => x"26",
          2760 => x"71",
          2761 => x"9a",
          2762 => x"71",
          2763 => x"9f",
          2764 => x"80",
          2765 => x"f4",
          2766 => x"39",
          2767 => x"51",
          2768 => x"82",
          2769 => x"80",
          2770 => x"a0",
          2771 => x"e4",
          2772 => x"b4",
          2773 => x"39",
          2774 => x"51",
          2775 => x"82",
          2776 => x"80",
          2777 => x"a0",
          2778 => x"c8",
          2779 => x"88",
          2780 => x"39",
          2781 => x"51",
          2782 => x"a1",
          2783 => x"39",
          2784 => x"51",
          2785 => x"a1",
          2786 => x"39",
          2787 => x"51",
          2788 => x"a2",
          2789 => x"39",
          2790 => x"51",
          2791 => x"a2",
          2792 => x"39",
          2793 => x"51",
          2794 => x"a3",
          2795 => x"39",
          2796 => x"51",
          2797 => x"83",
          2798 => x"fb",
          2799 => x"79",
          2800 => x"87",
          2801 => x"38",
          2802 => x"87",
          2803 => x"90",
          2804 => x"52",
          2805 => x"ab",
          2806 => x"dc",
          2807 => x"51",
          2808 => x"82",
          2809 => x"54",
          2810 => x"52",
          2811 => x"51",
          2812 => x"3f",
          2813 => x"04",
          2814 => x"66",
          2815 => x"80",
          2816 => x"5b",
          2817 => x"78",
          2818 => x"07",
          2819 => x"57",
          2820 => x"56",
          2821 => x"26",
          2822 => x"56",
          2823 => x"70",
          2824 => x"51",
          2825 => x"74",
          2826 => x"81",
          2827 => x"8c",
          2828 => x"56",
          2829 => x"3f",
          2830 => x"08",
          2831 => x"dc",
          2832 => x"82",
          2833 => x"87",
          2834 => x"0c",
          2835 => x"08",
          2836 => x"d4",
          2837 => x"80",
          2838 => x"75",
          2839 => x"f5",
          2840 => x"dc",
          2841 => x"bb",
          2842 => x"38",
          2843 => x"80",
          2844 => x"74",
          2845 => x"59",
          2846 => x"96",
          2847 => x"51",
          2848 => x"3f",
          2849 => x"78",
          2850 => x"7b",
          2851 => x"2a",
          2852 => x"57",
          2853 => x"80",
          2854 => x"82",
          2855 => x"87",
          2856 => x"08",
          2857 => x"fe",
          2858 => x"56",
          2859 => x"dc",
          2860 => x"0d",
          2861 => x"0d",
          2862 => x"05",
          2863 => x"58",
          2864 => x"80",
          2865 => x"7a",
          2866 => x"3f",
          2867 => x"08",
          2868 => x"80",
          2869 => x"76",
          2870 => x"38",
          2871 => x"d3",
          2872 => x"55",
          2873 => x"bb",
          2874 => x"52",
          2875 => x"2d",
          2876 => x"08",
          2877 => x"78",
          2878 => x"bb",
          2879 => x"3d",
          2880 => x"3d",
          2881 => x"63",
          2882 => x"80",
          2883 => x"73",
          2884 => x"41",
          2885 => x"5e",
          2886 => x"52",
          2887 => x"51",
          2888 => x"3f",
          2889 => x"51",
          2890 => x"3f",
          2891 => x"79",
          2892 => x"38",
          2893 => x"89",
          2894 => x"2e",
          2895 => x"c6",
          2896 => x"53",
          2897 => x"8e",
          2898 => x"52",
          2899 => x"51",
          2900 => x"3f",
          2901 => x"a3",
          2902 => x"b8",
          2903 => x"15",
          2904 => x"39",
          2905 => x"72",
          2906 => x"38",
          2907 => x"82",
          2908 => x"ff",
          2909 => x"89",
          2910 => x"dc",
          2911 => x"d8",
          2912 => x"55",
          2913 => x"18",
          2914 => x"27",
          2915 => x"33",
          2916 => x"e8",
          2917 => x"c0",
          2918 => x"82",
          2919 => x"ff",
          2920 => x"81",
          2921 => x"d3",
          2922 => x"a0",
          2923 => x"3f",
          2924 => x"82",
          2925 => x"ff",
          2926 => x"80",
          2927 => x"27",
          2928 => x"74",
          2929 => x"55",
          2930 => x"72",
          2931 => x"38",
          2932 => x"53",
          2933 => x"83",
          2934 => x"75",
          2935 => x"81",
          2936 => x"53",
          2937 => x"90",
          2938 => x"fe",
          2939 => x"82",
          2940 => x"52",
          2941 => x"39",
          2942 => x"08",
          2943 => x"d7",
          2944 => x"15",
          2945 => x"39",
          2946 => x"51",
          2947 => x"78",
          2948 => x"5c",
          2949 => x"3f",
          2950 => x"08",
          2951 => x"98",
          2952 => x"76",
          2953 => x"81",
          2954 => x"a0",
          2955 => x"bb",
          2956 => x"2b",
          2957 => x"70",
          2958 => x"30",
          2959 => x"70",
          2960 => x"07",
          2961 => x"06",
          2962 => x"59",
          2963 => x"80",
          2964 => x"38",
          2965 => x"09",
          2966 => x"38",
          2967 => x"39",
          2968 => x"72",
          2969 => x"b2",
          2970 => x"72",
          2971 => x"0c",
          2972 => x"04",
          2973 => x"02",
          2974 => x"82",
          2975 => x"82",
          2976 => x"55",
          2977 => x"3f",
          2978 => x"22",
          2979 => x"3f",
          2980 => x"54",
          2981 => x"53",
          2982 => x"33",
          2983 => x"a4",
          2984 => x"b4",
          2985 => x"2e",
          2986 => x"8b",
          2987 => x"0d",
          2988 => x"0d",
          2989 => x"80",
          2990 => x"b6",
          2991 => x"9c",
          2992 => x"a4",
          2993 => x"d6",
          2994 => x"9c",
          2995 => x"81",
          2996 => x"06",
          2997 => x"80",
          2998 => x"81",
          2999 => x"3f",
          3000 => x"51",
          3001 => x"80",
          3002 => x"3f",
          3003 => x"70",
          3004 => x"52",
          3005 => x"92",
          3006 => x"9c",
          3007 => x"a4",
          3008 => x"9a",
          3009 => x"9b",
          3010 => x"83",
          3011 => x"06",
          3012 => x"80",
          3013 => x"81",
          3014 => x"3f",
          3015 => x"51",
          3016 => x"80",
          3017 => x"3f",
          3018 => x"70",
          3019 => x"52",
          3020 => x"92",
          3021 => x"9b",
          3022 => x"a5",
          3023 => x"de",
          3024 => x"9b",
          3025 => x"85",
          3026 => x"06",
          3027 => x"80",
          3028 => x"81",
          3029 => x"3f",
          3030 => x"51",
          3031 => x"80",
          3032 => x"3f",
          3033 => x"70",
          3034 => x"52",
          3035 => x"92",
          3036 => x"9b",
          3037 => x"a5",
          3038 => x"a2",
          3039 => x"9b",
          3040 => x"87",
          3041 => x"06",
          3042 => x"80",
          3043 => x"81",
          3044 => x"3f",
          3045 => x"51",
          3046 => x"80",
          3047 => x"3f",
          3048 => x"70",
          3049 => x"52",
          3050 => x"92",
          3051 => x"9a",
          3052 => x"a5",
          3053 => x"e6",
          3054 => x"9a",
          3055 => x"ba",
          3056 => x"0d",
          3057 => x"0d",
          3058 => x"05",
          3059 => x"70",
          3060 => x"80",
          3061 => x"e3",
          3062 => x"0b",
          3063 => x"33",
          3064 => x"38",
          3065 => x"a6",
          3066 => x"d2",
          3067 => x"fc",
          3068 => x"bb",
          3069 => x"70",
          3070 => x"08",
          3071 => x"82",
          3072 => x"51",
          3073 => x"0b",
          3074 => x"34",
          3075 => x"b6",
          3076 => x"73",
          3077 => x"81",
          3078 => x"82",
          3079 => x"74",
          3080 => x"81",
          3081 => x"82",
          3082 => x"80",
          3083 => x"82",
          3084 => x"51",
          3085 => x"91",
          3086 => x"dc",
          3087 => x"a1",
          3088 => x"0b",
          3089 => x"d8",
          3090 => x"82",
          3091 => x"54",
          3092 => x"09",
          3093 => x"38",
          3094 => x"53",
          3095 => x"51",
          3096 => x"80",
          3097 => x"dc",
          3098 => x"0d",
          3099 => x"0d",
          3100 => x"82",
          3101 => x"5f",
          3102 => x"7c",
          3103 => x"cb",
          3104 => x"dc",
          3105 => x"06",
          3106 => x"2e",
          3107 => x"a3",
          3108 => x"59",
          3109 => x"a6",
          3110 => x"51",
          3111 => x"7c",
          3112 => x"82",
          3113 => x"80",
          3114 => x"82",
          3115 => x"7d",
          3116 => x"82",
          3117 => x"91",
          3118 => x"70",
          3119 => x"a6",
          3120 => x"b2",
          3121 => x"3d",
          3122 => x"80",
          3123 => x"51",
          3124 => x"b4",
          3125 => x"05",
          3126 => x"3f",
          3127 => x"08",
          3128 => x"90",
          3129 => x"78",
          3130 => x"89",
          3131 => x"80",
          3132 => x"d9",
          3133 => x"2e",
          3134 => x"78",
          3135 => x"38",
          3136 => x"81",
          3137 => x"82",
          3138 => x"78",
          3139 => x"ae",
          3140 => x"39",
          3141 => x"82",
          3142 => x"94",
          3143 => x"38",
          3144 => x"78",
          3145 => x"fc",
          3146 => x"24",
          3147 => x"b0",
          3148 => x"38",
          3149 => x"84",
          3150 => x"d7",
          3151 => x"2e",
          3152 => x"78",
          3153 => x"86",
          3154 => x"c7",
          3155 => x"d5",
          3156 => x"38",
          3157 => x"24",
          3158 => x"80",
          3159 => x"d9",
          3160 => x"d0",
          3161 => x"78",
          3162 => x"89",
          3163 => x"80",
          3164 => x"a5",
          3165 => x"39",
          3166 => x"2e",
          3167 => x"78",
          3168 => x"8c",
          3169 => x"8b",
          3170 => x"82",
          3171 => x"38",
          3172 => x"24",
          3173 => x"80",
          3174 => x"f4",
          3175 => x"f9",
          3176 => x"38",
          3177 => x"78",
          3178 => x"8d",
          3179 => x"81",
          3180 => x"d9",
          3181 => x"39",
          3182 => x"80",
          3183 => x"84",
          3184 => x"88",
          3185 => x"dc",
          3186 => x"82",
          3187 => x"8f",
          3188 => x"3d",
          3189 => x"53",
          3190 => x"51",
          3191 => x"82",
          3192 => x"80",
          3193 => x"81",
          3194 => x"38",
          3195 => x"80",
          3196 => x"52",
          3197 => x"05",
          3198 => x"c8",
          3199 => x"bb",
          3200 => x"ff",
          3201 => x"8d",
          3202 => x"84",
          3203 => x"3f",
          3204 => x"aa",
          3205 => x"94",
          3206 => x"39",
          3207 => x"80",
          3208 => x"84",
          3209 => x"a4",
          3210 => x"dc",
          3211 => x"fd",
          3212 => x"53",
          3213 => x"80",
          3214 => x"51",
          3215 => x"3f",
          3216 => x"08",
          3217 => x"ac",
          3218 => x"39",
          3219 => x"80",
          3220 => x"84",
          3221 => x"f4",
          3222 => x"dc",
          3223 => x"87",
          3224 => x"26",
          3225 => x"b4",
          3226 => x"11",
          3227 => x"05",
          3228 => x"3f",
          3229 => x"08",
          3230 => x"bb",
          3231 => x"63",
          3232 => x"b4",
          3233 => x"ff",
          3234 => x"02",
          3235 => x"33",
          3236 => x"63",
          3237 => x"82",
          3238 => x"51",
          3239 => x"3f",
          3240 => x"08",
          3241 => x"82",
          3242 => x"ca",
          3243 => x"5d",
          3244 => x"b4",
          3245 => x"05",
          3246 => x"3f",
          3247 => x"08",
          3248 => x"84",
          3249 => x"90",
          3250 => x"53",
          3251 => x"08",
          3252 => x"f2",
          3253 => x"d1",
          3254 => x"ff",
          3255 => x"8f",
          3256 => x"bb",
          3257 => x"3d",
          3258 => x"52",
          3259 => x"3f",
          3260 => x"08",
          3261 => x"84",
          3262 => x"90",
          3263 => x"bb",
          3264 => x"3d",
          3265 => x"52",
          3266 => x"3f",
          3267 => x"58",
          3268 => x"57",
          3269 => x"55",
          3270 => x"08",
          3271 => x"54",
          3272 => x"52",
          3273 => x"8d",
          3274 => x"dc",
          3275 => x"fb",
          3276 => x"bb",
          3277 => x"ef",
          3278 => x"82",
          3279 => x"ff",
          3280 => x"ff",
          3281 => x"e9",
          3282 => x"bb",
          3283 => x"2e",
          3284 => x"b4",
          3285 => x"11",
          3286 => x"05",
          3287 => x"3f",
          3288 => x"08",
          3289 => x"d6",
          3290 => x"fe",
          3291 => x"ff",
          3292 => x"e8",
          3293 => x"bb",
          3294 => x"38",
          3295 => x"08",
          3296 => x"b8",
          3297 => x"d0",
          3298 => x"5c",
          3299 => x"27",
          3300 => x"61",
          3301 => x"70",
          3302 => x"0c",
          3303 => x"f5",
          3304 => x"39",
          3305 => x"80",
          3306 => x"84",
          3307 => x"9c",
          3308 => x"dc",
          3309 => x"fa",
          3310 => x"3d",
          3311 => x"53",
          3312 => x"51",
          3313 => x"82",
          3314 => x"80",
          3315 => x"38",
          3316 => x"f8",
          3317 => x"84",
          3318 => x"f0",
          3319 => x"dc",
          3320 => x"f9",
          3321 => x"a7",
          3322 => x"ab",
          3323 => x"5a",
          3324 => x"81",
          3325 => x"59",
          3326 => x"05",
          3327 => x"34",
          3328 => x"42",
          3329 => x"3d",
          3330 => x"53",
          3331 => x"51",
          3332 => x"82",
          3333 => x"80",
          3334 => x"38",
          3335 => x"fc",
          3336 => x"84",
          3337 => x"a4",
          3338 => x"dc",
          3339 => x"f9",
          3340 => x"3d",
          3341 => x"53",
          3342 => x"51",
          3343 => x"82",
          3344 => x"80",
          3345 => x"38",
          3346 => x"51",
          3347 => x"3f",
          3348 => x"63",
          3349 => x"61",
          3350 => x"33",
          3351 => x"78",
          3352 => x"38",
          3353 => x"54",
          3354 => x"79",
          3355 => x"e4",
          3356 => x"e4",
          3357 => x"62",
          3358 => x"5a",
          3359 => x"51",
          3360 => x"f8",
          3361 => x"3d",
          3362 => x"53",
          3363 => x"51",
          3364 => x"82",
          3365 => x"80",
          3366 => x"ba",
          3367 => x"78",
          3368 => x"38",
          3369 => x"08",
          3370 => x"39",
          3371 => x"33",
          3372 => x"2e",
          3373 => x"ba",
          3374 => x"bc",
          3375 => x"ca",
          3376 => x"80",
          3377 => x"82",
          3378 => x"44",
          3379 => x"ba",
          3380 => x"78",
          3381 => x"38",
          3382 => x"08",
          3383 => x"82",
          3384 => x"59",
          3385 => x"88",
          3386 => x"a0",
          3387 => x"39",
          3388 => x"08",
          3389 => x"44",
          3390 => x"fc",
          3391 => x"84",
          3392 => x"c8",
          3393 => x"dc",
          3394 => x"38",
          3395 => x"33",
          3396 => x"2e",
          3397 => x"ba",
          3398 => x"80",
          3399 => x"ba",
          3400 => x"78",
          3401 => x"38",
          3402 => x"08",
          3403 => x"82",
          3404 => x"59",
          3405 => x"88",
          3406 => x"94",
          3407 => x"39",
          3408 => x"33",
          3409 => x"2e",
          3410 => x"ba",
          3411 => x"99",
          3412 => x"c6",
          3413 => x"80",
          3414 => x"82",
          3415 => x"43",
          3416 => x"ba",
          3417 => x"05",
          3418 => x"fe",
          3419 => x"ff",
          3420 => x"e4",
          3421 => x"bb",
          3422 => x"2e",
          3423 => x"62",
          3424 => x"88",
          3425 => x"81",
          3426 => x"32",
          3427 => x"72",
          3428 => x"70",
          3429 => x"51",
          3430 => x"80",
          3431 => x"7a",
          3432 => x"38",
          3433 => x"a8",
          3434 => x"b7",
          3435 => x"63",
          3436 => x"62",
          3437 => x"ee",
          3438 => x"a8",
          3439 => x"ce",
          3440 => x"ff",
          3441 => x"ff",
          3442 => x"e3",
          3443 => x"bb",
          3444 => x"2e",
          3445 => x"b4",
          3446 => x"11",
          3447 => x"05",
          3448 => x"3f",
          3449 => x"08",
          3450 => x"38",
          3451 => x"80",
          3452 => x"79",
          3453 => x"05",
          3454 => x"fe",
          3455 => x"ff",
          3456 => x"e3",
          3457 => x"bb",
          3458 => x"38",
          3459 => x"63",
          3460 => x"52",
          3461 => x"51",
          3462 => x"3f",
          3463 => x"08",
          3464 => x"52",
          3465 => x"a8",
          3466 => x"45",
          3467 => x"78",
          3468 => x"8a",
          3469 => x"27",
          3470 => x"3d",
          3471 => x"53",
          3472 => x"51",
          3473 => x"82",
          3474 => x"80",
          3475 => x"63",
          3476 => x"cb",
          3477 => x"34",
          3478 => x"44",
          3479 => x"82",
          3480 => x"c2",
          3481 => x"a7",
          3482 => x"fe",
          3483 => x"ff",
          3484 => x"dd",
          3485 => x"bb",
          3486 => x"2e",
          3487 => x"b4",
          3488 => x"11",
          3489 => x"05",
          3490 => x"3f",
          3491 => x"08",
          3492 => x"38",
          3493 => x"be",
          3494 => x"70",
          3495 => x"23",
          3496 => x"3d",
          3497 => x"53",
          3498 => x"51",
          3499 => x"82",
          3500 => x"e0",
          3501 => x"39",
          3502 => x"54",
          3503 => x"a8",
          3504 => x"94",
          3505 => x"ac",
          3506 => x"f8",
          3507 => x"ff",
          3508 => x"79",
          3509 => x"59",
          3510 => x"f3",
          3511 => x"9f",
          3512 => x"60",
          3513 => x"d0",
          3514 => x"fe",
          3515 => x"ff",
          3516 => x"dc",
          3517 => x"bb",
          3518 => x"2e",
          3519 => x"59",
          3520 => x"22",
          3521 => x"05",
          3522 => x"41",
          3523 => x"82",
          3524 => x"c1",
          3525 => x"a0",
          3526 => x"fe",
          3527 => x"ff",
          3528 => x"db",
          3529 => x"bb",
          3530 => x"2e",
          3531 => x"b4",
          3532 => x"11",
          3533 => x"05",
          3534 => x"3f",
          3535 => x"08",
          3536 => x"38",
          3537 => x"0c",
          3538 => x"05",
          3539 => x"fe",
          3540 => x"ff",
          3541 => x"db",
          3542 => x"bb",
          3543 => x"38",
          3544 => x"60",
          3545 => x"52",
          3546 => x"51",
          3547 => x"3f",
          3548 => x"08",
          3549 => x"52",
          3550 => x"a5",
          3551 => x"45",
          3552 => x"78",
          3553 => x"b6",
          3554 => x"27",
          3555 => x"3d",
          3556 => x"53",
          3557 => x"51",
          3558 => x"82",
          3559 => x"80",
          3560 => x"60",
          3561 => x"59",
          3562 => x"41",
          3563 => x"82",
          3564 => x"c0",
          3565 => x"ab",
          3566 => x"c4",
          3567 => x"3f",
          3568 => x"89",
          3569 => x"39",
          3570 => x"51",
          3571 => x"a2",
          3572 => x"3f",
          3573 => x"82",
          3574 => x"c0",
          3575 => x"80",
          3576 => x"c0",
          3577 => x"84",
          3578 => x"87",
          3579 => x"0c",
          3580 => x"82",
          3581 => x"ff",
          3582 => x"8c",
          3583 => x"87",
          3584 => x"0c",
          3585 => x"0b",
          3586 => x"94",
          3587 => x"39",
          3588 => x"80",
          3589 => x"84",
          3590 => x"b0",
          3591 => x"dc",
          3592 => x"f1",
          3593 => x"52",
          3594 => x"51",
          3595 => x"3f",
          3596 => x"04",
          3597 => x"80",
          3598 => x"84",
          3599 => x"8c",
          3600 => x"dc",
          3601 => x"f0",
          3602 => x"52",
          3603 => x"51",
          3604 => x"3f",
          3605 => x"2d",
          3606 => x"08",
          3607 => x"de",
          3608 => x"dc",
          3609 => x"a9",
          3610 => x"a2",
          3611 => x"ce",
          3612 => x"ec",
          3613 => x"eb",
          3614 => x"bd",
          3615 => x"39",
          3616 => x"51",
          3617 => x"3f",
          3618 => x"a6",
          3619 => x"3f",
          3620 => x"79",
          3621 => x"59",
          3622 => x"f0",
          3623 => x"7d",
          3624 => x"80",
          3625 => x"38",
          3626 => x"84",
          3627 => x"cb",
          3628 => x"dc",
          3629 => x"5c",
          3630 => x"b2",
          3631 => x"24",
          3632 => x"81",
          3633 => x"80",
          3634 => x"83",
          3635 => x"80",
          3636 => x"aa",
          3637 => x"55",
          3638 => x"54",
          3639 => x"aa",
          3640 => x"3d",
          3641 => x"51",
          3642 => x"3f",
          3643 => x"52",
          3644 => x"b0",
          3645 => x"fb",
          3646 => x"7a",
          3647 => x"a0",
          3648 => x"82",
          3649 => x"b4",
          3650 => x"05",
          3651 => x"b0",
          3652 => x"7a",
          3653 => x"82",
          3654 => x"b4",
          3655 => x"05",
          3656 => x"9c",
          3657 => x"80",
          3658 => x"8c",
          3659 => x"64",
          3660 => x"82",
          3661 => x"82",
          3662 => x"b4",
          3663 => x"05",
          3664 => x"3f",
          3665 => x"08",
          3666 => x"08",
          3667 => x"70",
          3668 => x"25",
          3669 => x"5f",
          3670 => x"83",
          3671 => x"81",
          3672 => x"06",
          3673 => x"2e",
          3674 => x"1c",
          3675 => x"06",
          3676 => x"fe",
          3677 => x"81",
          3678 => x"32",
          3679 => x"8a",
          3680 => x"2e",
          3681 => x"ee",
          3682 => x"aa",
          3683 => x"bc",
          3684 => x"aa",
          3685 => x"0d",
          3686 => x"bc",
          3687 => x"c0",
          3688 => x"08",
          3689 => x"84",
          3690 => x"51",
          3691 => x"82",
          3692 => x"90",
          3693 => x"55",
          3694 => x"80",
          3695 => x"d3",
          3696 => x"82",
          3697 => x"07",
          3698 => x"c0",
          3699 => x"08",
          3700 => x"84",
          3701 => x"51",
          3702 => x"82",
          3703 => x"90",
          3704 => x"55",
          3705 => x"80",
          3706 => x"d3",
          3707 => x"82",
          3708 => x"07",
          3709 => x"80",
          3710 => x"c0",
          3711 => x"8c",
          3712 => x"87",
          3713 => x"0c",
          3714 => x"5a",
          3715 => x"5b",
          3716 => x"05",
          3717 => x"80",
          3718 => x"ac",
          3719 => x"70",
          3720 => x"70",
          3721 => x"d3",
          3722 => x"89",
          3723 => x"c2",
          3724 => x"d8",
          3725 => x"ab",
          3726 => x"e4",
          3727 => x"a3",
          3728 => x"b1",
          3729 => x"3f",
          3730 => x"a8",
          3731 => x"3f",
          3732 => x"3d",
          3733 => x"83",
          3734 => x"2b",
          3735 => x"3f",
          3736 => x"08",
          3737 => x"72",
          3738 => x"54",
          3739 => x"25",
          3740 => x"82",
          3741 => x"84",
          3742 => x"fc",
          3743 => x"70",
          3744 => x"80",
          3745 => x"72",
          3746 => x"8a",
          3747 => x"51",
          3748 => x"09",
          3749 => x"38",
          3750 => x"f1",
          3751 => x"51",
          3752 => x"09",
          3753 => x"38",
          3754 => x"81",
          3755 => x"73",
          3756 => x"81",
          3757 => x"84",
          3758 => x"52",
          3759 => x"52",
          3760 => x"2e",
          3761 => x"54",
          3762 => x"9d",
          3763 => x"38",
          3764 => x"12",
          3765 => x"33",
          3766 => x"a0",
          3767 => x"81",
          3768 => x"2e",
          3769 => x"ea",
          3770 => x"33",
          3771 => x"a0",
          3772 => x"06",
          3773 => x"54",
          3774 => x"70",
          3775 => x"25",
          3776 => x"51",
          3777 => x"2e",
          3778 => x"72",
          3779 => x"54",
          3780 => x"0c",
          3781 => x"82",
          3782 => x"86",
          3783 => x"fc",
          3784 => x"53",
          3785 => x"2e",
          3786 => x"3d",
          3787 => x"72",
          3788 => x"3f",
          3789 => x"08",
          3790 => x"53",
          3791 => x"53",
          3792 => x"dc",
          3793 => x"0d",
          3794 => x"0d",
          3795 => x"33",
          3796 => x"53",
          3797 => x"8b",
          3798 => x"38",
          3799 => x"ff",
          3800 => x"52",
          3801 => x"81",
          3802 => x"13",
          3803 => x"52",
          3804 => x"80",
          3805 => x"13",
          3806 => x"52",
          3807 => x"80",
          3808 => x"13",
          3809 => x"52",
          3810 => x"80",
          3811 => x"13",
          3812 => x"52",
          3813 => x"26",
          3814 => x"8a",
          3815 => x"87",
          3816 => x"e7",
          3817 => x"38",
          3818 => x"c0",
          3819 => x"72",
          3820 => x"98",
          3821 => x"13",
          3822 => x"98",
          3823 => x"13",
          3824 => x"98",
          3825 => x"13",
          3826 => x"98",
          3827 => x"13",
          3828 => x"98",
          3829 => x"13",
          3830 => x"98",
          3831 => x"87",
          3832 => x"0c",
          3833 => x"98",
          3834 => x"0b",
          3835 => x"9c",
          3836 => x"71",
          3837 => x"0c",
          3838 => x"04",
          3839 => x"7f",
          3840 => x"98",
          3841 => x"7d",
          3842 => x"98",
          3843 => x"7d",
          3844 => x"c0",
          3845 => x"5a",
          3846 => x"34",
          3847 => x"b4",
          3848 => x"83",
          3849 => x"c0",
          3850 => x"5a",
          3851 => x"34",
          3852 => x"ac",
          3853 => x"85",
          3854 => x"c0",
          3855 => x"5a",
          3856 => x"34",
          3857 => x"a4",
          3858 => x"88",
          3859 => x"c0",
          3860 => x"5a",
          3861 => x"23",
          3862 => x"79",
          3863 => x"06",
          3864 => x"ff",
          3865 => x"86",
          3866 => x"85",
          3867 => x"84",
          3868 => x"83",
          3869 => x"82",
          3870 => x"7d",
          3871 => x"06",
          3872 => x"fc",
          3873 => x"d0",
          3874 => x"0d",
          3875 => x"0d",
          3876 => x"33",
          3877 => x"33",
          3878 => x"06",
          3879 => x"87",
          3880 => x"51",
          3881 => x"86",
          3882 => x"94",
          3883 => x"08",
          3884 => x"70",
          3885 => x"54",
          3886 => x"2e",
          3887 => x"91",
          3888 => x"06",
          3889 => x"d7",
          3890 => x"32",
          3891 => x"51",
          3892 => x"2e",
          3893 => x"93",
          3894 => x"06",
          3895 => x"ff",
          3896 => x"81",
          3897 => x"87",
          3898 => x"52",
          3899 => x"86",
          3900 => x"94",
          3901 => x"72",
          3902 => x"bb",
          3903 => x"3d",
          3904 => x"3d",
          3905 => x"05",
          3906 => x"70",
          3907 => x"52",
          3908 => x"b9",
          3909 => x"3d",
          3910 => x"3d",
          3911 => x"05",
          3912 => x"8a",
          3913 => x"06",
          3914 => x"52",
          3915 => x"3f",
          3916 => x"33",
          3917 => x"06",
          3918 => x"c0",
          3919 => x"76",
          3920 => x"38",
          3921 => x"94",
          3922 => x"70",
          3923 => x"81",
          3924 => x"54",
          3925 => x"8c",
          3926 => x"2a",
          3927 => x"51",
          3928 => x"38",
          3929 => x"70",
          3930 => x"53",
          3931 => x"8d",
          3932 => x"2a",
          3933 => x"51",
          3934 => x"be",
          3935 => x"ff",
          3936 => x"c0",
          3937 => x"72",
          3938 => x"38",
          3939 => x"90",
          3940 => x"0c",
          3941 => x"bb",
          3942 => x"3d",
          3943 => x"3d",
          3944 => x"80",
          3945 => x"81",
          3946 => x"53",
          3947 => x"2e",
          3948 => x"71",
          3949 => x"81",
          3950 => x"fc",
          3951 => x"ff",
          3952 => x"55",
          3953 => x"94",
          3954 => x"80",
          3955 => x"87",
          3956 => x"51",
          3957 => x"96",
          3958 => x"06",
          3959 => x"70",
          3960 => x"38",
          3961 => x"70",
          3962 => x"51",
          3963 => x"72",
          3964 => x"81",
          3965 => x"70",
          3966 => x"38",
          3967 => x"70",
          3968 => x"51",
          3969 => x"38",
          3970 => x"06",
          3971 => x"94",
          3972 => x"80",
          3973 => x"87",
          3974 => x"52",
          3975 => x"81",
          3976 => x"70",
          3977 => x"53",
          3978 => x"ff",
          3979 => x"82",
          3980 => x"89",
          3981 => x"fe",
          3982 => x"b9",
          3983 => x"81",
          3984 => x"52",
          3985 => x"84",
          3986 => x"2e",
          3987 => x"c0",
          3988 => x"70",
          3989 => x"2a",
          3990 => x"51",
          3991 => x"80",
          3992 => x"71",
          3993 => x"51",
          3994 => x"80",
          3995 => x"2e",
          3996 => x"c0",
          3997 => x"71",
          3998 => x"ff",
          3999 => x"dc",
          4000 => x"3d",
          4001 => x"af",
          4002 => x"dc",
          4003 => x"06",
          4004 => x"0c",
          4005 => x"0d",
          4006 => x"33",
          4007 => x"06",
          4008 => x"c0",
          4009 => x"70",
          4010 => x"38",
          4011 => x"94",
          4012 => x"70",
          4013 => x"81",
          4014 => x"51",
          4015 => x"80",
          4016 => x"72",
          4017 => x"51",
          4018 => x"80",
          4019 => x"2e",
          4020 => x"c0",
          4021 => x"71",
          4022 => x"2b",
          4023 => x"51",
          4024 => x"82",
          4025 => x"84",
          4026 => x"ff",
          4027 => x"c0",
          4028 => x"70",
          4029 => x"06",
          4030 => x"80",
          4031 => x"38",
          4032 => x"a4",
          4033 => x"80",
          4034 => x"9e",
          4035 => x"ba",
          4036 => x"c0",
          4037 => x"82",
          4038 => x"87",
          4039 => x"08",
          4040 => x"0c",
          4041 => x"9c",
          4042 => x"90",
          4043 => x"9e",
          4044 => x"ba",
          4045 => x"c0",
          4046 => x"82",
          4047 => x"87",
          4048 => x"08",
          4049 => x"0c",
          4050 => x"b4",
          4051 => x"a0",
          4052 => x"9e",
          4053 => x"ba",
          4054 => x"c0",
          4055 => x"82",
          4056 => x"87",
          4057 => x"08",
          4058 => x"0c",
          4059 => x"c4",
          4060 => x"b0",
          4061 => x"9e",
          4062 => x"70",
          4063 => x"23",
          4064 => x"84",
          4065 => x"b8",
          4066 => x"9e",
          4067 => x"ba",
          4068 => x"c0",
          4069 => x"82",
          4070 => x"81",
          4071 => x"c4",
          4072 => x"87",
          4073 => x"08",
          4074 => x"0a",
          4075 => x"52",
          4076 => x"83",
          4077 => x"71",
          4078 => x"34",
          4079 => x"c0",
          4080 => x"70",
          4081 => x"06",
          4082 => x"70",
          4083 => x"38",
          4084 => x"82",
          4085 => x"80",
          4086 => x"9e",
          4087 => x"90",
          4088 => x"51",
          4089 => x"80",
          4090 => x"81",
          4091 => x"ba",
          4092 => x"0b",
          4093 => x"90",
          4094 => x"80",
          4095 => x"52",
          4096 => x"2e",
          4097 => x"52",
          4098 => x"c8",
          4099 => x"87",
          4100 => x"08",
          4101 => x"80",
          4102 => x"52",
          4103 => x"83",
          4104 => x"71",
          4105 => x"34",
          4106 => x"c0",
          4107 => x"70",
          4108 => x"06",
          4109 => x"70",
          4110 => x"38",
          4111 => x"82",
          4112 => x"80",
          4113 => x"9e",
          4114 => x"84",
          4115 => x"51",
          4116 => x"80",
          4117 => x"81",
          4118 => x"ba",
          4119 => x"0b",
          4120 => x"90",
          4121 => x"80",
          4122 => x"52",
          4123 => x"2e",
          4124 => x"52",
          4125 => x"cc",
          4126 => x"87",
          4127 => x"08",
          4128 => x"80",
          4129 => x"52",
          4130 => x"83",
          4131 => x"71",
          4132 => x"34",
          4133 => x"c0",
          4134 => x"70",
          4135 => x"06",
          4136 => x"70",
          4137 => x"38",
          4138 => x"82",
          4139 => x"80",
          4140 => x"9e",
          4141 => x"a0",
          4142 => x"52",
          4143 => x"2e",
          4144 => x"52",
          4145 => x"cf",
          4146 => x"9e",
          4147 => x"98",
          4148 => x"8a",
          4149 => x"51",
          4150 => x"d0",
          4151 => x"87",
          4152 => x"08",
          4153 => x"06",
          4154 => x"70",
          4155 => x"38",
          4156 => x"82",
          4157 => x"87",
          4158 => x"08",
          4159 => x"06",
          4160 => x"51",
          4161 => x"82",
          4162 => x"80",
          4163 => x"9e",
          4164 => x"88",
          4165 => x"52",
          4166 => x"83",
          4167 => x"71",
          4168 => x"34",
          4169 => x"90",
          4170 => x"06",
          4171 => x"82",
          4172 => x"83",
          4173 => x"fb",
          4174 => x"ab",
          4175 => x"ad",
          4176 => x"ba",
          4177 => x"73",
          4178 => x"38",
          4179 => x"51",
          4180 => x"3f",
          4181 => x"51",
          4182 => x"3f",
          4183 => x"33",
          4184 => x"2e",
          4185 => x"ba",
          4186 => x"ba",
          4187 => x"54",
          4188 => x"d4",
          4189 => x"e0",
          4190 => x"cb",
          4191 => x"80",
          4192 => x"82",
          4193 => x"82",
          4194 => x"11",
          4195 => x"ab",
          4196 => x"90",
          4197 => x"ba",
          4198 => x"73",
          4199 => x"38",
          4200 => x"08",
          4201 => x"08",
          4202 => x"82",
          4203 => x"ff",
          4204 => x"82",
          4205 => x"54",
          4206 => x"94",
          4207 => x"88",
          4208 => x"8c",
          4209 => x"52",
          4210 => x"51",
          4211 => x"3f",
          4212 => x"33",
          4213 => x"2e",
          4214 => x"ba",
          4215 => x"ba",
          4216 => x"54",
          4217 => x"c4",
          4218 => x"ec",
          4219 => x"cf",
          4220 => x"80",
          4221 => x"82",
          4222 => x"52",
          4223 => x"51",
          4224 => x"3f",
          4225 => x"33",
          4226 => x"2e",
          4227 => x"ba",
          4228 => x"82",
          4229 => x"ff",
          4230 => x"82",
          4231 => x"54",
          4232 => x"8e",
          4233 => x"d2",
          4234 => x"ad",
          4235 => x"8f",
          4236 => x"ba",
          4237 => x"73",
          4238 => x"38",
          4239 => x"51",
          4240 => x"3f",
          4241 => x"33",
          4242 => x"2e",
          4243 => x"ad",
          4244 => x"ab",
          4245 => x"ba",
          4246 => x"73",
          4247 => x"38",
          4248 => x"51",
          4249 => x"3f",
          4250 => x"33",
          4251 => x"2e",
          4252 => x"ad",
          4253 => x"aa",
          4254 => x"ba",
          4255 => x"73",
          4256 => x"38",
          4257 => x"51",
          4258 => x"3f",
          4259 => x"51",
          4260 => x"3f",
          4261 => x"08",
          4262 => x"90",
          4263 => x"b8",
          4264 => x"ac",
          4265 => x"ae",
          4266 => x"8e",
          4267 => x"ba",
          4268 => x"82",
          4269 => x"ff",
          4270 => x"82",
          4271 => x"ff",
          4272 => x"82",
          4273 => x"52",
          4274 => x"51",
          4275 => x"3f",
          4276 => x"08",
          4277 => x"c0",
          4278 => x"c1",
          4279 => x"bb",
          4280 => x"84",
          4281 => x"71",
          4282 => x"82",
          4283 => x"52",
          4284 => x"51",
          4285 => x"3f",
          4286 => x"33",
          4287 => x"2e",
          4288 => x"ba",
          4289 => x"bd",
          4290 => x"75",
          4291 => x"3f",
          4292 => x"08",
          4293 => x"29",
          4294 => x"54",
          4295 => x"dc",
          4296 => x"af",
          4297 => x"8d",
          4298 => x"ba",
          4299 => x"73",
          4300 => x"38",
          4301 => x"08",
          4302 => x"c0",
          4303 => x"c0",
          4304 => x"bb",
          4305 => x"84",
          4306 => x"71",
          4307 => x"82",
          4308 => x"52",
          4309 => x"51",
          4310 => x"3f",
          4311 => x"51",
          4312 => x"3f",
          4313 => x"04",
          4314 => x"02",
          4315 => x"ff",
          4316 => x"84",
          4317 => x"71",
          4318 => x"9a",
          4319 => x"71",
          4320 => x"b0",
          4321 => x"39",
          4322 => x"51",
          4323 => x"b0",
          4324 => x"39",
          4325 => x"51",
          4326 => x"b0",
          4327 => x"39",
          4328 => x"51",
          4329 => x"3f",
          4330 => x"04",
          4331 => x"0c",
          4332 => x"0d",
          4333 => x"84",
          4334 => x"52",
          4335 => x"70",
          4336 => x"82",
          4337 => x"72",
          4338 => x"0d",
          4339 => x"0d",
          4340 => x"84",
          4341 => x"ba",
          4342 => x"80",
          4343 => x"09",
          4344 => x"d8",
          4345 => x"82",
          4346 => x"73",
          4347 => x"3d",
          4348 => x"0b",
          4349 => x"84",
          4350 => x"ba",
          4351 => x"c0",
          4352 => x"04",
          4353 => x"76",
          4354 => x"98",
          4355 => x"2b",
          4356 => x"72",
          4357 => x"82",
          4358 => x"51",
          4359 => x"80",
          4360 => x"ec",
          4361 => x"53",
          4362 => x"9c",
          4363 => x"e8",
          4364 => x"02",
          4365 => x"05",
          4366 => x"52",
          4367 => x"72",
          4368 => x"06",
          4369 => x"53",
          4370 => x"dc",
          4371 => x"0d",
          4372 => x"0d",
          4373 => x"05",
          4374 => x"71",
          4375 => x"54",
          4376 => x"b1",
          4377 => x"b0",
          4378 => x"51",
          4379 => x"3f",
          4380 => x"08",
          4381 => x"ff",
          4382 => x"82",
          4383 => x"52",
          4384 => x"aa",
          4385 => x"33",
          4386 => x"72",
          4387 => x"81",
          4388 => x"cc",
          4389 => x"ff",
          4390 => x"74",
          4391 => x"3d",
          4392 => x"3d",
          4393 => x"84",
          4394 => x"33",
          4395 => x"bb",
          4396 => x"bb",
          4397 => x"84",
          4398 => x"dc",
          4399 => x"51",
          4400 => x"58",
          4401 => x"2e",
          4402 => x"51",
          4403 => x"82",
          4404 => x"70",
          4405 => x"ba",
          4406 => x"19",
          4407 => x"56",
          4408 => x"3f",
          4409 => x"08",
          4410 => x"bb",
          4411 => x"84",
          4412 => x"dc",
          4413 => x"51",
          4414 => x"80",
          4415 => x"75",
          4416 => x"74",
          4417 => x"dd",
          4418 => x"b4",
          4419 => x"55",
          4420 => x"b4",
          4421 => x"ff",
          4422 => x"75",
          4423 => x"80",
          4424 => x"b4",
          4425 => x"2e",
          4426 => x"bb",
          4427 => x"75",
          4428 => x"38",
          4429 => x"33",
          4430 => x"38",
          4431 => x"05",
          4432 => x"78",
          4433 => x"80",
          4434 => x"82",
          4435 => x"52",
          4436 => x"8f",
          4437 => x"bb",
          4438 => x"80",
          4439 => x"8c",
          4440 => x"fd",
          4441 => x"ba",
          4442 => x"54",
          4443 => x"71",
          4444 => x"38",
          4445 => x"d0",
          4446 => x"0c",
          4447 => x"14",
          4448 => x"80",
          4449 => x"80",
          4450 => x"b4",
          4451 => x"b0",
          4452 => x"80",
          4453 => x"71",
          4454 => x"c5",
          4455 => x"b0",
          4456 => x"a4",
          4457 => x"82",
          4458 => x"85",
          4459 => x"dc",
          4460 => x"57",
          4461 => x"bb",
          4462 => x"80",
          4463 => x"82",
          4464 => x"80",
          4465 => x"bb",
          4466 => x"80",
          4467 => x"3d",
          4468 => x"81",
          4469 => x"82",
          4470 => x"80",
          4471 => x"75",
          4472 => x"a1",
          4473 => x"dc",
          4474 => x"0b",
          4475 => x"08",
          4476 => x"82",
          4477 => x"ff",
          4478 => x"55",
          4479 => x"34",
          4480 => x"52",
          4481 => x"b3",
          4482 => x"ff",
          4483 => x"74",
          4484 => x"81",
          4485 => x"38",
          4486 => x"04",
          4487 => x"aa",
          4488 => x"3d",
          4489 => x"81",
          4490 => x"80",
          4491 => x"b0",
          4492 => x"e2",
          4493 => x"bb",
          4494 => x"95",
          4495 => x"82",
          4496 => x"54",
          4497 => x"52",
          4498 => x"52",
          4499 => x"86",
          4500 => x"dc",
          4501 => x"a5",
          4502 => x"ff",
          4503 => x"82",
          4504 => x"81",
          4505 => x"80",
          4506 => x"dc",
          4507 => x"38",
          4508 => x"08",
          4509 => x"17",
          4510 => x"74",
          4511 => x"70",
          4512 => x"07",
          4513 => x"55",
          4514 => x"2e",
          4515 => x"ff",
          4516 => x"bb",
          4517 => x"11",
          4518 => x"80",
          4519 => x"82",
          4520 => x"80",
          4521 => x"82",
          4522 => x"ff",
          4523 => x"78",
          4524 => x"81",
          4525 => x"75",
          4526 => x"ff",
          4527 => x"79",
          4528 => x"c1",
          4529 => x"08",
          4530 => x"dc",
          4531 => x"80",
          4532 => x"bb",
          4533 => x"3d",
          4534 => x"3d",
          4535 => x"71",
          4536 => x"33",
          4537 => x"58",
          4538 => x"09",
          4539 => x"38",
          4540 => x"05",
          4541 => x"27",
          4542 => x"17",
          4543 => x"71",
          4544 => x"55",
          4545 => x"09",
          4546 => x"38",
          4547 => x"ea",
          4548 => x"73",
          4549 => x"bb",
          4550 => x"08",
          4551 => x"ad",
          4552 => x"bb",
          4553 => x"79",
          4554 => x"51",
          4555 => x"3f",
          4556 => x"08",
          4557 => x"84",
          4558 => x"74",
          4559 => x"38",
          4560 => x"88",
          4561 => x"fc",
          4562 => x"39",
          4563 => x"8c",
          4564 => x"53",
          4565 => x"c0",
          4566 => x"bb",
          4567 => x"2e",
          4568 => x"1b",
          4569 => x"77",
          4570 => x"3f",
          4571 => x"08",
          4572 => x"55",
          4573 => x"74",
          4574 => x"81",
          4575 => x"ff",
          4576 => x"82",
          4577 => x"8b",
          4578 => x"73",
          4579 => x"0c",
          4580 => x"04",
          4581 => x"b0",
          4582 => x"3d",
          4583 => x"08",
          4584 => x"80",
          4585 => x"34",
          4586 => x"33",
          4587 => x"08",
          4588 => x"81",
          4589 => x"82",
          4590 => x"55",
          4591 => x"38",
          4592 => x"80",
          4593 => x"38",
          4594 => x"06",
          4595 => x"80",
          4596 => x"38",
          4597 => x"86",
          4598 => x"dc",
          4599 => x"b0",
          4600 => x"dc",
          4601 => x"81",
          4602 => x"53",
          4603 => x"bb",
          4604 => x"80",
          4605 => x"82",
          4606 => x"80",
          4607 => x"82",
          4608 => x"ff",
          4609 => x"80",
          4610 => x"bb",
          4611 => x"82",
          4612 => x"53",
          4613 => x"90",
          4614 => x"54",
          4615 => x"3f",
          4616 => x"08",
          4617 => x"dc",
          4618 => x"09",
          4619 => x"d0",
          4620 => x"dc",
          4621 => x"ab",
          4622 => x"bb",
          4623 => x"80",
          4624 => x"dc",
          4625 => x"38",
          4626 => x"08",
          4627 => x"17",
          4628 => x"74",
          4629 => x"74",
          4630 => x"52",
          4631 => x"c2",
          4632 => x"70",
          4633 => x"5c",
          4634 => x"27",
          4635 => x"5b",
          4636 => x"09",
          4637 => x"97",
          4638 => x"75",
          4639 => x"34",
          4640 => x"82",
          4641 => x"80",
          4642 => x"f9",
          4643 => x"3d",
          4644 => x"3f",
          4645 => x"08",
          4646 => x"98",
          4647 => x"78",
          4648 => x"38",
          4649 => x"06",
          4650 => x"33",
          4651 => x"70",
          4652 => x"d3",
          4653 => x"98",
          4654 => x"2c",
          4655 => x"05",
          4656 => x"82",
          4657 => x"70",
          4658 => x"33",
          4659 => x"51",
          4660 => x"59",
          4661 => x"56",
          4662 => x"80",
          4663 => x"74",
          4664 => x"74",
          4665 => x"29",
          4666 => x"05",
          4667 => x"51",
          4668 => x"24",
          4669 => x"76",
          4670 => x"77",
          4671 => x"3f",
          4672 => x"08",
          4673 => x"54",
          4674 => x"d7",
          4675 => x"d3",
          4676 => x"56",
          4677 => x"81",
          4678 => x"81",
          4679 => x"70",
          4680 => x"81",
          4681 => x"51",
          4682 => x"26",
          4683 => x"53",
          4684 => x"51",
          4685 => x"82",
          4686 => x"81",
          4687 => x"73",
          4688 => x"39",
          4689 => x"80",
          4690 => x"38",
          4691 => x"74",
          4692 => x"34",
          4693 => x"70",
          4694 => x"d3",
          4695 => x"98",
          4696 => x"2c",
          4697 => x"70",
          4698 => x"b0",
          4699 => x"5e",
          4700 => x"57",
          4701 => x"74",
          4702 => x"81",
          4703 => x"38",
          4704 => x"14",
          4705 => x"80",
          4706 => x"88",
          4707 => x"82",
          4708 => x"92",
          4709 => x"d3",
          4710 => x"82",
          4711 => x"78",
          4712 => x"75",
          4713 => x"54",
          4714 => x"fd",
          4715 => x"84",
          4716 => x"80",
          4717 => x"08",
          4718 => x"90",
          4719 => x"7e",
          4720 => x"38",
          4721 => x"33",
          4722 => x"27",
          4723 => x"98",
          4724 => x"2c",
          4725 => x"75",
          4726 => x"74",
          4727 => x"33",
          4728 => x"74",
          4729 => x"29",
          4730 => x"05",
          4731 => x"82",
          4732 => x"56",
          4733 => x"39",
          4734 => x"33",
          4735 => x"54",
          4736 => x"90",
          4737 => x"54",
          4738 => x"74",
          4739 => x"8c",
          4740 => x"7e",
          4741 => x"81",
          4742 => x"82",
          4743 => x"82",
          4744 => x"70",
          4745 => x"29",
          4746 => x"05",
          4747 => x"82",
          4748 => x"5a",
          4749 => x"74",
          4750 => x"38",
          4751 => x"08",
          4752 => x"70",
          4753 => x"ff",
          4754 => x"74",
          4755 => x"29",
          4756 => x"05",
          4757 => x"82",
          4758 => x"56",
          4759 => x"75",
          4760 => x"82",
          4761 => x"70",
          4762 => x"98",
          4763 => x"8c",
          4764 => x"56",
          4765 => x"25",
          4766 => x"82",
          4767 => x"52",
          4768 => x"9e",
          4769 => x"81",
          4770 => x"81",
          4771 => x"70",
          4772 => x"d3",
          4773 => x"51",
          4774 => x"24",
          4775 => x"ee",
          4776 => x"34",
          4777 => x"1b",
          4778 => x"90",
          4779 => x"82",
          4780 => x"f3",
          4781 => x"fd",
          4782 => x"90",
          4783 => x"ff",
          4784 => x"73",
          4785 => x"c6",
          4786 => x"8c",
          4787 => x"54",
          4788 => x"8c",
          4789 => x"54",
          4790 => x"90",
          4791 => x"b0",
          4792 => x"51",
          4793 => x"3f",
          4794 => x"33",
          4795 => x"70",
          4796 => x"d3",
          4797 => x"51",
          4798 => x"74",
          4799 => x"74",
          4800 => x"14",
          4801 => x"82",
          4802 => x"52",
          4803 => x"ff",
          4804 => x"74",
          4805 => x"29",
          4806 => x"05",
          4807 => x"82",
          4808 => x"58",
          4809 => x"75",
          4810 => x"82",
          4811 => x"52",
          4812 => x"9c",
          4813 => x"d3",
          4814 => x"98",
          4815 => x"2c",
          4816 => x"33",
          4817 => x"57",
          4818 => x"fa",
          4819 => x"d3",
          4820 => x"88",
          4821 => x"da",
          4822 => x"80",
          4823 => x"80",
          4824 => x"98",
          4825 => x"8c",
          4826 => x"55",
          4827 => x"de",
          4828 => x"39",
          4829 => x"33",
          4830 => x"80",
          4831 => x"d3",
          4832 => x"8a",
          4833 => x"aa",
          4834 => x"8c",
          4835 => x"f6",
          4836 => x"bb",
          4837 => x"ff",
          4838 => x"96",
          4839 => x"8c",
          4840 => x"80",
          4841 => x"81",
          4842 => x"79",
          4843 => x"3f",
          4844 => x"7a",
          4845 => x"82",
          4846 => x"80",
          4847 => x"8c",
          4848 => x"bb",
          4849 => x"3d",
          4850 => x"d3",
          4851 => x"73",
          4852 => x"ba",
          4853 => x"b0",
          4854 => x"51",
          4855 => x"3f",
          4856 => x"33",
          4857 => x"73",
          4858 => x"34",
          4859 => x"06",
          4860 => x"82",
          4861 => x"82",
          4862 => x"55",
          4863 => x"2e",
          4864 => x"ff",
          4865 => x"82",
          4866 => x"74",
          4867 => x"98",
          4868 => x"ff",
          4869 => x"55",
          4870 => x"ad",
          4871 => x"54",
          4872 => x"74",
          4873 => x"b0",
          4874 => x"33",
          4875 => x"82",
          4876 => x"80",
          4877 => x"80",
          4878 => x"98",
          4879 => x"8c",
          4880 => x"55",
          4881 => x"d5",
          4882 => x"b0",
          4883 => x"51",
          4884 => x"3f",
          4885 => x"33",
          4886 => x"70",
          4887 => x"d3",
          4888 => x"51",
          4889 => x"74",
          4890 => x"38",
          4891 => x"08",
          4892 => x"ff",
          4893 => x"74",
          4894 => x"29",
          4895 => x"05",
          4896 => x"82",
          4897 => x"58",
          4898 => x"75",
          4899 => x"f7",
          4900 => x"d3",
          4901 => x"81",
          4902 => x"d3",
          4903 => x"56",
          4904 => x"27",
          4905 => x"82",
          4906 => x"52",
          4907 => x"73",
          4908 => x"34",
          4909 => x"33",
          4910 => x"99",
          4911 => x"d3",
          4912 => x"81",
          4913 => x"d3",
          4914 => x"56",
          4915 => x"26",
          4916 => x"ba",
          4917 => x"90",
          4918 => x"82",
          4919 => x"ee",
          4920 => x"0b",
          4921 => x"34",
          4922 => x"d3",
          4923 => x"9e",
          4924 => x"38",
          4925 => x"08",
          4926 => x"2e",
          4927 => x"51",
          4928 => x"3f",
          4929 => x"08",
          4930 => x"34",
          4931 => x"08",
          4932 => x"81",
          4933 => x"52",
          4934 => x"a3",
          4935 => x"5b",
          4936 => x"7a",
          4937 => x"ba",
          4938 => x"11",
          4939 => x"74",
          4940 => x"38",
          4941 => x"a1",
          4942 => x"bb",
          4943 => x"d3",
          4944 => x"bb",
          4945 => x"ff",
          4946 => x"53",
          4947 => x"51",
          4948 => x"3f",
          4949 => x"80",
          4950 => x"08",
          4951 => x"2e",
          4952 => x"74",
          4953 => x"9d",
          4954 => x"7a",
          4955 => x"81",
          4956 => x"82",
          4957 => x"55",
          4958 => x"a4",
          4959 => x"ff",
          4960 => x"82",
          4961 => x"82",
          4962 => x"82",
          4963 => x"81",
          4964 => x"05",
          4965 => x"79",
          4966 => x"c9",
          4967 => x"39",
          4968 => x"82",
          4969 => x"70",
          4970 => x"74",
          4971 => x"38",
          4972 => x"a0",
          4973 => x"bb",
          4974 => x"d3",
          4975 => x"bb",
          4976 => x"ff",
          4977 => x"53",
          4978 => x"51",
          4979 => x"3f",
          4980 => x"73",
          4981 => x"5b",
          4982 => x"82",
          4983 => x"74",
          4984 => x"d3",
          4985 => x"d3",
          4986 => x"79",
          4987 => x"3f",
          4988 => x"82",
          4989 => x"70",
          4990 => x"82",
          4991 => x"59",
          4992 => x"77",
          4993 => x"38",
          4994 => x"08",
          4995 => x"54",
          4996 => x"90",
          4997 => x"70",
          4998 => x"ff",
          4999 => x"f4",
          5000 => x"d3",
          5001 => x"73",
          5002 => x"e2",
          5003 => x"b0",
          5004 => x"51",
          5005 => x"3f",
          5006 => x"33",
          5007 => x"73",
          5008 => x"34",
          5009 => x"f9",
          5010 => x"c0",
          5011 => x"bb",
          5012 => x"80",
          5013 => x"d0",
          5014 => x"53",
          5015 => x"c0",
          5016 => x"a6",
          5017 => x"bb",
          5018 => x"80",
          5019 => x"34",
          5020 => x"81",
          5021 => x"bb",
          5022 => x"77",
          5023 => x"76",
          5024 => x"82",
          5025 => x"54",
          5026 => x"34",
          5027 => x"34",
          5028 => x"08",
          5029 => x"22",
          5030 => x"80",
          5031 => x"83",
          5032 => x"70",
          5033 => x"51",
          5034 => x"88",
          5035 => x"89",
          5036 => x"bb",
          5037 => x"88",
          5038 => x"d4",
          5039 => x"11",
          5040 => x"77",
          5041 => x"76",
          5042 => x"89",
          5043 => x"ff",
          5044 => x"52",
          5045 => x"72",
          5046 => x"fb",
          5047 => x"82",
          5048 => x"ff",
          5049 => x"51",
          5050 => x"bb",
          5051 => x"3d",
          5052 => x"3d",
          5053 => x"05",
          5054 => x"05",
          5055 => x"71",
          5056 => x"d4",
          5057 => x"2b",
          5058 => x"83",
          5059 => x"70",
          5060 => x"33",
          5061 => x"07",
          5062 => x"ae",
          5063 => x"81",
          5064 => x"07",
          5065 => x"53",
          5066 => x"54",
          5067 => x"53",
          5068 => x"77",
          5069 => x"18",
          5070 => x"d4",
          5071 => x"88",
          5072 => x"70",
          5073 => x"74",
          5074 => x"82",
          5075 => x"70",
          5076 => x"81",
          5077 => x"88",
          5078 => x"83",
          5079 => x"f8",
          5080 => x"56",
          5081 => x"73",
          5082 => x"06",
          5083 => x"54",
          5084 => x"82",
          5085 => x"81",
          5086 => x"72",
          5087 => x"82",
          5088 => x"16",
          5089 => x"34",
          5090 => x"34",
          5091 => x"04",
          5092 => x"82",
          5093 => x"02",
          5094 => x"05",
          5095 => x"2b",
          5096 => x"11",
          5097 => x"33",
          5098 => x"71",
          5099 => x"58",
          5100 => x"55",
          5101 => x"84",
          5102 => x"13",
          5103 => x"2b",
          5104 => x"2a",
          5105 => x"52",
          5106 => x"34",
          5107 => x"34",
          5108 => x"08",
          5109 => x"11",
          5110 => x"33",
          5111 => x"71",
          5112 => x"56",
          5113 => x"72",
          5114 => x"33",
          5115 => x"71",
          5116 => x"70",
          5117 => x"56",
          5118 => x"86",
          5119 => x"87",
          5120 => x"bb",
          5121 => x"70",
          5122 => x"33",
          5123 => x"07",
          5124 => x"ff",
          5125 => x"2a",
          5126 => x"53",
          5127 => x"34",
          5128 => x"34",
          5129 => x"04",
          5130 => x"02",
          5131 => x"82",
          5132 => x"71",
          5133 => x"11",
          5134 => x"12",
          5135 => x"2b",
          5136 => x"29",
          5137 => x"81",
          5138 => x"98",
          5139 => x"2b",
          5140 => x"53",
          5141 => x"56",
          5142 => x"71",
          5143 => x"f6",
          5144 => x"fe",
          5145 => x"bb",
          5146 => x"16",
          5147 => x"12",
          5148 => x"2b",
          5149 => x"07",
          5150 => x"33",
          5151 => x"71",
          5152 => x"70",
          5153 => x"ff",
          5154 => x"52",
          5155 => x"5a",
          5156 => x"05",
          5157 => x"54",
          5158 => x"13",
          5159 => x"13",
          5160 => x"d4",
          5161 => x"70",
          5162 => x"33",
          5163 => x"71",
          5164 => x"56",
          5165 => x"72",
          5166 => x"81",
          5167 => x"88",
          5168 => x"81",
          5169 => x"70",
          5170 => x"51",
          5171 => x"72",
          5172 => x"81",
          5173 => x"3d",
          5174 => x"3d",
          5175 => x"d4",
          5176 => x"05",
          5177 => x"70",
          5178 => x"11",
          5179 => x"83",
          5180 => x"8b",
          5181 => x"2b",
          5182 => x"59",
          5183 => x"73",
          5184 => x"81",
          5185 => x"88",
          5186 => x"8c",
          5187 => x"22",
          5188 => x"88",
          5189 => x"53",
          5190 => x"73",
          5191 => x"14",
          5192 => x"d4",
          5193 => x"70",
          5194 => x"33",
          5195 => x"71",
          5196 => x"56",
          5197 => x"72",
          5198 => x"33",
          5199 => x"71",
          5200 => x"70",
          5201 => x"55",
          5202 => x"82",
          5203 => x"83",
          5204 => x"bb",
          5205 => x"82",
          5206 => x"12",
          5207 => x"2b",
          5208 => x"dc",
          5209 => x"87",
          5210 => x"f7",
          5211 => x"82",
          5212 => x"31",
          5213 => x"83",
          5214 => x"70",
          5215 => x"fd",
          5216 => x"bb",
          5217 => x"83",
          5218 => x"82",
          5219 => x"12",
          5220 => x"2b",
          5221 => x"07",
          5222 => x"33",
          5223 => x"71",
          5224 => x"90",
          5225 => x"42",
          5226 => x"5b",
          5227 => x"54",
          5228 => x"8d",
          5229 => x"80",
          5230 => x"fe",
          5231 => x"84",
          5232 => x"33",
          5233 => x"71",
          5234 => x"83",
          5235 => x"11",
          5236 => x"53",
          5237 => x"55",
          5238 => x"34",
          5239 => x"06",
          5240 => x"14",
          5241 => x"d4",
          5242 => x"84",
          5243 => x"13",
          5244 => x"2b",
          5245 => x"2a",
          5246 => x"56",
          5247 => x"16",
          5248 => x"16",
          5249 => x"d4",
          5250 => x"80",
          5251 => x"34",
          5252 => x"14",
          5253 => x"d4",
          5254 => x"84",
          5255 => x"85",
          5256 => x"bb",
          5257 => x"70",
          5258 => x"33",
          5259 => x"07",
          5260 => x"80",
          5261 => x"2a",
          5262 => x"56",
          5263 => x"34",
          5264 => x"34",
          5265 => x"04",
          5266 => x"73",
          5267 => x"d4",
          5268 => x"f7",
          5269 => x"80",
          5270 => x"71",
          5271 => x"3f",
          5272 => x"04",
          5273 => x"80",
          5274 => x"f8",
          5275 => x"bb",
          5276 => x"ff",
          5277 => x"bb",
          5278 => x"11",
          5279 => x"33",
          5280 => x"07",
          5281 => x"56",
          5282 => x"ff",
          5283 => x"78",
          5284 => x"38",
          5285 => x"17",
          5286 => x"12",
          5287 => x"2b",
          5288 => x"ff",
          5289 => x"31",
          5290 => x"ff",
          5291 => x"27",
          5292 => x"56",
          5293 => x"79",
          5294 => x"73",
          5295 => x"38",
          5296 => x"5b",
          5297 => x"85",
          5298 => x"88",
          5299 => x"54",
          5300 => x"78",
          5301 => x"2e",
          5302 => x"79",
          5303 => x"76",
          5304 => x"bb",
          5305 => x"70",
          5306 => x"33",
          5307 => x"07",
          5308 => x"ff",
          5309 => x"5a",
          5310 => x"73",
          5311 => x"38",
          5312 => x"54",
          5313 => x"81",
          5314 => x"54",
          5315 => x"81",
          5316 => x"7a",
          5317 => x"06",
          5318 => x"51",
          5319 => x"81",
          5320 => x"80",
          5321 => x"52",
          5322 => x"c6",
          5323 => x"d4",
          5324 => x"86",
          5325 => x"12",
          5326 => x"2b",
          5327 => x"07",
          5328 => x"55",
          5329 => x"17",
          5330 => x"ff",
          5331 => x"2a",
          5332 => x"54",
          5333 => x"34",
          5334 => x"06",
          5335 => x"15",
          5336 => x"d4",
          5337 => x"2b",
          5338 => x"1e",
          5339 => x"87",
          5340 => x"88",
          5341 => x"88",
          5342 => x"5e",
          5343 => x"54",
          5344 => x"34",
          5345 => x"34",
          5346 => x"08",
          5347 => x"11",
          5348 => x"33",
          5349 => x"71",
          5350 => x"53",
          5351 => x"74",
          5352 => x"86",
          5353 => x"87",
          5354 => x"bb",
          5355 => x"16",
          5356 => x"11",
          5357 => x"33",
          5358 => x"07",
          5359 => x"53",
          5360 => x"56",
          5361 => x"16",
          5362 => x"16",
          5363 => x"d4",
          5364 => x"05",
          5365 => x"bb",
          5366 => x"3d",
          5367 => x"3d",
          5368 => x"82",
          5369 => x"84",
          5370 => x"3f",
          5371 => x"80",
          5372 => x"71",
          5373 => x"3f",
          5374 => x"08",
          5375 => x"bb",
          5376 => x"3d",
          5377 => x"3d",
          5378 => x"40",
          5379 => x"42",
          5380 => x"d4",
          5381 => x"09",
          5382 => x"38",
          5383 => x"7b",
          5384 => x"51",
          5385 => x"82",
          5386 => x"54",
          5387 => x"7e",
          5388 => x"51",
          5389 => x"7e",
          5390 => x"39",
          5391 => x"8f",
          5392 => x"dc",
          5393 => x"ff",
          5394 => x"d4",
          5395 => x"31",
          5396 => x"83",
          5397 => x"70",
          5398 => x"11",
          5399 => x"12",
          5400 => x"2b",
          5401 => x"31",
          5402 => x"ff",
          5403 => x"29",
          5404 => x"88",
          5405 => x"33",
          5406 => x"71",
          5407 => x"70",
          5408 => x"44",
          5409 => x"41",
          5410 => x"5b",
          5411 => x"5b",
          5412 => x"25",
          5413 => x"81",
          5414 => x"75",
          5415 => x"ff",
          5416 => x"54",
          5417 => x"83",
          5418 => x"88",
          5419 => x"88",
          5420 => x"33",
          5421 => x"71",
          5422 => x"90",
          5423 => x"47",
          5424 => x"54",
          5425 => x"8b",
          5426 => x"31",
          5427 => x"ff",
          5428 => x"77",
          5429 => x"fe",
          5430 => x"54",
          5431 => x"09",
          5432 => x"38",
          5433 => x"c0",
          5434 => x"ff",
          5435 => x"81",
          5436 => x"8e",
          5437 => x"24",
          5438 => x"51",
          5439 => x"81",
          5440 => x"18",
          5441 => x"24",
          5442 => x"79",
          5443 => x"33",
          5444 => x"71",
          5445 => x"53",
          5446 => x"f4",
          5447 => x"78",
          5448 => x"3f",
          5449 => x"08",
          5450 => x"06",
          5451 => x"53",
          5452 => x"82",
          5453 => x"11",
          5454 => x"55",
          5455 => x"db",
          5456 => x"d4",
          5457 => x"05",
          5458 => x"ff",
          5459 => x"81",
          5460 => x"15",
          5461 => x"24",
          5462 => x"78",
          5463 => x"3f",
          5464 => x"08",
          5465 => x"33",
          5466 => x"71",
          5467 => x"53",
          5468 => x"9c",
          5469 => x"78",
          5470 => x"3f",
          5471 => x"08",
          5472 => x"06",
          5473 => x"53",
          5474 => x"82",
          5475 => x"11",
          5476 => x"55",
          5477 => x"83",
          5478 => x"d4",
          5479 => x"05",
          5480 => x"19",
          5481 => x"83",
          5482 => x"58",
          5483 => x"7f",
          5484 => x"b0",
          5485 => x"dc",
          5486 => x"bb",
          5487 => x"2e",
          5488 => x"53",
          5489 => x"bb",
          5490 => x"ff",
          5491 => x"73",
          5492 => x"3f",
          5493 => x"78",
          5494 => x"80",
          5495 => x"78",
          5496 => x"3f",
          5497 => x"2b",
          5498 => x"08",
          5499 => x"51",
          5500 => x"7b",
          5501 => x"bb",
          5502 => x"3d",
          5503 => x"3d",
          5504 => x"29",
          5505 => x"fb",
          5506 => x"bb",
          5507 => x"82",
          5508 => x"80",
          5509 => x"73",
          5510 => x"82",
          5511 => x"51",
          5512 => x"3f",
          5513 => x"dc",
          5514 => x"0d",
          5515 => x"0d",
          5516 => x"33",
          5517 => x"70",
          5518 => x"38",
          5519 => x"11",
          5520 => x"82",
          5521 => x"83",
          5522 => x"fc",
          5523 => x"9b",
          5524 => x"84",
          5525 => x"33",
          5526 => x"51",
          5527 => x"80",
          5528 => x"84",
          5529 => x"92",
          5530 => x"51",
          5531 => x"80",
          5532 => x"81",
          5533 => x"72",
          5534 => x"92",
          5535 => x"81",
          5536 => x"0b",
          5537 => x"8c",
          5538 => x"71",
          5539 => x"06",
          5540 => x"80",
          5541 => x"87",
          5542 => x"08",
          5543 => x"38",
          5544 => x"80",
          5545 => x"71",
          5546 => x"c0",
          5547 => x"51",
          5548 => x"87",
          5549 => x"bb",
          5550 => x"82",
          5551 => x"33",
          5552 => x"bb",
          5553 => x"3d",
          5554 => x"3d",
          5555 => x"64",
          5556 => x"bf",
          5557 => x"40",
          5558 => x"74",
          5559 => x"cd",
          5560 => x"dc",
          5561 => x"7a",
          5562 => x"81",
          5563 => x"72",
          5564 => x"87",
          5565 => x"11",
          5566 => x"8c",
          5567 => x"92",
          5568 => x"5a",
          5569 => x"58",
          5570 => x"c0",
          5571 => x"76",
          5572 => x"76",
          5573 => x"70",
          5574 => x"81",
          5575 => x"54",
          5576 => x"8e",
          5577 => x"52",
          5578 => x"81",
          5579 => x"81",
          5580 => x"74",
          5581 => x"53",
          5582 => x"83",
          5583 => x"78",
          5584 => x"8f",
          5585 => x"2e",
          5586 => x"c0",
          5587 => x"52",
          5588 => x"87",
          5589 => x"08",
          5590 => x"2e",
          5591 => x"84",
          5592 => x"38",
          5593 => x"87",
          5594 => x"15",
          5595 => x"70",
          5596 => x"52",
          5597 => x"ff",
          5598 => x"39",
          5599 => x"81",
          5600 => x"ff",
          5601 => x"57",
          5602 => x"90",
          5603 => x"80",
          5604 => x"71",
          5605 => x"78",
          5606 => x"38",
          5607 => x"80",
          5608 => x"80",
          5609 => x"81",
          5610 => x"72",
          5611 => x"0c",
          5612 => x"04",
          5613 => x"60",
          5614 => x"8c",
          5615 => x"33",
          5616 => x"5b",
          5617 => x"74",
          5618 => x"e1",
          5619 => x"dc",
          5620 => x"79",
          5621 => x"78",
          5622 => x"06",
          5623 => x"77",
          5624 => x"87",
          5625 => x"11",
          5626 => x"8c",
          5627 => x"92",
          5628 => x"59",
          5629 => x"85",
          5630 => x"98",
          5631 => x"7d",
          5632 => x"0c",
          5633 => x"08",
          5634 => x"70",
          5635 => x"53",
          5636 => x"2e",
          5637 => x"70",
          5638 => x"33",
          5639 => x"18",
          5640 => x"2a",
          5641 => x"51",
          5642 => x"2e",
          5643 => x"c0",
          5644 => x"52",
          5645 => x"87",
          5646 => x"08",
          5647 => x"2e",
          5648 => x"84",
          5649 => x"38",
          5650 => x"87",
          5651 => x"15",
          5652 => x"70",
          5653 => x"52",
          5654 => x"ff",
          5655 => x"39",
          5656 => x"81",
          5657 => x"80",
          5658 => x"52",
          5659 => x"90",
          5660 => x"80",
          5661 => x"71",
          5662 => x"7a",
          5663 => x"38",
          5664 => x"80",
          5665 => x"80",
          5666 => x"81",
          5667 => x"72",
          5668 => x"0c",
          5669 => x"04",
          5670 => x"7a",
          5671 => x"a3",
          5672 => x"88",
          5673 => x"33",
          5674 => x"56",
          5675 => x"3f",
          5676 => x"08",
          5677 => x"83",
          5678 => x"fe",
          5679 => x"87",
          5680 => x"0c",
          5681 => x"76",
          5682 => x"38",
          5683 => x"93",
          5684 => x"2b",
          5685 => x"8c",
          5686 => x"71",
          5687 => x"38",
          5688 => x"71",
          5689 => x"c6",
          5690 => x"39",
          5691 => x"81",
          5692 => x"06",
          5693 => x"71",
          5694 => x"38",
          5695 => x"8c",
          5696 => x"e8",
          5697 => x"98",
          5698 => x"71",
          5699 => x"73",
          5700 => x"92",
          5701 => x"72",
          5702 => x"06",
          5703 => x"f7",
          5704 => x"80",
          5705 => x"88",
          5706 => x"0c",
          5707 => x"80",
          5708 => x"56",
          5709 => x"56",
          5710 => x"82",
          5711 => x"88",
          5712 => x"fe",
          5713 => x"81",
          5714 => x"33",
          5715 => x"07",
          5716 => x"0c",
          5717 => x"3d",
          5718 => x"3d",
          5719 => x"11",
          5720 => x"33",
          5721 => x"71",
          5722 => x"81",
          5723 => x"72",
          5724 => x"75",
          5725 => x"82",
          5726 => x"52",
          5727 => x"54",
          5728 => x"0d",
          5729 => x"0d",
          5730 => x"05",
          5731 => x"52",
          5732 => x"70",
          5733 => x"34",
          5734 => x"51",
          5735 => x"83",
          5736 => x"ff",
          5737 => x"75",
          5738 => x"72",
          5739 => x"54",
          5740 => x"2a",
          5741 => x"70",
          5742 => x"34",
          5743 => x"51",
          5744 => x"81",
          5745 => x"70",
          5746 => x"70",
          5747 => x"3d",
          5748 => x"3d",
          5749 => x"77",
          5750 => x"70",
          5751 => x"38",
          5752 => x"05",
          5753 => x"70",
          5754 => x"34",
          5755 => x"eb",
          5756 => x"0d",
          5757 => x"0d",
          5758 => x"54",
          5759 => x"72",
          5760 => x"54",
          5761 => x"51",
          5762 => x"84",
          5763 => x"fc",
          5764 => x"77",
          5765 => x"53",
          5766 => x"05",
          5767 => x"70",
          5768 => x"33",
          5769 => x"ff",
          5770 => x"52",
          5771 => x"2e",
          5772 => x"80",
          5773 => x"71",
          5774 => x"0c",
          5775 => x"04",
          5776 => x"74",
          5777 => x"89",
          5778 => x"2e",
          5779 => x"11",
          5780 => x"52",
          5781 => x"70",
          5782 => x"dc",
          5783 => x"0d",
          5784 => x"82",
          5785 => x"04",
          5786 => x"bb",
          5787 => x"f7",
          5788 => x"56",
          5789 => x"17",
          5790 => x"74",
          5791 => x"d6",
          5792 => x"b0",
          5793 => x"b4",
          5794 => x"81",
          5795 => x"59",
          5796 => x"82",
          5797 => x"7a",
          5798 => x"06",
          5799 => x"bb",
          5800 => x"17",
          5801 => x"08",
          5802 => x"08",
          5803 => x"08",
          5804 => x"74",
          5805 => x"38",
          5806 => x"55",
          5807 => x"09",
          5808 => x"38",
          5809 => x"18",
          5810 => x"81",
          5811 => x"f9",
          5812 => x"39",
          5813 => x"82",
          5814 => x"8b",
          5815 => x"fa",
          5816 => x"7a",
          5817 => x"57",
          5818 => x"08",
          5819 => x"75",
          5820 => x"3f",
          5821 => x"08",
          5822 => x"dc",
          5823 => x"81",
          5824 => x"b4",
          5825 => x"16",
          5826 => x"be",
          5827 => x"dc",
          5828 => x"85",
          5829 => x"81",
          5830 => x"17",
          5831 => x"bb",
          5832 => x"3d",
          5833 => x"3d",
          5834 => x"52",
          5835 => x"3f",
          5836 => x"08",
          5837 => x"dc",
          5838 => x"38",
          5839 => x"74",
          5840 => x"81",
          5841 => x"38",
          5842 => x"59",
          5843 => x"09",
          5844 => x"e3",
          5845 => x"53",
          5846 => x"08",
          5847 => x"70",
          5848 => x"91",
          5849 => x"d5",
          5850 => x"17",
          5851 => x"3f",
          5852 => x"a4",
          5853 => x"51",
          5854 => x"86",
          5855 => x"f2",
          5856 => x"17",
          5857 => x"3f",
          5858 => x"52",
          5859 => x"51",
          5860 => x"8c",
          5861 => x"84",
          5862 => x"fc",
          5863 => x"17",
          5864 => x"70",
          5865 => x"79",
          5866 => x"52",
          5867 => x"51",
          5868 => x"77",
          5869 => x"80",
          5870 => x"81",
          5871 => x"f9",
          5872 => x"bb",
          5873 => x"2e",
          5874 => x"58",
          5875 => x"dc",
          5876 => x"0d",
          5877 => x"0d",
          5878 => x"98",
          5879 => x"05",
          5880 => x"80",
          5881 => x"27",
          5882 => x"14",
          5883 => x"29",
          5884 => x"05",
          5885 => x"82",
          5886 => x"87",
          5887 => x"f9",
          5888 => x"7a",
          5889 => x"54",
          5890 => x"27",
          5891 => x"76",
          5892 => x"27",
          5893 => x"ff",
          5894 => x"58",
          5895 => x"80",
          5896 => x"82",
          5897 => x"72",
          5898 => x"38",
          5899 => x"72",
          5900 => x"8e",
          5901 => x"39",
          5902 => x"17",
          5903 => x"a4",
          5904 => x"53",
          5905 => x"fd",
          5906 => x"bb",
          5907 => x"9f",
          5908 => x"ff",
          5909 => x"11",
          5910 => x"70",
          5911 => x"18",
          5912 => x"76",
          5913 => x"53",
          5914 => x"82",
          5915 => x"80",
          5916 => x"83",
          5917 => x"b4",
          5918 => x"88",
          5919 => x"79",
          5920 => x"84",
          5921 => x"58",
          5922 => x"80",
          5923 => x"9f",
          5924 => x"80",
          5925 => x"88",
          5926 => x"08",
          5927 => x"51",
          5928 => x"82",
          5929 => x"80",
          5930 => x"10",
          5931 => x"74",
          5932 => x"51",
          5933 => x"82",
          5934 => x"83",
          5935 => x"58",
          5936 => x"87",
          5937 => x"08",
          5938 => x"51",
          5939 => x"82",
          5940 => x"9b",
          5941 => x"2b",
          5942 => x"74",
          5943 => x"51",
          5944 => x"82",
          5945 => x"f0",
          5946 => x"83",
          5947 => x"77",
          5948 => x"0c",
          5949 => x"04",
          5950 => x"7a",
          5951 => x"58",
          5952 => x"81",
          5953 => x"9e",
          5954 => x"17",
          5955 => x"96",
          5956 => x"53",
          5957 => x"81",
          5958 => x"79",
          5959 => x"72",
          5960 => x"38",
          5961 => x"72",
          5962 => x"b8",
          5963 => x"39",
          5964 => x"17",
          5965 => x"a4",
          5966 => x"53",
          5967 => x"fb",
          5968 => x"bb",
          5969 => x"82",
          5970 => x"81",
          5971 => x"83",
          5972 => x"b4",
          5973 => x"78",
          5974 => x"56",
          5975 => x"76",
          5976 => x"38",
          5977 => x"9f",
          5978 => x"33",
          5979 => x"07",
          5980 => x"74",
          5981 => x"83",
          5982 => x"89",
          5983 => x"08",
          5984 => x"51",
          5985 => x"82",
          5986 => x"59",
          5987 => x"08",
          5988 => x"74",
          5989 => x"16",
          5990 => x"84",
          5991 => x"76",
          5992 => x"88",
          5993 => x"81",
          5994 => x"8f",
          5995 => x"53",
          5996 => x"80",
          5997 => x"88",
          5998 => x"08",
          5999 => x"51",
          6000 => x"82",
          6001 => x"59",
          6002 => x"08",
          6003 => x"77",
          6004 => x"06",
          6005 => x"83",
          6006 => x"05",
          6007 => x"f7",
          6008 => x"39",
          6009 => x"a4",
          6010 => x"52",
          6011 => x"ef",
          6012 => x"dc",
          6013 => x"bb",
          6014 => x"38",
          6015 => x"06",
          6016 => x"83",
          6017 => x"18",
          6018 => x"54",
          6019 => x"f6",
          6020 => x"bb",
          6021 => x"0a",
          6022 => x"52",
          6023 => x"83",
          6024 => x"83",
          6025 => x"82",
          6026 => x"8a",
          6027 => x"f8",
          6028 => x"7c",
          6029 => x"59",
          6030 => x"81",
          6031 => x"38",
          6032 => x"08",
          6033 => x"73",
          6034 => x"38",
          6035 => x"52",
          6036 => x"a4",
          6037 => x"dc",
          6038 => x"bb",
          6039 => x"f2",
          6040 => x"82",
          6041 => x"39",
          6042 => x"e6",
          6043 => x"dc",
          6044 => x"de",
          6045 => x"78",
          6046 => x"3f",
          6047 => x"08",
          6048 => x"dc",
          6049 => x"80",
          6050 => x"bb",
          6051 => x"2e",
          6052 => x"bb",
          6053 => x"2e",
          6054 => x"53",
          6055 => x"51",
          6056 => x"82",
          6057 => x"c5",
          6058 => x"08",
          6059 => x"18",
          6060 => x"57",
          6061 => x"90",
          6062 => x"90",
          6063 => x"16",
          6064 => x"54",
          6065 => x"34",
          6066 => x"78",
          6067 => x"38",
          6068 => x"82",
          6069 => x"8a",
          6070 => x"f6",
          6071 => x"7e",
          6072 => x"5b",
          6073 => x"38",
          6074 => x"58",
          6075 => x"88",
          6076 => x"08",
          6077 => x"38",
          6078 => x"39",
          6079 => x"51",
          6080 => x"81",
          6081 => x"bb",
          6082 => x"82",
          6083 => x"bb",
          6084 => x"82",
          6085 => x"ff",
          6086 => x"38",
          6087 => x"82",
          6088 => x"26",
          6089 => x"79",
          6090 => x"08",
          6091 => x"73",
          6092 => x"b9",
          6093 => x"2e",
          6094 => x"80",
          6095 => x"1a",
          6096 => x"08",
          6097 => x"38",
          6098 => x"52",
          6099 => x"af",
          6100 => x"82",
          6101 => x"81",
          6102 => x"06",
          6103 => x"bb",
          6104 => x"82",
          6105 => x"09",
          6106 => x"72",
          6107 => x"70",
          6108 => x"bb",
          6109 => x"51",
          6110 => x"73",
          6111 => x"82",
          6112 => x"80",
          6113 => x"8c",
          6114 => x"81",
          6115 => x"38",
          6116 => x"08",
          6117 => x"73",
          6118 => x"75",
          6119 => x"77",
          6120 => x"56",
          6121 => x"76",
          6122 => x"82",
          6123 => x"26",
          6124 => x"75",
          6125 => x"f8",
          6126 => x"bb",
          6127 => x"2e",
          6128 => x"59",
          6129 => x"08",
          6130 => x"81",
          6131 => x"82",
          6132 => x"59",
          6133 => x"08",
          6134 => x"70",
          6135 => x"25",
          6136 => x"51",
          6137 => x"73",
          6138 => x"75",
          6139 => x"81",
          6140 => x"38",
          6141 => x"f5",
          6142 => x"75",
          6143 => x"f9",
          6144 => x"bb",
          6145 => x"bb",
          6146 => x"70",
          6147 => x"08",
          6148 => x"51",
          6149 => x"80",
          6150 => x"73",
          6151 => x"38",
          6152 => x"52",
          6153 => x"d0",
          6154 => x"dc",
          6155 => x"a5",
          6156 => x"18",
          6157 => x"08",
          6158 => x"18",
          6159 => x"74",
          6160 => x"38",
          6161 => x"18",
          6162 => x"33",
          6163 => x"73",
          6164 => x"97",
          6165 => x"74",
          6166 => x"38",
          6167 => x"55",
          6168 => x"bb",
          6169 => x"85",
          6170 => x"75",
          6171 => x"bb",
          6172 => x"3d",
          6173 => x"3d",
          6174 => x"52",
          6175 => x"3f",
          6176 => x"08",
          6177 => x"82",
          6178 => x"80",
          6179 => x"52",
          6180 => x"c1",
          6181 => x"dc",
          6182 => x"dc",
          6183 => x"0c",
          6184 => x"53",
          6185 => x"15",
          6186 => x"f2",
          6187 => x"56",
          6188 => x"16",
          6189 => x"22",
          6190 => x"27",
          6191 => x"54",
          6192 => x"76",
          6193 => x"33",
          6194 => x"3f",
          6195 => x"08",
          6196 => x"38",
          6197 => x"76",
          6198 => x"70",
          6199 => x"9f",
          6200 => x"56",
          6201 => x"bb",
          6202 => x"3d",
          6203 => x"3d",
          6204 => x"71",
          6205 => x"57",
          6206 => x"0a",
          6207 => x"38",
          6208 => x"53",
          6209 => x"38",
          6210 => x"0c",
          6211 => x"54",
          6212 => x"75",
          6213 => x"73",
          6214 => x"a8",
          6215 => x"73",
          6216 => x"85",
          6217 => x"0b",
          6218 => x"5a",
          6219 => x"27",
          6220 => x"a8",
          6221 => x"18",
          6222 => x"39",
          6223 => x"70",
          6224 => x"58",
          6225 => x"b2",
          6226 => x"76",
          6227 => x"3f",
          6228 => x"08",
          6229 => x"dc",
          6230 => x"bd",
          6231 => x"82",
          6232 => x"27",
          6233 => x"16",
          6234 => x"dc",
          6235 => x"38",
          6236 => x"39",
          6237 => x"55",
          6238 => x"52",
          6239 => x"d5",
          6240 => x"dc",
          6241 => x"0c",
          6242 => x"0c",
          6243 => x"53",
          6244 => x"80",
          6245 => x"85",
          6246 => x"94",
          6247 => x"2a",
          6248 => x"0c",
          6249 => x"06",
          6250 => x"9c",
          6251 => x"58",
          6252 => x"dc",
          6253 => x"0d",
          6254 => x"0d",
          6255 => x"90",
          6256 => x"05",
          6257 => x"f0",
          6258 => x"27",
          6259 => x"0b",
          6260 => x"98",
          6261 => x"84",
          6262 => x"2e",
          6263 => x"76",
          6264 => x"58",
          6265 => x"38",
          6266 => x"15",
          6267 => x"08",
          6268 => x"38",
          6269 => x"88",
          6270 => x"53",
          6271 => x"81",
          6272 => x"c0",
          6273 => x"22",
          6274 => x"89",
          6275 => x"72",
          6276 => x"74",
          6277 => x"f3",
          6278 => x"bb",
          6279 => x"82",
          6280 => x"82",
          6281 => x"27",
          6282 => x"81",
          6283 => x"dc",
          6284 => x"80",
          6285 => x"16",
          6286 => x"dc",
          6287 => x"ca",
          6288 => x"38",
          6289 => x"0c",
          6290 => x"dd",
          6291 => x"08",
          6292 => x"f9",
          6293 => x"bb",
          6294 => x"87",
          6295 => x"dc",
          6296 => x"80",
          6297 => x"55",
          6298 => x"08",
          6299 => x"38",
          6300 => x"bb",
          6301 => x"2e",
          6302 => x"bb",
          6303 => x"75",
          6304 => x"3f",
          6305 => x"08",
          6306 => x"94",
          6307 => x"52",
          6308 => x"c1",
          6309 => x"dc",
          6310 => x"0c",
          6311 => x"0c",
          6312 => x"05",
          6313 => x"80",
          6314 => x"bb",
          6315 => x"3d",
          6316 => x"3d",
          6317 => x"71",
          6318 => x"57",
          6319 => x"51",
          6320 => x"82",
          6321 => x"54",
          6322 => x"08",
          6323 => x"82",
          6324 => x"56",
          6325 => x"52",
          6326 => x"83",
          6327 => x"dc",
          6328 => x"bb",
          6329 => x"d2",
          6330 => x"dc",
          6331 => x"08",
          6332 => x"54",
          6333 => x"e5",
          6334 => x"06",
          6335 => x"58",
          6336 => x"08",
          6337 => x"38",
          6338 => x"75",
          6339 => x"80",
          6340 => x"81",
          6341 => x"7a",
          6342 => x"06",
          6343 => x"39",
          6344 => x"08",
          6345 => x"76",
          6346 => x"3f",
          6347 => x"08",
          6348 => x"dc",
          6349 => x"ff",
          6350 => x"84",
          6351 => x"06",
          6352 => x"54",
          6353 => x"dc",
          6354 => x"0d",
          6355 => x"0d",
          6356 => x"52",
          6357 => x"3f",
          6358 => x"08",
          6359 => x"06",
          6360 => x"51",
          6361 => x"83",
          6362 => x"06",
          6363 => x"14",
          6364 => x"3f",
          6365 => x"08",
          6366 => x"07",
          6367 => x"bb",
          6368 => x"3d",
          6369 => x"3d",
          6370 => x"70",
          6371 => x"06",
          6372 => x"53",
          6373 => x"ed",
          6374 => x"33",
          6375 => x"83",
          6376 => x"06",
          6377 => x"90",
          6378 => x"15",
          6379 => x"3f",
          6380 => x"04",
          6381 => x"7b",
          6382 => x"84",
          6383 => x"58",
          6384 => x"80",
          6385 => x"38",
          6386 => x"52",
          6387 => x"8f",
          6388 => x"dc",
          6389 => x"bb",
          6390 => x"f5",
          6391 => x"08",
          6392 => x"53",
          6393 => x"84",
          6394 => x"39",
          6395 => x"70",
          6396 => x"81",
          6397 => x"51",
          6398 => x"16",
          6399 => x"dc",
          6400 => x"81",
          6401 => x"38",
          6402 => x"ae",
          6403 => x"81",
          6404 => x"54",
          6405 => x"2e",
          6406 => x"8f",
          6407 => x"82",
          6408 => x"76",
          6409 => x"54",
          6410 => x"09",
          6411 => x"38",
          6412 => x"7a",
          6413 => x"80",
          6414 => x"fa",
          6415 => x"bb",
          6416 => x"82",
          6417 => x"89",
          6418 => x"08",
          6419 => x"86",
          6420 => x"98",
          6421 => x"82",
          6422 => x"8b",
          6423 => x"fb",
          6424 => x"70",
          6425 => x"81",
          6426 => x"fc",
          6427 => x"bb",
          6428 => x"82",
          6429 => x"b4",
          6430 => x"08",
          6431 => x"ec",
          6432 => x"bb",
          6433 => x"82",
          6434 => x"a0",
          6435 => x"82",
          6436 => x"52",
          6437 => x"51",
          6438 => x"8b",
          6439 => x"52",
          6440 => x"51",
          6441 => x"81",
          6442 => x"34",
          6443 => x"dc",
          6444 => x"0d",
          6445 => x"0d",
          6446 => x"98",
          6447 => x"70",
          6448 => x"ec",
          6449 => x"bb",
          6450 => x"38",
          6451 => x"53",
          6452 => x"81",
          6453 => x"34",
          6454 => x"04",
          6455 => x"78",
          6456 => x"80",
          6457 => x"34",
          6458 => x"80",
          6459 => x"38",
          6460 => x"18",
          6461 => x"9c",
          6462 => x"70",
          6463 => x"56",
          6464 => x"a0",
          6465 => x"71",
          6466 => x"81",
          6467 => x"81",
          6468 => x"89",
          6469 => x"06",
          6470 => x"73",
          6471 => x"55",
          6472 => x"55",
          6473 => x"81",
          6474 => x"81",
          6475 => x"74",
          6476 => x"75",
          6477 => x"52",
          6478 => x"13",
          6479 => x"08",
          6480 => x"33",
          6481 => x"9c",
          6482 => x"11",
          6483 => x"8a",
          6484 => x"dc",
          6485 => x"96",
          6486 => x"e7",
          6487 => x"dc",
          6488 => x"23",
          6489 => x"e7",
          6490 => x"bb",
          6491 => x"17",
          6492 => x"0d",
          6493 => x"0d",
          6494 => x"5e",
          6495 => x"70",
          6496 => x"55",
          6497 => x"83",
          6498 => x"73",
          6499 => x"91",
          6500 => x"2e",
          6501 => x"1d",
          6502 => x"0c",
          6503 => x"15",
          6504 => x"70",
          6505 => x"56",
          6506 => x"09",
          6507 => x"38",
          6508 => x"80",
          6509 => x"30",
          6510 => x"78",
          6511 => x"54",
          6512 => x"73",
          6513 => x"60",
          6514 => x"54",
          6515 => x"96",
          6516 => x"0b",
          6517 => x"80",
          6518 => x"f6",
          6519 => x"bb",
          6520 => x"85",
          6521 => x"3d",
          6522 => x"5c",
          6523 => x"53",
          6524 => x"51",
          6525 => x"80",
          6526 => x"88",
          6527 => x"5c",
          6528 => x"09",
          6529 => x"d4",
          6530 => x"70",
          6531 => x"71",
          6532 => x"30",
          6533 => x"73",
          6534 => x"51",
          6535 => x"57",
          6536 => x"38",
          6537 => x"75",
          6538 => x"17",
          6539 => x"75",
          6540 => x"30",
          6541 => x"51",
          6542 => x"80",
          6543 => x"38",
          6544 => x"87",
          6545 => x"26",
          6546 => x"77",
          6547 => x"a4",
          6548 => x"27",
          6549 => x"a0",
          6550 => x"39",
          6551 => x"33",
          6552 => x"57",
          6553 => x"27",
          6554 => x"75",
          6555 => x"30",
          6556 => x"32",
          6557 => x"80",
          6558 => x"25",
          6559 => x"56",
          6560 => x"80",
          6561 => x"84",
          6562 => x"58",
          6563 => x"70",
          6564 => x"55",
          6565 => x"09",
          6566 => x"38",
          6567 => x"80",
          6568 => x"30",
          6569 => x"77",
          6570 => x"54",
          6571 => x"81",
          6572 => x"ae",
          6573 => x"06",
          6574 => x"54",
          6575 => x"74",
          6576 => x"80",
          6577 => x"7b",
          6578 => x"30",
          6579 => x"70",
          6580 => x"25",
          6581 => x"07",
          6582 => x"51",
          6583 => x"a7",
          6584 => x"8b",
          6585 => x"39",
          6586 => x"54",
          6587 => x"8c",
          6588 => x"ff",
          6589 => x"a4",
          6590 => x"54",
          6591 => x"e1",
          6592 => x"dc",
          6593 => x"b2",
          6594 => x"70",
          6595 => x"71",
          6596 => x"54",
          6597 => x"82",
          6598 => x"80",
          6599 => x"38",
          6600 => x"76",
          6601 => x"df",
          6602 => x"54",
          6603 => x"81",
          6604 => x"55",
          6605 => x"34",
          6606 => x"52",
          6607 => x"51",
          6608 => x"82",
          6609 => x"bf",
          6610 => x"16",
          6611 => x"26",
          6612 => x"16",
          6613 => x"06",
          6614 => x"17",
          6615 => x"34",
          6616 => x"fd",
          6617 => x"19",
          6618 => x"80",
          6619 => x"79",
          6620 => x"81",
          6621 => x"81",
          6622 => x"85",
          6623 => x"54",
          6624 => x"8f",
          6625 => x"86",
          6626 => x"39",
          6627 => x"f3",
          6628 => x"73",
          6629 => x"80",
          6630 => x"52",
          6631 => x"ce",
          6632 => x"dc",
          6633 => x"bb",
          6634 => x"d7",
          6635 => x"08",
          6636 => x"e6",
          6637 => x"bb",
          6638 => x"82",
          6639 => x"80",
          6640 => x"1b",
          6641 => x"55",
          6642 => x"2e",
          6643 => x"8b",
          6644 => x"06",
          6645 => x"1c",
          6646 => x"33",
          6647 => x"70",
          6648 => x"55",
          6649 => x"38",
          6650 => x"52",
          6651 => x"9f",
          6652 => x"dc",
          6653 => x"8b",
          6654 => x"7a",
          6655 => x"3f",
          6656 => x"75",
          6657 => x"57",
          6658 => x"2e",
          6659 => x"84",
          6660 => x"06",
          6661 => x"75",
          6662 => x"81",
          6663 => x"2a",
          6664 => x"73",
          6665 => x"38",
          6666 => x"54",
          6667 => x"fb",
          6668 => x"80",
          6669 => x"34",
          6670 => x"c1",
          6671 => x"06",
          6672 => x"38",
          6673 => x"39",
          6674 => x"70",
          6675 => x"54",
          6676 => x"86",
          6677 => x"84",
          6678 => x"06",
          6679 => x"73",
          6680 => x"38",
          6681 => x"83",
          6682 => x"b4",
          6683 => x"51",
          6684 => x"82",
          6685 => x"88",
          6686 => x"ea",
          6687 => x"bb",
          6688 => x"3d",
          6689 => x"3d",
          6690 => x"ff",
          6691 => x"71",
          6692 => x"5c",
          6693 => x"80",
          6694 => x"38",
          6695 => x"05",
          6696 => x"a0",
          6697 => x"71",
          6698 => x"38",
          6699 => x"71",
          6700 => x"81",
          6701 => x"38",
          6702 => x"11",
          6703 => x"06",
          6704 => x"70",
          6705 => x"38",
          6706 => x"81",
          6707 => x"05",
          6708 => x"76",
          6709 => x"38",
          6710 => x"b5",
          6711 => x"77",
          6712 => x"57",
          6713 => x"05",
          6714 => x"70",
          6715 => x"33",
          6716 => x"53",
          6717 => x"99",
          6718 => x"e0",
          6719 => x"ff",
          6720 => x"ff",
          6721 => x"70",
          6722 => x"38",
          6723 => x"81",
          6724 => x"51",
          6725 => x"9f",
          6726 => x"72",
          6727 => x"81",
          6728 => x"70",
          6729 => x"72",
          6730 => x"32",
          6731 => x"72",
          6732 => x"73",
          6733 => x"53",
          6734 => x"70",
          6735 => x"38",
          6736 => x"19",
          6737 => x"75",
          6738 => x"38",
          6739 => x"83",
          6740 => x"74",
          6741 => x"59",
          6742 => x"39",
          6743 => x"33",
          6744 => x"bb",
          6745 => x"3d",
          6746 => x"3d",
          6747 => x"80",
          6748 => x"34",
          6749 => x"17",
          6750 => x"75",
          6751 => x"3f",
          6752 => x"bb",
          6753 => x"80",
          6754 => x"16",
          6755 => x"3f",
          6756 => x"08",
          6757 => x"06",
          6758 => x"73",
          6759 => x"2e",
          6760 => x"80",
          6761 => x"0b",
          6762 => x"56",
          6763 => x"e9",
          6764 => x"06",
          6765 => x"57",
          6766 => x"32",
          6767 => x"80",
          6768 => x"51",
          6769 => x"8a",
          6770 => x"e8",
          6771 => x"06",
          6772 => x"53",
          6773 => x"52",
          6774 => x"51",
          6775 => x"82",
          6776 => x"55",
          6777 => x"08",
          6778 => x"38",
          6779 => x"b4",
          6780 => x"86",
          6781 => x"97",
          6782 => x"dc",
          6783 => x"bb",
          6784 => x"2e",
          6785 => x"55",
          6786 => x"dc",
          6787 => x"0d",
          6788 => x"0d",
          6789 => x"05",
          6790 => x"33",
          6791 => x"75",
          6792 => x"fc",
          6793 => x"bb",
          6794 => x"8b",
          6795 => x"82",
          6796 => x"24",
          6797 => x"82",
          6798 => x"84",
          6799 => x"94",
          6800 => x"55",
          6801 => x"73",
          6802 => x"e6",
          6803 => x"0c",
          6804 => x"06",
          6805 => x"57",
          6806 => x"ae",
          6807 => x"33",
          6808 => x"3f",
          6809 => x"08",
          6810 => x"70",
          6811 => x"55",
          6812 => x"76",
          6813 => x"b8",
          6814 => x"2a",
          6815 => x"51",
          6816 => x"72",
          6817 => x"86",
          6818 => x"74",
          6819 => x"15",
          6820 => x"81",
          6821 => x"d7",
          6822 => x"bb",
          6823 => x"ff",
          6824 => x"06",
          6825 => x"56",
          6826 => x"38",
          6827 => x"8f",
          6828 => x"2a",
          6829 => x"51",
          6830 => x"72",
          6831 => x"80",
          6832 => x"52",
          6833 => x"3f",
          6834 => x"08",
          6835 => x"57",
          6836 => x"09",
          6837 => x"e2",
          6838 => x"74",
          6839 => x"56",
          6840 => x"33",
          6841 => x"72",
          6842 => x"38",
          6843 => x"51",
          6844 => x"82",
          6845 => x"57",
          6846 => x"84",
          6847 => x"ff",
          6848 => x"56",
          6849 => x"25",
          6850 => x"0b",
          6851 => x"56",
          6852 => x"05",
          6853 => x"83",
          6854 => x"2e",
          6855 => x"52",
          6856 => x"c6",
          6857 => x"dc",
          6858 => x"06",
          6859 => x"27",
          6860 => x"16",
          6861 => x"27",
          6862 => x"56",
          6863 => x"84",
          6864 => x"56",
          6865 => x"84",
          6866 => x"14",
          6867 => x"3f",
          6868 => x"08",
          6869 => x"06",
          6870 => x"80",
          6871 => x"06",
          6872 => x"80",
          6873 => x"db",
          6874 => x"bb",
          6875 => x"ff",
          6876 => x"77",
          6877 => x"d8",
          6878 => x"de",
          6879 => x"dc",
          6880 => x"9c",
          6881 => x"c4",
          6882 => x"15",
          6883 => x"14",
          6884 => x"70",
          6885 => x"51",
          6886 => x"56",
          6887 => x"84",
          6888 => x"81",
          6889 => x"71",
          6890 => x"16",
          6891 => x"53",
          6892 => x"23",
          6893 => x"8b",
          6894 => x"73",
          6895 => x"80",
          6896 => x"8d",
          6897 => x"39",
          6898 => x"51",
          6899 => x"82",
          6900 => x"53",
          6901 => x"08",
          6902 => x"72",
          6903 => x"8d",
          6904 => x"ce",
          6905 => x"14",
          6906 => x"3f",
          6907 => x"08",
          6908 => x"06",
          6909 => x"38",
          6910 => x"51",
          6911 => x"82",
          6912 => x"55",
          6913 => x"51",
          6914 => x"82",
          6915 => x"83",
          6916 => x"53",
          6917 => x"80",
          6918 => x"38",
          6919 => x"78",
          6920 => x"2a",
          6921 => x"78",
          6922 => x"86",
          6923 => x"22",
          6924 => x"31",
          6925 => x"cb",
          6926 => x"dc",
          6927 => x"bb",
          6928 => x"2e",
          6929 => x"82",
          6930 => x"80",
          6931 => x"f5",
          6932 => x"83",
          6933 => x"ff",
          6934 => x"38",
          6935 => x"9f",
          6936 => x"38",
          6937 => x"39",
          6938 => x"80",
          6939 => x"38",
          6940 => x"98",
          6941 => x"a0",
          6942 => x"1c",
          6943 => x"0c",
          6944 => x"17",
          6945 => x"76",
          6946 => x"81",
          6947 => x"80",
          6948 => x"d9",
          6949 => x"bb",
          6950 => x"ff",
          6951 => x"8d",
          6952 => x"8e",
          6953 => x"8a",
          6954 => x"14",
          6955 => x"3f",
          6956 => x"08",
          6957 => x"74",
          6958 => x"a2",
          6959 => x"79",
          6960 => x"ee",
          6961 => x"a8",
          6962 => x"15",
          6963 => x"2e",
          6964 => x"10",
          6965 => x"2a",
          6966 => x"05",
          6967 => x"ff",
          6968 => x"53",
          6969 => x"9c",
          6970 => x"81",
          6971 => x"0b",
          6972 => x"ff",
          6973 => x"0c",
          6974 => x"84",
          6975 => x"83",
          6976 => x"06",
          6977 => x"80",
          6978 => x"d8",
          6979 => x"bb",
          6980 => x"ff",
          6981 => x"72",
          6982 => x"81",
          6983 => x"38",
          6984 => x"73",
          6985 => x"3f",
          6986 => x"08",
          6987 => x"82",
          6988 => x"84",
          6989 => x"b2",
          6990 => x"87",
          6991 => x"dc",
          6992 => x"ff",
          6993 => x"82",
          6994 => x"09",
          6995 => x"c8",
          6996 => x"51",
          6997 => x"82",
          6998 => x"84",
          6999 => x"d2",
          7000 => x"06",
          7001 => x"98",
          7002 => x"ee",
          7003 => x"dc",
          7004 => x"85",
          7005 => x"09",
          7006 => x"38",
          7007 => x"51",
          7008 => x"82",
          7009 => x"90",
          7010 => x"a0",
          7011 => x"ca",
          7012 => x"dc",
          7013 => x"0c",
          7014 => x"82",
          7015 => x"81",
          7016 => x"82",
          7017 => x"72",
          7018 => x"80",
          7019 => x"0c",
          7020 => x"82",
          7021 => x"90",
          7022 => x"fb",
          7023 => x"54",
          7024 => x"80",
          7025 => x"73",
          7026 => x"80",
          7027 => x"72",
          7028 => x"80",
          7029 => x"86",
          7030 => x"15",
          7031 => x"71",
          7032 => x"81",
          7033 => x"81",
          7034 => x"d0",
          7035 => x"bb",
          7036 => x"06",
          7037 => x"38",
          7038 => x"54",
          7039 => x"80",
          7040 => x"71",
          7041 => x"82",
          7042 => x"87",
          7043 => x"fa",
          7044 => x"ab",
          7045 => x"58",
          7046 => x"05",
          7047 => x"e6",
          7048 => x"80",
          7049 => x"dc",
          7050 => x"38",
          7051 => x"08",
          7052 => x"d3",
          7053 => x"08",
          7054 => x"80",
          7055 => x"80",
          7056 => x"54",
          7057 => x"84",
          7058 => x"34",
          7059 => x"75",
          7060 => x"2e",
          7061 => x"53",
          7062 => x"53",
          7063 => x"f7",
          7064 => x"bb",
          7065 => x"73",
          7066 => x"0c",
          7067 => x"04",
          7068 => x"67",
          7069 => x"80",
          7070 => x"59",
          7071 => x"78",
          7072 => x"c8",
          7073 => x"06",
          7074 => x"3d",
          7075 => x"99",
          7076 => x"52",
          7077 => x"3f",
          7078 => x"08",
          7079 => x"dc",
          7080 => x"38",
          7081 => x"52",
          7082 => x"52",
          7083 => x"3f",
          7084 => x"08",
          7085 => x"dc",
          7086 => x"02",
          7087 => x"33",
          7088 => x"55",
          7089 => x"25",
          7090 => x"55",
          7091 => x"54",
          7092 => x"81",
          7093 => x"80",
          7094 => x"74",
          7095 => x"81",
          7096 => x"75",
          7097 => x"3f",
          7098 => x"08",
          7099 => x"02",
          7100 => x"91",
          7101 => x"81",
          7102 => x"82",
          7103 => x"06",
          7104 => x"80",
          7105 => x"88",
          7106 => x"39",
          7107 => x"58",
          7108 => x"38",
          7109 => x"70",
          7110 => x"54",
          7111 => x"81",
          7112 => x"52",
          7113 => x"a5",
          7114 => x"dc",
          7115 => x"88",
          7116 => x"62",
          7117 => x"d4",
          7118 => x"54",
          7119 => x"15",
          7120 => x"62",
          7121 => x"e8",
          7122 => x"52",
          7123 => x"51",
          7124 => x"7a",
          7125 => x"83",
          7126 => x"80",
          7127 => x"38",
          7128 => x"08",
          7129 => x"53",
          7130 => x"3d",
          7131 => x"dd",
          7132 => x"bb",
          7133 => x"82",
          7134 => x"82",
          7135 => x"39",
          7136 => x"38",
          7137 => x"33",
          7138 => x"70",
          7139 => x"55",
          7140 => x"2e",
          7141 => x"55",
          7142 => x"77",
          7143 => x"81",
          7144 => x"73",
          7145 => x"38",
          7146 => x"54",
          7147 => x"a0",
          7148 => x"82",
          7149 => x"52",
          7150 => x"a3",
          7151 => x"dc",
          7152 => x"18",
          7153 => x"55",
          7154 => x"dc",
          7155 => x"38",
          7156 => x"70",
          7157 => x"54",
          7158 => x"86",
          7159 => x"c0",
          7160 => x"b0",
          7161 => x"1b",
          7162 => x"1b",
          7163 => x"70",
          7164 => x"d9",
          7165 => x"dc",
          7166 => x"dc",
          7167 => x"0c",
          7168 => x"52",
          7169 => x"3f",
          7170 => x"08",
          7171 => x"08",
          7172 => x"77",
          7173 => x"86",
          7174 => x"1a",
          7175 => x"1a",
          7176 => x"91",
          7177 => x"0b",
          7178 => x"80",
          7179 => x"0c",
          7180 => x"70",
          7181 => x"54",
          7182 => x"81",
          7183 => x"bb",
          7184 => x"2e",
          7185 => x"82",
          7186 => x"94",
          7187 => x"17",
          7188 => x"2b",
          7189 => x"57",
          7190 => x"52",
          7191 => x"9f",
          7192 => x"dc",
          7193 => x"bb",
          7194 => x"26",
          7195 => x"55",
          7196 => x"08",
          7197 => x"81",
          7198 => x"79",
          7199 => x"31",
          7200 => x"70",
          7201 => x"25",
          7202 => x"76",
          7203 => x"81",
          7204 => x"55",
          7205 => x"38",
          7206 => x"0c",
          7207 => x"75",
          7208 => x"54",
          7209 => x"a2",
          7210 => x"7a",
          7211 => x"3f",
          7212 => x"08",
          7213 => x"55",
          7214 => x"89",
          7215 => x"dc",
          7216 => x"1a",
          7217 => x"80",
          7218 => x"54",
          7219 => x"dc",
          7220 => x"0d",
          7221 => x"0d",
          7222 => x"64",
          7223 => x"59",
          7224 => x"90",
          7225 => x"52",
          7226 => x"cf",
          7227 => x"dc",
          7228 => x"bb",
          7229 => x"38",
          7230 => x"55",
          7231 => x"86",
          7232 => x"82",
          7233 => x"19",
          7234 => x"55",
          7235 => x"80",
          7236 => x"38",
          7237 => x"0b",
          7238 => x"82",
          7239 => x"39",
          7240 => x"1a",
          7241 => x"82",
          7242 => x"19",
          7243 => x"08",
          7244 => x"7c",
          7245 => x"74",
          7246 => x"2e",
          7247 => x"94",
          7248 => x"83",
          7249 => x"56",
          7250 => x"38",
          7251 => x"22",
          7252 => x"89",
          7253 => x"55",
          7254 => x"75",
          7255 => x"19",
          7256 => x"39",
          7257 => x"52",
          7258 => x"93",
          7259 => x"dc",
          7260 => x"75",
          7261 => x"38",
          7262 => x"ff",
          7263 => x"98",
          7264 => x"19",
          7265 => x"51",
          7266 => x"82",
          7267 => x"80",
          7268 => x"38",
          7269 => x"08",
          7270 => x"2a",
          7271 => x"80",
          7272 => x"38",
          7273 => x"8a",
          7274 => x"5c",
          7275 => x"27",
          7276 => x"7a",
          7277 => x"54",
          7278 => x"52",
          7279 => x"51",
          7280 => x"82",
          7281 => x"fe",
          7282 => x"83",
          7283 => x"56",
          7284 => x"9f",
          7285 => x"08",
          7286 => x"74",
          7287 => x"38",
          7288 => x"b4",
          7289 => x"16",
          7290 => x"89",
          7291 => x"51",
          7292 => x"77",
          7293 => x"b9",
          7294 => x"1a",
          7295 => x"08",
          7296 => x"84",
          7297 => x"57",
          7298 => x"27",
          7299 => x"56",
          7300 => x"52",
          7301 => x"c7",
          7302 => x"dc",
          7303 => x"38",
          7304 => x"19",
          7305 => x"06",
          7306 => x"52",
          7307 => x"a2",
          7308 => x"31",
          7309 => x"7f",
          7310 => x"94",
          7311 => x"94",
          7312 => x"5c",
          7313 => x"80",
          7314 => x"bb",
          7315 => x"3d",
          7316 => x"3d",
          7317 => x"65",
          7318 => x"5d",
          7319 => x"0c",
          7320 => x"05",
          7321 => x"f6",
          7322 => x"bb",
          7323 => x"82",
          7324 => x"8a",
          7325 => x"33",
          7326 => x"2e",
          7327 => x"56",
          7328 => x"90",
          7329 => x"81",
          7330 => x"06",
          7331 => x"87",
          7332 => x"2e",
          7333 => x"95",
          7334 => x"91",
          7335 => x"56",
          7336 => x"81",
          7337 => x"34",
          7338 => x"8e",
          7339 => x"08",
          7340 => x"56",
          7341 => x"84",
          7342 => x"5c",
          7343 => x"82",
          7344 => x"18",
          7345 => x"ff",
          7346 => x"74",
          7347 => x"7e",
          7348 => x"ff",
          7349 => x"2a",
          7350 => x"7a",
          7351 => x"8c",
          7352 => x"08",
          7353 => x"38",
          7354 => x"39",
          7355 => x"52",
          7356 => x"e7",
          7357 => x"dc",
          7358 => x"bb",
          7359 => x"2e",
          7360 => x"74",
          7361 => x"91",
          7362 => x"2e",
          7363 => x"74",
          7364 => x"88",
          7365 => x"38",
          7366 => x"0c",
          7367 => x"15",
          7368 => x"08",
          7369 => x"06",
          7370 => x"51",
          7371 => x"82",
          7372 => x"fe",
          7373 => x"18",
          7374 => x"51",
          7375 => x"82",
          7376 => x"80",
          7377 => x"38",
          7378 => x"08",
          7379 => x"2a",
          7380 => x"80",
          7381 => x"38",
          7382 => x"8a",
          7383 => x"5b",
          7384 => x"27",
          7385 => x"7b",
          7386 => x"54",
          7387 => x"52",
          7388 => x"51",
          7389 => x"82",
          7390 => x"fe",
          7391 => x"b0",
          7392 => x"31",
          7393 => x"79",
          7394 => x"84",
          7395 => x"16",
          7396 => x"89",
          7397 => x"52",
          7398 => x"cc",
          7399 => x"55",
          7400 => x"16",
          7401 => x"2b",
          7402 => x"39",
          7403 => x"94",
          7404 => x"93",
          7405 => x"cd",
          7406 => x"bb",
          7407 => x"e3",
          7408 => x"b0",
          7409 => x"76",
          7410 => x"94",
          7411 => x"ff",
          7412 => x"71",
          7413 => x"7b",
          7414 => x"38",
          7415 => x"18",
          7416 => x"51",
          7417 => x"82",
          7418 => x"fd",
          7419 => x"53",
          7420 => x"18",
          7421 => x"06",
          7422 => x"51",
          7423 => x"7e",
          7424 => x"83",
          7425 => x"76",
          7426 => x"17",
          7427 => x"1e",
          7428 => x"18",
          7429 => x"0c",
          7430 => x"58",
          7431 => x"74",
          7432 => x"38",
          7433 => x"8c",
          7434 => x"90",
          7435 => x"33",
          7436 => x"55",
          7437 => x"34",
          7438 => x"82",
          7439 => x"90",
          7440 => x"f8",
          7441 => x"8b",
          7442 => x"53",
          7443 => x"f2",
          7444 => x"bb",
          7445 => x"82",
          7446 => x"80",
          7447 => x"16",
          7448 => x"2a",
          7449 => x"51",
          7450 => x"80",
          7451 => x"38",
          7452 => x"52",
          7453 => x"e7",
          7454 => x"dc",
          7455 => x"bb",
          7456 => x"d4",
          7457 => x"08",
          7458 => x"a0",
          7459 => x"73",
          7460 => x"88",
          7461 => x"74",
          7462 => x"51",
          7463 => x"8c",
          7464 => x"9c",
          7465 => x"fb",
          7466 => x"b2",
          7467 => x"15",
          7468 => x"3f",
          7469 => x"15",
          7470 => x"3f",
          7471 => x"0b",
          7472 => x"78",
          7473 => x"3f",
          7474 => x"08",
          7475 => x"81",
          7476 => x"57",
          7477 => x"34",
          7478 => x"dc",
          7479 => x"0d",
          7480 => x"0d",
          7481 => x"54",
          7482 => x"82",
          7483 => x"53",
          7484 => x"08",
          7485 => x"3d",
          7486 => x"73",
          7487 => x"3f",
          7488 => x"08",
          7489 => x"dc",
          7490 => x"82",
          7491 => x"74",
          7492 => x"bb",
          7493 => x"3d",
          7494 => x"3d",
          7495 => x"51",
          7496 => x"8b",
          7497 => x"82",
          7498 => x"24",
          7499 => x"bb",
          7500 => x"d3",
          7501 => x"52",
          7502 => x"dc",
          7503 => x"0d",
          7504 => x"0d",
          7505 => x"3d",
          7506 => x"94",
          7507 => x"c1",
          7508 => x"dc",
          7509 => x"bb",
          7510 => x"e0",
          7511 => x"63",
          7512 => x"d4",
          7513 => x"8d",
          7514 => x"dc",
          7515 => x"bb",
          7516 => x"38",
          7517 => x"05",
          7518 => x"2b",
          7519 => x"80",
          7520 => x"76",
          7521 => x"0c",
          7522 => x"02",
          7523 => x"70",
          7524 => x"81",
          7525 => x"56",
          7526 => x"9e",
          7527 => x"53",
          7528 => x"db",
          7529 => x"bb",
          7530 => x"15",
          7531 => x"82",
          7532 => x"84",
          7533 => x"06",
          7534 => x"55",
          7535 => x"dc",
          7536 => x"0d",
          7537 => x"0d",
          7538 => x"5b",
          7539 => x"80",
          7540 => x"ff",
          7541 => x"9f",
          7542 => x"b5",
          7543 => x"dc",
          7544 => x"bb",
          7545 => x"fc",
          7546 => x"7a",
          7547 => x"08",
          7548 => x"64",
          7549 => x"2e",
          7550 => x"a0",
          7551 => x"70",
          7552 => x"ea",
          7553 => x"dc",
          7554 => x"bb",
          7555 => x"d4",
          7556 => x"7b",
          7557 => x"3f",
          7558 => x"08",
          7559 => x"dc",
          7560 => x"38",
          7561 => x"51",
          7562 => x"82",
          7563 => x"45",
          7564 => x"51",
          7565 => x"82",
          7566 => x"57",
          7567 => x"08",
          7568 => x"80",
          7569 => x"da",
          7570 => x"bb",
          7571 => x"82",
          7572 => x"a4",
          7573 => x"7b",
          7574 => x"3f",
          7575 => x"dc",
          7576 => x"38",
          7577 => x"51",
          7578 => x"82",
          7579 => x"57",
          7580 => x"08",
          7581 => x"38",
          7582 => x"09",
          7583 => x"38",
          7584 => x"e0",
          7585 => x"dc",
          7586 => x"ff",
          7587 => x"74",
          7588 => x"3f",
          7589 => x"78",
          7590 => x"33",
          7591 => x"56",
          7592 => x"91",
          7593 => x"05",
          7594 => x"81",
          7595 => x"56",
          7596 => x"f5",
          7597 => x"54",
          7598 => x"81",
          7599 => x"80",
          7600 => x"78",
          7601 => x"55",
          7602 => x"11",
          7603 => x"18",
          7604 => x"58",
          7605 => x"34",
          7606 => x"ff",
          7607 => x"55",
          7608 => x"34",
          7609 => x"77",
          7610 => x"81",
          7611 => x"ff",
          7612 => x"55",
          7613 => x"34",
          7614 => x"d3",
          7615 => x"84",
          7616 => x"94",
          7617 => x"70",
          7618 => x"56",
          7619 => x"76",
          7620 => x"81",
          7621 => x"70",
          7622 => x"56",
          7623 => x"82",
          7624 => x"78",
          7625 => x"80",
          7626 => x"27",
          7627 => x"19",
          7628 => x"7a",
          7629 => x"5c",
          7630 => x"55",
          7631 => x"7a",
          7632 => x"5c",
          7633 => x"2e",
          7634 => x"85",
          7635 => x"94",
          7636 => x"81",
          7637 => x"73",
          7638 => x"81",
          7639 => x"7a",
          7640 => x"38",
          7641 => x"76",
          7642 => x"0c",
          7643 => x"04",
          7644 => x"7b",
          7645 => x"fc",
          7646 => x"53",
          7647 => x"bb",
          7648 => x"dc",
          7649 => x"bb",
          7650 => x"fa",
          7651 => x"33",
          7652 => x"f2",
          7653 => x"08",
          7654 => x"27",
          7655 => x"15",
          7656 => x"2a",
          7657 => x"51",
          7658 => x"83",
          7659 => x"94",
          7660 => x"80",
          7661 => x"0c",
          7662 => x"2e",
          7663 => x"79",
          7664 => x"70",
          7665 => x"51",
          7666 => x"2e",
          7667 => x"52",
          7668 => x"fe",
          7669 => x"82",
          7670 => x"ff",
          7671 => x"70",
          7672 => x"fe",
          7673 => x"82",
          7674 => x"73",
          7675 => x"76",
          7676 => x"06",
          7677 => x"0c",
          7678 => x"98",
          7679 => x"58",
          7680 => x"39",
          7681 => x"54",
          7682 => x"73",
          7683 => x"cd",
          7684 => x"bb",
          7685 => x"82",
          7686 => x"81",
          7687 => x"38",
          7688 => x"08",
          7689 => x"9b",
          7690 => x"dc",
          7691 => x"0c",
          7692 => x"0c",
          7693 => x"81",
          7694 => x"76",
          7695 => x"38",
          7696 => x"94",
          7697 => x"94",
          7698 => x"16",
          7699 => x"2a",
          7700 => x"51",
          7701 => x"72",
          7702 => x"38",
          7703 => x"51",
          7704 => x"82",
          7705 => x"54",
          7706 => x"08",
          7707 => x"bb",
          7708 => x"a7",
          7709 => x"74",
          7710 => x"3f",
          7711 => x"08",
          7712 => x"2e",
          7713 => x"74",
          7714 => x"79",
          7715 => x"14",
          7716 => x"38",
          7717 => x"0c",
          7718 => x"94",
          7719 => x"94",
          7720 => x"83",
          7721 => x"72",
          7722 => x"38",
          7723 => x"51",
          7724 => x"82",
          7725 => x"94",
          7726 => x"91",
          7727 => x"53",
          7728 => x"81",
          7729 => x"34",
          7730 => x"39",
          7731 => x"82",
          7732 => x"05",
          7733 => x"08",
          7734 => x"08",
          7735 => x"38",
          7736 => x"0c",
          7737 => x"80",
          7738 => x"72",
          7739 => x"73",
          7740 => x"53",
          7741 => x"8c",
          7742 => x"16",
          7743 => x"38",
          7744 => x"0c",
          7745 => x"82",
          7746 => x"8b",
          7747 => x"f9",
          7748 => x"56",
          7749 => x"80",
          7750 => x"38",
          7751 => x"3d",
          7752 => x"8a",
          7753 => x"51",
          7754 => x"82",
          7755 => x"55",
          7756 => x"08",
          7757 => x"77",
          7758 => x"52",
          7759 => x"b5",
          7760 => x"dc",
          7761 => x"bb",
          7762 => x"c3",
          7763 => x"33",
          7764 => x"55",
          7765 => x"24",
          7766 => x"16",
          7767 => x"2a",
          7768 => x"51",
          7769 => x"80",
          7770 => x"9c",
          7771 => x"77",
          7772 => x"3f",
          7773 => x"08",
          7774 => x"77",
          7775 => x"22",
          7776 => x"74",
          7777 => x"ce",
          7778 => x"bb",
          7779 => x"74",
          7780 => x"81",
          7781 => x"85",
          7782 => x"74",
          7783 => x"38",
          7784 => x"74",
          7785 => x"bb",
          7786 => x"3d",
          7787 => x"3d",
          7788 => x"3d",
          7789 => x"70",
          7790 => x"ff",
          7791 => x"dc",
          7792 => x"82",
          7793 => x"73",
          7794 => x"0d",
          7795 => x"0d",
          7796 => x"3d",
          7797 => x"71",
          7798 => x"e7",
          7799 => x"bb",
          7800 => x"82",
          7801 => x"80",
          7802 => x"93",
          7803 => x"dc",
          7804 => x"51",
          7805 => x"82",
          7806 => x"53",
          7807 => x"82",
          7808 => x"52",
          7809 => x"ac",
          7810 => x"dc",
          7811 => x"bb",
          7812 => x"2e",
          7813 => x"85",
          7814 => x"87",
          7815 => x"dc",
          7816 => x"74",
          7817 => x"d5",
          7818 => x"52",
          7819 => x"89",
          7820 => x"dc",
          7821 => x"70",
          7822 => x"07",
          7823 => x"82",
          7824 => x"06",
          7825 => x"54",
          7826 => x"dc",
          7827 => x"0d",
          7828 => x"0d",
          7829 => x"53",
          7830 => x"53",
          7831 => x"56",
          7832 => x"82",
          7833 => x"55",
          7834 => x"08",
          7835 => x"52",
          7836 => x"81",
          7837 => x"dc",
          7838 => x"bb",
          7839 => x"38",
          7840 => x"05",
          7841 => x"2b",
          7842 => x"80",
          7843 => x"86",
          7844 => x"76",
          7845 => x"38",
          7846 => x"51",
          7847 => x"74",
          7848 => x"0c",
          7849 => x"04",
          7850 => x"63",
          7851 => x"80",
          7852 => x"ec",
          7853 => x"3d",
          7854 => x"3f",
          7855 => x"08",
          7856 => x"dc",
          7857 => x"38",
          7858 => x"73",
          7859 => x"08",
          7860 => x"13",
          7861 => x"58",
          7862 => x"26",
          7863 => x"7c",
          7864 => x"39",
          7865 => x"cc",
          7866 => x"81",
          7867 => x"bb",
          7868 => x"33",
          7869 => x"81",
          7870 => x"06",
          7871 => x"75",
          7872 => x"52",
          7873 => x"05",
          7874 => x"3f",
          7875 => x"08",
          7876 => x"38",
          7877 => x"08",
          7878 => x"38",
          7879 => x"08",
          7880 => x"bb",
          7881 => x"80",
          7882 => x"81",
          7883 => x"59",
          7884 => x"14",
          7885 => x"ca",
          7886 => x"39",
          7887 => x"82",
          7888 => x"57",
          7889 => x"38",
          7890 => x"18",
          7891 => x"ff",
          7892 => x"82",
          7893 => x"5b",
          7894 => x"08",
          7895 => x"7c",
          7896 => x"12",
          7897 => x"52",
          7898 => x"82",
          7899 => x"06",
          7900 => x"14",
          7901 => x"cb",
          7902 => x"dc",
          7903 => x"ff",
          7904 => x"70",
          7905 => x"82",
          7906 => x"51",
          7907 => x"b4",
          7908 => x"bb",
          7909 => x"bb",
          7910 => x"0a",
          7911 => x"70",
          7912 => x"84",
          7913 => x"51",
          7914 => x"ff",
          7915 => x"56",
          7916 => x"38",
          7917 => x"7c",
          7918 => x"0c",
          7919 => x"81",
          7920 => x"74",
          7921 => x"7a",
          7922 => x"0c",
          7923 => x"04",
          7924 => x"79",
          7925 => x"05",
          7926 => x"57",
          7927 => x"82",
          7928 => x"56",
          7929 => x"08",
          7930 => x"91",
          7931 => x"75",
          7932 => x"90",
          7933 => x"81",
          7934 => x"06",
          7935 => x"87",
          7936 => x"2e",
          7937 => x"94",
          7938 => x"73",
          7939 => x"27",
          7940 => x"73",
          7941 => x"bb",
          7942 => x"88",
          7943 => x"76",
          7944 => x"3f",
          7945 => x"08",
          7946 => x"0c",
          7947 => x"39",
          7948 => x"52",
          7949 => x"bf",
          7950 => x"bb",
          7951 => x"2e",
          7952 => x"83",
          7953 => x"82",
          7954 => x"81",
          7955 => x"06",
          7956 => x"56",
          7957 => x"a0",
          7958 => x"82",
          7959 => x"98",
          7960 => x"94",
          7961 => x"08",
          7962 => x"dc",
          7963 => x"51",
          7964 => x"82",
          7965 => x"56",
          7966 => x"8c",
          7967 => x"17",
          7968 => x"07",
          7969 => x"18",
          7970 => x"2e",
          7971 => x"91",
          7972 => x"55",
          7973 => x"dc",
          7974 => x"0d",
          7975 => x"0d",
          7976 => x"3d",
          7977 => x"52",
          7978 => x"da",
          7979 => x"bb",
          7980 => x"82",
          7981 => x"81",
          7982 => x"45",
          7983 => x"52",
          7984 => x"52",
          7985 => x"3f",
          7986 => x"08",
          7987 => x"dc",
          7988 => x"38",
          7989 => x"05",
          7990 => x"2a",
          7991 => x"51",
          7992 => x"55",
          7993 => x"38",
          7994 => x"54",
          7995 => x"81",
          7996 => x"80",
          7997 => x"70",
          7998 => x"54",
          7999 => x"81",
          8000 => x"52",
          8001 => x"c5",
          8002 => x"dc",
          8003 => x"2a",
          8004 => x"51",
          8005 => x"80",
          8006 => x"38",
          8007 => x"bb",
          8008 => x"15",
          8009 => x"86",
          8010 => x"82",
          8011 => x"5c",
          8012 => x"3d",
          8013 => x"c7",
          8014 => x"bb",
          8015 => x"82",
          8016 => x"80",
          8017 => x"bb",
          8018 => x"73",
          8019 => x"3f",
          8020 => x"08",
          8021 => x"dc",
          8022 => x"87",
          8023 => x"39",
          8024 => x"08",
          8025 => x"38",
          8026 => x"08",
          8027 => x"77",
          8028 => x"3f",
          8029 => x"08",
          8030 => x"08",
          8031 => x"bb",
          8032 => x"80",
          8033 => x"55",
          8034 => x"94",
          8035 => x"2e",
          8036 => x"53",
          8037 => x"51",
          8038 => x"82",
          8039 => x"55",
          8040 => x"78",
          8041 => x"fe",
          8042 => x"dc",
          8043 => x"82",
          8044 => x"a0",
          8045 => x"e9",
          8046 => x"53",
          8047 => x"05",
          8048 => x"51",
          8049 => x"82",
          8050 => x"54",
          8051 => x"08",
          8052 => x"78",
          8053 => x"8e",
          8054 => x"58",
          8055 => x"82",
          8056 => x"54",
          8057 => x"08",
          8058 => x"54",
          8059 => x"82",
          8060 => x"84",
          8061 => x"06",
          8062 => x"02",
          8063 => x"33",
          8064 => x"81",
          8065 => x"86",
          8066 => x"f6",
          8067 => x"74",
          8068 => x"70",
          8069 => x"c3",
          8070 => x"dc",
          8071 => x"56",
          8072 => x"08",
          8073 => x"54",
          8074 => x"08",
          8075 => x"81",
          8076 => x"82",
          8077 => x"dc",
          8078 => x"09",
          8079 => x"38",
          8080 => x"b4",
          8081 => x"b0",
          8082 => x"dc",
          8083 => x"51",
          8084 => x"82",
          8085 => x"54",
          8086 => x"08",
          8087 => x"8b",
          8088 => x"b4",
          8089 => x"b7",
          8090 => x"54",
          8091 => x"15",
          8092 => x"90",
          8093 => x"34",
          8094 => x"0a",
          8095 => x"19",
          8096 => x"9f",
          8097 => x"78",
          8098 => x"51",
          8099 => x"a0",
          8100 => x"11",
          8101 => x"05",
          8102 => x"b6",
          8103 => x"ae",
          8104 => x"15",
          8105 => x"78",
          8106 => x"53",
          8107 => x"3f",
          8108 => x"0b",
          8109 => x"77",
          8110 => x"3f",
          8111 => x"08",
          8112 => x"dc",
          8113 => x"82",
          8114 => x"52",
          8115 => x"51",
          8116 => x"3f",
          8117 => x"52",
          8118 => x"aa",
          8119 => x"90",
          8120 => x"34",
          8121 => x"0b",
          8122 => x"78",
          8123 => x"b6",
          8124 => x"dc",
          8125 => x"39",
          8126 => x"52",
          8127 => x"be",
          8128 => x"82",
          8129 => x"99",
          8130 => x"da",
          8131 => x"3d",
          8132 => x"d2",
          8133 => x"53",
          8134 => x"84",
          8135 => x"3d",
          8136 => x"3f",
          8137 => x"08",
          8138 => x"dc",
          8139 => x"38",
          8140 => x"3d",
          8141 => x"3d",
          8142 => x"cc",
          8143 => x"bb",
          8144 => x"82",
          8145 => x"82",
          8146 => x"81",
          8147 => x"81",
          8148 => x"86",
          8149 => x"aa",
          8150 => x"a4",
          8151 => x"a8",
          8152 => x"05",
          8153 => x"ea",
          8154 => x"77",
          8155 => x"70",
          8156 => x"b4",
          8157 => x"3d",
          8158 => x"51",
          8159 => x"82",
          8160 => x"55",
          8161 => x"08",
          8162 => x"6f",
          8163 => x"06",
          8164 => x"a2",
          8165 => x"92",
          8166 => x"81",
          8167 => x"bb",
          8168 => x"2e",
          8169 => x"81",
          8170 => x"51",
          8171 => x"82",
          8172 => x"55",
          8173 => x"08",
          8174 => x"68",
          8175 => x"a8",
          8176 => x"05",
          8177 => x"51",
          8178 => x"3f",
          8179 => x"33",
          8180 => x"8b",
          8181 => x"84",
          8182 => x"06",
          8183 => x"73",
          8184 => x"a0",
          8185 => x"8b",
          8186 => x"54",
          8187 => x"15",
          8188 => x"33",
          8189 => x"70",
          8190 => x"55",
          8191 => x"2e",
          8192 => x"6e",
          8193 => x"df",
          8194 => x"78",
          8195 => x"3f",
          8196 => x"08",
          8197 => x"ff",
          8198 => x"82",
          8199 => x"dc",
          8200 => x"80",
          8201 => x"bb",
          8202 => x"78",
          8203 => x"af",
          8204 => x"dc",
          8205 => x"d4",
          8206 => x"55",
          8207 => x"08",
          8208 => x"81",
          8209 => x"73",
          8210 => x"81",
          8211 => x"63",
          8212 => x"76",
          8213 => x"3f",
          8214 => x"0b",
          8215 => x"87",
          8216 => x"dc",
          8217 => x"77",
          8218 => x"3f",
          8219 => x"08",
          8220 => x"dc",
          8221 => x"78",
          8222 => x"aa",
          8223 => x"dc",
          8224 => x"82",
          8225 => x"a8",
          8226 => x"ed",
          8227 => x"80",
          8228 => x"02",
          8229 => x"df",
          8230 => x"57",
          8231 => x"3d",
          8232 => x"96",
          8233 => x"e9",
          8234 => x"dc",
          8235 => x"bb",
          8236 => x"cf",
          8237 => x"65",
          8238 => x"d4",
          8239 => x"b5",
          8240 => x"dc",
          8241 => x"bb",
          8242 => x"38",
          8243 => x"05",
          8244 => x"06",
          8245 => x"73",
          8246 => x"a7",
          8247 => x"09",
          8248 => x"71",
          8249 => x"06",
          8250 => x"55",
          8251 => x"15",
          8252 => x"81",
          8253 => x"34",
          8254 => x"b4",
          8255 => x"bb",
          8256 => x"74",
          8257 => x"0c",
          8258 => x"04",
          8259 => x"64",
          8260 => x"93",
          8261 => x"52",
          8262 => x"d1",
          8263 => x"bb",
          8264 => x"82",
          8265 => x"80",
          8266 => x"58",
          8267 => x"3d",
          8268 => x"c8",
          8269 => x"bb",
          8270 => x"82",
          8271 => x"b4",
          8272 => x"c7",
          8273 => x"a0",
          8274 => x"55",
          8275 => x"84",
          8276 => x"17",
          8277 => x"2b",
          8278 => x"96",
          8279 => x"b0",
          8280 => x"54",
          8281 => x"15",
          8282 => x"ff",
          8283 => x"82",
          8284 => x"55",
          8285 => x"dc",
          8286 => x"0d",
          8287 => x"0d",
          8288 => x"5a",
          8289 => x"3d",
          8290 => x"99",
          8291 => x"81",
          8292 => x"dc",
          8293 => x"dc",
          8294 => x"82",
          8295 => x"07",
          8296 => x"55",
          8297 => x"2e",
          8298 => x"81",
          8299 => x"55",
          8300 => x"2e",
          8301 => x"7b",
          8302 => x"80",
          8303 => x"70",
          8304 => x"be",
          8305 => x"bb",
          8306 => x"82",
          8307 => x"80",
          8308 => x"52",
          8309 => x"dc",
          8310 => x"dc",
          8311 => x"bb",
          8312 => x"38",
          8313 => x"08",
          8314 => x"08",
          8315 => x"56",
          8316 => x"19",
          8317 => x"59",
          8318 => x"74",
          8319 => x"56",
          8320 => x"ec",
          8321 => x"75",
          8322 => x"74",
          8323 => x"2e",
          8324 => x"16",
          8325 => x"33",
          8326 => x"73",
          8327 => x"38",
          8328 => x"84",
          8329 => x"06",
          8330 => x"7a",
          8331 => x"76",
          8332 => x"07",
          8333 => x"54",
          8334 => x"80",
          8335 => x"80",
          8336 => x"7b",
          8337 => x"53",
          8338 => x"93",
          8339 => x"dc",
          8340 => x"bb",
          8341 => x"38",
          8342 => x"55",
          8343 => x"56",
          8344 => x"8b",
          8345 => x"56",
          8346 => x"83",
          8347 => x"75",
          8348 => x"51",
          8349 => x"3f",
          8350 => x"08",
          8351 => x"82",
          8352 => x"98",
          8353 => x"e6",
          8354 => x"53",
          8355 => x"b8",
          8356 => x"3d",
          8357 => x"3f",
          8358 => x"08",
          8359 => x"08",
          8360 => x"bb",
          8361 => x"98",
          8362 => x"a0",
          8363 => x"70",
          8364 => x"ae",
          8365 => x"6d",
          8366 => x"81",
          8367 => x"57",
          8368 => x"74",
          8369 => x"38",
          8370 => x"81",
          8371 => x"81",
          8372 => x"52",
          8373 => x"89",
          8374 => x"dc",
          8375 => x"a5",
          8376 => x"33",
          8377 => x"54",
          8378 => x"3f",
          8379 => x"08",
          8380 => x"38",
          8381 => x"76",
          8382 => x"05",
          8383 => x"39",
          8384 => x"08",
          8385 => x"15",
          8386 => x"ff",
          8387 => x"73",
          8388 => x"38",
          8389 => x"83",
          8390 => x"56",
          8391 => x"75",
          8392 => x"82",
          8393 => x"33",
          8394 => x"2e",
          8395 => x"52",
          8396 => x"51",
          8397 => x"3f",
          8398 => x"08",
          8399 => x"ff",
          8400 => x"38",
          8401 => x"88",
          8402 => x"8a",
          8403 => x"38",
          8404 => x"ec",
          8405 => x"75",
          8406 => x"74",
          8407 => x"73",
          8408 => x"05",
          8409 => x"17",
          8410 => x"70",
          8411 => x"34",
          8412 => x"70",
          8413 => x"ff",
          8414 => x"55",
          8415 => x"26",
          8416 => x"8b",
          8417 => x"86",
          8418 => x"e5",
          8419 => x"38",
          8420 => x"99",
          8421 => x"05",
          8422 => x"70",
          8423 => x"73",
          8424 => x"81",
          8425 => x"ff",
          8426 => x"ed",
          8427 => x"80",
          8428 => x"91",
          8429 => x"55",
          8430 => x"3f",
          8431 => x"08",
          8432 => x"dc",
          8433 => x"38",
          8434 => x"51",
          8435 => x"3f",
          8436 => x"08",
          8437 => x"dc",
          8438 => x"76",
          8439 => x"67",
          8440 => x"34",
          8441 => x"82",
          8442 => x"84",
          8443 => x"06",
          8444 => x"80",
          8445 => x"2e",
          8446 => x"81",
          8447 => x"ff",
          8448 => x"82",
          8449 => x"54",
          8450 => x"08",
          8451 => x"53",
          8452 => x"08",
          8453 => x"ff",
          8454 => x"67",
          8455 => x"8b",
          8456 => x"53",
          8457 => x"51",
          8458 => x"3f",
          8459 => x"0b",
          8460 => x"79",
          8461 => x"ee",
          8462 => x"dc",
          8463 => x"55",
          8464 => x"dc",
          8465 => x"0d",
          8466 => x"0d",
          8467 => x"88",
          8468 => x"05",
          8469 => x"fc",
          8470 => x"54",
          8471 => x"d2",
          8472 => x"bb",
          8473 => x"82",
          8474 => x"82",
          8475 => x"1a",
          8476 => x"82",
          8477 => x"80",
          8478 => x"8c",
          8479 => x"78",
          8480 => x"1a",
          8481 => x"2a",
          8482 => x"51",
          8483 => x"90",
          8484 => x"82",
          8485 => x"58",
          8486 => x"81",
          8487 => x"39",
          8488 => x"22",
          8489 => x"70",
          8490 => x"56",
          8491 => x"bd",
          8492 => x"14",
          8493 => x"30",
          8494 => x"9f",
          8495 => x"dc",
          8496 => x"19",
          8497 => x"5a",
          8498 => x"81",
          8499 => x"38",
          8500 => x"77",
          8501 => x"82",
          8502 => x"56",
          8503 => x"74",
          8504 => x"ff",
          8505 => x"81",
          8506 => x"55",
          8507 => x"75",
          8508 => x"82",
          8509 => x"dc",
          8510 => x"ff",
          8511 => x"bb",
          8512 => x"2e",
          8513 => x"82",
          8514 => x"8e",
          8515 => x"56",
          8516 => x"09",
          8517 => x"38",
          8518 => x"59",
          8519 => x"77",
          8520 => x"06",
          8521 => x"87",
          8522 => x"39",
          8523 => x"ba",
          8524 => x"55",
          8525 => x"2e",
          8526 => x"15",
          8527 => x"2e",
          8528 => x"83",
          8529 => x"75",
          8530 => x"7e",
          8531 => x"a8",
          8532 => x"dc",
          8533 => x"bb",
          8534 => x"ce",
          8535 => x"16",
          8536 => x"56",
          8537 => x"38",
          8538 => x"19",
          8539 => x"8c",
          8540 => x"7d",
          8541 => x"38",
          8542 => x"0c",
          8543 => x"0c",
          8544 => x"80",
          8545 => x"73",
          8546 => x"98",
          8547 => x"05",
          8548 => x"57",
          8549 => x"26",
          8550 => x"7b",
          8551 => x"0c",
          8552 => x"81",
          8553 => x"84",
          8554 => x"54",
          8555 => x"dc",
          8556 => x"0d",
          8557 => x"0d",
          8558 => x"88",
          8559 => x"05",
          8560 => x"54",
          8561 => x"c5",
          8562 => x"56",
          8563 => x"bb",
          8564 => x"8b",
          8565 => x"bb",
          8566 => x"29",
          8567 => x"05",
          8568 => x"55",
          8569 => x"84",
          8570 => x"34",
          8571 => x"08",
          8572 => x"5f",
          8573 => x"51",
          8574 => x"3f",
          8575 => x"08",
          8576 => x"70",
          8577 => x"57",
          8578 => x"8b",
          8579 => x"82",
          8580 => x"06",
          8581 => x"56",
          8582 => x"38",
          8583 => x"05",
          8584 => x"7e",
          8585 => x"f0",
          8586 => x"dc",
          8587 => x"67",
          8588 => x"2e",
          8589 => x"82",
          8590 => x"8b",
          8591 => x"75",
          8592 => x"80",
          8593 => x"81",
          8594 => x"2e",
          8595 => x"80",
          8596 => x"38",
          8597 => x"0a",
          8598 => x"ff",
          8599 => x"55",
          8600 => x"86",
          8601 => x"8a",
          8602 => x"89",
          8603 => x"2a",
          8604 => x"77",
          8605 => x"59",
          8606 => x"81",
          8607 => x"70",
          8608 => x"07",
          8609 => x"56",
          8610 => x"38",
          8611 => x"05",
          8612 => x"7e",
          8613 => x"80",
          8614 => x"82",
          8615 => x"8a",
          8616 => x"83",
          8617 => x"06",
          8618 => x"08",
          8619 => x"74",
          8620 => x"41",
          8621 => x"56",
          8622 => x"8a",
          8623 => x"61",
          8624 => x"55",
          8625 => x"27",
          8626 => x"93",
          8627 => x"80",
          8628 => x"38",
          8629 => x"70",
          8630 => x"43",
          8631 => x"95",
          8632 => x"06",
          8633 => x"2e",
          8634 => x"77",
          8635 => x"74",
          8636 => x"83",
          8637 => x"06",
          8638 => x"82",
          8639 => x"2e",
          8640 => x"78",
          8641 => x"2e",
          8642 => x"80",
          8643 => x"ae",
          8644 => x"2a",
          8645 => x"82",
          8646 => x"56",
          8647 => x"2e",
          8648 => x"77",
          8649 => x"82",
          8650 => x"79",
          8651 => x"70",
          8652 => x"5a",
          8653 => x"86",
          8654 => x"27",
          8655 => x"52",
          8656 => x"b8",
          8657 => x"bb",
          8658 => x"29",
          8659 => x"70",
          8660 => x"55",
          8661 => x"0b",
          8662 => x"08",
          8663 => x"05",
          8664 => x"ff",
          8665 => x"27",
          8666 => x"88",
          8667 => x"ae",
          8668 => x"2a",
          8669 => x"82",
          8670 => x"56",
          8671 => x"2e",
          8672 => x"77",
          8673 => x"82",
          8674 => x"79",
          8675 => x"70",
          8676 => x"5a",
          8677 => x"86",
          8678 => x"27",
          8679 => x"52",
          8680 => x"b7",
          8681 => x"bb",
          8682 => x"84",
          8683 => x"bb",
          8684 => x"f5",
          8685 => x"81",
          8686 => x"dc",
          8687 => x"bb",
          8688 => x"71",
          8689 => x"83",
          8690 => x"5e",
          8691 => x"89",
          8692 => x"5c",
          8693 => x"1c",
          8694 => x"05",
          8695 => x"ff",
          8696 => x"70",
          8697 => x"31",
          8698 => x"57",
          8699 => x"83",
          8700 => x"06",
          8701 => x"1c",
          8702 => x"5c",
          8703 => x"1d",
          8704 => x"29",
          8705 => x"31",
          8706 => x"55",
          8707 => x"87",
          8708 => x"7c",
          8709 => x"7a",
          8710 => x"31",
          8711 => x"b6",
          8712 => x"bb",
          8713 => x"7d",
          8714 => x"81",
          8715 => x"82",
          8716 => x"83",
          8717 => x"80",
          8718 => x"87",
          8719 => x"81",
          8720 => x"fd",
          8721 => x"f8",
          8722 => x"2e",
          8723 => x"80",
          8724 => x"ff",
          8725 => x"bb",
          8726 => x"a0",
          8727 => x"38",
          8728 => x"74",
          8729 => x"86",
          8730 => x"fd",
          8731 => x"81",
          8732 => x"80",
          8733 => x"83",
          8734 => x"39",
          8735 => x"08",
          8736 => x"92",
          8737 => x"b8",
          8738 => x"59",
          8739 => x"27",
          8740 => x"86",
          8741 => x"55",
          8742 => x"09",
          8743 => x"38",
          8744 => x"f5",
          8745 => x"38",
          8746 => x"55",
          8747 => x"86",
          8748 => x"80",
          8749 => x"7a",
          8750 => x"b9",
          8751 => x"82",
          8752 => x"7a",
          8753 => x"8a",
          8754 => x"52",
          8755 => x"ff",
          8756 => x"79",
          8757 => x"7b",
          8758 => x"06",
          8759 => x"51",
          8760 => x"3f",
          8761 => x"1c",
          8762 => x"32",
          8763 => x"96",
          8764 => x"06",
          8765 => x"91",
          8766 => x"a1",
          8767 => x"55",
          8768 => x"ff",
          8769 => x"74",
          8770 => x"06",
          8771 => x"51",
          8772 => x"3f",
          8773 => x"52",
          8774 => x"ff",
          8775 => x"f8",
          8776 => x"34",
          8777 => x"1b",
          8778 => x"d9",
          8779 => x"52",
          8780 => x"ff",
          8781 => x"60",
          8782 => x"51",
          8783 => x"3f",
          8784 => x"09",
          8785 => x"cb",
          8786 => x"b2",
          8787 => x"c3",
          8788 => x"a0",
          8789 => x"52",
          8790 => x"ff",
          8791 => x"82",
          8792 => x"51",
          8793 => x"3f",
          8794 => x"1b",
          8795 => x"95",
          8796 => x"b2",
          8797 => x"a0",
          8798 => x"80",
          8799 => x"1c",
          8800 => x"80",
          8801 => x"93",
          8802 => x"ec",
          8803 => x"1b",
          8804 => x"82",
          8805 => x"52",
          8806 => x"ff",
          8807 => x"7c",
          8808 => x"06",
          8809 => x"51",
          8810 => x"3f",
          8811 => x"a4",
          8812 => x"0b",
          8813 => x"93",
          8814 => x"80",
          8815 => x"51",
          8816 => x"3f",
          8817 => x"52",
          8818 => x"70",
          8819 => x"9f",
          8820 => x"54",
          8821 => x"52",
          8822 => x"9b",
          8823 => x"56",
          8824 => x"08",
          8825 => x"7d",
          8826 => x"81",
          8827 => x"38",
          8828 => x"86",
          8829 => x"52",
          8830 => x"9b",
          8831 => x"80",
          8832 => x"7a",
          8833 => x"ed",
          8834 => x"85",
          8835 => x"7a",
          8836 => x"8f",
          8837 => x"85",
          8838 => x"83",
          8839 => x"ff",
          8840 => x"ff",
          8841 => x"e8",
          8842 => x"9e",
          8843 => x"52",
          8844 => x"51",
          8845 => x"3f",
          8846 => x"52",
          8847 => x"9e",
          8848 => x"54",
          8849 => x"53",
          8850 => x"51",
          8851 => x"3f",
          8852 => x"16",
          8853 => x"7e",
          8854 => x"d8",
          8855 => x"80",
          8856 => x"ff",
          8857 => x"7f",
          8858 => x"7d",
          8859 => x"81",
          8860 => x"f8",
          8861 => x"ff",
          8862 => x"ff",
          8863 => x"51",
          8864 => x"3f",
          8865 => x"88",
          8866 => x"39",
          8867 => x"f8",
          8868 => x"2e",
          8869 => x"55",
          8870 => x"51",
          8871 => x"3f",
          8872 => x"57",
          8873 => x"83",
          8874 => x"76",
          8875 => x"7a",
          8876 => x"ff",
          8877 => x"82",
          8878 => x"82",
          8879 => x"80",
          8880 => x"dc",
          8881 => x"51",
          8882 => x"3f",
          8883 => x"78",
          8884 => x"74",
          8885 => x"18",
          8886 => x"2e",
          8887 => x"79",
          8888 => x"2e",
          8889 => x"55",
          8890 => x"62",
          8891 => x"74",
          8892 => x"75",
          8893 => x"7e",
          8894 => x"b8",
          8895 => x"dc",
          8896 => x"38",
          8897 => x"78",
          8898 => x"74",
          8899 => x"56",
          8900 => x"93",
          8901 => x"66",
          8902 => x"26",
          8903 => x"56",
          8904 => x"83",
          8905 => x"64",
          8906 => x"77",
          8907 => x"84",
          8908 => x"52",
          8909 => x"9d",
          8910 => x"d4",
          8911 => x"51",
          8912 => x"3f",
          8913 => x"55",
          8914 => x"81",
          8915 => x"34",
          8916 => x"16",
          8917 => x"16",
          8918 => x"16",
          8919 => x"05",
          8920 => x"c1",
          8921 => x"fe",
          8922 => x"fe",
          8923 => x"34",
          8924 => x"08",
          8925 => x"07",
          8926 => x"16",
          8927 => x"dc",
          8928 => x"34",
          8929 => x"c6",
          8930 => x"9c",
          8931 => x"52",
          8932 => x"51",
          8933 => x"3f",
          8934 => x"53",
          8935 => x"51",
          8936 => x"3f",
          8937 => x"bb",
          8938 => x"38",
          8939 => x"52",
          8940 => x"99",
          8941 => x"56",
          8942 => x"08",
          8943 => x"39",
          8944 => x"39",
          8945 => x"39",
          8946 => x"08",
          8947 => x"bb",
          8948 => x"3d",
          8949 => x"3d",
          8950 => x"5b",
          8951 => x"60",
          8952 => x"57",
          8953 => x"25",
          8954 => x"3d",
          8955 => x"55",
          8956 => x"15",
          8957 => x"c9",
          8958 => x"81",
          8959 => x"06",
          8960 => x"3d",
          8961 => x"8d",
          8962 => x"74",
          8963 => x"05",
          8964 => x"17",
          8965 => x"2e",
          8966 => x"c9",
          8967 => x"34",
          8968 => x"83",
          8969 => x"74",
          8970 => x"0c",
          8971 => x"04",
          8972 => x"7b",
          8973 => x"b3",
          8974 => x"57",
          8975 => x"09",
          8976 => x"38",
          8977 => x"51",
          8978 => x"17",
          8979 => x"76",
          8980 => x"88",
          8981 => x"17",
          8982 => x"59",
          8983 => x"81",
          8984 => x"76",
          8985 => x"8b",
          8986 => x"54",
          8987 => x"17",
          8988 => x"51",
          8989 => x"79",
          8990 => x"30",
          8991 => x"9f",
          8992 => x"53",
          8993 => x"75",
          8994 => x"81",
          8995 => x"0c",
          8996 => x"04",
          8997 => x"79",
          8998 => x"56",
          8999 => x"24",
          9000 => x"3d",
          9001 => x"74",
          9002 => x"52",
          9003 => x"cb",
          9004 => x"bb",
          9005 => x"38",
          9006 => x"78",
          9007 => x"06",
          9008 => x"16",
          9009 => x"39",
          9010 => x"82",
          9011 => x"89",
          9012 => x"fd",
          9013 => x"54",
          9014 => x"80",
          9015 => x"ff",
          9016 => x"76",
          9017 => x"3d",
          9018 => x"3d",
          9019 => x"e3",
          9020 => x"53",
          9021 => x"53",
          9022 => x"3f",
          9023 => x"51",
          9024 => x"72",
          9025 => x"3f",
          9026 => x"04",
          9027 => x"ff",
          9028 => x"ff",
          9029 => x"ff",
          9030 => x"00",
          9031 => x"aa",
          9032 => x"2e",
          9033 => x"35",
          9034 => x"3c",
          9035 => x"43",
          9036 => x"4a",
          9037 => x"51",
          9038 => x"58",
          9039 => x"5f",
          9040 => x"66",
          9041 => x"6d",
          9042 => x"74",
          9043 => x"7a",
          9044 => x"80",
          9045 => x"86",
          9046 => x"8c",
          9047 => x"92",
          9048 => x"98",
          9049 => x"9e",
          9050 => x"a4",
          9051 => x"82",
          9052 => x"88",
          9053 => x"8e",
          9054 => x"94",
          9055 => x"9a",
          9056 => x"b9",
          9057 => x"b9",
          9058 => x"ca",
          9059 => x"22",
          9060 => x"a1",
          9061 => x"8e",
          9062 => x"92",
          9063 => x"f3",
          9064 => x"d5",
          9065 => x"6b",
          9066 => x"f1",
          9067 => x"74",
          9068 => x"8e",
          9069 => x"ca",
          9070 => x"f3",
          9071 => x"92",
          9072 => x"8e",
          9073 => x"8e",
          9074 => x"f1",
          9075 => x"6b",
          9076 => x"f3",
          9077 => x"22",
          9078 => x"31",
          9079 => x"1a",
          9080 => x"1a",
          9081 => x"60",
          9082 => x"1a",
          9083 => x"1a",
          9084 => x"1a",
          9085 => x"1a",
          9086 => x"1a",
          9087 => x"1a",
          9088 => x"1a",
          9089 => x"1d",
          9090 => x"1a",
          9091 => x"48",
          9092 => x"78",
          9093 => x"1a",
          9094 => x"1a",
          9095 => x"1a",
          9096 => x"1a",
          9097 => x"1a",
          9098 => x"1a",
          9099 => x"1a",
          9100 => x"1a",
          9101 => x"1a",
          9102 => x"1a",
          9103 => x"1a",
          9104 => x"1a",
          9105 => x"1a",
          9106 => x"1a",
          9107 => x"1a",
          9108 => x"1a",
          9109 => x"1a",
          9110 => x"1a",
          9111 => x"1a",
          9112 => x"1a",
          9113 => x"1a",
          9114 => x"1a",
          9115 => x"1a",
          9116 => x"1a",
          9117 => x"1a",
          9118 => x"1a",
          9119 => x"1a",
          9120 => x"1a",
          9121 => x"1a",
          9122 => x"1a",
          9123 => x"1a",
          9124 => x"1a",
          9125 => x"1a",
          9126 => x"1a",
          9127 => x"1a",
          9128 => x"1a",
          9129 => x"a8",
          9130 => x"1a",
          9131 => x"1a",
          9132 => x"1a",
          9133 => x"1a",
          9134 => x"16",
          9135 => x"1a",
          9136 => x"1a",
          9137 => x"1a",
          9138 => x"1a",
          9139 => x"1a",
          9140 => x"1a",
          9141 => x"1a",
          9142 => x"1a",
          9143 => x"1a",
          9144 => x"1a",
          9145 => x"d8",
          9146 => x"3f",
          9147 => x"af",
          9148 => x"af",
          9149 => x"af",
          9150 => x"1a",
          9151 => x"3f",
          9152 => x"1a",
          9153 => x"1a",
          9154 => x"98",
          9155 => x"1a",
          9156 => x"1a",
          9157 => x"ec",
          9158 => x"f7",
          9159 => x"1a",
          9160 => x"1a",
          9161 => x"11",
          9162 => x"1a",
          9163 => x"1f",
          9164 => x"1a",
          9165 => x"1a",
          9166 => x"16",
          9167 => x"69",
          9168 => x"00",
          9169 => x"63",
          9170 => x"00",
          9171 => x"69",
          9172 => x"00",
          9173 => x"61",
          9174 => x"00",
          9175 => x"65",
          9176 => x"00",
          9177 => x"65",
          9178 => x"00",
          9179 => x"70",
          9180 => x"00",
          9181 => x"66",
          9182 => x"00",
          9183 => x"6d",
          9184 => x"00",
          9185 => x"00",
          9186 => x"00",
          9187 => x"00",
          9188 => x"00",
          9189 => x"00",
          9190 => x"00",
          9191 => x"00",
          9192 => x"6c",
          9193 => x"00",
          9194 => x"00",
          9195 => x"74",
          9196 => x"00",
          9197 => x"65",
          9198 => x"00",
          9199 => x"6f",
          9200 => x"00",
          9201 => x"74",
          9202 => x"00",
          9203 => x"73",
          9204 => x"00",
          9205 => x"73",
          9206 => x"00",
          9207 => x"6f",
          9208 => x"00",
          9209 => x"00",
          9210 => x"6b",
          9211 => x"72",
          9212 => x"00",
          9213 => x"65",
          9214 => x"6c",
          9215 => x"72",
          9216 => x"00",
          9217 => x"6b",
          9218 => x"74",
          9219 => x"61",
          9220 => x"00",
          9221 => x"66",
          9222 => x"20",
          9223 => x"6e",
          9224 => x"00",
          9225 => x"70",
          9226 => x"20",
          9227 => x"6e",
          9228 => x"00",
          9229 => x"61",
          9230 => x"20",
          9231 => x"65",
          9232 => x"65",
          9233 => x"00",
          9234 => x"65",
          9235 => x"64",
          9236 => x"65",
          9237 => x"00",
          9238 => x"65",
          9239 => x"72",
          9240 => x"79",
          9241 => x"69",
          9242 => x"2e",
          9243 => x"00",
          9244 => x"65",
          9245 => x"6e",
          9246 => x"20",
          9247 => x"61",
          9248 => x"2e",
          9249 => x"00",
          9250 => x"69",
          9251 => x"72",
          9252 => x"20",
          9253 => x"74",
          9254 => x"65",
          9255 => x"00",
          9256 => x"76",
          9257 => x"75",
          9258 => x"72",
          9259 => x"20",
          9260 => x"61",
          9261 => x"2e",
          9262 => x"00",
          9263 => x"6b",
          9264 => x"74",
          9265 => x"61",
          9266 => x"64",
          9267 => x"00",
          9268 => x"63",
          9269 => x"61",
          9270 => x"6c",
          9271 => x"69",
          9272 => x"79",
          9273 => x"6d",
          9274 => x"75",
          9275 => x"6f",
          9276 => x"69",
          9277 => x"00",
          9278 => x"6d",
          9279 => x"61",
          9280 => x"74",
          9281 => x"00",
          9282 => x"65",
          9283 => x"2c",
          9284 => x"65",
          9285 => x"69",
          9286 => x"63",
          9287 => x"65",
          9288 => x"64",
          9289 => x"00",
          9290 => x"65",
          9291 => x"20",
          9292 => x"6b",
          9293 => x"00",
          9294 => x"75",
          9295 => x"63",
          9296 => x"74",
          9297 => x"6d",
          9298 => x"2e",
          9299 => x"00",
          9300 => x"20",
          9301 => x"79",
          9302 => x"65",
          9303 => x"69",
          9304 => x"2e",
          9305 => x"00",
          9306 => x"61",
          9307 => x"65",
          9308 => x"69",
          9309 => x"72",
          9310 => x"74",
          9311 => x"00",
          9312 => x"63",
          9313 => x"2e",
          9314 => x"00",
          9315 => x"6e",
          9316 => x"20",
          9317 => x"6f",
          9318 => x"00",
          9319 => x"75",
          9320 => x"74",
          9321 => x"25",
          9322 => x"74",
          9323 => x"75",
          9324 => x"74",
          9325 => x"73",
          9326 => x"0a",
          9327 => x"00",
          9328 => x"64",
          9329 => x"00",
          9330 => x"6c",
          9331 => x"00",
          9332 => x"00",
          9333 => x"58",
          9334 => x"00",
          9335 => x"20",
          9336 => x"20",
          9337 => x"00",
          9338 => x"58",
          9339 => x"00",
          9340 => x"00",
          9341 => x"00",
          9342 => x"00",
          9343 => x"54",
          9344 => x"00",
          9345 => x"20",
          9346 => x"28",
          9347 => x"00",
          9348 => x"30",
          9349 => x"30",
          9350 => x"00",
          9351 => x"35",
          9352 => x"00",
          9353 => x"55",
          9354 => x"65",
          9355 => x"30",
          9356 => x"20",
          9357 => x"25",
          9358 => x"2a",
          9359 => x"00",
          9360 => x"54",
          9361 => x"6e",
          9362 => x"72",
          9363 => x"20",
          9364 => x"64",
          9365 => x"00",
          9366 => x"65",
          9367 => x"6e",
          9368 => x"72",
          9369 => x"00",
          9370 => x"20",
          9371 => x"65",
          9372 => x"70",
          9373 => x"00",
          9374 => x"54",
          9375 => x"44",
          9376 => x"74",
          9377 => x"75",
          9378 => x"00",
          9379 => x"54",
          9380 => x"52",
          9381 => x"74",
          9382 => x"75",
          9383 => x"00",
          9384 => x"54",
          9385 => x"58",
          9386 => x"74",
          9387 => x"75",
          9388 => x"00",
          9389 => x"54",
          9390 => x"58",
          9391 => x"74",
          9392 => x"75",
          9393 => x"00",
          9394 => x"54",
          9395 => x"58",
          9396 => x"74",
          9397 => x"75",
          9398 => x"00",
          9399 => x"54",
          9400 => x"58",
          9401 => x"74",
          9402 => x"75",
          9403 => x"00",
          9404 => x"74",
          9405 => x"20",
          9406 => x"74",
          9407 => x"72",
          9408 => x"00",
          9409 => x"62",
          9410 => x"67",
          9411 => x"6d",
          9412 => x"2e",
          9413 => x"00",
          9414 => x"6f",
          9415 => x"63",
          9416 => x"74",
          9417 => x"00",
          9418 => x"74",
          9419 => x"73",
          9420 => x"00",
          9421 => x"00",
          9422 => x"6c",
          9423 => x"74",
          9424 => x"6e",
          9425 => x"61",
          9426 => x"65",
          9427 => x"20",
          9428 => x"64",
          9429 => x"20",
          9430 => x"61",
          9431 => x"69",
          9432 => x"20",
          9433 => x"75",
          9434 => x"79",
          9435 => x"00",
          9436 => x"00",
          9437 => x"20",
          9438 => x"6b",
          9439 => x"21",
          9440 => x"00",
          9441 => x"74",
          9442 => x"69",
          9443 => x"2e",
          9444 => x"00",
          9445 => x"6c",
          9446 => x"74",
          9447 => x"6e",
          9448 => x"61",
          9449 => x"65",
          9450 => x"00",
          9451 => x"25",
          9452 => x"00",
          9453 => x"00",
          9454 => x"61",
          9455 => x"67",
          9456 => x"2e",
          9457 => x"00",
          9458 => x"79",
          9459 => x"2e",
          9460 => x"00",
          9461 => x"70",
          9462 => x"6e",
          9463 => x"2e",
          9464 => x"00",
          9465 => x"6c",
          9466 => x"30",
          9467 => x"2d",
          9468 => x"38",
          9469 => x"25",
          9470 => x"29",
          9471 => x"00",
          9472 => x"70",
          9473 => x"6d",
          9474 => x"00",
          9475 => x"6d",
          9476 => x"74",
          9477 => x"00",
          9478 => x"6c",
          9479 => x"30",
          9480 => x"00",
          9481 => x"00",
          9482 => x"6c",
          9483 => x"30",
          9484 => x"00",
          9485 => x"6c",
          9486 => x"30",
          9487 => x"2d",
          9488 => x"00",
          9489 => x"61",
          9490 => x"6e",
          9491 => x"6e",
          9492 => x"72",
          9493 => x"73",
          9494 => x"00",
          9495 => x"62",
          9496 => x"67",
          9497 => x"74",
          9498 => x"75",
          9499 => x"00",
          9500 => x"61",
          9501 => x"64",
          9502 => x"72",
          9503 => x"69",
          9504 => x"00",
          9505 => x"62",
          9506 => x"67",
          9507 => x"72",
          9508 => x"69",
          9509 => x"00",
          9510 => x"63",
          9511 => x"6e",
          9512 => x"6f",
          9513 => x"40",
          9514 => x"38",
          9515 => x"2e",
          9516 => x"00",
          9517 => x"6c",
          9518 => x"20",
          9519 => x"65",
          9520 => x"25",
          9521 => x"78",
          9522 => x"2e",
          9523 => x"00",
          9524 => x"6c",
          9525 => x"74",
          9526 => x"65",
          9527 => x"6f",
          9528 => x"28",
          9529 => x"2e",
          9530 => x"00",
          9531 => x"74",
          9532 => x"69",
          9533 => x"61",
          9534 => x"69",
          9535 => x"69",
          9536 => x"2e",
          9537 => x"00",
          9538 => x"64",
          9539 => x"62",
          9540 => x"69",
          9541 => x"2e",
          9542 => x"00",
          9543 => x"00",
          9544 => x"00",
          9545 => x"5c",
          9546 => x"25",
          9547 => x"73",
          9548 => x"00",
          9549 => x"5c",
          9550 => x"25",
          9551 => x"00",
          9552 => x"5c",
          9553 => x"00",
          9554 => x"20",
          9555 => x"6d",
          9556 => x"2e",
          9557 => x"00",
          9558 => x"6e",
          9559 => x"2e",
          9560 => x"00",
          9561 => x"62",
          9562 => x"67",
          9563 => x"74",
          9564 => x"75",
          9565 => x"2e",
          9566 => x"00",
          9567 => x"25",
          9568 => x"64",
          9569 => x"3a",
          9570 => x"25",
          9571 => x"64",
          9572 => x"00",
          9573 => x"20",
          9574 => x"66",
          9575 => x"72",
          9576 => x"6f",
          9577 => x"00",
          9578 => x"72",
          9579 => x"53",
          9580 => x"63",
          9581 => x"69",
          9582 => x"00",
          9583 => x"65",
          9584 => x"65",
          9585 => x"6d",
          9586 => x"6d",
          9587 => x"65",
          9588 => x"00",
          9589 => x"20",
          9590 => x"53",
          9591 => x"4d",
          9592 => x"25",
          9593 => x"3a",
          9594 => x"58",
          9595 => x"00",
          9596 => x"20",
          9597 => x"41",
          9598 => x"20",
          9599 => x"25",
          9600 => x"3a",
          9601 => x"58",
          9602 => x"00",
          9603 => x"20",
          9604 => x"4e",
          9605 => x"41",
          9606 => x"25",
          9607 => x"3a",
          9608 => x"58",
          9609 => x"00",
          9610 => x"20",
          9611 => x"4d",
          9612 => x"20",
          9613 => x"25",
          9614 => x"3a",
          9615 => x"58",
          9616 => x"00",
          9617 => x"20",
          9618 => x"20",
          9619 => x"20",
          9620 => x"25",
          9621 => x"3a",
          9622 => x"58",
          9623 => x"00",
          9624 => x"20",
          9625 => x"43",
          9626 => x"20",
          9627 => x"44",
          9628 => x"63",
          9629 => x"3d",
          9630 => x"64",
          9631 => x"00",
          9632 => x"20",
          9633 => x"45",
          9634 => x"20",
          9635 => x"54",
          9636 => x"72",
          9637 => x"3d",
          9638 => x"64",
          9639 => x"00",
          9640 => x"20",
          9641 => x"52",
          9642 => x"52",
          9643 => x"43",
          9644 => x"6e",
          9645 => x"3d",
          9646 => x"64",
          9647 => x"00",
          9648 => x"20",
          9649 => x"48",
          9650 => x"45",
          9651 => x"53",
          9652 => x"00",
          9653 => x"20",
          9654 => x"49",
          9655 => x"00",
          9656 => x"20",
          9657 => x"54",
          9658 => x"00",
          9659 => x"20",
          9660 => x"0a",
          9661 => x"00",
          9662 => x"20",
          9663 => x"0a",
          9664 => x"00",
          9665 => x"72",
          9666 => x"65",
          9667 => x"00",
          9668 => x"20",
          9669 => x"20",
          9670 => x"65",
          9671 => x"65",
          9672 => x"72",
          9673 => x"64",
          9674 => x"73",
          9675 => x"25",
          9676 => x"0a",
          9677 => x"00",
          9678 => x"20",
          9679 => x"20",
          9680 => x"6f",
          9681 => x"53",
          9682 => x"74",
          9683 => x"64",
          9684 => x"73",
          9685 => x"25",
          9686 => x"0a",
          9687 => x"00",
          9688 => x"20",
          9689 => x"63",
          9690 => x"74",
          9691 => x"20",
          9692 => x"72",
          9693 => x"20",
          9694 => x"20",
          9695 => x"25",
          9696 => x"0a",
          9697 => x"00",
          9698 => x"63",
          9699 => x"00",
          9700 => x"20",
          9701 => x"20",
          9702 => x"20",
          9703 => x"20",
          9704 => x"20",
          9705 => x"20",
          9706 => x"20",
          9707 => x"25",
          9708 => x"0a",
          9709 => x"00",
          9710 => x"20",
          9711 => x"74",
          9712 => x"43",
          9713 => x"6b",
          9714 => x"65",
          9715 => x"20",
          9716 => x"20",
          9717 => x"25",
          9718 => x"30",
          9719 => x"48",
          9720 => x"00",
          9721 => x"20",
          9722 => x"41",
          9723 => x"6c",
          9724 => x"20",
          9725 => x"71",
          9726 => x"20",
          9727 => x"20",
          9728 => x"25",
          9729 => x"30",
          9730 => x"48",
          9731 => x"00",
          9732 => x"20",
          9733 => x"68",
          9734 => x"65",
          9735 => x"52",
          9736 => x"43",
          9737 => x"6b",
          9738 => x"65",
          9739 => x"25",
          9740 => x"30",
          9741 => x"48",
          9742 => x"00",
          9743 => x"6c",
          9744 => x"00",
          9745 => x"69",
          9746 => x"00",
          9747 => x"78",
          9748 => x"00",
          9749 => x"00",
          9750 => x"6d",
          9751 => x"00",
          9752 => x"6e",
          9753 => x"00",
          9754 => x"c4",
          9755 => x"00",
          9756 => x"02",
          9757 => x"c0",
          9758 => x"00",
          9759 => x"03",
          9760 => x"bc",
          9761 => x"00",
          9762 => x"04",
          9763 => x"b8",
          9764 => x"00",
          9765 => x"05",
          9766 => x"b4",
          9767 => x"00",
          9768 => x"06",
          9769 => x"b0",
          9770 => x"00",
          9771 => x"07",
          9772 => x"ac",
          9773 => x"00",
          9774 => x"01",
          9775 => x"a8",
          9776 => x"00",
          9777 => x"08",
          9778 => x"a4",
          9779 => x"00",
          9780 => x"0b",
          9781 => x"a0",
          9782 => x"00",
          9783 => x"09",
          9784 => x"9c",
          9785 => x"00",
          9786 => x"0a",
          9787 => x"98",
          9788 => x"00",
          9789 => x"0d",
          9790 => x"94",
          9791 => x"00",
          9792 => x"0c",
          9793 => x"90",
          9794 => x"00",
          9795 => x"0e",
          9796 => x"8c",
          9797 => x"00",
          9798 => x"0f",
          9799 => x"88",
          9800 => x"00",
          9801 => x"0f",
          9802 => x"84",
          9803 => x"00",
          9804 => x"10",
          9805 => x"80",
          9806 => x"00",
          9807 => x"11",
          9808 => x"7c",
          9809 => x"00",
          9810 => x"12",
          9811 => x"78",
          9812 => x"00",
          9813 => x"13",
          9814 => x"74",
          9815 => x"00",
          9816 => x"14",
          9817 => x"70",
          9818 => x"00",
          9819 => x"15",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"00",
          9824 => x"7e",
          9825 => x"7e",
          9826 => x"7e",
          9827 => x"00",
          9828 => x"7e",
          9829 => x"7e",
          9830 => x"7e",
          9831 => x"00",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"00",
          9836 => x"00",
          9837 => x"00",
          9838 => x"00",
          9839 => x"00",
          9840 => x"00",
          9841 => x"00",
          9842 => x"74",
          9843 => x"00",
          9844 => x"74",
          9845 => x"00",
          9846 => x"00",
          9847 => x"6c",
          9848 => x"25",
          9849 => x"00",
          9850 => x"6c",
          9851 => x"74",
          9852 => x"65",
          9853 => x"20",
          9854 => x"20",
          9855 => x"74",
          9856 => x"20",
          9857 => x"65",
          9858 => x"20",
          9859 => x"2e",
          9860 => x"00",
          9861 => x"6e",
          9862 => x"6f",
          9863 => x"2f",
          9864 => x"61",
          9865 => x"68",
          9866 => x"6f",
          9867 => x"66",
          9868 => x"2c",
          9869 => x"73",
          9870 => x"69",
          9871 => x"00",
          9872 => x"00",
          9873 => x"2c",
          9874 => x"3d",
          9875 => x"5d",
          9876 => x"00",
          9877 => x"00",
          9878 => x"33",
          9879 => x"00",
          9880 => x"4d",
          9881 => x"53",
          9882 => x"00",
          9883 => x"4e",
          9884 => x"20",
          9885 => x"46",
          9886 => x"32",
          9887 => x"00",
          9888 => x"4e",
          9889 => x"20",
          9890 => x"46",
          9891 => x"20",
          9892 => x"00",
          9893 => x"40",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"41",
          9898 => x"80",
          9899 => x"49",
          9900 => x"8f",
          9901 => x"4f",
          9902 => x"55",
          9903 => x"9b",
          9904 => x"9f",
          9905 => x"55",
          9906 => x"a7",
          9907 => x"ab",
          9908 => x"af",
          9909 => x"b3",
          9910 => x"b7",
          9911 => x"bb",
          9912 => x"bf",
          9913 => x"c3",
          9914 => x"c7",
          9915 => x"cb",
          9916 => x"cf",
          9917 => x"d3",
          9918 => x"d7",
          9919 => x"db",
          9920 => x"df",
          9921 => x"e3",
          9922 => x"e7",
          9923 => x"eb",
          9924 => x"ef",
          9925 => x"f3",
          9926 => x"f7",
          9927 => x"fb",
          9928 => x"ff",
          9929 => x"3b",
          9930 => x"2f",
          9931 => x"3a",
          9932 => x"7c",
          9933 => x"00",
          9934 => x"04",
          9935 => x"40",
          9936 => x"00",
          9937 => x"00",
          9938 => x"02",
          9939 => x"08",
          9940 => x"20",
          9941 => x"00",
          9942 => x"00",
          9943 => x"3c",
          9944 => x"00",
          9945 => x"00",
          9946 => x"00",
          9947 => x"44",
          9948 => x"00",
          9949 => x"00",
          9950 => x"00",
          9951 => x"4c",
          9952 => x"00",
          9953 => x"00",
          9954 => x"00",
          9955 => x"54",
          9956 => x"00",
          9957 => x"00",
          9958 => x"00",
          9959 => x"5c",
          9960 => x"00",
          9961 => x"00",
          9962 => x"00",
          9963 => x"64",
          9964 => x"00",
          9965 => x"00",
          9966 => x"00",
          9967 => x"6c",
          9968 => x"00",
          9969 => x"00",
          9970 => x"00",
          9971 => x"74",
          9972 => x"00",
          9973 => x"00",
          9974 => x"00",
          9975 => x"7c",
          9976 => x"00",
          9977 => x"00",
          9978 => x"00",
          9979 => x"84",
          9980 => x"00",
          9981 => x"00",
          9982 => x"00",
          9983 => x"88",
          9984 => x"00",
          9985 => x"00",
          9986 => x"00",
          9987 => x"8c",
          9988 => x"00",
          9989 => x"00",
          9990 => x"00",
          9991 => x"90",
          9992 => x"00",
          9993 => x"00",
          9994 => x"00",
          9995 => x"94",
          9996 => x"00",
          9997 => x"00",
          9998 => x"00",
          9999 => x"98",
         10000 => x"00",
         10001 => x"00",
         10002 => x"00",
         10003 => x"9c",
         10004 => x"00",
         10005 => x"00",
         10006 => x"00",
         10007 => x"a0",
         10008 => x"00",
         10009 => x"00",
         10010 => x"00",
         10011 => x"a8",
         10012 => x"00",
         10013 => x"00",
         10014 => x"00",
         10015 => x"ac",
         10016 => x"00",
         10017 => x"00",
         10018 => x"00",
         10019 => x"b4",
         10020 => x"00",
         10021 => x"00",
         10022 => x"00",
         10023 => x"bc",
         10024 => x"00",
         10025 => x"00",
         10026 => x"00",
         10027 => x"c4",
         10028 => x"00",
         10029 => x"00",
         10030 => x"00",
         10031 => x"cc",
         10032 => x"00",
         10033 => x"00",
         10034 => x"00",
         10035 => x"d4",
         10036 => x"00",
         10037 => x"00",
         10038 => x"00",
         10039 => x"dc",
         10040 => x"00",
         10041 => x"00",
         10042 => x"00",
         10043 => x"e4",
         10044 => x"00",
         10045 => x"00",
         10046 => x"00",
         10047 => x"00",
         10048 => x"00",
         10049 => x"ff",
         10050 => x"00",
         10051 => x"ff",
         10052 => x"00",
         10053 => x"ff",
         10054 => x"00",
         10055 => x"00",
         10056 => x"00",
         10057 => x"ff",
         10058 => x"00",
         10059 => x"00",
         10060 => x"00",
         10061 => x"00",
         10062 => x"00",
         10063 => x"00",
         10064 => x"00",
         10065 => x"00",
         10066 => x"01",
         10067 => x"01",
         10068 => x"01",
         10069 => x"00",
         10070 => x"00",
         10071 => x"00",
         10072 => x"00",
         10073 => x"00",
         10074 => x"00",
         10075 => x"00",
         10076 => x"00",
         10077 => x"00",
         10078 => x"00",
         10079 => x"00",
         10080 => x"00",
         10081 => x"00",
         10082 => x"00",
         10083 => x"00",
         10084 => x"00",
         10085 => x"00",
         10086 => x"00",
         10087 => x"00",
         10088 => x"00",
         10089 => x"00",
         10090 => x"00",
         10091 => x"00",
         10092 => x"00",
         10093 => x"00",
         10094 => x"c8",
         10095 => x"00",
         10096 => x"d0",
         10097 => x"00",
         10098 => x"d8",
         10099 => x"00",
         10100 => x"00",
         10101 => x"00",
         10102 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"83",
             1 => x"0b",
             2 => x"b9",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"82",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"80",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"80",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a4",
           270 => x"0b",
           271 => x"0b",
           272 => x"c2",
           273 => x"0b",
           274 => x"0b",
           275 => x"e0",
           276 => x"0b",
           277 => x"0b",
           278 => x"80",
           279 => x"0b",
           280 => x"0b",
           281 => x"9e",
           282 => x"0b",
           283 => x"0b",
           284 => x"bd",
           285 => x"0b",
           286 => x"0b",
           287 => x"dd",
           288 => x"0b",
           289 => x"0b",
           290 => x"fd",
           291 => x"0b",
           292 => x"0b",
           293 => x"9d",
           294 => x"0b",
           295 => x"0b",
           296 => x"bd",
           297 => x"0b",
           298 => x"0b",
           299 => x"dd",
           300 => x"0b",
           301 => x"0b",
           302 => x"fd",
           303 => x"0b",
           304 => x"0b",
           305 => x"9d",
           306 => x"0b",
           307 => x"0b",
           308 => x"bd",
           309 => x"0b",
           310 => x"0b",
           311 => x"dd",
           312 => x"0b",
           313 => x"0b",
           314 => x"fd",
           315 => x"0b",
           316 => x"0b",
           317 => x"9d",
           318 => x"0b",
           319 => x"0b",
           320 => x"bd",
           321 => x"0b",
           322 => x"0b",
           323 => x"dd",
           324 => x"0b",
           325 => x"0b",
           326 => x"fd",
           327 => x"0b",
           328 => x"0b",
           329 => x"9d",
           330 => x"0b",
           331 => x"0b",
           332 => x"bd",
           333 => x"0b",
           334 => x"0b",
           335 => x"dd",
           336 => x"0b",
           337 => x"0b",
           338 => x"fd",
           339 => x"0b",
           340 => x"0b",
           341 => x"9d",
           342 => x"0b",
           343 => x"0b",
           344 => x"bd",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"bb",
           386 => x"f9",
           387 => x"bb",
           388 => x"d8",
           389 => x"bb",
           390 => x"b2",
           391 => x"e8",
           392 => x"90",
           393 => x"e8",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"82",
           399 => x"82",
           400 => x"82",
           401 => x"94",
           402 => x"bb",
           403 => x"d8",
           404 => x"bb",
           405 => x"c2",
           406 => x"e8",
           407 => x"90",
           408 => x"e8",
           409 => x"cc",
           410 => x"e8",
           411 => x"90",
           412 => x"e8",
           413 => x"fb",
           414 => x"e8",
           415 => x"90",
           416 => x"e8",
           417 => x"2d",
           418 => x"08",
           419 => x"04",
           420 => x"0c",
           421 => x"82",
           422 => x"82",
           423 => x"82",
           424 => x"97",
           425 => x"bb",
           426 => x"d8",
           427 => x"bb",
           428 => x"fc",
           429 => x"bb",
           430 => x"d8",
           431 => x"bb",
           432 => x"fd",
           433 => x"bb",
           434 => x"d8",
           435 => x"bb",
           436 => x"f4",
           437 => x"bb",
           438 => x"d8",
           439 => x"bb",
           440 => x"f6",
           441 => x"bb",
           442 => x"d8",
           443 => x"bb",
           444 => x"f7",
           445 => x"bb",
           446 => x"d8",
           447 => x"bb",
           448 => x"dc",
           449 => x"bb",
           450 => x"d8",
           451 => x"bb",
           452 => x"e9",
           453 => x"bb",
           454 => x"d8",
           455 => x"bb",
           456 => x"e1",
           457 => x"bb",
           458 => x"d8",
           459 => x"bb",
           460 => x"e4",
           461 => x"bb",
           462 => x"d8",
           463 => x"bb",
           464 => x"ee",
           465 => x"bb",
           466 => x"d8",
           467 => x"bb",
           468 => x"f7",
           469 => x"bb",
           470 => x"d8",
           471 => x"bb",
           472 => x"e8",
           473 => x"bb",
           474 => x"d8",
           475 => x"bb",
           476 => x"f2",
           477 => x"bb",
           478 => x"d8",
           479 => x"bb",
           480 => x"f3",
           481 => x"bb",
           482 => x"d8",
           483 => x"bb",
           484 => x"f3",
           485 => x"bb",
           486 => x"d8",
           487 => x"bb",
           488 => x"fb",
           489 => x"bb",
           490 => x"d8",
           491 => x"bb",
           492 => x"f9",
           493 => x"bb",
           494 => x"d8",
           495 => x"bb",
           496 => x"fe",
           497 => x"bb",
           498 => x"d8",
           499 => x"bb",
           500 => x"f4",
           501 => x"bb",
           502 => x"d8",
           503 => x"bb",
           504 => x"81",
           505 => x"bb",
           506 => x"d8",
           507 => x"bb",
           508 => x"82",
           509 => x"bb",
           510 => x"d8",
           511 => x"bb",
           512 => x"ea",
           513 => x"bb",
           514 => x"d8",
           515 => x"bb",
           516 => x"ea",
           517 => x"bb",
           518 => x"d8",
           519 => x"bb",
           520 => x"eb",
           521 => x"bb",
           522 => x"d8",
           523 => x"bb",
           524 => x"f5",
           525 => x"bb",
           526 => x"d8",
           527 => x"bb",
           528 => x"82",
           529 => x"bb",
           530 => x"d8",
           531 => x"bb",
           532 => x"85",
           533 => x"bb",
           534 => x"d8",
           535 => x"bb",
           536 => x"88",
           537 => x"bb",
           538 => x"d8",
           539 => x"bb",
           540 => x"dc",
           541 => x"bb",
           542 => x"d8",
           543 => x"bb",
           544 => x"8b",
           545 => x"bb",
           546 => x"d8",
           547 => x"bb",
           548 => x"99",
           549 => x"bb",
           550 => x"d8",
           551 => x"bb",
           552 => x"97",
           553 => x"bb",
           554 => x"d8",
           555 => x"bb",
           556 => x"ad",
           557 => x"bb",
           558 => x"d8",
           559 => x"bb",
           560 => x"af",
           561 => x"bb",
           562 => x"d8",
           563 => x"bb",
           564 => x"b1",
           565 => x"bb",
           566 => x"d8",
           567 => x"bb",
           568 => x"f4",
           569 => x"bb",
           570 => x"d8",
           571 => x"bb",
           572 => x"f6",
           573 => x"bb",
           574 => x"d8",
           575 => x"bb",
           576 => x"fa",
           577 => x"bb",
           578 => x"d8",
           579 => x"bb",
           580 => x"d6",
           581 => x"bb",
           582 => x"d8",
           583 => x"bb",
           584 => x"a7",
           585 => x"bb",
           586 => x"d8",
           587 => x"bb",
           588 => x"a8",
           589 => x"bb",
           590 => x"d8",
           591 => x"bb",
           592 => x"ab",
           593 => x"bb",
           594 => x"d8",
           595 => x"bb",
           596 => x"a4",
           597 => x"bb",
           598 => x"d8",
           599 => x"04",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"04",
           609 => x"81",
           610 => x"83",
           611 => x"05",
           612 => x"10",
           613 => x"72",
           614 => x"51",
           615 => x"72",
           616 => x"06",
           617 => x"72",
           618 => x"10",
           619 => x"10",
           620 => x"ed",
           621 => x"53",
           622 => x"bb",
           623 => x"d3",
           624 => x"38",
           625 => x"84",
           626 => x"0b",
           627 => x"bc",
           628 => x"51",
           629 => x"04",
           630 => x"e8",
           631 => x"bb",
           632 => x"3d",
           633 => x"e8",
           634 => x"70",
           635 => x"08",
           636 => x"82",
           637 => x"fc",
           638 => x"82",
           639 => x"88",
           640 => x"82",
           641 => x"52",
           642 => x"3f",
           643 => x"08",
           644 => x"e8",
           645 => x"0c",
           646 => x"08",
           647 => x"70",
           648 => x"0c",
           649 => x"3d",
           650 => x"e8",
           651 => x"bb",
           652 => x"82",
           653 => x"fb",
           654 => x"bb",
           655 => x"05",
           656 => x"33",
           657 => x"70",
           658 => x"51",
           659 => x"8f",
           660 => x"82",
           661 => x"8c",
           662 => x"83",
           663 => x"80",
           664 => x"e8",
           665 => x"0c",
           666 => x"82",
           667 => x"8c",
           668 => x"05",
           669 => x"08",
           670 => x"80",
           671 => x"e8",
           672 => x"0c",
           673 => x"08",
           674 => x"82",
           675 => x"fc",
           676 => x"bb",
           677 => x"05",
           678 => x"80",
           679 => x"0b",
           680 => x"08",
           681 => x"25",
           682 => x"82",
           683 => x"90",
           684 => x"a0",
           685 => x"bb",
           686 => x"82",
           687 => x"f8",
           688 => x"82",
           689 => x"f8",
           690 => x"2e",
           691 => x"8d",
           692 => x"82",
           693 => x"f4",
           694 => x"d2",
           695 => x"e8",
           696 => x"08",
           697 => x"08",
           698 => x"53",
           699 => x"34",
           700 => x"08",
           701 => x"ff",
           702 => x"e8",
           703 => x"0c",
           704 => x"08",
           705 => x"81",
           706 => x"e8",
           707 => x"0c",
           708 => x"82",
           709 => x"fc",
           710 => x"80",
           711 => x"bb",
           712 => x"05",
           713 => x"bb",
           714 => x"05",
           715 => x"bb",
           716 => x"05",
           717 => x"dc",
           718 => x"0d",
           719 => x"0c",
           720 => x"e8",
           721 => x"bb",
           722 => x"3d",
           723 => x"82",
           724 => x"e5",
           725 => x"bb",
           726 => x"05",
           727 => x"e8",
           728 => x"0c",
           729 => x"82",
           730 => x"e8",
           731 => x"bb",
           732 => x"05",
           733 => x"e8",
           734 => x"0c",
           735 => x"08",
           736 => x"54",
           737 => x"08",
           738 => x"53",
           739 => x"08",
           740 => x"53",
           741 => x"8d",
           742 => x"dc",
           743 => x"bb",
           744 => x"05",
           745 => x"e8",
           746 => x"08",
           747 => x"08",
           748 => x"05",
           749 => x"74",
           750 => x"e8",
           751 => x"08",
           752 => x"dc",
           753 => x"3d",
           754 => x"e8",
           755 => x"bb",
           756 => x"82",
           757 => x"fb",
           758 => x"bb",
           759 => x"05",
           760 => x"e8",
           761 => x"0c",
           762 => x"08",
           763 => x"54",
           764 => x"08",
           765 => x"53",
           766 => x"08",
           767 => x"52",
           768 => x"82",
           769 => x"70",
           770 => x"08",
           771 => x"82",
           772 => x"f8",
           773 => x"82",
           774 => x"51",
           775 => x"0d",
           776 => x"0c",
           777 => x"e8",
           778 => x"bb",
           779 => x"3d",
           780 => x"82",
           781 => x"e4",
           782 => x"bb",
           783 => x"05",
           784 => x"0b",
           785 => x"82",
           786 => x"88",
           787 => x"11",
           788 => x"2a",
           789 => x"70",
           790 => x"51",
           791 => x"72",
           792 => x"38",
           793 => x"bb",
           794 => x"05",
           795 => x"39",
           796 => x"08",
           797 => x"53",
           798 => x"72",
           799 => x"08",
           800 => x"72",
           801 => x"53",
           802 => x"95",
           803 => x"bb",
           804 => x"05",
           805 => x"82",
           806 => x"8c",
           807 => x"bb",
           808 => x"05",
           809 => x"06",
           810 => x"80",
           811 => x"38",
           812 => x"08",
           813 => x"53",
           814 => x"81",
           815 => x"bb",
           816 => x"05",
           817 => x"b9",
           818 => x"38",
           819 => x"08",
           820 => x"53",
           821 => x"09",
           822 => x"c5",
           823 => x"e8",
           824 => x"33",
           825 => x"70",
           826 => x"51",
           827 => x"38",
           828 => x"08",
           829 => x"70",
           830 => x"81",
           831 => x"06",
           832 => x"53",
           833 => x"99",
           834 => x"e8",
           835 => x"22",
           836 => x"07",
           837 => x"82",
           838 => x"e4",
           839 => x"d0",
           840 => x"e8",
           841 => x"33",
           842 => x"70",
           843 => x"70",
           844 => x"11",
           845 => x"51",
           846 => x"55",
           847 => x"bb",
           848 => x"05",
           849 => x"e8",
           850 => x"33",
           851 => x"e8",
           852 => x"33",
           853 => x"11",
           854 => x"72",
           855 => x"08",
           856 => x"82",
           857 => x"e8",
           858 => x"98",
           859 => x"2c",
           860 => x"72",
           861 => x"38",
           862 => x"82",
           863 => x"e8",
           864 => x"bb",
           865 => x"05",
           866 => x"2a",
           867 => x"51",
           868 => x"fd",
           869 => x"bb",
           870 => x"05",
           871 => x"2b",
           872 => x"70",
           873 => x"88",
           874 => x"51",
           875 => x"82",
           876 => x"ec",
           877 => x"b8",
           878 => x"e8",
           879 => x"22",
           880 => x"70",
           881 => x"51",
           882 => x"2e",
           883 => x"bb",
           884 => x"05",
           885 => x"2b",
           886 => x"51",
           887 => x"8a",
           888 => x"82",
           889 => x"e8",
           890 => x"bb",
           891 => x"05",
           892 => x"82",
           893 => x"c4",
           894 => x"82",
           895 => x"c4",
           896 => x"d8",
           897 => x"38",
           898 => x"08",
           899 => x"70",
           900 => x"9b",
           901 => x"08",
           902 => x"53",
           903 => x"bb",
           904 => x"05",
           905 => x"07",
           906 => x"82",
           907 => x"e4",
           908 => x"bb",
           909 => x"05",
           910 => x"07",
           911 => x"82",
           912 => x"e4",
           913 => x"a8",
           914 => x"e8",
           915 => x"22",
           916 => x"07",
           917 => x"82",
           918 => x"e4",
           919 => x"90",
           920 => x"e8",
           921 => x"22",
           922 => x"07",
           923 => x"82",
           924 => x"e4",
           925 => x"f8",
           926 => x"e8",
           927 => x"22",
           928 => x"51",
           929 => x"bb",
           930 => x"05",
           931 => x"82",
           932 => x"e8",
           933 => x"d8",
           934 => x"e8",
           935 => x"22",
           936 => x"51",
           937 => x"bb",
           938 => x"05",
           939 => x"39",
           940 => x"bb",
           941 => x"05",
           942 => x"e8",
           943 => x"22",
           944 => x"53",
           945 => x"e8",
           946 => x"23",
           947 => x"82",
           948 => x"f8",
           949 => x"a8",
           950 => x"e8",
           951 => x"08",
           952 => x"08",
           953 => x"84",
           954 => x"e8",
           955 => x"0c",
           956 => x"53",
           957 => x"e8",
           958 => x"34",
           959 => x"08",
           960 => x"ff",
           961 => x"72",
           962 => x"08",
           963 => x"8c",
           964 => x"bb",
           965 => x"05",
           966 => x"e8",
           967 => x"08",
           968 => x"bb",
           969 => x"05",
           970 => x"82",
           971 => x"fc",
           972 => x"bb",
           973 => x"05",
           974 => x"2a",
           975 => x"51",
           976 => x"72",
           977 => x"38",
           978 => x"08",
           979 => x"70",
           980 => x"72",
           981 => x"82",
           982 => x"fc",
           983 => x"53",
           984 => x"82",
           985 => x"53",
           986 => x"e8",
           987 => x"23",
           988 => x"bb",
           989 => x"05",
           990 => x"8a",
           991 => x"dc",
           992 => x"82",
           993 => x"f4",
           994 => x"bb",
           995 => x"05",
           996 => x"bb",
           997 => x"05",
           998 => x"31",
           999 => x"82",
          1000 => x"ec",
          1001 => x"d8",
          1002 => x"e8",
          1003 => x"08",
          1004 => x"08",
          1005 => x"84",
          1006 => x"e8",
          1007 => x"0c",
          1008 => x"bb",
          1009 => x"05",
          1010 => x"e8",
          1011 => x"22",
          1012 => x"70",
          1013 => x"51",
          1014 => x"80",
          1015 => x"82",
          1016 => x"e8",
          1017 => x"98",
          1018 => x"98",
          1019 => x"bb",
          1020 => x"05",
          1021 => x"a1",
          1022 => x"bb",
          1023 => x"72",
          1024 => x"08",
          1025 => x"99",
          1026 => x"e8",
          1027 => x"08",
          1028 => x"3f",
          1029 => x"08",
          1030 => x"bb",
          1031 => x"05",
          1032 => x"e8",
          1033 => x"22",
          1034 => x"e8",
          1035 => x"22",
          1036 => x"54",
          1037 => x"bb",
          1038 => x"05",
          1039 => x"39",
          1040 => x"08",
          1041 => x"70",
          1042 => x"81",
          1043 => x"53",
          1044 => x"a4",
          1045 => x"e8",
          1046 => x"08",
          1047 => x"08",
          1048 => x"84",
          1049 => x"e8",
          1050 => x"0c",
          1051 => x"bb",
          1052 => x"05",
          1053 => x"39",
          1054 => x"08",
          1055 => x"82",
          1056 => x"90",
          1057 => x"05",
          1058 => x"08",
          1059 => x"70",
          1060 => x"e8",
          1061 => x"0c",
          1062 => x"e8",
          1063 => x"08",
          1064 => x"08",
          1065 => x"82",
          1066 => x"fc",
          1067 => x"25",
          1068 => x"bb",
          1069 => x"05",
          1070 => x"07",
          1071 => x"82",
          1072 => x"e4",
          1073 => x"bb",
          1074 => x"05",
          1075 => x"bb",
          1076 => x"05",
          1077 => x"e8",
          1078 => x"22",
          1079 => x"06",
          1080 => x"82",
          1081 => x"e4",
          1082 => x"af",
          1083 => x"82",
          1084 => x"f4",
          1085 => x"39",
          1086 => x"08",
          1087 => x"70",
          1088 => x"51",
          1089 => x"bb",
          1090 => x"05",
          1091 => x"0b",
          1092 => x"08",
          1093 => x"90",
          1094 => x"e8",
          1095 => x"23",
          1096 => x"08",
          1097 => x"70",
          1098 => x"81",
          1099 => x"53",
          1100 => x"a4",
          1101 => x"e8",
          1102 => x"08",
          1103 => x"08",
          1104 => x"84",
          1105 => x"e8",
          1106 => x"0c",
          1107 => x"bb",
          1108 => x"05",
          1109 => x"39",
          1110 => x"08",
          1111 => x"82",
          1112 => x"90",
          1113 => x"05",
          1114 => x"08",
          1115 => x"70",
          1116 => x"e8",
          1117 => x"0c",
          1118 => x"e8",
          1119 => x"08",
          1120 => x"08",
          1121 => x"82",
          1122 => x"e4",
          1123 => x"cf",
          1124 => x"72",
          1125 => x"08",
          1126 => x"82",
          1127 => x"82",
          1128 => x"f0",
          1129 => x"bb",
          1130 => x"05",
          1131 => x"e8",
          1132 => x"22",
          1133 => x"08",
          1134 => x"71",
          1135 => x"56",
          1136 => x"f3",
          1137 => x"dc",
          1138 => x"75",
          1139 => x"e8",
          1140 => x"08",
          1141 => x"08",
          1142 => x"82",
          1143 => x"f0",
          1144 => x"33",
          1145 => x"73",
          1146 => x"82",
          1147 => x"f0",
          1148 => x"72",
          1149 => x"bb",
          1150 => x"05",
          1151 => x"df",
          1152 => x"53",
          1153 => x"e8",
          1154 => x"34",
          1155 => x"bb",
          1156 => x"05",
          1157 => x"33",
          1158 => x"53",
          1159 => x"e8",
          1160 => x"34",
          1161 => x"08",
          1162 => x"53",
          1163 => x"08",
          1164 => x"73",
          1165 => x"e8",
          1166 => x"08",
          1167 => x"bb",
          1168 => x"05",
          1169 => x"e8",
          1170 => x"22",
          1171 => x"bb",
          1172 => x"05",
          1173 => x"a2",
          1174 => x"bb",
          1175 => x"82",
          1176 => x"fc",
          1177 => x"82",
          1178 => x"fc",
          1179 => x"2e",
          1180 => x"b2",
          1181 => x"e8",
          1182 => x"08",
          1183 => x"54",
          1184 => x"74",
          1185 => x"51",
          1186 => x"bb",
          1187 => x"05",
          1188 => x"e8",
          1189 => x"22",
          1190 => x"51",
          1191 => x"2e",
          1192 => x"bb",
          1193 => x"05",
          1194 => x"51",
          1195 => x"bb",
          1196 => x"05",
          1197 => x"e8",
          1198 => x"22",
          1199 => x"70",
          1200 => x"51",
          1201 => x"2e",
          1202 => x"82",
          1203 => x"ec",
          1204 => x"90",
          1205 => x"e8",
          1206 => x"0c",
          1207 => x"08",
          1208 => x"90",
          1209 => x"e8",
          1210 => x"0c",
          1211 => x"08",
          1212 => x"51",
          1213 => x"2e",
          1214 => x"95",
          1215 => x"e8",
          1216 => x"08",
          1217 => x"72",
          1218 => x"08",
          1219 => x"93",
          1220 => x"e8",
          1221 => x"08",
          1222 => x"72",
          1223 => x"08",
          1224 => x"82",
          1225 => x"c8",
          1226 => x"bb",
          1227 => x"05",
          1228 => x"e8",
          1229 => x"22",
          1230 => x"70",
          1231 => x"51",
          1232 => x"2e",
          1233 => x"82",
          1234 => x"e8",
          1235 => x"98",
          1236 => x"2c",
          1237 => x"08",
          1238 => x"57",
          1239 => x"72",
          1240 => x"38",
          1241 => x"08",
          1242 => x"70",
          1243 => x"53",
          1244 => x"e8",
          1245 => x"23",
          1246 => x"bb",
          1247 => x"05",
          1248 => x"bb",
          1249 => x"05",
          1250 => x"31",
          1251 => x"82",
          1252 => x"e8",
          1253 => x"bb",
          1254 => x"05",
          1255 => x"2a",
          1256 => x"51",
          1257 => x"80",
          1258 => x"82",
          1259 => x"e8",
          1260 => x"88",
          1261 => x"2b",
          1262 => x"70",
          1263 => x"51",
          1264 => x"72",
          1265 => x"e8",
          1266 => x"22",
          1267 => x"51",
          1268 => x"bb",
          1269 => x"05",
          1270 => x"82",
          1271 => x"fc",
          1272 => x"88",
          1273 => x"2b",
          1274 => x"70",
          1275 => x"51",
          1276 => x"72",
          1277 => x"e8",
          1278 => x"22",
          1279 => x"51",
          1280 => x"bb",
          1281 => x"05",
          1282 => x"e8",
          1283 => x"22",
          1284 => x"06",
          1285 => x"b0",
          1286 => x"e8",
          1287 => x"22",
          1288 => x"54",
          1289 => x"e8",
          1290 => x"23",
          1291 => x"70",
          1292 => x"53",
          1293 => x"90",
          1294 => x"e8",
          1295 => x"08",
          1296 => x"8a",
          1297 => x"39",
          1298 => x"08",
          1299 => x"70",
          1300 => x"81",
          1301 => x"53",
          1302 => x"91",
          1303 => x"e8",
          1304 => x"08",
          1305 => x"8a",
          1306 => x"c7",
          1307 => x"e8",
          1308 => x"22",
          1309 => x"70",
          1310 => x"51",
          1311 => x"2e",
          1312 => x"bb",
          1313 => x"05",
          1314 => x"51",
          1315 => x"a3",
          1316 => x"e8",
          1317 => x"22",
          1318 => x"70",
          1319 => x"51",
          1320 => x"2e",
          1321 => x"bb",
          1322 => x"05",
          1323 => x"51",
          1324 => x"82",
          1325 => x"e4",
          1326 => x"86",
          1327 => x"06",
          1328 => x"72",
          1329 => x"38",
          1330 => x"08",
          1331 => x"52",
          1332 => x"df",
          1333 => x"e8",
          1334 => x"22",
          1335 => x"2e",
          1336 => x"94",
          1337 => x"e8",
          1338 => x"08",
          1339 => x"e8",
          1340 => x"33",
          1341 => x"3f",
          1342 => x"08",
          1343 => x"70",
          1344 => x"81",
          1345 => x"53",
          1346 => x"b0",
          1347 => x"e8",
          1348 => x"22",
          1349 => x"54",
          1350 => x"e8",
          1351 => x"23",
          1352 => x"70",
          1353 => x"53",
          1354 => x"90",
          1355 => x"e8",
          1356 => x"08",
          1357 => x"88",
          1358 => x"39",
          1359 => x"08",
          1360 => x"70",
          1361 => x"81",
          1362 => x"53",
          1363 => x"b0",
          1364 => x"e8",
          1365 => x"33",
          1366 => x"54",
          1367 => x"e8",
          1368 => x"34",
          1369 => x"70",
          1370 => x"53",
          1371 => x"90",
          1372 => x"e8",
          1373 => x"08",
          1374 => x"88",
          1375 => x"39",
          1376 => x"08",
          1377 => x"70",
          1378 => x"81",
          1379 => x"53",
          1380 => x"82",
          1381 => x"ec",
          1382 => x"11",
          1383 => x"82",
          1384 => x"ec",
          1385 => x"90",
          1386 => x"2c",
          1387 => x"73",
          1388 => x"82",
          1389 => x"88",
          1390 => x"a0",
          1391 => x"3f",
          1392 => x"bb",
          1393 => x"05",
          1394 => x"80",
          1395 => x"81",
          1396 => x"82",
          1397 => x"88",
          1398 => x"82",
          1399 => x"fc",
          1400 => x"87",
          1401 => x"ee",
          1402 => x"e8",
          1403 => x"33",
          1404 => x"f3",
          1405 => x"06",
          1406 => x"82",
          1407 => x"f4",
          1408 => x"11",
          1409 => x"82",
          1410 => x"f4",
          1411 => x"83",
          1412 => x"53",
          1413 => x"ff",
          1414 => x"38",
          1415 => x"08",
          1416 => x"52",
          1417 => x"08",
          1418 => x"70",
          1419 => x"bb",
          1420 => x"05",
          1421 => x"82",
          1422 => x"fc",
          1423 => x"86",
          1424 => x"b7",
          1425 => x"e8",
          1426 => x"33",
          1427 => x"d3",
          1428 => x"06",
          1429 => x"82",
          1430 => x"f4",
          1431 => x"11",
          1432 => x"82",
          1433 => x"f4",
          1434 => x"83",
          1435 => x"53",
          1436 => x"ff",
          1437 => x"38",
          1438 => x"08",
          1439 => x"52",
          1440 => x"08",
          1441 => x"70",
          1442 => x"86",
          1443 => x"bb",
          1444 => x"05",
          1445 => x"82",
          1446 => x"fc",
          1447 => x"b7",
          1448 => x"e8",
          1449 => x"08",
          1450 => x"2e",
          1451 => x"bb",
          1452 => x"05",
          1453 => x"bb",
          1454 => x"05",
          1455 => x"82",
          1456 => x"f0",
          1457 => x"bb",
          1458 => x"05",
          1459 => x"52",
          1460 => x"3f",
          1461 => x"bb",
          1462 => x"05",
          1463 => x"2a",
          1464 => x"51",
          1465 => x"80",
          1466 => x"38",
          1467 => x"08",
          1468 => x"ff",
          1469 => x"72",
          1470 => x"08",
          1471 => x"73",
          1472 => x"90",
          1473 => x"80",
          1474 => x"38",
          1475 => x"08",
          1476 => x"52",
          1477 => x"9b",
          1478 => x"82",
          1479 => x"88",
          1480 => x"82",
          1481 => x"f8",
          1482 => x"85",
          1483 => x"0b",
          1484 => x"08",
          1485 => x"ea",
          1486 => x"bb",
          1487 => x"05",
          1488 => x"a5",
          1489 => x"06",
          1490 => x"0b",
          1491 => x"08",
          1492 => x"80",
          1493 => x"e8",
          1494 => x"23",
          1495 => x"bb",
          1496 => x"05",
          1497 => x"82",
          1498 => x"f4",
          1499 => x"80",
          1500 => x"e8",
          1501 => x"08",
          1502 => x"e8",
          1503 => x"33",
          1504 => x"3f",
          1505 => x"82",
          1506 => x"88",
          1507 => x"11",
          1508 => x"bb",
          1509 => x"05",
          1510 => x"82",
          1511 => x"e0",
          1512 => x"bb",
          1513 => x"3d",
          1514 => x"e8",
          1515 => x"bb",
          1516 => x"82",
          1517 => x"fd",
          1518 => x"d3",
          1519 => x"82",
          1520 => x"8c",
          1521 => x"82",
          1522 => x"88",
          1523 => x"e4",
          1524 => x"bb",
          1525 => x"82",
          1526 => x"54",
          1527 => x"82",
          1528 => x"04",
          1529 => x"08",
          1530 => x"e8",
          1531 => x"0d",
          1532 => x"bb",
          1533 => x"05",
          1534 => x"b0",
          1535 => x"33",
          1536 => x"70",
          1537 => x"81",
          1538 => x"51",
          1539 => x"80",
          1540 => x"ff",
          1541 => x"e8",
          1542 => x"0c",
          1543 => x"82",
          1544 => x"88",
          1545 => x"72",
          1546 => x"e8",
          1547 => x"08",
          1548 => x"bb",
          1549 => x"05",
          1550 => x"82",
          1551 => x"fc",
          1552 => x"81",
          1553 => x"72",
          1554 => x"38",
          1555 => x"08",
          1556 => x"08",
          1557 => x"e8",
          1558 => x"33",
          1559 => x"08",
          1560 => x"2d",
          1561 => x"08",
          1562 => x"2e",
          1563 => x"ff",
          1564 => x"e8",
          1565 => x"0c",
          1566 => x"82",
          1567 => x"82",
          1568 => x"53",
          1569 => x"90",
          1570 => x"72",
          1571 => x"dc",
          1572 => x"80",
          1573 => x"ff",
          1574 => x"e8",
          1575 => x"0c",
          1576 => x"08",
          1577 => x"70",
          1578 => x"08",
          1579 => x"53",
          1580 => x"08",
          1581 => x"82",
          1582 => x"87",
          1583 => x"bb",
          1584 => x"82",
          1585 => x"02",
          1586 => x"0c",
          1587 => x"80",
          1588 => x"e8",
          1589 => x"0c",
          1590 => x"08",
          1591 => x"85",
          1592 => x"81",
          1593 => x"32",
          1594 => x"51",
          1595 => x"53",
          1596 => x"8d",
          1597 => x"82",
          1598 => x"f4",
          1599 => x"f3",
          1600 => x"e8",
          1601 => x"08",
          1602 => x"82",
          1603 => x"88",
          1604 => x"05",
          1605 => x"08",
          1606 => x"53",
          1607 => x"e8",
          1608 => x"34",
          1609 => x"06",
          1610 => x"2e",
          1611 => x"bb",
          1612 => x"05",
          1613 => x"e8",
          1614 => x"08",
          1615 => x"e8",
          1616 => x"33",
          1617 => x"08",
          1618 => x"2d",
          1619 => x"08",
          1620 => x"2e",
          1621 => x"ff",
          1622 => x"e8",
          1623 => x"0c",
          1624 => x"82",
          1625 => x"f8",
          1626 => x"82",
          1627 => x"f4",
          1628 => x"82",
          1629 => x"f4",
          1630 => x"bb",
          1631 => x"3d",
          1632 => x"e8",
          1633 => x"bb",
          1634 => x"82",
          1635 => x"fe",
          1636 => x"d3",
          1637 => x"82",
          1638 => x"88",
          1639 => x"93",
          1640 => x"dc",
          1641 => x"bb",
          1642 => x"84",
          1643 => x"bb",
          1644 => x"82",
          1645 => x"02",
          1646 => x"0c",
          1647 => x"82",
          1648 => x"8c",
          1649 => x"11",
          1650 => x"2a",
          1651 => x"70",
          1652 => x"51",
          1653 => x"72",
          1654 => x"38",
          1655 => x"bb",
          1656 => x"05",
          1657 => x"39",
          1658 => x"08",
          1659 => x"85",
          1660 => x"82",
          1661 => x"06",
          1662 => x"53",
          1663 => x"80",
          1664 => x"bb",
          1665 => x"05",
          1666 => x"e8",
          1667 => x"08",
          1668 => x"14",
          1669 => x"08",
          1670 => x"82",
          1671 => x"8c",
          1672 => x"08",
          1673 => x"e8",
          1674 => x"08",
          1675 => x"54",
          1676 => x"73",
          1677 => x"74",
          1678 => x"e8",
          1679 => x"08",
          1680 => x"81",
          1681 => x"0c",
          1682 => x"08",
          1683 => x"70",
          1684 => x"08",
          1685 => x"51",
          1686 => x"39",
          1687 => x"08",
          1688 => x"82",
          1689 => x"8c",
          1690 => x"82",
          1691 => x"88",
          1692 => x"81",
          1693 => x"90",
          1694 => x"54",
          1695 => x"82",
          1696 => x"53",
          1697 => x"82",
          1698 => x"8c",
          1699 => x"11",
          1700 => x"8c",
          1701 => x"bb",
          1702 => x"05",
          1703 => x"bb",
          1704 => x"05",
          1705 => x"8a",
          1706 => x"82",
          1707 => x"fc",
          1708 => x"bb",
          1709 => x"05",
          1710 => x"dc",
          1711 => x"0d",
          1712 => x"0c",
          1713 => x"e8",
          1714 => x"bb",
          1715 => x"3d",
          1716 => x"e8",
          1717 => x"08",
          1718 => x"70",
          1719 => x"81",
          1720 => x"51",
          1721 => x"2e",
          1722 => x"0b",
          1723 => x"08",
          1724 => x"83",
          1725 => x"bb",
          1726 => x"05",
          1727 => x"33",
          1728 => x"70",
          1729 => x"51",
          1730 => x"80",
          1731 => x"38",
          1732 => x"08",
          1733 => x"82",
          1734 => x"88",
          1735 => x"53",
          1736 => x"70",
          1737 => x"51",
          1738 => x"14",
          1739 => x"e8",
          1740 => x"08",
          1741 => x"81",
          1742 => x"0c",
          1743 => x"08",
          1744 => x"84",
          1745 => x"82",
          1746 => x"f8",
          1747 => x"51",
          1748 => x"39",
          1749 => x"08",
          1750 => x"85",
          1751 => x"82",
          1752 => x"06",
          1753 => x"52",
          1754 => x"80",
          1755 => x"bb",
          1756 => x"05",
          1757 => x"70",
          1758 => x"e8",
          1759 => x"0c",
          1760 => x"bb",
          1761 => x"05",
          1762 => x"82",
          1763 => x"88",
          1764 => x"bb",
          1765 => x"05",
          1766 => x"85",
          1767 => x"a0",
          1768 => x"71",
          1769 => x"ff",
          1770 => x"e8",
          1771 => x"0c",
          1772 => x"82",
          1773 => x"88",
          1774 => x"08",
          1775 => x"0c",
          1776 => x"39",
          1777 => x"08",
          1778 => x"82",
          1779 => x"88",
          1780 => x"94",
          1781 => x"52",
          1782 => x"bb",
          1783 => x"82",
          1784 => x"fc",
          1785 => x"82",
          1786 => x"fc",
          1787 => x"25",
          1788 => x"82",
          1789 => x"88",
          1790 => x"bb",
          1791 => x"05",
          1792 => x"e8",
          1793 => x"08",
          1794 => x"82",
          1795 => x"f0",
          1796 => x"82",
          1797 => x"fc",
          1798 => x"2e",
          1799 => x"95",
          1800 => x"e8",
          1801 => x"08",
          1802 => x"71",
          1803 => x"08",
          1804 => x"93",
          1805 => x"e8",
          1806 => x"08",
          1807 => x"71",
          1808 => x"08",
          1809 => x"82",
          1810 => x"f4",
          1811 => x"82",
          1812 => x"ec",
          1813 => x"13",
          1814 => x"82",
          1815 => x"f8",
          1816 => x"39",
          1817 => x"08",
          1818 => x"8c",
          1819 => x"05",
          1820 => x"82",
          1821 => x"fc",
          1822 => x"81",
          1823 => x"82",
          1824 => x"f8",
          1825 => x"51",
          1826 => x"e8",
          1827 => x"08",
          1828 => x"0c",
          1829 => x"82",
          1830 => x"04",
          1831 => x"08",
          1832 => x"e8",
          1833 => x"0d",
          1834 => x"08",
          1835 => x"82",
          1836 => x"fc",
          1837 => x"bb",
          1838 => x"05",
          1839 => x"e8",
          1840 => x"0c",
          1841 => x"08",
          1842 => x"80",
          1843 => x"38",
          1844 => x"08",
          1845 => x"82",
          1846 => x"fc",
          1847 => x"81",
          1848 => x"bb",
          1849 => x"05",
          1850 => x"e8",
          1851 => x"08",
          1852 => x"bb",
          1853 => x"05",
          1854 => x"81",
          1855 => x"bb",
          1856 => x"05",
          1857 => x"e8",
          1858 => x"08",
          1859 => x"e8",
          1860 => x"0c",
          1861 => x"08",
          1862 => x"82",
          1863 => x"90",
          1864 => x"82",
          1865 => x"f8",
          1866 => x"bb",
          1867 => x"05",
          1868 => x"82",
          1869 => x"90",
          1870 => x"bb",
          1871 => x"05",
          1872 => x"82",
          1873 => x"90",
          1874 => x"bb",
          1875 => x"05",
          1876 => x"81",
          1877 => x"bb",
          1878 => x"05",
          1879 => x"82",
          1880 => x"fc",
          1881 => x"bb",
          1882 => x"05",
          1883 => x"82",
          1884 => x"f8",
          1885 => x"bb",
          1886 => x"05",
          1887 => x"e8",
          1888 => x"08",
          1889 => x"33",
          1890 => x"ae",
          1891 => x"e8",
          1892 => x"08",
          1893 => x"bb",
          1894 => x"05",
          1895 => x"e8",
          1896 => x"08",
          1897 => x"bb",
          1898 => x"05",
          1899 => x"e8",
          1900 => x"08",
          1901 => x"38",
          1902 => x"08",
          1903 => x"51",
          1904 => x"bb",
          1905 => x"05",
          1906 => x"82",
          1907 => x"f8",
          1908 => x"bb",
          1909 => x"05",
          1910 => x"71",
          1911 => x"bb",
          1912 => x"05",
          1913 => x"82",
          1914 => x"fc",
          1915 => x"ad",
          1916 => x"e8",
          1917 => x"08",
          1918 => x"dc",
          1919 => x"3d",
          1920 => x"e8",
          1921 => x"bb",
          1922 => x"82",
          1923 => x"fe",
          1924 => x"bb",
          1925 => x"05",
          1926 => x"e8",
          1927 => x"0c",
          1928 => x"08",
          1929 => x"52",
          1930 => x"bb",
          1931 => x"05",
          1932 => x"82",
          1933 => x"fc",
          1934 => x"81",
          1935 => x"51",
          1936 => x"83",
          1937 => x"82",
          1938 => x"fc",
          1939 => x"05",
          1940 => x"08",
          1941 => x"82",
          1942 => x"fc",
          1943 => x"bb",
          1944 => x"05",
          1945 => x"82",
          1946 => x"51",
          1947 => x"82",
          1948 => x"04",
          1949 => x"08",
          1950 => x"e8",
          1951 => x"0d",
          1952 => x"08",
          1953 => x"82",
          1954 => x"fc",
          1955 => x"bb",
          1956 => x"05",
          1957 => x"33",
          1958 => x"08",
          1959 => x"81",
          1960 => x"e8",
          1961 => x"0c",
          1962 => x"08",
          1963 => x"53",
          1964 => x"34",
          1965 => x"08",
          1966 => x"81",
          1967 => x"e8",
          1968 => x"0c",
          1969 => x"06",
          1970 => x"2e",
          1971 => x"be",
          1972 => x"e8",
          1973 => x"08",
          1974 => x"dc",
          1975 => x"3d",
          1976 => x"e8",
          1977 => x"bb",
          1978 => x"82",
          1979 => x"fd",
          1980 => x"bb",
          1981 => x"05",
          1982 => x"e8",
          1983 => x"0c",
          1984 => x"08",
          1985 => x"82",
          1986 => x"f8",
          1987 => x"bb",
          1988 => x"05",
          1989 => x"80",
          1990 => x"bb",
          1991 => x"05",
          1992 => x"82",
          1993 => x"90",
          1994 => x"bb",
          1995 => x"05",
          1996 => x"82",
          1997 => x"90",
          1998 => x"bb",
          1999 => x"05",
          2000 => x"ba",
          2001 => x"e8",
          2002 => x"08",
          2003 => x"82",
          2004 => x"f8",
          2005 => x"05",
          2006 => x"08",
          2007 => x"82",
          2008 => x"fc",
          2009 => x"52",
          2010 => x"82",
          2011 => x"fc",
          2012 => x"05",
          2013 => x"08",
          2014 => x"ff",
          2015 => x"bb",
          2016 => x"05",
          2017 => x"bb",
          2018 => x"85",
          2019 => x"bb",
          2020 => x"82",
          2021 => x"02",
          2022 => x"0c",
          2023 => x"82",
          2024 => x"90",
          2025 => x"2e",
          2026 => x"82",
          2027 => x"8c",
          2028 => x"71",
          2029 => x"e8",
          2030 => x"08",
          2031 => x"bb",
          2032 => x"05",
          2033 => x"e8",
          2034 => x"08",
          2035 => x"81",
          2036 => x"54",
          2037 => x"71",
          2038 => x"80",
          2039 => x"bb",
          2040 => x"05",
          2041 => x"33",
          2042 => x"08",
          2043 => x"81",
          2044 => x"e8",
          2045 => x"0c",
          2046 => x"06",
          2047 => x"8d",
          2048 => x"82",
          2049 => x"fc",
          2050 => x"9b",
          2051 => x"e8",
          2052 => x"08",
          2053 => x"bb",
          2054 => x"05",
          2055 => x"e8",
          2056 => x"08",
          2057 => x"38",
          2058 => x"82",
          2059 => x"90",
          2060 => x"2e",
          2061 => x"82",
          2062 => x"88",
          2063 => x"33",
          2064 => x"8d",
          2065 => x"82",
          2066 => x"fc",
          2067 => x"d7",
          2068 => x"e8",
          2069 => x"08",
          2070 => x"bb",
          2071 => x"05",
          2072 => x"e8",
          2073 => x"08",
          2074 => x"52",
          2075 => x"81",
          2076 => x"e8",
          2077 => x"0c",
          2078 => x"bb",
          2079 => x"05",
          2080 => x"82",
          2081 => x"8c",
          2082 => x"33",
          2083 => x"70",
          2084 => x"08",
          2085 => x"53",
          2086 => x"53",
          2087 => x"0b",
          2088 => x"08",
          2089 => x"82",
          2090 => x"fc",
          2091 => x"bb",
          2092 => x"3d",
          2093 => x"e8",
          2094 => x"bb",
          2095 => x"82",
          2096 => x"fd",
          2097 => x"bb",
          2098 => x"05",
          2099 => x"e8",
          2100 => x"0c",
          2101 => x"08",
          2102 => x"8d",
          2103 => x"82",
          2104 => x"fc",
          2105 => x"ec",
          2106 => x"e8",
          2107 => x"08",
          2108 => x"82",
          2109 => x"f8",
          2110 => x"05",
          2111 => x"08",
          2112 => x"70",
          2113 => x"51",
          2114 => x"2e",
          2115 => x"bb",
          2116 => x"05",
          2117 => x"82",
          2118 => x"8c",
          2119 => x"bb",
          2120 => x"05",
          2121 => x"84",
          2122 => x"39",
          2123 => x"08",
          2124 => x"ff",
          2125 => x"e8",
          2126 => x"0c",
          2127 => x"08",
          2128 => x"82",
          2129 => x"88",
          2130 => x"70",
          2131 => x"08",
          2132 => x"51",
          2133 => x"08",
          2134 => x"82",
          2135 => x"85",
          2136 => x"bb",
          2137 => x"82",
          2138 => x"02",
          2139 => x"0c",
          2140 => x"82",
          2141 => x"88",
          2142 => x"bb",
          2143 => x"05",
          2144 => x"e8",
          2145 => x"08",
          2146 => x"d4",
          2147 => x"e8",
          2148 => x"08",
          2149 => x"bb",
          2150 => x"05",
          2151 => x"e8",
          2152 => x"08",
          2153 => x"bb",
          2154 => x"05",
          2155 => x"e8",
          2156 => x"08",
          2157 => x"38",
          2158 => x"08",
          2159 => x"51",
          2160 => x"e8",
          2161 => x"08",
          2162 => x"71",
          2163 => x"e8",
          2164 => x"08",
          2165 => x"bb",
          2166 => x"05",
          2167 => x"39",
          2168 => x"08",
          2169 => x"70",
          2170 => x"0c",
          2171 => x"0d",
          2172 => x"0c",
          2173 => x"e8",
          2174 => x"bb",
          2175 => x"3d",
          2176 => x"82",
          2177 => x"fc",
          2178 => x"bb",
          2179 => x"05",
          2180 => x"b9",
          2181 => x"e8",
          2182 => x"08",
          2183 => x"e8",
          2184 => x"0c",
          2185 => x"bb",
          2186 => x"05",
          2187 => x"e8",
          2188 => x"08",
          2189 => x"0b",
          2190 => x"08",
          2191 => x"82",
          2192 => x"f4",
          2193 => x"bb",
          2194 => x"05",
          2195 => x"e8",
          2196 => x"08",
          2197 => x"38",
          2198 => x"08",
          2199 => x"30",
          2200 => x"08",
          2201 => x"80",
          2202 => x"e8",
          2203 => x"0c",
          2204 => x"08",
          2205 => x"8a",
          2206 => x"82",
          2207 => x"f0",
          2208 => x"bb",
          2209 => x"05",
          2210 => x"e8",
          2211 => x"0c",
          2212 => x"bb",
          2213 => x"05",
          2214 => x"bb",
          2215 => x"05",
          2216 => x"c5",
          2217 => x"dc",
          2218 => x"bb",
          2219 => x"05",
          2220 => x"bb",
          2221 => x"05",
          2222 => x"90",
          2223 => x"e8",
          2224 => x"08",
          2225 => x"e8",
          2226 => x"0c",
          2227 => x"08",
          2228 => x"70",
          2229 => x"0c",
          2230 => x"0d",
          2231 => x"0c",
          2232 => x"e8",
          2233 => x"bb",
          2234 => x"3d",
          2235 => x"82",
          2236 => x"fc",
          2237 => x"bb",
          2238 => x"05",
          2239 => x"99",
          2240 => x"e8",
          2241 => x"08",
          2242 => x"e8",
          2243 => x"0c",
          2244 => x"bb",
          2245 => x"05",
          2246 => x"e8",
          2247 => x"08",
          2248 => x"38",
          2249 => x"08",
          2250 => x"30",
          2251 => x"08",
          2252 => x"81",
          2253 => x"e8",
          2254 => x"08",
          2255 => x"e8",
          2256 => x"08",
          2257 => x"3f",
          2258 => x"08",
          2259 => x"e8",
          2260 => x"0c",
          2261 => x"e8",
          2262 => x"08",
          2263 => x"38",
          2264 => x"08",
          2265 => x"30",
          2266 => x"08",
          2267 => x"82",
          2268 => x"f8",
          2269 => x"82",
          2270 => x"54",
          2271 => x"82",
          2272 => x"04",
          2273 => x"08",
          2274 => x"e8",
          2275 => x"0d",
          2276 => x"bb",
          2277 => x"05",
          2278 => x"bb",
          2279 => x"05",
          2280 => x"c5",
          2281 => x"dc",
          2282 => x"bb",
          2283 => x"85",
          2284 => x"bb",
          2285 => x"82",
          2286 => x"02",
          2287 => x"0c",
          2288 => x"81",
          2289 => x"e8",
          2290 => x"08",
          2291 => x"e8",
          2292 => x"08",
          2293 => x"82",
          2294 => x"70",
          2295 => x"0c",
          2296 => x"0d",
          2297 => x"0c",
          2298 => x"e8",
          2299 => x"bb",
          2300 => x"3d",
          2301 => x"82",
          2302 => x"fc",
          2303 => x"0b",
          2304 => x"08",
          2305 => x"82",
          2306 => x"8c",
          2307 => x"bb",
          2308 => x"05",
          2309 => x"38",
          2310 => x"08",
          2311 => x"80",
          2312 => x"80",
          2313 => x"e8",
          2314 => x"08",
          2315 => x"82",
          2316 => x"8c",
          2317 => x"82",
          2318 => x"8c",
          2319 => x"bb",
          2320 => x"05",
          2321 => x"bb",
          2322 => x"05",
          2323 => x"39",
          2324 => x"08",
          2325 => x"80",
          2326 => x"38",
          2327 => x"08",
          2328 => x"82",
          2329 => x"88",
          2330 => x"ad",
          2331 => x"e8",
          2332 => x"08",
          2333 => x"08",
          2334 => x"31",
          2335 => x"08",
          2336 => x"82",
          2337 => x"f8",
          2338 => x"bb",
          2339 => x"05",
          2340 => x"bb",
          2341 => x"05",
          2342 => x"e8",
          2343 => x"08",
          2344 => x"bb",
          2345 => x"05",
          2346 => x"e8",
          2347 => x"08",
          2348 => x"bb",
          2349 => x"05",
          2350 => x"39",
          2351 => x"08",
          2352 => x"80",
          2353 => x"82",
          2354 => x"88",
          2355 => x"82",
          2356 => x"f4",
          2357 => x"91",
          2358 => x"e8",
          2359 => x"08",
          2360 => x"e8",
          2361 => x"0c",
          2362 => x"e8",
          2363 => x"08",
          2364 => x"0c",
          2365 => x"82",
          2366 => x"04",
          2367 => x"08",
          2368 => x"e8",
          2369 => x"0d",
          2370 => x"bb",
          2371 => x"05",
          2372 => x"e8",
          2373 => x"08",
          2374 => x"0c",
          2375 => x"08",
          2376 => x"70",
          2377 => x"72",
          2378 => x"82",
          2379 => x"f8",
          2380 => x"81",
          2381 => x"72",
          2382 => x"81",
          2383 => x"82",
          2384 => x"88",
          2385 => x"08",
          2386 => x"0c",
          2387 => x"82",
          2388 => x"f8",
          2389 => x"72",
          2390 => x"81",
          2391 => x"81",
          2392 => x"e8",
          2393 => x"34",
          2394 => x"08",
          2395 => x"70",
          2396 => x"71",
          2397 => x"51",
          2398 => x"82",
          2399 => x"f8",
          2400 => x"bb",
          2401 => x"05",
          2402 => x"b0",
          2403 => x"06",
          2404 => x"82",
          2405 => x"88",
          2406 => x"08",
          2407 => x"0c",
          2408 => x"53",
          2409 => x"bb",
          2410 => x"05",
          2411 => x"e8",
          2412 => x"33",
          2413 => x"08",
          2414 => x"82",
          2415 => x"e8",
          2416 => x"e2",
          2417 => x"82",
          2418 => x"e8",
          2419 => x"f8",
          2420 => x"80",
          2421 => x"0b",
          2422 => x"08",
          2423 => x"82",
          2424 => x"88",
          2425 => x"08",
          2426 => x"0c",
          2427 => x"53",
          2428 => x"bb",
          2429 => x"05",
          2430 => x"39",
          2431 => x"bb",
          2432 => x"05",
          2433 => x"e8",
          2434 => x"08",
          2435 => x"05",
          2436 => x"08",
          2437 => x"33",
          2438 => x"08",
          2439 => x"80",
          2440 => x"bb",
          2441 => x"05",
          2442 => x"a0",
          2443 => x"81",
          2444 => x"e8",
          2445 => x"0c",
          2446 => x"82",
          2447 => x"f8",
          2448 => x"af",
          2449 => x"38",
          2450 => x"08",
          2451 => x"53",
          2452 => x"83",
          2453 => x"80",
          2454 => x"e8",
          2455 => x"0c",
          2456 => x"88",
          2457 => x"e8",
          2458 => x"34",
          2459 => x"bb",
          2460 => x"05",
          2461 => x"73",
          2462 => x"82",
          2463 => x"f8",
          2464 => x"72",
          2465 => x"38",
          2466 => x"0b",
          2467 => x"08",
          2468 => x"82",
          2469 => x"0b",
          2470 => x"08",
          2471 => x"80",
          2472 => x"e8",
          2473 => x"0c",
          2474 => x"08",
          2475 => x"53",
          2476 => x"81",
          2477 => x"bb",
          2478 => x"05",
          2479 => x"e0",
          2480 => x"38",
          2481 => x"08",
          2482 => x"e0",
          2483 => x"72",
          2484 => x"08",
          2485 => x"82",
          2486 => x"f8",
          2487 => x"11",
          2488 => x"82",
          2489 => x"f8",
          2490 => x"bb",
          2491 => x"05",
          2492 => x"73",
          2493 => x"82",
          2494 => x"f8",
          2495 => x"11",
          2496 => x"82",
          2497 => x"f8",
          2498 => x"bb",
          2499 => x"05",
          2500 => x"89",
          2501 => x"80",
          2502 => x"e8",
          2503 => x"0c",
          2504 => x"82",
          2505 => x"f8",
          2506 => x"bb",
          2507 => x"05",
          2508 => x"72",
          2509 => x"38",
          2510 => x"bb",
          2511 => x"05",
          2512 => x"39",
          2513 => x"08",
          2514 => x"70",
          2515 => x"08",
          2516 => x"29",
          2517 => x"08",
          2518 => x"70",
          2519 => x"e8",
          2520 => x"0c",
          2521 => x"08",
          2522 => x"70",
          2523 => x"71",
          2524 => x"51",
          2525 => x"53",
          2526 => x"bb",
          2527 => x"05",
          2528 => x"39",
          2529 => x"08",
          2530 => x"53",
          2531 => x"90",
          2532 => x"e8",
          2533 => x"08",
          2534 => x"e8",
          2535 => x"0c",
          2536 => x"08",
          2537 => x"82",
          2538 => x"fc",
          2539 => x"0c",
          2540 => x"82",
          2541 => x"ec",
          2542 => x"bb",
          2543 => x"05",
          2544 => x"dc",
          2545 => x"0d",
          2546 => x"0c",
          2547 => x"e8",
          2548 => x"bb",
          2549 => x"3d",
          2550 => x"82",
          2551 => x"f0",
          2552 => x"bb",
          2553 => x"05",
          2554 => x"73",
          2555 => x"e8",
          2556 => x"08",
          2557 => x"53",
          2558 => x"72",
          2559 => x"08",
          2560 => x"72",
          2561 => x"53",
          2562 => x"09",
          2563 => x"38",
          2564 => x"08",
          2565 => x"70",
          2566 => x"71",
          2567 => x"39",
          2568 => x"08",
          2569 => x"53",
          2570 => x"09",
          2571 => x"38",
          2572 => x"bb",
          2573 => x"05",
          2574 => x"e8",
          2575 => x"08",
          2576 => x"05",
          2577 => x"08",
          2578 => x"33",
          2579 => x"08",
          2580 => x"82",
          2581 => x"f8",
          2582 => x"72",
          2583 => x"81",
          2584 => x"38",
          2585 => x"08",
          2586 => x"70",
          2587 => x"71",
          2588 => x"51",
          2589 => x"82",
          2590 => x"f8",
          2591 => x"bb",
          2592 => x"05",
          2593 => x"e8",
          2594 => x"0c",
          2595 => x"08",
          2596 => x"80",
          2597 => x"38",
          2598 => x"08",
          2599 => x"80",
          2600 => x"38",
          2601 => x"90",
          2602 => x"e8",
          2603 => x"34",
          2604 => x"08",
          2605 => x"70",
          2606 => x"71",
          2607 => x"51",
          2608 => x"82",
          2609 => x"f8",
          2610 => x"a4",
          2611 => x"82",
          2612 => x"f4",
          2613 => x"bb",
          2614 => x"05",
          2615 => x"81",
          2616 => x"70",
          2617 => x"72",
          2618 => x"e8",
          2619 => x"34",
          2620 => x"82",
          2621 => x"f8",
          2622 => x"72",
          2623 => x"38",
          2624 => x"bb",
          2625 => x"05",
          2626 => x"39",
          2627 => x"08",
          2628 => x"53",
          2629 => x"90",
          2630 => x"e8",
          2631 => x"33",
          2632 => x"26",
          2633 => x"39",
          2634 => x"bb",
          2635 => x"05",
          2636 => x"39",
          2637 => x"bb",
          2638 => x"05",
          2639 => x"82",
          2640 => x"f8",
          2641 => x"af",
          2642 => x"38",
          2643 => x"08",
          2644 => x"53",
          2645 => x"83",
          2646 => x"80",
          2647 => x"e8",
          2648 => x"0c",
          2649 => x"8a",
          2650 => x"e8",
          2651 => x"34",
          2652 => x"bb",
          2653 => x"05",
          2654 => x"e8",
          2655 => x"33",
          2656 => x"27",
          2657 => x"82",
          2658 => x"f8",
          2659 => x"80",
          2660 => x"94",
          2661 => x"e8",
          2662 => x"33",
          2663 => x"53",
          2664 => x"e8",
          2665 => x"34",
          2666 => x"08",
          2667 => x"d0",
          2668 => x"72",
          2669 => x"08",
          2670 => x"82",
          2671 => x"f8",
          2672 => x"90",
          2673 => x"38",
          2674 => x"08",
          2675 => x"f9",
          2676 => x"72",
          2677 => x"08",
          2678 => x"82",
          2679 => x"f8",
          2680 => x"72",
          2681 => x"38",
          2682 => x"bb",
          2683 => x"05",
          2684 => x"39",
          2685 => x"08",
          2686 => x"82",
          2687 => x"f4",
          2688 => x"54",
          2689 => x"8d",
          2690 => x"82",
          2691 => x"ec",
          2692 => x"f7",
          2693 => x"e8",
          2694 => x"33",
          2695 => x"e8",
          2696 => x"08",
          2697 => x"e8",
          2698 => x"33",
          2699 => x"bb",
          2700 => x"05",
          2701 => x"e8",
          2702 => x"08",
          2703 => x"05",
          2704 => x"08",
          2705 => x"55",
          2706 => x"82",
          2707 => x"f8",
          2708 => x"a5",
          2709 => x"e8",
          2710 => x"33",
          2711 => x"2e",
          2712 => x"bb",
          2713 => x"05",
          2714 => x"bb",
          2715 => x"05",
          2716 => x"e8",
          2717 => x"08",
          2718 => x"08",
          2719 => x"71",
          2720 => x"0b",
          2721 => x"08",
          2722 => x"82",
          2723 => x"ec",
          2724 => x"bb",
          2725 => x"3d",
          2726 => x"e8",
          2727 => x"3d",
          2728 => x"08",
          2729 => x"58",
          2730 => x"80",
          2731 => x"39",
          2732 => x"e6",
          2733 => x"bb",
          2734 => x"78",
          2735 => x"33",
          2736 => x"39",
          2737 => x"73",
          2738 => x"81",
          2739 => x"81",
          2740 => x"39",
          2741 => x"90",
          2742 => x"dc",
          2743 => x"52",
          2744 => x"3f",
          2745 => x"08",
          2746 => x"75",
          2747 => x"a3",
          2748 => x"dc",
          2749 => x"84",
          2750 => x"73",
          2751 => x"b0",
          2752 => x"70",
          2753 => x"58",
          2754 => x"27",
          2755 => x"54",
          2756 => x"dc",
          2757 => x"0d",
          2758 => x"0d",
          2759 => x"93",
          2760 => x"38",
          2761 => x"82",
          2762 => x"52",
          2763 => x"82",
          2764 => x"81",
          2765 => x"9f",
          2766 => x"f9",
          2767 => x"84",
          2768 => x"39",
          2769 => x"51",
          2770 => x"82",
          2771 => x"80",
          2772 => x"a0",
          2773 => x"dd",
          2774 => x"c8",
          2775 => x"39",
          2776 => x"51",
          2777 => x"82",
          2778 => x"80",
          2779 => x"a1",
          2780 => x"c1",
          2781 => x"a0",
          2782 => x"82",
          2783 => x"b5",
          2784 => x"d0",
          2785 => x"82",
          2786 => x"a9",
          2787 => x"88",
          2788 => x"82",
          2789 => x"9d",
          2790 => x"b8",
          2791 => x"82",
          2792 => x"91",
          2793 => x"e8",
          2794 => x"82",
          2795 => x"85",
          2796 => x"8c",
          2797 => x"3f",
          2798 => x"04",
          2799 => x"77",
          2800 => x"74",
          2801 => x"8a",
          2802 => x"75",
          2803 => x"51",
          2804 => x"e8",
          2805 => x"ef",
          2806 => x"bb",
          2807 => x"75",
          2808 => x"3f",
          2809 => x"08",
          2810 => x"75",
          2811 => x"9c",
          2812 => x"e5",
          2813 => x"0d",
          2814 => x"0d",
          2815 => x"05",
          2816 => x"33",
          2817 => x"68",
          2818 => x"7a",
          2819 => x"51",
          2820 => x"78",
          2821 => x"ff",
          2822 => x"81",
          2823 => x"07",
          2824 => x"06",
          2825 => x"56",
          2826 => x"38",
          2827 => x"52",
          2828 => x"52",
          2829 => x"b9",
          2830 => x"dc",
          2831 => x"bb",
          2832 => x"38",
          2833 => x"08",
          2834 => x"88",
          2835 => x"dc",
          2836 => x"3d",
          2837 => x"84",
          2838 => x"52",
          2839 => x"88",
          2840 => x"bb",
          2841 => x"82",
          2842 => x"90",
          2843 => x"74",
          2844 => x"38",
          2845 => x"19",
          2846 => x"39",
          2847 => x"05",
          2848 => x"de",
          2849 => x"70",
          2850 => x"25",
          2851 => x"9f",
          2852 => x"51",
          2853 => x"74",
          2854 => x"38",
          2855 => x"53",
          2856 => x"88",
          2857 => x"51",
          2858 => x"76",
          2859 => x"bb",
          2860 => x"3d",
          2861 => x"3d",
          2862 => x"84",
          2863 => x"33",
          2864 => x"58",
          2865 => x"52",
          2866 => x"ad",
          2867 => x"dc",
          2868 => x"76",
          2869 => x"38",
          2870 => x"9c",
          2871 => x"82",
          2872 => x"61",
          2873 => x"82",
          2874 => x"7f",
          2875 => x"78",
          2876 => x"dc",
          2877 => x"39",
          2878 => x"82",
          2879 => x"8a",
          2880 => x"f3",
          2881 => x"61",
          2882 => x"05",
          2883 => x"33",
          2884 => x"68",
          2885 => x"5c",
          2886 => x"7a",
          2887 => x"c8",
          2888 => x"b5",
          2889 => x"d0",
          2890 => x"ad",
          2891 => x"74",
          2892 => x"80",
          2893 => x"2e",
          2894 => x"a0",
          2895 => x"80",
          2896 => x"18",
          2897 => x"27",
          2898 => x"22",
          2899 => x"d4",
          2900 => x"85",
          2901 => x"82",
          2902 => x"ff",
          2903 => x"82",
          2904 => x"c3",
          2905 => x"53",
          2906 => x"8e",
          2907 => x"52",
          2908 => x"51",
          2909 => x"3f",
          2910 => x"a3",
          2911 => x"b8",
          2912 => x"15",
          2913 => x"74",
          2914 => x"7a",
          2915 => x"72",
          2916 => x"a3",
          2917 => x"b8",
          2918 => x"39",
          2919 => x"51",
          2920 => x"3f",
          2921 => x"82",
          2922 => x"52",
          2923 => x"83",
          2924 => x"39",
          2925 => x"51",
          2926 => x"3f",
          2927 => x"79",
          2928 => x"38",
          2929 => x"33",
          2930 => x"56",
          2931 => x"83",
          2932 => x"80",
          2933 => x"27",
          2934 => x"53",
          2935 => x"70",
          2936 => x"51",
          2937 => x"2e",
          2938 => x"80",
          2939 => x"38",
          2940 => x"08",
          2941 => x"88",
          2942 => x"b0",
          2943 => x"51",
          2944 => x"81",
          2945 => x"b6",
          2946 => x"f8",
          2947 => x"3f",
          2948 => x"1c",
          2949 => x"fe",
          2950 => x"dc",
          2951 => x"70",
          2952 => x"57",
          2953 => x"09",
          2954 => x"38",
          2955 => x"82",
          2956 => x"98",
          2957 => x"2c",
          2958 => x"70",
          2959 => x"32",
          2960 => x"72",
          2961 => x"07",
          2962 => x"58",
          2963 => x"57",
          2964 => x"d8",
          2965 => x"2e",
          2966 => x"85",
          2967 => x"8c",
          2968 => x"53",
          2969 => x"fd",
          2970 => x"53",
          2971 => x"dc",
          2972 => x"0d",
          2973 => x"0d",
          2974 => x"33",
          2975 => x"53",
          2976 => x"52",
          2977 => x"d1",
          2978 => x"b4",
          2979 => x"d9",
          2980 => x"90",
          2981 => x"9c",
          2982 => x"b5",
          2983 => x"a4",
          2984 => x"b6",
          2985 => x"80",
          2986 => x"a5",
          2987 => x"3d",
          2988 => x"3d",
          2989 => x"96",
          2990 => x"aa",
          2991 => x"51",
          2992 => x"82",
          2993 => x"9d",
          2994 => x"51",
          2995 => x"72",
          2996 => x"81",
          2997 => x"71",
          2998 => x"38",
          2999 => x"a3",
          3000 => x"d8",
          3001 => x"3f",
          3002 => x"97",
          3003 => x"2a",
          3004 => x"51",
          3005 => x"2e",
          3006 => x"51",
          3007 => x"82",
          3008 => x"9d",
          3009 => x"51",
          3010 => x"72",
          3011 => x"81",
          3012 => x"71",
          3013 => x"38",
          3014 => x"e7",
          3015 => x"f8",
          3016 => x"3f",
          3017 => x"db",
          3018 => x"2a",
          3019 => x"51",
          3020 => x"2e",
          3021 => x"51",
          3022 => x"82",
          3023 => x"9c",
          3024 => x"51",
          3025 => x"72",
          3026 => x"81",
          3027 => x"71",
          3028 => x"38",
          3029 => x"ab",
          3030 => x"a0",
          3031 => x"3f",
          3032 => x"9f",
          3033 => x"2a",
          3034 => x"51",
          3035 => x"2e",
          3036 => x"51",
          3037 => x"82",
          3038 => x"9c",
          3039 => x"51",
          3040 => x"72",
          3041 => x"81",
          3042 => x"71",
          3043 => x"38",
          3044 => x"ef",
          3045 => x"c8",
          3046 => x"3f",
          3047 => x"e3",
          3048 => x"2a",
          3049 => x"51",
          3050 => x"2e",
          3051 => x"51",
          3052 => x"82",
          3053 => x"9b",
          3054 => x"51",
          3055 => x"a8",
          3056 => x"3d",
          3057 => x"3d",
          3058 => x"84",
          3059 => x"33",
          3060 => x"56",
          3061 => x"51",
          3062 => x"0b",
          3063 => x"d8",
          3064 => x"a9",
          3065 => x"82",
          3066 => x"82",
          3067 => x"80",
          3068 => x"82",
          3069 => x"30",
          3070 => x"dc",
          3071 => x"25",
          3072 => x"51",
          3073 => x"0b",
          3074 => x"d8",
          3075 => x"82",
          3076 => x"54",
          3077 => x"09",
          3078 => x"38",
          3079 => x"53",
          3080 => x"51",
          3081 => x"3f",
          3082 => x"08",
          3083 => x"38",
          3084 => x"08",
          3085 => x"3f",
          3086 => x"d2",
          3087 => x"89",
          3088 => x"0b",
          3089 => x"b6",
          3090 => x"0b",
          3091 => x"33",
          3092 => x"2e",
          3093 => x"8c",
          3094 => x"a8",
          3095 => x"75",
          3096 => x"3f",
          3097 => x"bb",
          3098 => x"3d",
          3099 => x"3d",
          3100 => x"71",
          3101 => x"0c",
          3102 => x"52",
          3103 => x"cb",
          3104 => x"bb",
          3105 => x"ff",
          3106 => x"7d",
          3107 => x"06",
          3108 => x"3d",
          3109 => x"82",
          3110 => x"78",
          3111 => x"3f",
          3112 => x"52",
          3113 => x"51",
          3114 => x"3f",
          3115 => x"08",
          3116 => x"38",
          3117 => x"51",
          3118 => x"81",
          3119 => x"82",
          3120 => x"ff",
          3121 => x"96",
          3122 => x"5a",
          3123 => x"79",
          3124 => x"3f",
          3125 => x"84",
          3126 => x"c2",
          3127 => x"dc",
          3128 => x"70",
          3129 => x"59",
          3130 => x"2e",
          3131 => x"78",
          3132 => x"80",
          3133 => x"ab",
          3134 => x"38",
          3135 => x"a4",
          3136 => x"2e",
          3137 => x"78",
          3138 => x"38",
          3139 => x"ff",
          3140 => x"80",
          3141 => x"2e",
          3142 => x"78",
          3143 => x"ad",
          3144 => x"39",
          3145 => x"84",
          3146 => x"bd",
          3147 => x"78",
          3148 => x"a6",
          3149 => x"2e",
          3150 => x"8e",
          3151 => x"bf",
          3152 => x"38",
          3153 => x"2e",
          3154 => x"8e",
          3155 => x"80",
          3156 => x"a0",
          3157 => x"d5",
          3158 => x"78",
          3159 => x"8c",
          3160 => x"80",
          3161 => x"38",
          3162 => x"2e",
          3163 => x"78",
          3164 => x"8b",
          3165 => x"9c",
          3166 => x"d1",
          3167 => x"38",
          3168 => x"2e",
          3169 => x"8e",
          3170 => x"81",
          3171 => x"e2",
          3172 => x"82",
          3173 => x"78",
          3174 => x"8c",
          3175 => x"80",
          3176 => x"91",
          3177 => x"39",
          3178 => x"2e",
          3179 => x"78",
          3180 => x"8d",
          3181 => x"dc",
          3182 => x"ff",
          3183 => x"ff",
          3184 => x"ec",
          3185 => x"bb",
          3186 => x"38",
          3187 => x"51",
          3188 => x"b4",
          3189 => x"11",
          3190 => x"05",
          3191 => x"3f",
          3192 => x"08",
          3193 => x"38",
          3194 => x"83",
          3195 => x"02",
          3196 => x"33",
          3197 => x"cf",
          3198 => x"80",
          3199 => x"82",
          3200 => x"81",
          3201 => x"78",
          3202 => x"a7",
          3203 => x"d4",
          3204 => x"fd",
          3205 => x"a7",
          3206 => x"f3",
          3207 => x"ff",
          3208 => x"ff",
          3209 => x"eb",
          3210 => x"bb",
          3211 => x"2e",
          3212 => x"80",
          3213 => x"02",
          3214 => x"33",
          3215 => x"d9",
          3216 => x"dc",
          3217 => x"a7",
          3218 => x"9f",
          3219 => x"ff",
          3220 => x"ff",
          3221 => x"ea",
          3222 => x"bb",
          3223 => x"2e",
          3224 => x"89",
          3225 => x"38",
          3226 => x"fc",
          3227 => x"84",
          3228 => x"d9",
          3229 => x"dc",
          3230 => x"82",
          3231 => x"43",
          3232 => x"a7",
          3233 => x"51",
          3234 => x"3f",
          3235 => x"05",
          3236 => x"52",
          3237 => x"29",
          3238 => x"05",
          3239 => x"f0",
          3240 => x"dc",
          3241 => x"38",
          3242 => x"51",
          3243 => x"81",
          3244 => x"39",
          3245 => x"84",
          3246 => x"c0",
          3247 => x"dc",
          3248 => x"ff",
          3249 => x"5b",
          3250 => x"81",
          3251 => x"dc",
          3252 => x"51",
          3253 => x"80",
          3254 => x"3d",
          3255 => x"51",
          3256 => x"82",
          3257 => x"b5",
          3258 => x"05",
          3259 => x"b0",
          3260 => x"dc",
          3261 => x"ff",
          3262 => x"5a",
          3263 => x"82",
          3264 => x"b5",
          3265 => x"05",
          3266 => x"94",
          3267 => x"80",
          3268 => x"8c",
          3269 => x"80",
          3270 => x"dc",
          3271 => x"06",
          3272 => x"79",
          3273 => x"f3",
          3274 => x"bb",
          3275 => x"2e",
          3276 => x"82",
          3277 => x"51",
          3278 => x"fb",
          3279 => x"3d",
          3280 => x"53",
          3281 => x"51",
          3282 => x"82",
          3283 => x"80",
          3284 => x"38",
          3285 => x"fc",
          3286 => x"84",
          3287 => x"ed",
          3288 => x"dc",
          3289 => x"fa",
          3290 => x"3d",
          3291 => x"53",
          3292 => x"51",
          3293 => x"82",
          3294 => x"86",
          3295 => x"dc",
          3296 => x"a7",
          3297 => x"ac",
          3298 => x"63",
          3299 => x"7b",
          3300 => x"38",
          3301 => x"7a",
          3302 => x"5c",
          3303 => x"26",
          3304 => x"db",
          3305 => x"ff",
          3306 => x"ff",
          3307 => x"e8",
          3308 => x"bb",
          3309 => x"2e",
          3310 => x"b4",
          3311 => x"11",
          3312 => x"05",
          3313 => x"3f",
          3314 => x"08",
          3315 => x"ef",
          3316 => x"fe",
          3317 => x"ff",
          3318 => x"e7",
          3319 => x"bb",
          3320 => x"2e",
          3321 => x"82",
          3322 => x"ff",
          3323 => x"63",
          3324 => x"27",
          3325 => x"61",
          3326 => x"81",
          3327 => x"79",
          3328 => x"05",
          3329 => x"b4",
          3330 => x"11",
          3331 => x"05",
          3332 => x"3f",
          3333 => x"08",
          3334 => x"a3",
          3335 => x"fe",
          3336 => x"ff",
          3337 => x"e7",
          3338 => x"bb",
          3339 => x"2e",
          3340 => x"b4",
          3341 => x"11",
          3342 => x"05",
          3343 => x"3f",
          3344 => x"08",
          3345 => x"f7",
          3346 => x"d4",
          3347 => x"89",
          3348 => x"79",
          3349 => x"38",
          3350 => x"7b",
          3351 => x"5b",
          3352 => x"92",
          3353 => x"7a",
          3354 => x"53",
          3355 => x"a7",
          3356 => x"aa",
          3357 => x"1a",
          3358 => x"43",
          3359 => x"8a",
          3360 => x"3f",
          3361 => x"b4",
          3362 => x"11",
          3363 => x"05",
          3364 => x"3f",
          3365 => x"08",
          3366 => x"82",
          3367 => x"59",
          3368 => x"89",
          3369 => x"80",
          3370 => x"cd",
          3371 => x"c9",
          3372 => x"80",
          3373 => x"82",
          3374 => x"44",
          3375 => x"ba",
          3376 => x"78",
          3377 => x"38",
          3378 => x"08",
          3379 => x"82",
          3380 => x"59",
          3381 => x"88",
          3382 => x"98",
          3383 => x"39",
          3384 => x"33",
          3385 => x"2e",
          3386 => x"ba",
          3387 => x"89",
          3388 => x"b0",
          3389 => x"05",
          3390 => x"fe",
          3391 => x"ff",
          3392 => x"e5",
          3393 => x"bb",
          3394 => x"de",
          3395 => x"c8",
          3396 => x"80",
          3397 => x"82",
          3398 => x"43",
          3399 => x"82",
          3400 => x"59",
          3401 => x"88",
          3402 => x"8c",
          3403 => x"39",
          3404 => x"33",
          3405 => x"2e",
          3406 => x"ba",
          3407 => x"aa",
          3408 => x"cb",
          3409 => x"80",
          3410 => x"82",
          3411 => x"43",
          3412 => x"ba",
          3413 => x"78",
          3414 => x"38",
          3415 => x"08",
          3416 => x"82",
          3417 => x"88",
          3418 => x"3d",
          3419 => x"53",
          3420 => x"51",
          3421 => x"82",
          3422 => x"80",
          3423 => x"80",
          3424 => x"7a",
          3425 => x"38",
          3426 => x"90",
          3427 => x"70",
          3428 => x"2a",
          3429 => x"51",
          3430 => x"78",
          3431 => x"38",
          3432 => x"83",
          3433 => x"82",
          3434 => x"c4",
          3435 => x"55",
          3436 => x"53",
          3437 => x"51",
          3438 => x"82",
          3439 => x"87",
          3440 => x"3d",
          3441 => x"53",
          3442 => x"51",
          3443 => x"82",
          3444 => x"80",
          3445 => x"38",
          3446 => x"fc",
          3447 => x"84",
          3448 => x"e9",
          3449 => x"dc",
          3450 => x"a4",
          3451 => x"02",
          3452 => x"33",
          3453 => x"81",
          3454 => x"3d",
          3455 => x"53",
          3456 => x"51",
          3457 => x"82",
          3458 => x"e1",
          3459 => x"39",
          3460 => x"54",
          3461 => x"98",
          3462 => x"bd",
          3463 => x"ac",
          3464 => x"f8",
          3465 => x"ff",
          3466 => x"79",
          3467 => x"59",
          3468 => x"f5",
          3469 => x"79",
          3470 => x"b4",
          3471 => x"11",
          3472 => x"05",
          3473 => x"3f",
          3474 => x"08",
          3475 => x"38",
          3476 => x"80",
          3477 => x"79",
          3478 => x"05",
          3479 => x"39",
          3480 => x"51",
          3481 => x"ff",
          3482 => x"3d",
          3483 => x"53",
          3484 => x"51",
          3485 => x"82",
          3486 => x"80",
          3487 => x"38",
          3488 => x"f0",
          3489 => x"84",
          3490 => x"f0",
          3491 => x"dc",
          3492 => x"a5",
          3493 => x"02",
          3494 => x"79",
          3495 => x"5b",
          3496 => x"b4",
          3497 => x"11",
          3498 => x"05",
          3499 => x"3f",
          3500 => x"08",
          3501 => x"87",
          3502 => x"22",
          3503 => x"a8",
          3504 => x"a6",
          3505 => x"d3",
          3506 => x"80",
          3507 => x"51",
          3508 => x"3f",
          3509 => x"33",
          3510 => x"2e",
          3511 => x"78",
          3512 => x"38",
          3513 => x"41",
          3514 => x"3d",
          3515 => x"53",
          3516 => x"51",
          3517 => x"82",
          3518 => x"80",
          3519 => x"60",
          3520 => x"05",
          3521 => x"82",
          3522 => x"78",
          3523 => x"39",
          3524 => x"51",
          3525 => x"ff",
          3526 => x"3d",
          3527 => x"53",
          3528 => x"51",
          3529 => x"82",
          3530 => x"80",
          3531 => x"38",
          3532 => x"f0",
          3533 => x"84",
          3534 => x"c0",
          3535 => x"dc",
          3536 => x"a0",
          3537 => x"71",
          3538 => x"84",
          3539 => x"3d",
          3540 => x"53",
          3541 => x"51",
          3542 => x"82",
          3543 => x"e5",
          3544 => x"39",
          3545 => x"54",
          3546 => x"b4",
          3547 => x"e9",
          3548 => x"ac",
          3549 => x"f8",
          3550 => x"ff",
          3551 => x"79",
          3552 => x"59",
          3553 => x"f2",
          3554 => x"79",
          3555 => x"b4",
          3556 => x"11",
          3557 => x"05",
          3558 => x"3f",
          3559 => x"08",
          3560 => x"38",
          3561 => x"0c",
          3562 => x"05",
          3563 => x"39",
          3564 => x"51",
          3565 => x"ff",
          3566 => x"a8",
          3567 => x"a4",
          3568 => x"98",
          3569 => x"f7",
          3570 => x"dc",
          3571 => x"3f",
          3572 => x"de",
          3573 => x"39",
          3574 => x"51",
          3575 => x"84",
          3576 => x"87",
          3577 => x"0c",
          3578 => x"0b",
          3579 => x"94",
          3580 => x"39",
          3581 => x"51",
          3582 => x"3f",
          3583 => x"0b",
          3584 => x"84",
          3585 => x"83",
          3586 => x"94",
          3587 => x"af",
          3588 => x"ff",
          3589 => x"ff",
          3590 => x"df",
          3591 => x"bb",
          3592 => x"2e",
          3593 => x"63",
          3594 => x"98",
          3595 => x"a9",
          3596 => x"78",
          3597 => x"ff",
          3598 => x"ff",
          3599 => x"df",
          3600 => x"bb",
          3601 => x"2e",
          3602 => x"63",
          3603 => x"b4",
          3604 => x"85",
          3605 => x"78",
          3606 => x"dc",
          3607 => x"f0",
          3608 => x"bb",
          3609 => x"82",
          3610 => x"ff",
          3611 => x"f0",
          3612 => x"a9",
          3613 => x"be",
          3614 => x"a2",
          3615 => x"bf",
          3616 => x"88",
          3617 => x"dc",
          3618 => x"ff",
          3619 => x"a8",
          3620 => x"39",
          3621 => x"33",
          3622 => x"2e",
          3623 => x"7d",
          3624 => x"78",
          3625 => x"cf",
          3626 => x"ff",
          3627 => x"83",
          3628 => x"bb",
          3629 => x"81",
          3630 => x"2e",
          3631 => x"82",
          3632 => x"7b",
          3633 => x"38",
          3634 => x"7b",
          3635 => x"38",
          3636 => x"82",
          3637 => x"7a",
          3638 => x"a0",
          3639 => x"82",
          3640 => x"b4",
          3641 => x"05",
          3642 => x"d5",
          3643 => x"7a",
          3644 => x"ff",
          3645 => x"ca",
          3646 => x"39",
          3647 => x"aa",
          3648 => x"53",
          3649 => x"52",
          3650 => x"b0",
          3651 => x"a4",
          3652 => x"39",
          3653 => x"53",
          3654 => x"52",
          3655 => x"b0",
          3656 => x"a4",
          3657 => x"ba",
          3658 => x"bc",
          3659 => x"56",
          3660 => x"54",
          3661 => x"53",
          3662 => x"52",
          3663 => x"b0",
          3664 => x"f2",
          3665 => x"dc",
          3666 => x"dc",
          3667 => x"30",
          3668 => x"80",
          3669 => x"5b",
          3670 => x"7b",
          3671 => x"38",
          3672 => x"7a",
          3673 => x"80",
          3674 => x"81",
          3675 => x"ff",
          3676 => x"7b",
          3677 => x"7d",
          3678 => x"81",
          3679 => x"78",
          3680 => x"ff",
          3681 => x"06",
          3682 => x"82",
          3683 => x"ff",
          3684 => x"ee",
          3685 => x"3d",
          3686 => x"82",
          3687 => x"87",
          3688 => x"70",
          3689 => x"87",
          3690 => x"72",
          3691 => x"3f",
          3692 => x"08",
          3693 => x"08",
          3694 => x"84",
          3695 => x"51",
          3696 => x"72",
          3697 => x"08",
          3698 => x"87",
          3699 => x"70",
          3700 => x"87",
          3701 => x"72",
          3702 => x"3f",
          3703 => x"08",
          3704 => x"08",
          3705 => x"84",
          3706 => x"51",
          3707 => x"72",
          3708 => x"08",
          3709 => x"8c",
          3710 => x"87",
          3711 => x"0c",
          3712 => x"0b",
          3713 => x"94",
          3714 => x"9a",
          3715 => x"86",
          3716 => x"84",
          3717 => x"34",
          3718 => x"d3",
          3719 => x"3d",
          3720 => x"0c",
          3721 => x"82",
          3722 => x"54",
          3723 => x"93",
          3724 => x"aa",
          3725 => x"bb",
          3726 => x"aa",
          3727 => x"bb",
          3728 => x"dd",
          3729 => x"e5",
          3730 => x"e8",
          3731 => x"9e",
          3732 => x"fe",
          3733 => x"52",
          3734 => x"88",
          3735 => x"d8",
          3736 => x"dc",
          3737 => x"06",
          3738 => x"14",
          3739 => x"80",
          3740 => x"71",
          3741 => x"0c",
          3742 => x"04",
          3743 => x"76",
          3744 => x"55",
          3745 => x"54",
          3746 => x"81",
          3747 => x"33",
          3748 => x"2e",
          3749 => x"86",
          3750 => x"53",
          3751 => x"33",
          3752 => x"2e",
          3753 => x"86",
          3754 => x"53",
          3755 => x"52",
          3756 => x"09",
          3757 => x"38",
          3758 => x"12",
          3759 => x"33",
          3760 => x"a2",
          3761 => x"81",
          3762 => x"2e",
          3763 => x"ea",
          3764 => x"81",
          3765 => x"72",
          3766 => x"70",
          3767 => x"38",
          3768 => x"80",
          3769 => x"73",
          3770 => x"72",
          3771 => x"70",
          3772 => x"81",
          3773 => x"81",
          3774 => x"32",
          3775 => x"80",
          3776 => x"51",
          3777 => x"80",
          3778 => x"80",
          3779 => x"05",
          3780 => x"75",
          3781 => x"70",
          3782 => x"0c",
          3783 => x"04",
          3784 => x"76",
          3785 => x"80",
          3786 => x"86",
          3787 => x"52",
          3788 => x"c8",
          3789 => x"dc",
          3790 => x"80",
          3791 => x"74",
          3792 => x"bb",
          3793 => x"3d",
          3794 => x"3d",
          3795 => x"11",
          3796 => x"52",
          3797 => x"70",
          3798 => x"98",
          3799 => x"33",
          3800 => x"82",
          3801 => x"26",
          3802 => x"84",
          3803 => x"83",
          3804 => x"26",
          3805 => x"85",
          3806 => x"84",
          3807 => x"26",
          3808 => x"86",
          3809 => x"85",
          3810 => x"26",
          3811 => x"88",
          3812 => x"86",
          3813 => x"e7",
          3814 => x"38",
          3815 => x"54",
          3816 => x"87",
          3817 => x"cc",
          3818 => x"87",
          3819 => x"0c",
          3820 => x"c0",
          3821 => x"82",
          3822 => x"c0",
          3823 => x"83",
          3824 => x"c0",
          3825 => x"84",
          3826 => x"c0",
          3827 => x"85",
          3828 => x"c0",
          3829 => x"86",
          3830 => x"c0",
          3831 => x"74",
          3832 => x"a4",
          3833 => x"c0",
          3834 => x"80",
          3835 => x"98",
          3836 => x"52",
          3837 => x"dc",
          3838 => x"0d",
          3839 => x"0d",
          3840 => x"c0",
          3841 => x"81",
          3842 => x"c0",
          3843 => x"5e",
          3844 => x"87",
          3845 => x"08",
          3846 => x"1c",
          3847 => x"98",
          3848 => x"79",
          3849 => x"87",
          3850 => x"08",
          3851 => x"1c",
          3852 => x"98",
          3853 => x"79",
          3854 => x"87",
          3855 => x"08",
          3856 => x"1c",
          3857 => x"98",
          3858 => x"7b",
          3859 => x"87",
          3860 => x"08",
          3861 => x"1c",
          3862 => x"0c",
          3863 => x"ff",
          3864 => x"83",
          3865 => x"58",
          3866 => x"57",
          3867 => x"56",
          3868 => x"55",
          3869 => x"54",
          3870 => x"53",
          3871 => x"ff",
          3872 => x"aa",
          3873 => x"9a",
          3874 => x"3d",
          3875 => x"3d",
          3876 => x"05",
          3877 => x"fc",
          3878 => x"ff",
          3879 => x"55",
          3880 => x"84",
          3881 => x"2e",
          3882 => x"c0",
          3883 => x"70",
          3884 => x"2a",
          3885 => x"53",
          3886 => x"80",
          3887 => x"71",
          3888 => x"81",
          3889 => x"70",
          3890 => x"81",
          3891 => x"06",
          3892 => x"80",
          3893 => x"71",
          3894 => x"81",
          3895 => x"70",
          3896 => x"73",
          3897 => x"51",
          3898 => x"80",
          3899 => x"2e",
          3900 => x"c0",
          3901 => x"74",
          3902 => x"82",
          3903 => x"87",
          3904 => x"ff",
          3905 => x"8f",
          3906 => x"30",
          3907 => x"51",
          3908 => x"82",
          3909 => x"83",
          3910 => x"f9",
          3911 => x"a7",
          3912 => x"77",
          3913 => x"81",
          3914 => x"7a",
          3915 => x"eb",
          3916 => x"fc",
          3917 => x"ff",
          3918 => x"87",
          3919 => x"53",
          3920 => x"86",
          3921 => x"94",
          3922 => x"08",
          3923 => x"70",
          3924 => x"56",
          3925 => x"2e",
          3926 => x"91",
          3927 => x"06",
          3928 => x"d7",
          3929 => x"32",
          3930 => x"51",
          3931 => x"2e",
          3932 => x"93",
          3933 => x"06",
          3934 => x"ff",
          3935 => x"81",
          3936 => x"87",
          3937 => x"54",
          3938 => x"86",
          3939 => x"94",
          3940 => x"74",
          3941 => x"82",
          3942 => x"89",
          3943 => x"f9",
          3944 => x"54",
          3945 => x"70",
          3946 => x"53",
          3947 => x"77",
          3948 => x"38",
          3949 => x"06",
          3950 => x"b9",
          3951 => x"81",
          3952 => x"57",
          3953 => x"c0",
          3954 => x"75",
          3955 => x"38",
          3956 => x"94",
          3957 => x"70",
          3958 => x"81",
          3959 => x"52",
          3960 => x"8c",
          3961 => x"2a",
          3962 => x"51",
          3963 => x"38",
          3964 => x"70",
          3965 => x"51",
          3966 => x"8d",
          3967 => x"2a",
          3968 => x"51",
          3969 => x"be",
          3970 => x"ff",
          3971 => x"c0",
          3972 => x"70",
          3973 => x"38",
          3974 => x"90",
          3975 => x"0c",
          3976 => x"33",
          3977 => x"06",
          3978 => x"70",
          3979 => x"76",
          3980 => x"0c",
          3981 => x"04",
          3982 => x"82",
          3983 => x"70",
          3984 => x"54",
          3985 => x"94",
          3986 => x"80",
          3987 => x"87",
          3988 => x"51",
          3989 => x"82",
          3990 => x"06",
          3991 => x"70",
          3992 => x"38",
          3993 => x"06",
          3994 => x"94",
          3995 => x"80",
          3996 => x"87",
          3997 => x"52",
          3998 => x"81",
          3999 => x"bb",
          4000 => x"84",
          4001 => x"ff",
          4002 => x"bb",
          4003 => x"ff",
          4004 => x"dc",
          4005 => x"3d",
          4006 => x"fc",
          4007 => x"ff",
          4008 => x"87",
          4009 => x"52",
          4010 => x"86",
          4011 => x"94",
          4012 => x"08",
          4013 => x"70",
          4014 => x"51",
          4015 => x"70",
          4016 => x"38",
          4017 => x"06",
          4018 => x"94",
          4019 => x"80",
          4020 => x"87",
          4021 => x"52",
          4022 => x"98",
          4023 => x"2c",
          4024 => x"71",
          4025 => x"0c",
          4026 => x"04",
          4027 => x"87",
          4028 => x"08",
          4029 => x"8a",
          4030 => x"70",
          4031 => x"b4",
          4032 => x"9e",
          4033 => x"ba",
          4034 => x"c0",
          4035 => x"82",
          4036 => x"87",
          4037 => x"08",
          4038 => x"0c",
          4039 => x"98",
          4040 => x"8c",
          4041 => x"9e",
          4042 => x"ba",
          4043 => x"c0",
          4044 => x"82",
          4045 => x"87",
          4046 => x"08",
          4047 => x"0c",
          4048 => x"b0",
          4049 => x"9c",
          4050 => x"9e",
          4051 => x"ba",
          4052 => x"c0",
          4053 => x"82",
          4054 => x"87",
          4055 => x"08",
          4056 => x"0c",
          4057 => x"c0",
          4058 => x"ac",
          4059 => x"9e",
          4060 => x"ba",
          4061 => x"c0",
          4062 => x"51",
          4063 => x"b4",
          4064 => x"9e",
          4065 => x"ba",
          4066 => x"c0",
          4067 => x"82",
          4068 => x"87",
          4069 => x"08",
          4070 => x"0c",
          4071 => x"ba",
          4072 => x"0b",
          4073 => x"90",
          4074 => x"80",
          4075 => x"52",
          4076 => x"2e",
          4077 => x"52",
          4078 => x"c5",
          4079 => x"87",
          4080 => x"08",
          4081 => x"0a",
          4082 => x"52",
          4083 => x"83",
          4084 => x"71",
          4085 => x"34",
          4086 => x"c0",
          4087 => x"70",
          4088 => x"06",
          4089 => x"70",
          4090 => x"38",
          4091 => x"82",
          4092 => x"80",
          4093 => x"9e",
          4094 => x"88",
          4095 => x"51",
          4096 => x"80",
          4097 => x"81",
          4098 => x"ba",
          4099 => x"0b",
          4100 => x"90",
          4101 => x"80",
          4102 => x"52",
          4103 => x"2e",
          4104 => x"52",
          4105 => x"c9",
          4106 => x"87",
          4107 => x"08",
          4108 => x"80",
          4109 => x"52",
          4110 => x"83",
          4111 => x"71",
          4112 => x"34",
          4113 => x"c0",
          4114 => x"70",
          4115 => x"06",
          4116 => x"70",
          4117 => x"38",
          4118 => x"82",
          4119 => x"80",
          4120 => x"9e",
          4121 => x"82",
          4122 => x"51",
          4123 => x"80",
          4124 => x"81",
          4125 => x"ba",
          4126 => x"0b",
          4127 => x"90",
          4128 => x"80",
          4129 => x"52",
          4130 => x"2e",
          4131 => x"52",
          4132 => x"cd",
          4133 => x"87",
          4134 => x"08",
          4135 => x"80",
          4136 => x"52",
          4137 => x"83",
          4138 => x"71",
          4139 => x"34",
          4140 => x"c0",
          4141 => x"70",
          4142 => x"51",
          4143 => x"80",
          4144 => x"81",
          4145 => x"ba",
          4146 => x"c0",
          4147 => x"70",
          4148 => x"70",
          4149 => x"51",
          4150 => x"ba",
          4151 => x"0b",
          4152 => x"90",
          4153 => x"80",
          4154 => x"52",
          4155 => x"83",
          4156 => x"71",
          4157 => x"34",
          4158 => x"90",
          4159 => x"f0",
          4160 => x"2a",
          4161 => x"70",
          4162 => x"34",
          4163 => x"c0",
          4164 => x"70",
          4165 => x"52",
          4166 => x"2e",
          4167 => x"52",
          4168 => x"d3",
          4169 => x"9e",
          4170 => x"87",
          4171 => x"70",
          4172 => x"34",
          4173 => x"04",
          4174 => x"82",
          4175 => x"ff",
          4176 => x"82",
          4177 => x"54",
          4178 => x"89",
          4179 => x"a8",
          4180 => x"90",
          4181 => x"bc",
          4182 => x"88",
          4183 => x"c6",
          4184 => x"80",
          4185 => x"82",
          4186 => x"82",
          4187 => x"11",
          4188 => x"ab",
          4189 => x"90",
          4190 => x"ba",
          4191 => x"73",
          4192 => x"38",
          4193 => x"08",
          4194 => x"08",
          4195 => x"82",
          4196 => x"ff",
          4197 => x"82",
          4198 => x"54",
          4199 => x"94",
          4200 => x"80",
          4201 => x"84",
          4202 => x"52",
          4203 => x"51",
          4204 => x"3f",
          4205 => x"33",
          4206 => x"2e",
          4207 => x"ba",
          4208 => x"ba",
          4209 => x"54",
          4210 => x"a8",
          4211 => x"89",
          4212 => x"ca",
          4213 => x"80",
          4214 => x"82",
          4215 => x"82",
          4216 => x"11",
          4217 => x"ac",
          4218 => x"8f",
          4219 => x"ba",
          4220 => x"73",
          4221 => x"38",
          4222 => x"33",
          4223 => x"e0",
          4224 => x"d5",
          4225 => x"d3",
          4226 => x"80",
          4227 => x"82",
          4228 => x"52",
          4229 => x"51",
          4230 => x"3f",
          4231 => x"33",
          4232 => x"2e",
          4233 => x"ba",
          4234 => x"82",
          4235 => x"ff",
          4236 => x"82",
          4237 => x"54",
          4238 => x"89",
          4239 => x"c0",
          4240 => x"a0",
          4241 => x"c7",
          4242 => x"80",
          4243 => x"82",
          4244 => x"ff",
          4245 => x"82",
          4246 => x"54",
          4247 => x"89",
          4248 => x"e0",
          4249 => x"fc",
          4250 => x"cd",
          4251 => x"80",
          4252 => x"82",
          4253 => x"ff",
          4254 => x"82",
          4255 => x"54",
          4256 => x"89",
          4257 => x"f8",
          4258 => x"d8",
          4259 => x"84",
          4260 => x"d0",
          4261 => x"a8",
          4262 => x"ae",
          4263 => x"8e",
          4264 => x"ba",
          4265 => x"82",
          4266 => x"ff",
          4267 => x"82",
          4268 => x"52",
          4269 => x"51",
          4270 => x"3f",
          4271 => x"51",
          4272 => x"3f",
          4273 => x"22",
          4274 => x"90",
          4275 => x"89",
          4276 => x"b8",
          4277 => x"84",
          4278 => x"51",
          4279 => x"82",
          4280 => x"bd",
          4281 => x"76",
          4282 => x"54",
          4283 => x"08",
          4284 => x"b8",
          4285 => x"e1",
          4286 => x"cb",
          4287 => x"80",
          4288 => x"82",
          4289 => x"56",
          4290 => x"52",
          4291 => x"f4",
          4292 => x"dc",
          4293 => x"c0",
          4294 => x"31",
          4295 => x"bb",
          4296 => x"82",
          4297 => x"ff",
          4298 => x"82",
          4299 => x"54",
          4300 => x"a9",
          4301 => x"c0",
          4302 => x"84",
          4303 => x"51",
          4304 => x"82",
          4305 => x"bd",
          4306 => x"76",
          4307 => x"54",
          4308 => x"08",
          4309 => x"90",
          4310 => x"fd",
          4311 => x"fc",
          4312 => x"80",
          4313 => x"0d",
          4314 => x"0d",
          4315 => x"33",
          4316 => x"71",
          4317 => x"38",
          4318 => x"82",
          4319 => x"52",
          4320 => x"82",
          4321 => x"9d",
          4322 => x"c4",
          4323 => x"82",
          4324 => x"91",
          4325 => x"d4",
          4326 => x"82",
          4327 => x"85",
          4328 => x"e0",
          4329 => x"bc",
          4330 => x"0d",
          4331 => x"80",
          4332 => x"3d",
          4333 => x"96",
          4334 => x"52",
          4335 => x"0c",
          4336 => x"70",
          4337 => x"0c",
          4338 => x"3d",
          4339 => x"3d",
          4340 => x"96",
          4341 => x"82",
          4342 => x"52",
          4343 => x"73",
          4344 => x"ba",
          4345 => x"70",
          4346 => x"0c",
          4347 => x"83",
          4348 => x"80",
          4349 => x"96",
          4350 => x"82",
          4351 => x"87",
          4352 => x"0c",
          4353 => x"0d",
          4354 => x"70",
          4355 => x"98",
          4356 => x"2c",
          4357 => x"70",
          4358 => x"53",
          4359 => x"51",
          4360 => x"b0",
          4361 => x"55",
          4362 => x"25",
          4363 => x"b0",
          4364 => x"12",
          4365 => x"97",
          4366 => x"33",
          4367 => x"70",
          4368 => x"81",
          4369 => x"81",
          4370 => x"bb",
          4371 => x"3d",
          4372 => x"3d",
          4373 => x"84",
          4374 => x"33",
          4375 => x"56",
          4376 => x"2e",
          4377 => x"d3",
          4378 => x"88",
          4379 => x"c3",
          4380 => x"b0",
          4381 => x"51",
          4382 => x"3f",
          4383 => x"08",
          4384 => x"ff",
          4385 => x"73",
          4386 => x"53",
          4387 => x"72",
          4388 => x"53",
          4389 => x"51",
          4390 => x"3f",
          4391 => x"87",
          4392 => x"f6",
          4393 => x"02",
          4394 => x"05",
          4395 => x"05",
          4396 => x"82",
          4397 => x"70",
          4398 => x"ba",
          4399 => x"08",
          4400 => x"5a",
          4401 => x"80",
          4402 => x"74",
          4403 => x"3f",
          4404 => x"33",
          4405 => x"82",
          4406 => x"81",
          4407 => x"58",
          4408 => x"fb",
          4409 => x"dc",
          4410 => x"82",
          4411 => x"70",
          4412 => x"ba",
          4413 => x"08",
          4414 => x"74",
          4415 => x"38",
          4416 => x"52",
          4417 => x"b3",
          4418 => x"bb",
          4419 => x"05",
          4420 => x"bb",
          4421 => x"81",
          4422 => x"93",
          4423 => x"38",
          4424 => x"bb",
          4425 => x"80",
          4426 => x"82",
          4427 => x"56",
          4428 => x"ac",
          4429 => x"ac",
          4430 => x"a4",
          4431 => x"fc",
          4432 => x"53",
          4433 => x"51",
          4434 => x"3f",
          4435 => x"08",
          4436 => x"81",
          4437 => x"82",
          4438 => x"51",
          4439 => x"3f",
          4440 => x"04",
          4441 => x"82",
          4442 => x"93",
          4443 => x"52",
          4444 => x"89",
          4445 => x"99",
          4446 => x"73",
          4447 => x"84",
          4448 => x"73",
          4449 => x"38",
          4450 => x"bb",
          4451 => x"bb",
          4452 => x"71",
          4453 => x"38",
          4454 => x"de",
          4455 => x"bb",
          4456 => x"99",
          4457 => x"0b",
          4458 => x"0c",
          4459 => x"04",
          4460 => x"81",
          4461 => x"82",
          4462 => x"51",
          4463 => x"3f",
          4464 => x"08",
          4465 => x"82",
          4466 => x"53",
          4467 => x"88",
          4468 => x"56",
          4469 => x"3f",
          4470 => x"08",
          4471 => x"38",
          4472 => x"b0",
          4473 => x"bb",
          4474 => x"80",
          4475 => x"dc",
          4476 => x"38",
          4477 => x"08",
          4478 => x"17",
          4479 => x"74",
          4480 => x"76",
          4481 => x"82",
          4482 => x"57",
          4483 => x"3f",
          4484 => x"09",
          4485 => x"af",
          4486 => x"0d",
          4487 => x"0d",
          4488 => x"ad",
          4489 => x"5a",
          4490 => x"58",
          4491 => x"bb",
          4492 => x"80",
          4493 => x"82",
          4494 => x"81",
          4495 => x"0b",
          4496 => x"08",
          4497 => x"f8",
          4498 => x"70",
          4499 => x"8b",
          4500 => x"bb",
          4501 => x"2e",
          4502 => x"51",
          4503 => x"3f",
          4504 => x"08",
          4505 => x"55",
          4506 => x"bb",
          4507 => x"8e",
          4508 => x"dc",
          4509 => x"70",
          4510 => x"80",
          4511 => x"09",
          4512 => x"72",
          4513 => x"51",
          4514 => x"77",
          4515 => x"73",
          4516 => x"82",
          4517 => x"8c",
          4518 => x"51",
          4519 => x"3f",
          4520 => x"08",
          4521 => x"38",
          4522 => x"51",
          4523 => x"3f",
          4524 => x"09",
          4525 => x"38",
          4526 => x"51",
          4527 => x"3f",
          4528 => x"ae",
          4529 => x"3d",
          4530 => x"bb",
          4531 => x"34",
          4532 => x"82",
          4533 => x"a9",
          4534 => x"f6",
          4535 => x"7e",
          4536 => x"72",
          4537 => x"5a",
          4538 => x"2e",
          4539 => x"a2",
          4540 => x"78",
          4541 => x"76",
          4542 => x"81",
          4543 => x"70",
          4544 => x"58",
          4545 => x"2e",
          4546 => x"86",
          4547 => x"26",
          4548 => x"54",
          4549 => x"82",
          4550 => x"70",
          4551 => x"ff",
          4552 => x"82",
          4553 => x"53",
          4554 => x"08",
          4555 => x"e3",
          4556 => x"dc",
          4557 => x"38",
          4558 => x"55",
          4559 => x"88",
          4560 => x"2e",
          4561 => x"39",
          4562 => x"ac",
          4563 => x"5a",
          4564 => x"11",
          4565 => x"51",
          4566 => x"82",
          4567 => x"80",
          4568 => x"ff",
          4569 => x"52",
          4570 => x"b1",
          4571 => x"dc",
          4572 => x"06",
          4573 => x"38",
          4574 => x"39",
          4575 => x"81",
          4576 => x"54",
          4577 => x"ff",
          4578 => x"54",
          4579 => x"dc",
          4580 => x"0d",
          4581 => x"0d",
          4582 => x"b2",
          4583 => x"3d",
          4584 => x"5a",
          4585 => x"3d",
          4586 => x"b4",
          4587 => x"b0",
          4588 => x"73",
          4589 => x"73",
          4590 => x"33",
          4591 => x"83",
          4592 => x"76",
          4593 => x"bc",
          4594 => x"76",
          4595 => x"73",
          4596 => x"ad",
          4597 => x"98",
          4598 => x"bb",
          4599 => x"bb",
          4600 => x"bb",
          4601 => x"2e",
          4602 => x"93",
          4603 => x"82",
          4604 => x"51",
          4605 => x"3f",
          4606 => x"08",
          4607 => x"38",
          4608 => x"51",
          4609 => x"3f",
          4610 => x"82",
          4611 => x"5b",
          4612 => x"08",
          4613 => x"52",
          4614 => x"52",
          4615 => x"b7",
          4616 => x"dc",
          4617 => x"bb",
          4618 => x"2e",
          4619 => x"80",
          4620 => x"bb",
          4621 => x"ff",
          4622 => x"82",
          4623 => x"55",
          4624 => x"bb",
          4625 => x"a9",
          4626 => x"dc",
          4627 => x"70",
          4628 => x"80",
          4629 => x"53",
          4630 => x"06",
          4631 => x"f8",
          4632 => x"1b",
          4633 => x"06",
          4634 => x"7b",
          4635 => x"80",
          4636 => x"2e",
          4637 => x"ff",
          4638 => x"39",
          4639 => x"ac",
          4640 => x"38",
          4641 => x"08",
          4642 => x"38",
          4643 => x"8f",
          4644 => x"82",
          4645 => x"dc",
          4646 => x"70",
          4647 => x"59",
          4648 => x"ee",
          4649 => x"ff",
          4650 => x"88",
          4651 => x"2b",
          4652 => x"82",
          4653 => x"70",
          4654 => x"97",
          4655 => x"2c",
          4656 => x"29",
          4657 => x"05",
          4658 => x"70",
          4659 => x"51",
          4660 => x"51",
          4661 => x"81",
          4662 => x"2e",
          4663 => x"77",
          4664 => x"38",
          4665 => x"0a",
          4666 => x"0a",
          4667 => x"2c",
          4668 => x"75",
          4669 => x"38",
          4670 => x"52",
          4671 => x"85",
          4672 => x"dc",
          4673 => x"06",
          4674 => x"2e",
          4675 => x"82",
          4676 => x"81",
          4677 => x"74",
          4678 => x"29",
          4679 => x"05",
          4680 => x"70",
          4681 => x"56",
          4682 => x"95",
          4683 => x"76",
          4684 => x"77",
          4685 => x"3f",
          4686 => x"08",
          4687 => x"54",
          4688 => x"d3",
          4689 => x"75",
          4690 => x"ca",
          4691 => x"55",
          4692 => x"88",
          4693 => x"2b",
          4694 => x"82",
          4695 => x"70",
          4696 => x"98",
          4697 => x"11",
          4698 => x"82",
          4699 => x"33",
          4700 => x"51",
          4701 => x"55",
          4702 => x"09",
          4703 => x"92",
          4704 => x"f0",
          4705 => x"0c",
          4706 => x"d3",
          4707 => x"0b",
          4708 => x"34",
          4709 => x"82",
          4710 => x"75",
          4711 => x"34",
          4712 => x"34",
          4713 => x"7e",
          4714 => x"26",
          4715 => x"73",
          4716 => x"9b",
          4717 => x"73",
          4718 => x"d3",
          4719 => x"73",
          4720 => x"cb",
          4721 => x"8c",
          4722 => x"75",
          4723 => x"74",
          4724 => x"98",
          4725 => x"73",
          4726 => x"38",
          4727 => x"73",
          4728 => x"34",
          4729 => x"0a",
          4730 => x"0a",
          4731 => x"2c",
          4732 => x"33",
          4733 => x"df",
          4734 => x"90",
          4735 => x"56",
          4736 => x"d3",
          4737 => x"1a",
          4738 => x"33",
          4739 => x"d3",
          4740 => x"73",
          4741 => x"38",
          4742 => x"73",
          4743 => x"34",
          4744 => x"33",
          4745 => x"0a",
          4746 => x"0a",
          4747 => x"2c",
          4748 => x"33",
          4749 => x"56",
          4750 => x"a8",
          4751 => x"b0",
          4752 => x"1a",
          4753 => x"54",
          4754 => x"3f",
          4755 => x"0a",
          4756 => x"0a",
          4757 => x"2c",
          4758 => x"33",
          4759 => x"73",
          4760 => x"38",
          4761 => x"33",
          4762 => x"70",
          4763 => x"d3",
          4764 => x"51",
          4765 => x"77",
          4766 => x"38",
          4767 => x"08",
          4768 => x"ff",
          4769 => x"74",
          4770 => x"29",
          4771 => x"05",
          4772 => x"82",
          4773 => x"56",
          4774 => x"75",
          4775 => x"fb",
          4776 => x"7a",
          4777 => x"81",
          4778 => x"d3",
          4779 => x"52",
          4780 => x"51",
          4781 => x"81",
          4782 => x"d3",
          4783 => x"81",
          4784 => x"55",
          4785 => x"fb",
          4786 => x"d3",
          4787 => x"05",
          4788 => x"d3",
          4789 => x"15",
          4790 => x"d3",
          4791 => x"d3",
          4792 => x"88",
          4793 => x"cb",
          4794 => x"90",
          4795 => x"2b",
          4796 => x"82",
          4797 => x"57",
          4798 => x"74",
          4799 => x"38",
          4800 => x"81",
          4801 => x"34",
          4802 => x"08",
          4803 => x"51",
          4804 => x"3f",
          4805 => x"0a",
          4806 => x"0a",
          4807 => x"2c",
          4808 => x"33",
          4809 => x"75",
          4810 => x"38",
          4811 => x"08",
          4812 => x"ff",
          4813 => x"82",
          4814 => x"70",
          4815 => x"98",
          4816 => x"8c",
          4817 => x"56",
          4818 => x"24",
          4819 => x"82",
          4820 => x"52",
          4821 => x"9c",
          4822 => x"81",
          4823 => x"81",
          4824 => x"70",
          4825 => x"d3",
          4826 => x"51",
          4827 => x"25",
          4828 => x"9b",
          4829 => x"8c",
          4830 => x"54",
          4831 => x"82",
          4832 => x"52",
          4833 => x"9c",
          4834 => x"d3",
          4835 => x"51",
          4836 => x"82",
          4837 => x"81",
          4838 => x"73",
          4839 => x"d3",
          4840 => x"73",
          4841 => x"38",
          4842 => x"52",
          4843 => x"f3",
          4844 => x"80",
          4845 => x"0b",
          4846 => x"34",
          4847 => x"d3",
          4848 => x"82",
          4849 => x"af",
          4850 => x"82",
          4851 => x"54",
          4852 => x"f9",
          4853 => x"d3",
          4854 => x"88",
          4855 => x"d3",
          4856 => x"90",
          4857 => x"54",
          4858 => x"90",
          4859 => x"ff",
          4860 => x"39",
          4861 => x"33",
          4862 => x"33",
          4863 => x"75",
          4864 => x"38",
          4865 => x"73",
          4866 => x"34",
          4867 => x"70",
          4868 => x"81",
          4869 => x"51",
          4870 => x"25",
          4871 => x"1a",
          4872 => x"33",
          4873 => x"d3",
          4874 => x"73",
          4875 => x"9b",
          4876 => x"81",
          4877 => x"81",
          4878 => x"70",
          4879 => x"d3",
          4880 => x"51",
          4881 => x"24",
          4882 => x"d3",
          4883 => x"a0",
          4884 => x"df",
          4885 => x"90",
          4886 => x"2b",
          4887 => x"82",
          4888 => x"57",
          4889 => x"74",
          4890 => x"a3",
          4891 => x"b0",
          4892 => x"51",
          4893 => x"3f",
          4894 => x"0a",
          4895 => x"0a",
          4896 => x"2c",
          4897 => x"33",
          4898 => x"75",
          4899 => x"38",
          4900 => x"82",
          4901 => x"70",
          4902 => x"82",
          4903 => x"59",
          4904 => x"77",
          4905 => x"38",
          4906 => x"08",
          4907 => x"54",
          4908 => x"90",
          4909 => x"70",
          4910 => x"ff",
          4911 => x"82",
          4912 => x"70",
          4913 => x"82",
          4914 => x"58",
          4915 => x"75",
          4916 => x"f7",
          4917 => x"d3",
          4918 => x"52",
          4919 => x"51",
          4920 => x"80",
          4921 => x"90",
          4922 => x"82",
          4923 => x"f7",
          4924 => x"b0",
          4925 => x"a8",
          4926 => x"80",
          4927 => x"74",
          4928 => x"82",
          4929 => x"dc",
          4930 => x"8c",
          4931 => x"dc",
          4932 => x"06",
          4933 => x"74",
          4934 => x"ff",
          4935 => x"93",
          4936 => x"39",
          4937 => x"82",
          4938 => x"fc",
          4939 => x"54",
          4940 => x"a7",
          4941 => x"ff",
          4942 => x"82",
          4943 => x"82",
          4944 => x"82",
          4945 => x"81",
          4946 => x"05",
          4947 => x"79",
          4948 => x"92",
          4949 => x"54",
          4950 => x"73",
          4951 => x"80",
          4952 => x"38",
          4953 => x"a1",
          4954 => x"39",
          4955 => x"09",
          4956 => x"38",
          4957 => x"08",
          4958 => x"2e",
          4959 => x"51",
          4960 => x"3f",
          4961 => x"08",
          4962 => x"34",
          4963 => x"08",
          4964 => x"81",
          4965 => x"52",
          4966 => x"a2",
          4967 => x"c3",
          4968 => x"29",
          4969 => x"05",
          4970 => x"54",
          4971 => x"ab",
          4972 => x"ff",
          4973 => x"82",
          4974 => x"82",
          4975 => x"82",
          4976 => x"81",
          4977 => x"05",
          4978 => x"79",
          4979 => x"96",
          4980 => x"54",
          4981 => x"06",
          4982 => x"74",
          4983 => x"34",
          4984 => x"82",
          4985 => x"82",
          4986 => x"52",
          4987 => x"e2",
          4988 => x"39",
          4989 => x"33",
          4990 => x"06",
          4991 => x"33",
          4992 => x"74",
          4993 => x"87",
          4994 => x"b0",
          4995 => x"14",
          4996 => x"d3",
          4997 => x"1a",
          4998 => x"54",
          4999 => x"3f",
          5000 => x"82",
          5001 => x"54",
          5002 => x"f4",
          5003 => x"d3",
          5004 => x"88",
          5005 => x"fb",
          5006 => x"90",
          5007 => x"54",
          5008 => x"90",
          5009 => x"39",
          5010 => x"83",
          5011 => x"82",
          5012 => x"84",
          5013 => x"bb",
          5014 => x"80",
          5015 => x"83",
          5016 => x"ff",
          5017 => x"82",
          5018 => x"54",
          5019 => x"74",
          5020 => x"76",
          5021 => x"82",
          5022 => x"54",
          5023 => x"34",
          5024 => x"34",
          5025 => x"08",
          5026 => x"15",
          5027 => x"15",
          5028 => x"d4",
          5029 => x"d0",
          5030 => x"fe",
          5031 => x"70",
          5032 => x"06",
          5033 => x"58",
          5034 => x"74",
          5035 => x"73",
          5036 => x"82",
          5037 => x"70",
          5038 => x"bb",
          5039 => x"f8",
          5040 => x"55",
          5041 => x"34",
          5042 => x"34",
          5043 => x"04",
          5044 => x"73",
          5045 => x"84",
          5046 => x"38",
          5047 => x"2a",
          5048 => x"83",
          5049 => x"51",
          5050 => x"82",
          5051 => x"83",
          5052 => x"f9",
          5053 => x"a6",
          5054 => x"84",
          5055 => x"22",
          5056 => x"bb",
          5057 => x"83",
          5058 => x"74",
          5059 => x"11",
          5060 => x"12",
          5061 => x"2b",
          5062 => x"05",
          5063 => x"71",
          5064 => x"06",
          5065 => x"2a",
          5066 => x"59",
          5067 => x"57",
          5068 => x"71",
          5069 => x"81",
          5070 => x"bb",
          5071 => x"75",
          5072 => x"54",
          5073 => x"34",
          5074 => x"34",
          5075 => x"08",
          5076 => x"33",
          5077 => x"71",
          5078 => x"70",
          5079 => x"ff",
          5080 => x"52",
          5081 => x"05",
          5082 => x"ff",
          5083 => x"2a",
          5084 => x"71",
          5085 => x"72",
          5086 => x"53",
          5087 => x"34",
          5088 => x"08",
          5089 => x"76",
          5090 => x"17",
          5091 => x"0d",
          5092 => x"0d",
          5093 => x"08",
          5094 => x"9e",
          5095 => x"83",
          5096 => x"86",
          5097 => x"12",
          5098 => x"2b",
          5099 => x"07",
          5100 => x"52",
          5101 => x"05",
          5102 => x"85",
          5103 => x"88",
          5104 => x"88",
          5105 => x"56",
          5106 => x"13",
          5107 => x"13",
          5108 => x"d4",
          5109 => x"84",
          5110 => x"12",
          5111 => x"2b",
          5112 => x"07",
          5113 => x"52",
          5114 => x"12",
          5115 => x"33",
          5116 => x"07",
          5117 => x"54",
          5118 => x"70",
          5119 => x"73",
          5120 => x"82",
          5121 => x"13",
          5122 => x"12",
          5123 => x"2b",
          5124 => x"ff",
          5125 => x"88",
          5126 => x"53",
          5127 => x"73",
          5128 => x"14",
          5129 => x"0d",
          5130 => x"0d",
          5131 => x"22",
          5132 => x"08",
          5133 => x"71",
          5134 => x"81",
          5135 => x"88",
          5136 => x"88",
          5137 => x"33",
          5138 => x"71",
          5139 => x"90",
          5140 => x"5f",
          5141 => x"5a",
          5142 => x"54",
          5143 => x"80",
          5144 => x"51",
          5145 => x"82",
          5146 => x"70",
          5147 => x"81",
          5148 => x"8b",
          5149 => x"2b",
          5150 => x"70",
          5151 => x"33",
          5152 => x"07",
          5153 => x"8f",
          5154 => x"51",
          5155 => x"53",
          5156 => x"72",
          5157 => x"2a",
          5158 => x"82",
          5159 => x"83",
          5160 => x"bb",
          5161 => x"16",
          5162 => x"12",
          5163 => x"2b",
          5164 => x"07",
          5165 => x"55",
          5166 => x"33",
          5167 => x"71",
          5168 => x"70",
          5169 => x"06",
          5170 => x"57",
          5171 => x"52",
          5172 => x"71",
          5173 => x"88",
          5174 => x"fb",
          5175 => x"bb",
          5176 => x"84",
          5177 => x"22",
          5178 => x"72",
          5179 => x"33",
          5180 => x"71",
          5181 => x"83",
          5182 => x"5b",
          5183 => x"52",
          5184 => x"33",
          5185 => x"71",
          5186 => x"02",
          5187 => x"05",
          5188 => x"70",
          5189 => x"51",
          5190 => x"71",
          5191 => x"81",
          5192 => x"bb",
          5193 => x"15",
          5194 => x"12",
          5195 => x"2b",
          5196 => x"07",
          5197 => x"52",
          5198 => x"12",
          5199 => x"33",
          5200 => x"07",
          5201 => x"54",
          5202 => x"70",
          5203 => x"72",
          5204 => x"82",
          5205 => x"14",
          5206 => x"83",
          5207 => x"88",
          5208 => x"bb",
          5209 => x"54",
          5210 => x"04",
          5211 => x"7b",
          5212 => x"08",
          5213 => x"70",
          5214 => x"06",
          5215 => x"53",
          5216 => x"82",
          5217 => x"76",
          5218 => x"11",
          5219 => x"83",
          5220 => x"8b",
          5221 => x"2b",
          5222 => x"70",
          5223 => x"33",
          5224 => x"71",
          5225 => x"53",
          5226 => x"53",
          5227 => x"59",
          5228 => x"25",
          5229 => x"80",
          5230 => x"51",
          5231 => x"81",
          5232 => x"14",
          5233 => x"33",
          5234 => x"71",
          5235 => x"76",
          5236 => x"2a",
          5237 => x"58",
          5238 => x"14",
          5239 => x"ff",
          5240 => x"87",
          5241 => x"bb",
          5242 => x"19",
          5243 => x"85",
          5244 => x"88",
          5245 => x"88",
          5246 => x"5b",
          5247 => x"84",
          5248 => x"85",
          5249 => x"bb",
          5250 => x"53",
          5251 => x"14",
          5252 => x"87",
          5253 => x"bb",
          5254 => x"76",
          5255 => x"75",
          5256 => x"82",
          5257 => x"18",
          5258 => x"12",
          5259 => x"2b",
          5260 => x"80",
          5261 => x"88",
          5262 => x"55",
          5263 => x"74",
          5264 => x"15",
          5265 => x"0d",
          5266 => x"0d",
          5267 => x"bb",
          5268 => x"38",
          5269 => x"71",
          5270 => x"38",
          5271 => x"8c",
          5272 => x"0d",
          5273 => x"0d",
          5274 => x"58",
          5275 => x"82",
          5276 => x"83",
          5277 => x"82",
          5278 => x"84",
          5279 => x"12",
          5280 => x"2b",
          5281 => x"59",
          5282 => x"81",
          5283 => x"75",
          5284 => x"cb",
          5285 => x"29",
          5286 => x"81",
          5287 => x"88",
          5288 => x"81",
          5289 => x"79",
          5290 => x"ff",
          5291 => x"7f",
          5292 => x"51",
          5293 => x"77",
          5294 => x"38",
          5295 => x"85",
          5296 => x"5a",
          5297 => x"33",
          5298 => x"71",
          5299 => x"57",
          5300 => x"38",
          5301 => x"ff",
          5302 => x"7a",
          5303 => x"80",
          5304 => x"82",
          5305 => x"11",
          5306 => x"12",
          5307 => x"2b",
          5308 => x"ff",
          5309 => x"52",
          5310 => x"55",
          5311 => x"83",
          5312 => x"80",
          5313 => x"26",
          5314 => x"74",
          5315 => x"2e",
          5316 => x"77",
          5317 => x"81",
          5318 => x"75",
          5319 => x"3f",
          5320 => x"82",
          5321 => x"79",
          5322 => x"f7",
          5323 => x"bb",
          5324 => x"1c",
          5325 => x"87",
          5326 => x"8b",
          5327 => x"2b",
          5328 => x"5e",
          5329 => x"7a",
          5330 => x"ff",
          5331 => x"88",
          5332 => x"56",
          5333 => x"15",
          5334 => x"ff",
          5335 => x"85",
          5336 => x"bb",
          5337 => x"83",
          5338 => x"72",
          5339 => x"33",
          5340 => x"71",
          5341 => x"70",
          5342 => x"5b",
          5343 => x"56",
          5344 => x"19",
          5345 => x"19",
          5346 => x"d4",
          5347 => x"84",
          5348 => x"12",
          5349 => x"2b",
          5350 => x"07",
          5351 => x"55",
          5352 => x"78",
          5353 => x"76",
          5354 => x"82",
          5355 => x"70",
          5356 => x"84",
          5357 => x"12",
          5358 => x"2b",
          5359 => x"2a",
          5360 => x"52",
          5361 => x"84",
          5362 => x"85",
          5363 => x"bb",
          5364 => x"84",
          5365 => x"82",
          5366 => x"8d",
          5367 => x"fe",
          5368 => x"52",
          5369 => x"08",
          5370 => x"dc",
          5371 => x"71",
          5372 => x"38",
          5373 => x"ed",
          5374 => x"dc",
          5375 => x"82",
          5376 => x"84",
          5377 => x"ee",
          5378 => x"66",
          5379 => x"70",
          5380 => x"bb",
          5381 => x"2e",
          5382 => x"84",
          5383 => x"3f",
          5384 => x"7e",
          5385 => x"3f",
          5386 => x"08",
          5387 => x"39",
          5388 => x"7b",
          5389 => x"3f",
          5390 => x"ba",
          5391 => x"f5",
          5392 => x"bb",
          5393 => x"ff",
          5394 => x"bb",
          5395 => x"71",
          5396 => x"70",
          5397 => x"06",
          5398 => x"73",
          5399 => x"81",
          5400 => x"88",
          5401 => x"75",
          5402 => x"ff",
          5403 => x"88",
          5404 => x"73",
          5405 => x"70",
          5406 => x"33",
          5407 => x"07",
          5408 => x"53",
          5409 => x"48",
          5410 => x"54",
          5411 => x"56",
          5412 => x"80",
          5413 => x"76",
          5414 => x"06",
          5415 => x"83",
          5416 => x"42",
          5417 => x"33",
          5418 => x"71",
          5419 => x"70",
          5420 => x"70",
          5421 => x"33",
          5422 => x"71",
          5423 => x"53",
          5424 => x"56",
          5425 => x"25",
          5426 => x"75",
          5427 => x"ff",
          5428 => x"54",
          5429 => x"81",
          5430 => x"18",
          5431 => x"2e",
          5432 => x"8f",
          5433 => x"f6",
          5434 => x"83",
          5435 => x"58",
          5436 => x"7f",
          5437 => x"74",
          5438 => x"78",
          5439 => x"3f",
          5440 => x"7f",
          5441 => x"75",
          5442 => x"38",
          5443 => x"11",
          5444 => x"33",
          5445 => x"07",
          5446 => x"f4",
          5447 => x"52",
          5448 => x"b7",
          5449 => x"dc",
          5450 => x"ff",
          5451 => x"7c",
          5452 => x"2b",
          5453 => x"08",
          5454 => x"53",
          5455 => x"8e",
          5456 => x"bb",
          5457 => x"84",
          5458 => x"ff",
          5459 => x"5c",
          5460 => x"60",
          5461 => x"74",
          5462 => x"38",
          5463 => x"c9",
          5464 => x"d4",
          5465 => x"11",
          5466 => x"33",
          5467 => x"07",
          5468 => x"f4",
          5469 => x"52",
          5470 => x"df",
          5471 => x"dc",
          5472 => x"ff",
          5473 => x"7c",
          5474 => x"2b",
          5475 => x"08",
          5476 => x"53",
          5477 => x"8e",
          5478 => x"bb",
          5479 => x"84",
          5480 => x"05",
          5481 => x"73",
          5482 => x"06",
          5483 => x"7b",
          5484 => x"f9",
          5485 => x"bb",
          5486 => x"82",
          5487 => x"80",
          5488 => x"7d",
          5489 => x"82",
          5490 => x"51",
          5491 => x"3f",
          5492 => x"98",
          5493 => x"7a",
          5494 => x"38",
          5495 => x"52",
          5496 => x"8f",
          5497 => x"83",
          5498 => x"d4",
          5499 => x"05",
          5500 => x"3f",
          5501 => x"82",
          5502 => x"94",
          5503 => x"fc",
          5504 => x"77",
          5505 => x"54",
          5506 => x"82",
          5507 => x"55",
          5508 => x"08",
          5509 => x"38",
          5510 => x"52",
          5511 => x"08",
          5512 => x"c3",
          5513 => x"bb",
          5514 => x"3d",
          5515 => x"3d",
          5516 => x"05",
          5517 => x"52",
          5518 => x"87",
          5519 => x"d8",
          5520 => x"71",
          5521 => x"0c",
          5522 => x"04",
          5523 => x"02",
          5524 => x"02",
          5525 => x"05",
          5526 => x"83",
          5527 => x"26",
          5528 => x"72",
          5529 => x"c0",
          5530 => x"53",
          5531 => x"74",
          5532 => x"38",
          5533 => x"73",
          5534 => x"c0",
          5535 => x"51",
          5536 => x"85",
          5537 => x"98",
          5538 => x"52",
          5539 => x"82",
          5540 => x"70",
          5541 => x"38",
          5542 => x"8c",
          5543 => x"ec",
          5544 => x"fc",
          5545 => x"52",
          5546 => x"87",
          5547 => x"08",
          5548 => x"2e",
          5549 => x"82",
          5550 => x"34",
          5551 => x"13",
          5552 => x"82",
          5553 => x"86",
          5554 => x"f3",
          5555 => x"62",
          5556 => x"05",
          5557 => x"57",
          5558 => x"83",
          5559 => x"fe",
          5560 => x"bb",
          5561 => x"06",
          5562 => x"71",
          5563 => x"71",
          5564 => x"2b",
          5565 => x"80",
          5566 => x"92",
          5567 => x"c0",
          5568 => x"41",
          5569 => x"5a",
          5570 => x"87",
          5571 => x"0c",
          5572 => x"84",
          5573 => x"08",
          5574 => x"70",
          5575 => x"53",
          5576 => x"2e",
          5577 => x"08",
          5578 => x"70",
          5579 => x"34",
          5580 => x"80",
          5581 => x"53",
          5582 => x"2e",
          5583 => x"53",
          5584 => x"26",
          5585 => x"80",
          5586 => x"87",
          5587 => x"08",
          5588 => x"38",
          5589 => x"8c",
          5590 => x"80",
          5591 => x"78",
          5592 => x"99",
          5593 => x"0c",
          5594 => x"8c",
          5595 => x"08",
          5596 => x"51",
          5597 => x"38",
          5598 => x"8d",
          5599 => x"17",
          5600 => x"81",
          5601 => x"53",
          5602 => x"2e",
          5603 => x"fc",
          5604 => x"52",
          5605 => x"7d",
          5606 => x"ed",
          5607 => x"80",
          5608 => x"71",
          5609 => x"38",
          5610 => x"53",
          5611 => x"dc",
          5612 => x"0d",
          5613 => x"0d",
          5614 => x"02",
          5615 => x"05",
          5616 => x"58",
          5617 => x"80",
          5618 => x"fc",
          5619 => x"bb",
          5620 => x"06",
          5621 => x"71",
          5622 => x"81",
          5623 => x"38",
          5624 => x"2b",
          5625 => x"80",
          5626 => x"92",
          5627 => x"c0",
          5628 => x"40",
          5629 => x"5a",
          5630 => x"c0",
          5631 => x"76",
          5632 => x"76",
          5633 => x"75",
          5634 => x"2a",
          5635 => x"51",
          5636 => x"80",
          5637 => x"7a",
          5638 => x"5c",
          5639 => x"81",
          5640 => x"81",
          5641 => x"06",
          5642 => x"80",
          5643 => x"87",
          5644 => x"08",
          5645 => x"38",
          5646 => x"8c",
          5647 => x"80",
          5648 => x"77",
          5649 => x"99",
          5650 => x"0c",
          5651 => x"8c",
          5652 => x"08",
          5653 => x"51",
          5654 => x"38",
          5655 => x"8d",
          5656 => x"70",
          5657 => x"84",
          5658 => x"5b",
          5659 => x"2e",
          5660 => x"fc",
          5661 => x"52",
          5662 => x"7d",
          5663 => x"f8",
          5664 => x"80",
          5665 => x"71",
          5666 => x"38",
          5667 => x"53",
          5668 => x"dc",
          5669 => x"0d",
          5670 => x"0d",
          5671 => x"05",
          5672 => x"02",
          5673 => x"05",
          5674 => x"54",
          5675 => x"fe",
          5676 => x"dc",
          5677 => x"53",
          5678 => x"80",
          5679 => x"0b",
          5680 => x"8c",
          5681 => x"71",
          5682 => x"dc",
          5683 => x"24",
          5684 => x"84",
          5685 => x"92",
          5686 => x"54",
          5687 => x"8d",
          5688 => x"39",
          5689 => x"80",
          5690 => x"cb",
          5691 => x"70",
          5692 => x"81",
          5693 => x"52",
          5694 => x"8a",
          5695 => x"98",
          5696 => x"71",
          5697 => x"c0",
          5698 => x"52",
          5699 => x"81",
          5700 => x"c0",
          5701 => x"53",
          5702 => x"82",
          5703 => x"71",
          5704 => x"39",
          5705 => x"39",
          5706 => x"77",
          5707 => x"81",
          5708 => x"72",
          5709 => x"84",
          5710 => x"73",
          5711 => x"0c",
          5712 => x"04",
          5713 => x"74",
          5714 => x"71",
          5715 => x"2b",
          5716 => x"dc",
          5717 => x"84",
          5718 => x"fd",
          5719 => x"83",
          5720 => x"12",
          5721 => x"2b",
          5722 => x"07",
          5723 => x"70",
          5724 => x"2b",
          5725 => x"07",
          5726 => x"0c",
          5727 => x"56",
          5728 => x"3d",
          5729 => x"3d",
          5730 => x"84",
          5731 => x"22",
          5732 => x"72",
          5733 => x"54",
          5734 => x"2a",
          5735 => x"34",
          5736 => x"04",
          5737 => x"73",
          5738 => x"70",
          5739 => x"05",
          5740 => x"88",
          5741 => x"72",
          5742 => x"54",
          5743 => x"2a",
          5744 => x"70",
          5745 => x"34",
          5746 => x"51",
          5747 => x"83",
          5748 => x"fe",
          5749 => x"75",
          5750 => x"51",
          5751 => x"92",
          5752 => x"81",
          5753 => x"73",
          5754 => x"55",
          5755 => x"51",
          5756 => x"3d",
          5757 => x"3d",
          5758 => x"76",
          5759 => x"72",
          5760 => x"05",
          5761 => x"11",
          5762 => x"38",
          5763 => x"04",
          5764 => x"78",
          5765 => x"56",
          5766 => x"81",
          5767 => x"74",
          5768 => x"56",
          5769 => x"31",
          5770 => x"52",
          5771 => x"80",
          5772 => x"71",
          5773 => x"38",
          5774 => x"dc",
          5775 => x"0d",
          5776 => x"0d",
          5777 => x"51",
          5778 => x"73",
          5779 => x"81",
          5780 => x"33",
          5781 => x"38",
          5782 => x"bb",
          5783 => x"3d",
          5784 => x"0b",
          5785 => x"0c",
          5786 => x"82",
          5787 => x"04",
          5788 => x"7b",
          5789 => x"83",
          5790 => x"5a",
          5791 => x"80",
          5792 => x"54",
          5793 => x"53",
          5794 => x"53",
          5795 => x"52",
          5796 => x"3f",
          5797 => x"08",
          5798 => x"81",
          5799 => x"82",
          5800 => x"83",
          5801 => x"16",
          5802 => x"18",
          5803 => x"18",
          5804 => x"58",
          5805 => x"9f",
          5806 => x"33",
          5807 => x"2e",
          5808 => x"93",
          5809 => x"76",
          5810 => x"52",
          5811 => x"51",
          5812 => x"83",
          5813 => x"79",
          5814 => x"0c",
          5815 => x"04",
          5816 => x"78",
          5817 => x"80",
          5818 => x"17",
          5819 => x"38",
          5820 => x"fc",
          5821 => x"dc",
          5822 => x"bb",
          5823 => x"38",
          5824 => x"53",
          5825 => x"81",
          5826 => x"f7",
          5827 => x"bb",
          5828 => x"2e",
          5829 => x"55",
          5830 => x"b0",
          5831 => x"82",
          5832 => x"88",
          5833 => x"f8",
          5834 => x"70",
          5835 => x"c0",
          5836 => x"dc",
          5837 => x"bb",
          5838 => x"91",
          5839 => x"55",
          5840 => x"09",
          5841 => x"f0",
          5842 => x"33",
          5843 => x"2e",
          5844 => x"80",
          5845 => x"80",
          5846 => x"dc",
          5847 => x"17",
          5848 => x"fd",
          5849 => x"d4",
          5850 => x"b2",
          5851 => x"96",
          5852 => x"85",
          5853 => x"75",
          5854 => x"3f",
          5855 => x"e4",
          5856 => x"98",
          5857 => x"9c",
          5858 => x"08",
          5859 => x"17",
          5860 => x"3f",
          5861 => x"52",
          5862 => x"51",
          5863 => x"a0",
          5864 => x"05",
          5865 => x"0c",
          5866 => x"75",
          5867 => x"33",
          5868 => x"3f",
          5869 => x"34",
          5870 => x"52",
          5871 => x"51",
          5872 => x"82",
          5873 => x"80",
          5874 => x"81",
          5875 => x"bb",
          5876 => x"3d",
          5877 => x"3d",
          5878 => x"1a",
          5879 => x"fe",
          5880 => x"54",
          5881 => x"73",
          5882 => x"8a",
          5883 => x"71",
          5884 => x"08",
          5885 => x"75",
          5886 => x"0c",
          5887 => x"04",
          5888 => x"7a",
          5889 => x"56",
          5890 => x"77",
          5891 => x"38",
          5892 => x"08",
          5893 => x"38",
          5894 => x"54",
          5895 => x"2e",
          5896 => x"72",
          5897 => x"38",
          5898 => x"8d",
          5899 => x"39",
          5900 => x"81",
          5901 => x"b6",
          5902 => x"2a",
          5903 => x"2a",
          5904 => x"05",
          5905 => x"55",
          5906 => x"82",
          5907 => x"81",
          5908 => x"83",
          5909 => x"b4",
          5910 => x"17",
          5911 => x"a4",
          5912 => x"55",
          5913 => x"57",
          5914 => x"3f",
          5915 => x"08",
          5916 => x"74",
          5917 => x"14",
          5918 => x"70",
          5919 => x"07",
          5920 => x"71",
          5921 => x"52",
          5922 => x"72",
          5923 => x"75",
          5924 => x"58",
          5925 => x"76",
          5926 => x"15",
          5927 => x"73",
          5928 => x"3f",
          5929 => x"08",
          5930 => x"76",
          5931 => x"06",
          5932 => x"05",
          5933 => x"3f",
          5934 => x"08",
          5935 => x"06",
          5936 => x"76",
          5937 => x"15",
          5938 => x"73",
          5939 => x"3f",
          5940 => x"08",
          5941 => x"82",
          5942 => x"06",
          5943 => x"05",
          5944 => x"3f",
          5945 => x"08",
          5946 => x"58",
          5947 => x"58",
          5948 => x"dc",
          5949 => x"0d",
          5950 => x"0d",
          5951 => x"5a",
          5952 => x"59",
          5953 => x"82",
          5954 => x"98",
          5955 => x"82",
          5956 => x"33",
          5957 => x"2e",
          5958 => x"72",
          5959 => x"38",
          5960 => x"8d",
          5961 => x"39",
          5962 => x"81",
          5963 => x"f7",
          5964 => x"2a",
          5965 => x"2a",
          5966 => x"05",
          5967 => x"55",
          5968 => x"82",
          5969 => x"59",
          5970 => x"08",
          5971 => x"74",
          5972 => x"16",
          5973 => x"16",
          5974 => x"59",
          5975 => x"53",
          5976 => x"8f",
          5977 => x"2b",
          5978 => x"74",
          5979 => x"71",
          5980 => x"72",
          5981 => x"0b",
          5982 => x"74",
          5983 => x"17",
          5984 => x"75",
          5985 => x"3f",
          5986 => x"08",
          5987 => x"dc",
          5988 => x"38",
          5989 => x"06",
          5990 => x"78",
          5991 => x"54",
          5992 => x"77",
          5993 => x"33",
          5994 => x"71",
          5995 => x"51",
          5996 => x"34",
          5997 => x"76",
          5998 => x"17",
          5999 => x"75",
          6000 => x"3f",
          6001 => x"08",
          6002 => x"dc",
          6003 => x"38",
          6004 => x"ff",
          6005 => x"10",
          6006 => x"76",
          6007 => x"51",
          6008 => x"be",
          6009 => x"2a",
          6010 => x"05",
          6011 => x"f9",
          6012 => x"bb",
          6013 => x"82",
          6014 => x"ab",
          6015 => x"0a",
          6016 => x"2b",
          6017 => x"70",
          6018 => x"70",
          6019 => x"54",
          6020 => x"82",
          6021 => x"8f",
          6022 => x"07",
          6023 => x"f7",
          6024 => x"0b",
          6025 => x"78",
          6026 => x"0c",
          6027 => x"04",
          6028 => x"7a",
          6029 => x"08",
          6030 => x"59",
          6031 => x"a4",
          6032 => x"17",
          6033 => x"38",
          6034 => x"aa",
          6035 => x"73",
          6036 => x"fd",
          6037 => x"bb",
          6038 => x"82",
          6039 => x"80",
          6040 => x"39",
          6041 => x"eb",
          6042 => x"80",
          6043 => x"bb",
          6044 => x"80",
          6045 => x"52",
          6046 => x"84",
          6047 => x"dc",
          6048 => x"bb",
          6049 => x"2e",
          6050 => x"82",
          6051 => x"81",
          6052 => x"82",
          6053 => x"ff",
          6054 => x"80",
          6055 => x"75",
          6056 => x"3f",
          6057 => x"08",
          6058 => x"16",
          6059 => x"90",
          6060 => x"55",
          6061 => x"27",
          6062 => x"15",
          6063 => x"84",
          6064 => x"07",
          6065 => x"17",
          6066 => x"76",
          6067 => x"a6",
          6068 => x"73",
          6069 => x"0c",
          6070 => x"04",
          6071 => x"7c",
          6072 => x"59",
          6073 => x"95",
          6074 => x"08",
          6075 => x"2e",
          6076 => x"17",
          6077 => x"b2",
          6078 => x"ae",
          6079 => x"7a",
          6080 => x"3f",
          6081 => x"82",
          6082 => x"27",
          6083 => x"82",
          6084 => x"55",
          6085 => x"08",
          6086 => x"d2",
          6087 => x"08",
          6088 => x"08",
          6089 => x"38",
          6090 => x"17",
          6091 => x"54",
          6092 => x"82",
          6093 => x"7a",
          6094 => x"06",
          6095 => x"81",
          6096 => x"17",
          6097 => x"83",
          6098 => x"75",
          6099 => x"f9",
          6100 => x"59",
          6101 => x"08",
          6102 => x"81",
          6103 => x"82",
          6104 => x"59",
          6105 => x"08",
          6106 => x"70",
          6107 => x"25",
          6108 => x"82",
          6109 => x"54",
          6110 => x"55",
          6111 => x"38",
          6112 => x"08",
          6113 => x"38",
          6114 => x"54",
          6115 => x"90",
          6116 => x"18",
          6117 => x"38",
          6118 => x"39",
          6119 => x"38",
          6120 => x"16",
          6121 => x"08",
          6122 => x"38",
          6123 => x"78",
          6124 => x"38",
          6125 => x"51",
          6126 => x"82",
          6127 => x"80",
          6128 => x"80",
          6129 => x"dc",
          6130 => x"09",
          6131 => x"38",
          6132 => x"08",
          6133 => x"dc",
          6134 => x"30",
          6135 => x"80",
          6136 => x"07",
          6137 => x"55",
          6138 => x"38",
          6139 => x"09",
          6140 => x"ae",
          6141 => x"80",
          6142 => x"53",
          6143 => x"51",
          6144 => x"82",
          6145 => x"82",
          6146 => x"30",
          6147 => x"dc",
          6148 => x"25",
          6149 => x"79",
          6150 => x"38",
          6151 => x"8f",
          6152 => x"79",
          6153 => x"f9",
          6154 => x"bb",
          6155 => x"74",
          6156 => x"8c",
          6157 => x"17",
          6158 => x"90",
          6159 => x"54",
          6160 => x"86",
          6161 => x"90",
          6162 => x"17",
          6163 => x"54",
          6164 => x"34",
          6165 => x"56",
          6166 => x"90",
          6167 => x"80",
          6168 => x"82",
          6169 => x"55",
          6170 => x"56",
          6171 => x"82",
          6172 => x"8c",
          6173 => x"f8",
          6174 => x"70",
          6175 => x"f0",
          6176 => x"dc",
          6177 => x"56",
          6178 => x"08",
          6179 => x"7b",
          6180 => x"f6",
          6181 => x"bb",
          6182 => x"bb",
          6183 => x"17",
          6184 => x"80",
          6185 => x"b4",
          6186 => x"57",
          6187 => x"77",
          6188 => x"81",
          6189 => x"15",
          6190 => x"78",
          6191 => x"81",
          6192 => x"53",
          6193 => x"15",
          6194 => x"e9",
          6195 => x"dc",
          6196 => x"df",
          6197 => x"22",
          6198 => x"30",
          6199 => x"70",
          6200 => x"51",
          6201 => x"82",
          6202 => x"8a",
          6203 => x"f8",
          6204 => x"7c",
          6205 => x"56",
          6206 => x"80",
          6207 => x"f1",
          6208 => x"06",
          6209 => x"e9",
          6210 => x"18",
          6211 => x"08",
          6212 => x"38",
          6213 => x"82",
          6214 => x"38",
          6215 => x"54",
          6216 => x"74",
          6217 => x"82",
          6218 => x"22",
          6219 => x"79",
          6220 => x"38",
          6221 => x"98",
          6222 => x"cd",
          6223 => x"22",
          6224 => x"54",
          6225 => x"26",
          6226 => x"52",
          6227 => x"b0",
          6228 => x"dc",
          6229 => x"bb",
          6230 => x"2e",
          6231 => x"0b",
          6232 => x"08",
          6233 => x"98",
          6234 => x"bb",
          6235 => x"85",
          6236 => x"bd",
          6237 => x"31",
          6238 => x"73",
          6239 => x"f4",
          6240 => x"bb",
          6241 => x"18",
          6242 => x"18",
          6243 => x"08",
          6244 => x"72",
          6245 => x"38",
          6246 => x"58",
          6247 => x"89",
          6248 => x"18",
          6249 => x"ff",
          6250 => x"05",
          6251 => x"80",
          6252 => x"bb",
          6253 => x"3d",
          6254 => x"3d",
          6255 => x"08",
          6256 => x"a0",
          6257 => x"54",
          6258 => x"77",
          6259 => x"80",
          6260 => x"0c",
          6261 => x"53",
          6262 => x"80",
          6263 => x"38",
          6264 => x"06",
          6265 => x"b5",
          6266 => x"98",
          6267 => x"14",
          6268 => x"92",
          6269 => x"2a",
          6270 => x"56",
          6271 => x"26",
          6272 => x"80",
          6273 => x"16",
          6274 => x"77",
          6275 => x"53",
          6276 => x"38",
          6277 => x"51",
          6278 => x"82",
          6279 => x"53",
          6280 => x"0b",
          6281 => x"08",
          6282 => x"38",
          6283 => x"bb",
          6284 => x"2e",
          6285 => x"98",
          6286 => x"bb",
          6287 => x"80",
          6288 => x"8a",
          6289 => x"15",
          6290 => x"80",
          6291 => x"14",
          6292 => x"51",
          6293 => x"82",
          6294 => x"53",
          6295 => x"bb",
          6296 => x"2e",
          6297 => x"82",
          6298 => x"dc",
          6299 => x"ba",
          6300 => x"82",
          6301 => x"ff",
          6302 => x"82",
          6303 => x"52",
          6304 => x"f3",
          6305 => x"dc",
          6306 => x"72",
          6307 => x"72",
          6308 => x"f2",
          6309 => x"bb",
          6310 => x"15",
          6311 => x"15",
          6312 => x"b4",
          6313 => x"0c",
          6314 => x"82",
          6315 => x"8a",
          6316 => x"f7",
          6317 => x"7d",
          6318 => x"5b",
          6319 => x"76",
          6320 => x"3f",
          6321 => x"08",
          6322 => x"dc",
          6323 => x"38",
          6324 => x"08",
          6325 => x"08",
          6326 => x"f0",
          6327 => x"bb",
          6328 => x"82",
          6329 => x"80",
          6330 => x"bb",
          6331 => x"18",
          6332 => x"51",
          6333 => x"81",
          6334 => x"81",
          6335 => x"81",
          6336 => x"dc",
          6337 => x"83",
          6338 => x"77",
          6339 => x"72",
          6340 => x"38",
          6341 => x"75",
          6342 => x"81",
          6343 => x"a5",
          6344 => x"dc",
          6345 => x"52",
          6346 => x"8e",
          6347 => x"dc",
          6348 => x"bb",
          6349 => x"2e",
          6350 => x"73",
          6351 => x"81",
          6352 => x"87",
          6353 => x"bb",
          6354 => x"3d",
          6355 => x"3d",
          6356 => x"11",
          6357 => x"ec",
          6358 => x"dc",
          6359 => x"ff",
          6360 => x"33",
          6361 => x"71",
          6362 => x"81",
          6363 => x"94",
          6364 => x"d0",
          6365 => x"dc",
          6366 => x"73",
          6367 => x"82",
          6368 => x"85",
          6369 => x"fc",
          6370 => x"79",
          6371 => x"ff",
          6372 => x"12",
          6373 => x"eb",
          6374 => x"70",
          6375 => x"72",
          6376 => x"81",
          6377 => x"73",
          6378 => x"94",
          6379 => x"d6",
          6380 => x"0d",
          6381 => x"0d",
          6382 => x"55",
          6383 => x"5a",
          6384 => x"08",
          6385 => x"8a",
          6386 => x"08",
          6387 => x"ee",
          6388 => x"bb",
          6389 => x"82",
          6390 => x"80",
          6391 => x"15",
          6392 => x"55",
          6393 => x"38",
          6394 => x"e6",
          6395 => x"33",
          6396 => x"70",
          6397 => x"58",
          6398 => x"86",
          6399 => x"bb",
          6400 => x"73",
          6401 => x"83",
          6402 => x"73",
          6403 => x"38",
          6404 => x"06",
          6405 => x"80",
          6406 => x"75",
          6407 => x"38",
          6408 => x"08",
          6409 => x"54",
          6410 => x"2e",
          6411 => x"83",
          6412 => x"73",
          6413 => x"38",
          6414 => x"51",
          6415 => x"82",
          6416 => x"58",
          6417 => x"08",
          6418 => x"15",
          6419 => x"38",
          6420 => x"0b",
          6421 => x"77",
          6422 => x"0c",
          6423 => x"04",
          6424 => x"77",
          6425 => x"54",
          6426 => x"51",
          6427 => x"82",
          6428 => x"55",
          6429 => x"08",
          6430 => x"14",
          6431 => x"51",
          6432 => x"82",
          6433 => x"55",
          6434 => x"08",
          6435 => x"53",
          6436 => x"08",
          6437 => x"08",
          6438 => x"3f",
          6439 => x"14",
          6440 => x"08",
          6441 => x"3f",
          6442 => x"17",
          6443 => x"bb",
          6444 => x"3d",
          6445 => x"3d",
          6446 => x"08",
          6447 => x"54",
          6448 => x"53",
          6449 => x"82",
          6450 => x"8d",
          6451 => x"08",
          6452 => x"34",
          6453 => x"15",
          6454 => x"0d",
          6455 => x"0d",
          6456 => x"57",
          6457 => x"17",
          6458 => x"08",
          6459 => x"82",
          6460 => x"89",
          6461 => x"55",
          6462 => x"14",
          6463 => x"16",
          6464 => x"71",
          6465 => x"38",
          6466 => x"09",
          6467 => x"38",
          6468 => x"73",
          6469 => x"81",
          6470 => x"ae",
          6471 => x"05",
          6472 => x"15",
          6473 => x"70",
          6474 => x"34",
          6475 => x"8a",
          6476 => x"38",
          6477 => x"05",
          6478 => x"81",
          6479 => x"17",
          6480 => x"12",
          6481 => x"34",
          6482 => x"9c",
          6483 => x"e8",
          6484 => x"bb",
          6485 => x"0c",
          6486 => x"e7",
          6487 => x"bb",
          6488 => x"17",
          6489 => x"51",
          6490 => x"82",
          6491 => x"84",
          6492 => x"3d",
          6493 => x"3d",
          6494 => x"08",
          6495 => x"61",
          6496 => x"55",
          6497 => x"2e",
          6498 => x"55",
          6499 => x"2e",
          6500 => x"80",
          6501 => x"94",
          6502 => x"1c",
          6503 => x"81",
          6504 => x"61",
          6505 => x"56",
          6506 => x"2e",
          6507 => x"83",
          6508 => x"73",
          6509 => x"70",
          6510 => x"25",
          6511 => x"51",
          6512 => x"38",
          6513 => x"0c",
          6514 => x"51",
          6515 => x"26",
          6516 => x"80",
          6517 => x"34",
          6518 => x"51",
          6519 => x"82",
          6520 => x"55",
          6521 => x"91",
          6522 => x"1d",
          6523 => x"8b",
          6524 => x"79",
          6525 => x"3f",
          6526 => x"57",
          6527 => x"55",
          6528 => x"2e",
          6529 => x"80",
          6530 => x"18",
          6531 => x"1a",
          6532 => x"70",
          6533 => x"2a",
          6534 => x"07",
          6535 => x"5a",
          6536 => x"8c",
          6537 => x"54",
          6538 => x"81",
          6539 => x"39",
          6540 => x"70",
          6541 => x"2a",
          6542 => x"75",
          6543 => x"8c",
          6544 => x"2e",
          6545 => x"a0",
          6546 => x"38",
          6547 => x"0c",
          6548 => x"76",
          6549 => x"38",
          6550 => x"b8",
          6551 => x"70",
          6552 => x"5a",
          6553 => x"76",
          6554 => x"38",
          6555 => x"70",
          6556 => x"dc",
          6557 => x"72",
          6558 => x"80",
          6559 => x"51",
          6560 => x"73",
          6561 => x"38",
          6562 => x"18",
          6563 => x"1a",
          6564 => x"55",
          6565 => x"2e",
          6566 => x"83",
          6567 => x"73",
          6568 => x"70",
          6569 => x"25",
          6570 => x"51",
          6571 => x"38",
          6572 => x"75",
          6573 => x"81",
          6574 => x"81",
          6575 => x"27",
          6576 => x"73",
          6577 => x"38",
          6578 => x"70",
          6579 => x"32",
          6580 => x"80",
          6581 => x"2a",
          6582 => x"56",
          6583 => x"81",
          6584 => x"57",
          6585 => x"f5",
          6586 => x"2b",
          6587 => x"25",
          6588 => x"80",
          6589 => x"b5",
          6590 => x"57",
          6591 => x"e6",
          6592 => x"bb",
          6593 => x"2e",
          6594 => x"18",
          6595 => x"1a",
          6596 => x"56",
          6597 => x"3f",
          6598 => x"08",
          6599 => x"e8",
          6600 => x"54",
          6601 => x"80",
          6602 => x"17",
          6603 => x"34",
          6604 => x"11",
          6605 => x"74",
          6606 => x"75",
          6607 => x"c4",
          6608 => x"3f",
          6609 => x"08",
          6610 => x"9f",
          6611 => x"99",
          6612 => x"e0",
          6613 => x"ff",
          6614 => x"79",
          6615 => x"74",
          6616 => x"57",
          6617 => x"77",
          6618 => x"76",
          6619 => x"38",
          6620 => x"73",
          6621 => x"09",
          6622 => x"38",
          6623 => x"84",
          6624 => x"27",
          6625 => x"39",
          6626 => x"f2",
          6627 => x"80",
          6628 => x"54",
          6629 => x"34",
          6630 => x"58",
          6631 => x"f2",
          6632 => x"bb",
          6633 => x"82",
          6634 => x"80",
          6635 => x"1b",
          6636 => x"51",
          6637 => x"82",
          6638 => x"56",
          6639 => x"08",
          6640 => x"9c",
          6641 => x"33",
          6642 => x"80",
          6643 => x"38",
          6644 => x"bf",
          6645 => x"86",
          6646 => x"15",
          6647 => x"2a",
          6648 => x"51",
          6649 => x"92",
          6650 => x"79",
          6651 => x"e4",
          6652 => x"bb",
          6653 => x"2e",
          6654 => x"52",
          6655 => x"ba",
          6656 => x"39",
          6657 => x"33",
          6658 => x"80",
          6659 => x"74",
          6660 => x"81",
          6661 => x"38",
          6662 => x"70",
          6663 => x"82",
          6664 => x"54",
          6665 => x"96",
          6666 => x"06",
          6667 => x"2e",
          6668 => x"ff",
          6669 => x"1c",
          6670 => x"80",
          6671 => x"81",
          6672 => x"ba",
          6673 => x"b6",
          6674 => x"2a",
          6675 => x"51",
          6676 => x"38",
          6677 => x"70",
          6678 => x"81",
          6679 => x"55",
          6680 => x"e1",
          6681 => x"08",
          6682 => x"1d",
          6683 => x"7c",
          6684 => x"3f",
          6685 => x"08",
          6686 => x"fa",
          6687 => x"82",
          6688 => x"8f",
          6689 => x"f6",
          6690 => x"5b",
          6691 => x"70",
          6692 => x"59",
          6693 => x"73",
          6694 => x"c6",
          6695 => x"81",
          6696 => x"70",
          6697 => x"52",
          6698 => x"8d",
          6699 => x"38",
          6700 => x"09",
          6701 => x"a5",
          6702 => x"d0",
          6703 => x"ff",
          6704 => x"53",
          6705 => x"91",
          6706 => x"73",
          6707 => x"d0",
          6708 => x"71",
          6709 => x"f7",
          6710 => x"82",
          6711 => x"55",
          6712 => x"55",
          6713 => x"81",
          6714 => x"74",
          6715 => x"56",
          6716 => x"12",
          6717 => x"70",
          6718 => x"38",
          6719 => x"81",
          6720 => x"51",
          6721 => x"51",
          6722 => x"89",
          6723 => x"70",
          6724 => x"53",
          6725 => x"70",
          6726 => x"51",
          6727 => x"09",
          6728 => x"38",
          6729 => x"38",
          6730 => x"77",
          6731 => x"70",
          6732 => x"2a",
          6733 => x"07",
          6734 => x"51",
          6735 => x"8f",
          6736 => x"84",
          6737 => x"83",
          6738 => x"94",
          6739 => x"74",
          6740 => x"38",
          6741 => x"0c",
          6742 => x"86",
          6743 => x"a8",
          6744 => x"82",
          6745 => x"8c",
          6746 => x"fa",
          6747 => x"56",
          6748 => x"17",
          6749 => x"b0",
          6750 => x"52",
          6751 => x"e0",
          6752 => x"82",
          6753 => x"81",
          6754 => x"b2",
          6755 => x"b4",
          6756 => x"dc",
          6757 => x"ff",
          6758 => x"55",
          6759 => x"d5",
          6760 => x"06",
          6761 => x"80",
          6762 => x"33",
          6763 => x"81",
          6764 => x"81",
          6765 => x"81",
          6766 => x"eb",
          6767 => x"70",
          6768 => x"07",
          6769 => x"73",
          6770 => x"81",
          6771 => x"81",
          6772 => x"83",
          6773 => x"d4",
          6774 => x"16",
          6775 => x"3f",
          6776 => x"08",
          6777 => x"dc",
          6778 => x"9d",
          6779 => x"82",
          6780 => x"81",
          6781 => x"e0",
          6782 => x"bb",
          6783 => x"82",
          6784 => x"80",
          6785 => x"82",
          6786 => x"bb",
          6787 => x"3d",
          6788 => x"3d",
          6789 => x"84",
          6790 => x"05",
          6791 => x"80",
          6792 => x"51",
          6793 => x"82",
          6794 => x"58",
          6795 => x"0b",
          6796 => x"08",
          6797 => x"38",
          6798 => x"08",
          6799 => x"d3",
          6800 => x"08",
          6801 => x"56",
          6802 => x"86",
          6803 => x"75",
          6804 => x"fe",
          6805 => x"54",
          6806 => x"2e",
          6807 => x"14",
          6808 => x"ca",
          6809 => x"dc",
          6810 => x"06",
          6811 => x"54",
          6812 => x"38",
          6813 => x"86",
          6814 => x"82",
          6815 => x"06",
          6816 => x"56",
          6817 => x"38",
          6818 => x"80",
          6819 => x"81",
          6820 => x"52",
          6821 => x"51",
          6822 => x"82",
          6823 => x"81",
          6824 => x"81",
          6825 => x"83",
          6826 => x"87",
          6827 => x"2e",
          6828 => x"82",
          6829 => x"06",
          6830 => x"56",
          6831 => x"38",
          6832 => x"74",
          6833 => x"a3",
          6834 => x"dc",
          6835 => x"06",
          6836 => x"2e",
          6837 => x"80",
          6838 => x"3d",
          6839 => x"83",
          6840 => x"15",
          6841 => x"53",
          6842 => x"8d",
          6843 => x"15",
          6844 => x"3f",
          6845 => x"08",
          6846 => x"70",
          6847 => x"0c",
          6848 => x"16",
          6849 => x"80",
          6850 => x"80",
          6851 => x"54",
          6852 => x"84",
          6853 => x"5b",
          6854 => x"80",
          6855 => x"7a",
          6856 => x"fc",
          6857 => x"bb",
          6858 => x"ff",
          6859 => x"77",
          6860 => x"81",
          6861 => x"76",
          6862 => x"81",
          6863 => x"2e",
          6864 => x"8d",
          6865 => x"26",
          6866 => x"bf",
          6867 => x"f4",
          6868 => x"dc",
          6869 => x"ff",
          6870 => x"84",
          6871 => x"81",
          6872 => x"38",
          6873 => x"51",
          6874 => x"82",
          6875 => x"83",
          6876 => x"58",
          6877 => x"80",
          6878 => x"db",
          6879 => x"bb",
          6880 => x"77",
          6881 => x"80",
          6882 => x"82",
          6883 => x"c4",
          6884 => x"11",
          6885 => x"06",
          6886 => x"8d",
          6887 => x"26",
          6888 => x"74",
          6889 => x"78",
          6890 => x"c1",
          6891 => x"59",
          6892 => x"15",
          6893 => x"2e",
          6894 => x"13",
          6895 => x"72",
          6896 => x"38",
          6897 => x"eb",
          6898 => x"14",
          6899 => x"3f",
          6900 => x"08",
          6901 => x"dc",
          6902 => x"23",
          6903 => x"57",
          6904 => x"83",
          6905 => x"c7",
          6906 => x"d8",
          6907 => x"dc",
          6908 => x"ff",
          6909 => x"8d",
          6910 => x"14",
          6911 => x"3f",
          6912 => x"08",
          6913 => x"14",
          6914 => x"3f",
          6915 => x"08",
          6916 => x"06",
          6917 => x"72",
          6918 => x"97",
          6919 => x"22",
          6920 => x"84",
          6921 => x"5a",
          6922 => x"83",
          6923 => x"14",
          6924 => x"79",
          6925 => x"ee",
          6926 => x"bb",
          6927 => x"82",
          6928 => x"80",
          6929 => x"38",
          6930 => x"08",
          6931 => x"ff",
          6932 => x"38",
          6933 => x"83",
          6934 => x"83",
          6935 => x"74",
          6936 => x"85",
          6937 => x"89",
          6938 => x"76",
          6939 => x"c3",
          6940 => x"70",
          6941 => x"7b",
          6942 => x"73",
          6943 => x"17",
          6944 => x"ac",
          6945 => x"55",
          6946 => x"09",
          6947 => x"38",
          6948 => x"51",
          6949 => x"82",
          6950 => x"83",
          6951 => x"53",
          6952 => x"82",
          6953 => x"82",
          6954 => x"e0",
          6955 => x"ab",
          6956 => x"dc",
          6957 => x"0c",
          6958 => x"53",
          6959 => x"56",
          6960 => x"81",
          6961 => x"13",
          6962 => x"74",
          6963 => x"82",
          6964 => x"74",
          6965 => x"81",
          6966 => x"06",
          6967 => x"83",
          6968 => x"2a",
          6969 => x"72",
          6970 => x"26",
          6971 => x"ff",
          6972 => x"0c",
          6973 => x"15",
          6974 => x"0b",
          6975 => x"76",
          6976 => x"81",
          6977 => x"38",
          6978 => x"51",
          6979 => x"82",
          6980 => x"83",
          6981 => x"53",
          6982 => x"09",
          6983 => x"f9",
          6984 => x"52",
          6985 => x"b8",
          6986 => x"dc",
          6987 => x"38",
          6988 => x"08",
          6989 => x"84",
          6990 => x"d8",
          6991 => x"bb",
          6992 => x"ff",
          6993 => x"72",
          6994 => x"2e",
          6995 => x"80",
          6996 => x"14",
          6997 => x"3f",
          6998 => x"08",
          6999 => x"a4",
          7000 => x"81",
          7001 => x"84",
          7002 => x"d7",
          7003 => x"bb",
          7004 => x"8a",
          7005 => x"2e",
          7006 => x"9d",
          7007 => x"14",
          7008 => x"3f",
          7009 => x"08",
          7010 => x"84",
          7011 => x"d7",
          7012 => x"bb",
          7013 => x"15",
          7014 => x"34",
          7015 => x"22",
          7016 => x"72",
          7017 => x"23",
          7018 => x"23",
          7019 => x"15",
          7020 => x"75",
          7021 => x"0c",
          7022 => x"04",
          7023 => x"77",
          7024 => x"73",
          7025 => x"38",
          7026 => x"72",
          7027 => x"38",
          7028 => x"71",
          7029 => x"38",
          7030 => x"84",
          7031 => x"52",
          7032 => x"09",
          7033 => x"38",
          7034 => x"51",
          7035 => x"82",
          7036 => x"81",
          7037 => x"88",
          7038 => x"08",
          7039 => x"39",
          7040 => x"73",
          7041 => x"74",
          7042 => x"0c",
          7043 => x"04",
          7044 => x"02",
          7045 => x"7a",
          7046 => x"fc",
          7047 => x"f4",
          7048 => x"54",
          7049 => x"bb",
          7050 => x"bc",
          7051 => x"dc",
          7052 => x"82",
          7053 => x"70",
          7054 => x"73",
          7055 => x"38",
          7056 => x"78",
          7057 => x"2e",
          7058 => x"74",
          7059 => x"0c",
          7060 => x"80",
          7061 => x"80",
          7062 => x"70",
          7063 => x"51",
          7064 => x"82",
          7065 => x"54",
          7066 => x"dc",
          7067 => x"0d",
          7068 => x"0d",
          7069 => x"05",
          7070 => x"33",
          7071 => x"54",
          7072 => x"84",
          7073 => x"bf",
          7074 => x"98",
          7075 => x"53",
          7076 => x"05",
          7077 => x"fa",
          7078 => x"dc",
          7079 => x"bb",
          7080 => x"a4",
          7081 => x"68",
          7082 => x"70",
          7083 => x"c6",
          7084 => x"dc",
          7085 => x"bb",
          7086 => x"38",
          7087 => x"05",
          7088 => x"2b",
          7089 => x"80",
          7090 => x"86",
          7091 => x"06",
          7092 => x"2e",
          7093 => x"74",
          7094 => x"38",
          7095 => x"09",
          7096 => x"38",
          7097 => x"f8",
          7098 => x"dc",
          7099 => x"39",
          7100 => x"33",
          7101 => x"73",
          7102 => x"77",
          7103 => x"81",
          7104 => x"73",
          7105 => x"38",
          7106 => x"bc",
          7107 => x"07",
          7108 => x"b4",
          7109 => x"2a",
          7110 => x"51",
          7111 => x"2e",
          7112 => x"62",
          7113 => x"e8",
          7114 => x"bb",
          7115 => x"82",
          7116 => x"52",
          7117 => x"51",
          7118 => x"62",
          7119 => x"8b",
          7120 => x"53",
          7121 => x"51",
          7122 => x"80",
          7123 => x"05",
          7124 => x"3f",
          7125 => x"0b",
          7126 => x"75",
          7127 => x"f1",
          7128 => x"11",
          7129 => x"80",
          7130 => x"97",
          7131 => x"51",
          7132 => x"82",
          7133 => x"55",
          7134 => x"08",
          7135 => x"b7",
          7136 => x"c4",
          7137 => x"05",
          7138 => x"2a",
          7139 => x"51",
          7140 => x"80",
          7141 => x"84",
          7142 => x"39",
          7143 => x"70",
          7144 => x"54",
          7145 => x"a9",
          7146 => x"06",
          7147 => x"2e",
          7148 => x"55",
          7149 => x"73",
          7150 => x"d6",
          7151 => x"bb",
          7152 => x"ff",
          7153 => x"0c",
          7154 => x"bb",
          7155 => x"f8",
          7156 => x"2a",
          7157 => x"51",
          7158 => x"2e",
          7159 => x"80",
          7160 => x"7a",
          7161 => x"a0",
          7162 => x"a4",
          7163 => x"53",
          7164 => x"e6",
          7165 => x"bb",
          7166 => x"bb",
          7167 => x"1b",
          7168 => x"05",
          7169 => x"d3",
          7170 => x"dc",
          7171 => x"dc",
          7172 => x"0c",
          7173 => x"56",
          7174 => x"84",
          7175 => x"90",
          7176 => x"0b",
          7177 => x"80",
          7178 => x"0c",
          7179 => x"1a",
          7180 => x"2a",
          7181 => x"51",
          7182 => x"2e",
          7183 => x"82",
          7184 => x"80",
          7185 => x"38",
          7186 => x"08",
          7187 => x"8a",
          7188 => x"89",
          7189 => x"59",
          7190 => x"76",
          7191 => x"d7",
          7192 => x"bb",
          7193 => x"82",
          7194 => x"81",
          7195 => x"82",
          7196 => x"dc",
          7197 => x"09",
          7198 => x"38",
          7199 => x"78",
          7200 => x"30",
          7201 => x"80",
          7202 => x"77",
          7203 => x"38",
          7204 => x"06",
          7205 => x"c3",
          7206 => x"1a",
          7207 => x"38",
          7208 => x"06",
          7209 => x"2e",
          7210 => x"52",
          7211 => x"a6",
          7212 => x"dc",
          7213 => x"82",
          7214 => x"75",
          7215 => x"bb",
          7216 => x"9c",
          7217 => x"39",
          7218 => x"74",
          7219 => x"bb",
          7220 => x"3d",
          7221 => x"3d",
          7222 => x"65",
          7223 => x"5d",
          7224 => x"0c",
          7225 => x"05",
          7226 => x"f9",
          7227 => x"bb",
          7228 => x"82",
          7229 => x"8a",
          7230 => x"33",
          7231 => x"2e",
          7232 => x"56",
          7233 => x"90",
          7234 => x"06",
          7235 => x"74",
          7236 => x"b6",
          7237 => x"82",
          7238 => x"34",
          7239 => x"aa",
          7240 => x"91",
          7241 => x"56",
          7242 => x"8c",
          7243 => x"1a",
          7244 => x"74",
          7245 => x"38",
          7246 => x"80",
          7247 => x"38",
          7248 => x"70",
          7249 => x"56",
          7250 => x"b2",
          7251 => x"11",
          7252 => x"77",
          7253 => x"5b",
          7254 => x"38",
          7255 => x"88",
          7256 => x"8f",
          7257 => x"08",
          7258 => x"d5",
          7259 => x"bb",
          7260 => x"81",
          7261 => x"9f",
          7262 => x"2e",
          7263 => x"74",
          7264 => x"98",
          7265 => x"7e",
          7266 => x"3f",
          7267 => x"08",
          7268 => x"83",
          7269 => x"dc",
          7270 => x"89",
          7271 => x"77",
          7272 => x"d6",
          7273 => x"7f",
          7274 => x"58",
          7275 => x"75",
          7276 => x"75",
          7277 => x"77",
          7278 => x"7c",
          7279 => x"33",
          7280 => x"3f",
          7281 => x"08",
          7282 => x"7e",
          7283 => x"56",
          7284 => x"2e",
          7285 => x"16",
          7286 => x"55",
          7287 => x"94",
          7288 => x"53",
          7289 => x"b0",
          7290 => x"31",
          7291 => x"05",
          7292 => x"3f",
          7293 => x"56",
          7294 => x"9c",
          7295 => x"19",
          7296 => x"06",
          7297 => x"31",
          7298 => x"76",
          7299 => x"7b",
          7300 => x"08",
          7301 => x"d1",
          7302 => x"bb",
          7303 => x"81",
          7304 => x"94",
          7305 => x"ff",
          7306 => x"05",
          7307 => x"cf",
          7308 => x"76",
          7309 => x"17",
          7310 => x"1e",
          7311 => x"18",
          7312 => x"5e",
          7313 => x"39",
          7314 => x"82",
          7315 => x"90",
          7316 => x"f2",
          7317 => x"63",
          7318 => x"40",
          7319 => x"7e",
          7320 => x"fc",
          7321 => x"51",
          7322 => x"82",
          7323 => x"55",
          7324 => x"08",
          7325 => x"18",
          7326 => x"80",
          7327 => x"74",
          7328 => x"39",
          7329 => x"70",
          7330 => x"81",
          7331 => x"56",
          7332 => x"80",
          7333 => x"38",
          7334 => x"0b",
          7335 => x"82",
          7336 => x"39",
          7337 => x"19",
          7338 => x"83",
          7339 => x"18",
          7340 => x"56",
          7341 => x"27",
          7342 => x"09",
          7343 => x"2e",
          7344 => x"94",
          7345 => x"83",
          7346 => x"56",
          7347 => x"38",
          7348 => x"22",
          7349 => x"89",
          7350 => x"55",
          7351 => x"75",
          7352 => x"18",
          7353 => x"9c",
          7354 => x"85",
          7355 => x"08",
          7356 => x"d7",
          7357 => x"bb",
          7358 => x"82",
          7359 => x"80",
          7360 => x"38",
          7361 => x"ff",
          7362 => x"ff",
          7363 => x"38",
          7364 => x"0c",
          7365 => x"85",
          7366 => x"19",
          7367 => x"b0",
          7368 => x"19",
          7369 => x"81",
          7370 => x"74",
          7371 => x"3f",
          7372 => x"08",
          7373 => x"98",
          7374 => x"7e",
          7375 => x"3f",
          7376 => x"08",
          7377 => x"d2",
          7378 => x"dc",
          7379 => x"89",
          7380 => x"78",
          7381 => x"d5",
          7382 => x"7f",
          7383 => x"58",
          7384 => x"75",
          7385 => x"75",
          7386 => x"78",
          7387 => x"7c",
          7388 => x"33",
          7389 => x"3f",
          7390 => x"08",
          7391 => x"7e",
          7392 => x"78",
          7393 => x"74",
          7394 => x"38",
          7395 => x"b0",
          7396 => x"31",
          7397 => x"05",
          7398 => x"51",
          7399 => x"7e",
          7400 => x"83",
          7401 => x"89",
          7402 => x"db",
          7403 => x"08",
          7404 => x"26",
          7405 => x"51",
          7406 => x"82",
          7407 => x"fd",
          7408 => x"77",
          7409 => x"55",
          7410 => x"0c",
          7411 => x"83",
          7412 => x"80",
          7413 => x"55",
          7414 => x"83",
          7415 => x"9c",
          7416 => x"7e",
          7417 => x"3f",
          7418 => x"08",
          7419 => x"75",
          7420 => x"94",
          7421 => x"ff",
          7422 => x"05",
          7423 => x"3f",
          7424 => x"0b",
          7425 => x"7b",
          7426 => x"08",
          7427 => x"76",
          7428 => x"08",
          7429 => x"1c",
          7430 => x"08",
          7431 => x"5c",
          7432 => x"83",
          7433 => x"74",
          7434 => x"fd",
          7435 => x"18",
          7436 => x"07",
          7437 => x"19",
          7438 => x"75",
          7439 => x"0c",
          7440 => x"04",
          7441 => x"7a",
          7442 => x"05",
          7443 => x"56",
          7444 => x"82",
          7445 => x"57",
          7446 => x"08",
          7447 => x"90",
          7448 => x"86",
          7449 => x"06",
          7450 => x"73",
          7451 => x"e9",
          7452 => x"08",
          7453 => x"cc",
          7454 => x"bb",
          7455 => x"82",
          7456 => x"80",
          7457 => x"16",
          7458 => x"33",
          7459 => x"55",
          7460 => x"34",
          7461 => x"53",
          7462 => x"08",
          7463 => x"3f",
          7464 => x"52",
          7465 => x"c9",
          7466 => x"88",
          7467 => x"96",
          7468 => x"f0",
          7469 => x"92",
          7470 => x"ca",
          7471 => x"81",
          7472 => x"34",
          7473 => x"df",
          7474 => x"dc",
          7475 => x"33",
          7476 => x"55",
          7477 => x"17",
          7478 => x"bb",
          7479 => x"3d",
          7480 => x"3d",
          7481 => x"52",
          7482 => x"3f",
          7483 => x"08",
          7484 => x"dc",
          7485 => x"86",
          7486 => x"52",
          7487 => x"bc",
          7488 => x"dc",
          7489 => x"bb",
          7490 => x"38",
          7491 => x"08",
          7492 => x"82",
          7493 => x"86",
          7494 => x"ff",
          7495 => x"3d",
          7496 => x"3f",
          7497 => x"0b",
          7498 => x"08",
          7499 => x"82",
          7500 => x"82",
          7501 => x"80",
          7502 => x"bb",
          7503 => x"3d",
          7504 => x"3d",
          7505 => x"93",
          7506 => x"52",
          7507 => x"e9",
          7508 => x"bb",
          7509 => x"82",
          7510 => x"80",
          7511 => x"58",
          7512 => x"3d",
          7513 => x"e0",
          7514 => x"bb",
          7515 => x"82",
          7516 => x"bc",
          7517 => x"c7",
          7518 => x"98",
          7519 => x"73",
          7520 => x"38",
          7521 => x"12",
          7522 => x"39",
          7523 => x"33",
          7524 => x"70",
          7525 => x"55",
          7526 => x"2e",
          7527 => x"7f",
          7528 => x"54",
          7529 => x"82",
          7530 => x"94",
          7531 => x"39",
          7532 => x"08",
          7533 => x"81",
          7534 => x"85",
          7535 => x"bb",
          7536 => x"3d",
          7537 => x"3d",
          7538 => x"5b",
          7539 => x"34",
          7540 => x"3d",
          7541 => x"52",
          7542 => x"e8",
          7543 => x"bb",
          7544 => x"82",
          7545 => x"82",
          7546 => x"43",
          7547 => x"11",
          7548 => x"58",
          7549 => x"80",
          7550 => x"38",
          7551 => x"3d",
          7552 => x"d5",
          7553 => x"bb",
          7554 => x"82",
          7555 => x"82",
          7556 => x"52",
          7557 => x"c8",
          7558 => x"dc",
          7559 => x"bb",
          7560 => x"c1",
          7561 => x"7b",
          7562 => x"3f",
          7563 => x"08",
          7564 => x"74",
          7565 => x"3f",
          7566 => x"08",
          7567 => x"dc",
          7568 => x"38",
          7569 => x"51",
          7570 => x"82",
          7571 => x"57",
          7572 => x"08",
          7573 => x"52",
          7574 => x"f2",
          7575 => x"bb",
          7576 => x"a6",
          7577 => x"74",
          7578 => x"3f",
          7579 => x"08",
          7580 => x"dc",
          7581 => x"cc",
          7582 => x"2e",
          7583 => x"86",
          7584 => x"81",
          7585 => x"81",
          7586 => x"3d",
          7587 => x"52",
          7588 => x"c9",
          7589 => x"3d",
          7590 => x"11",
          7591 => x"5a",
          7592 => x"2e",
          7593 => x"b9",
          7594 => x"16",
          7595 => x"33",
          7596 => x"73",
          7597 => x"16",
          7598 => x"26",
          7599 => x"75",
          7600 => x"38",
          7601 => x"05",
          7602 => x"6f",
          7603 => x"ff",
          7604 => x"55",
          7605 => x"74",
          7606 => x"38",
          7607 => x"11",
          7608 => x"74",
          7609 => x"39",
          7610 => x"09",
          7611 => x"38",
          7612 => x"11",
          7613 => x"74",
          7614 => x"82",
          7615 => x"70",
          7616 => x"b5",
          7617 => x"08",
          7618 => x"5c",
          7619 => x"73",
          7620 => x"38",
          7621 => x"1a",
          7622 => x"55",
          7623 => x"38",
          7624 => x"73",
          7625 => x"38",
          7626 => x"76",
          7627 => x"74",
          7628 => x"33",
          7629 => x"05",
          7630 => x"15",
          7631 => x"ba",
          7632 => x"05",
          7633 => x"ff",
          7634 => x"06",
          7635 => x"57",
          7636 => x"18",
          7637 => x"54",
          7638 => x"70",
          7639 => x"34",
          7640 => x"ee",
          7641 => x"34",
          7642 => x"dc",
          7643 => x"0d",
          7644 => x"0d",
          7645 => x"3d",
          7646 => x"71",
          7647 => x"ec",
          7648 => x"bb",
          7649 => x"82",
          7650 => x"82",
          7651 => x"15",
          7652 => x"82",
          7653 => x"15",
          7654 => x"76",
          7655 => x"90",
          7656 => x"81",
          7657 => x"06",
          7658 => x"72",
          7659 => x"56",
          7660 => x"54",
          7661 => x"17",
          7662 => x"78",
          7663 => x"38",
          7664 => x"22",
          7665 => x"59",
          7666 => x"78",
          7667 => x"76",
          7668 => x"51",
          7669 => x"3f",
          7670 => x"08",
          7671 => x"54",
          7672 => x"53",
          7673 => x"3f",
          7674 => x"08",
          7675 => x"38",
          7676 => x"75",
          7677 => x"18",
          7678 => x"31",
          7679 => x"57",
          7680 => x"b1",
          7681 => x"08",
          7682 => x"38",
          7683 => x"51",
          7684 => x"82",
          7685 => x"54",
          7686 => x"08",
          7687 => x"9a",
          7688 => x"dc",
          7689 => x"81",
          7690 => x"bb",
          7691 => x"16",
          7692 => x"16",
          7693 => x"2e",
          7694 => x"76",
          7695 => x"dc",
          7696 => x"31",
          7697 => x"18",
          7698 => x"90",
          7699 => x"81",
          7700 => x"06",
          7701 => x"56",
          7702 => x"9a",
          7703 => x"74",
          7704 => x"3f",
          7705 => x"08",
          7706 => x"dc",
          7707 => x"82",
          7708 => x"56",
          7709 => x"52",
          7710 => x"84",
          7711 => x"dc",
          7712 => x"ff",
          7713 => x"81",
          7714 => x"38",
          7715 => x"98",
          7716 => x"a6",
          7717 => x"16",
          7718 => x"39",
          7719 => x"16",
          7720 => x"75",
          7721 => x"53",
          7722 => x"aa",
          7723 => x"79",
          7724 => x"3f",
          7725 => x"08",
          7726 => x"0b",
          7727 => x"82",
          7728 => x"39",
          7729 => x"16",
          7730 => x"bb",
          7731 => x"2a",
          7732 => x"08",
          7733 => x"15",
          7734 => x"15",
          7735 => x"90",
          7736 => x"16",
          7737 => x"33",
          7738 => x"53",
          7739 => x"34",
          7740 => x"06",
          7741 => x"2e",
          7742 => x"9c",
          7743 => x"85",
          7744 => x"16",
          7745 => x"72",
          7746 => x"0c",
          7747 => x"04",
          7748 => x"79",
          7749 => x"75",
          7750 => x"8a",
          7751 => x"89",
          7752 => x"52",
          7753 => x"05",
          7754 => x"3f",
          7755 => x"08",
          7756 => x"dc",
          7757 => x"38",
          7758 => x"7a",
          7759 => x"d8",
          7760 => x"bb",
          7761 => x"82",
          7762 => x"80",
          7763 => x"16",
          7764 => x"2b",
          7765 => x"74",
          7766 => x"86",
          7767 => x"84",
          7768 => x"06",
          7769 => x"73",
          7770 => x"38",
          7771 => x"52",
          7772 => x"da",
          7773 => x"dc",
          7774 => x"0c",
          7775 => x"14",
          7776 => x"23",
          7777 => x"51",
          7778 => x"82",
          7779 => x"55",
          7780 => x"09",
          7781 => x"38",
          7782 => x"39",
          7783 => x"84",
          7784 => x"0c",
          7785 => x"82",
          7786 => x"89",
          7787 => x"fc",
          7788 => x"87",
          7789 => x"53",
          7790 => x"e7",
          7791 => x"bb",
          7792 => x"38",
          7793 => x"08",
          7794 => x"3d",
          7795 => x"3d",
          7796 => x"89",
          7797 => x"54",
          7798 => x"54",
          7799 => x"82",
          7800 => x"53",
          7801 => x"08",
          7802 => x"74",
          7803 => x"bb",
          7804 => x"73",
          7805 => x"3f",
          7806 => x"08",
          7807 => x"39",
          7808 => x"08",
          7809 => x"d3",
          7810 => x"bb",
          7811 => x"82",
          7812 => x"84",
          7813 => x"06",
          7814 => x"53",
          7815 => x"bb",
          7816 => x"38",
          7817 => x"51",
          7818 => x"72",
          7819 => x"cf",
          7820 => x"bb",
          7821 => x"32",
          7822 => x"72",
          7823 => x"70",
          7824 => x"08",
          7825 => x"54",
          7826 => x"bb",
          7827 => x"3d",
          7828 => x"3d",
          7829 => x"80",
          7830 => x"70",
          7831 => x"52",
          7832 => x"3f",
          7833 => x"08",
          7834 => x"dc",
          7835 => x"64",
          7836 => x"d6",
          7837 => x"bb",
          7838 => x"82",
          7839 => x"a0",
          7840 => x"cb",
          7841 => x"98",
          7842 => x"73",
          7843 => x"38",
          7844 => x"39",
          7845 => x"88",
          7846 => x"75",
          7847 => x"3f",
          7848 => x"dc",
          7849 => x"0d",
          7850 => x"0d",
          7851 => x"5c",
          7852 => x"3d",
          7853 => x"93",
          7854 => x"d6",
          7855 => x"dc",
          7856 => x"bb",
          7857 => x"80",
          7858 => x"0c",
          7859 => x"11",
          7860 => x"90",
          7861 => x"56",
          7862 => x"74",
          7863 => x"75",
          7864 => x"e4",
          7865 => x"81",
          7866 => x"5b",
          7867 => x"82",
          7868 => x"75",
          7869 => x"73",
          7870 => x"81",
          7871 => x"82",
          7872 => x"76",
          7873 => x"f0",
          7874 => x"f4",
          7875 => x"dc",
          7876 => x"d1",
          7877 => x"dc",
          7878 => x"ce",
          7879 => x"dc",
          7880 => x"82",
          7881 => x"07",
          7882 => x"05",
          7883 => x"53",
          7884 => x"98",
          7885 => x"26",
          7886 => x"f9",
          7887 => x"08",
          7888 => x"08",
          7889 => x"98",
          7890 => x"81",
          7891 => x"58",
          7892 => x"3f",
          7893 => x"08",
          7894 => x"dc",
          7895 => x"38",
          7896 => x"77",
          7897 => x"5d",
          7898 => x"74",
          7899 => x"81",
          7900 => x"b4",
          7901 => x"bb",
          7902 => x"bb",
          7903 => x"ff",
          7904 => x"30",
          7905 => x"1b",
          7906 => x"5b",
          7907 => x"39",
          7908 => x"ff",
          7909 => x"82",
          7910 => x"f0",
          7911 => x"30",
          7912 => x"1b",
          7913 => x"5b",
          7914 => x"83",
          7915 => x"58",
          7916 => x"92",
          7917 => x"0c",
          7918 => x"12",
          7919 => x"33",
          7920 => x"54",
          7921 => x"34",
          7922 => x"dc",
          7923 => x"0d",
          7924 => x"0d",
          7925 => x"fc",
          7926 => x"52",
          7927 => x"3f",
          7928 => x"08",
          7929 => x"dc",
          7930 => x"38",
          7931 => x"56",
          7932 => x"38",
          7933 => x"70",
          7934 => x"81",
          7935 => x"55",
          7936 => x"80",
          7937 => x"38",
          7938 => x"54",
          7939 => x"08",
          7940 => x"38",
          7941 => x"82",
          7942 => x"53",
          7943 => x"52",
          7944 => x"8c",
          7945 => x"dc",
          7946 => x"19",
          7947 => x"c9",
          7948 => x"08",
          7949 => x"ff",
          7950 => x"82",
          7951 => x"ff",
          7952 => x"06",
          7953 => x"56",
          7954 => x"08",
          7955 => x"81",
          7956 => x"82",
          7957 => x"75",
          7958 => x"54",
          7959 => x"08",
          7960 => x"27",
          7961 => x"17",
          7962 => x"bb",
          7963 => x"76",
          7964 => x"3f",
          7965 => x"08",
          7966 => x"08",
          7967 => x"90",
          7968 => x"c0",
          7969 => x"90",
          7970 => x"80",
          7971 => x"75",
          7972 => x"75",
          7973 => x"bb",
          7974 => x"3d",
          7975 => x"3d",
          7976 => x"a0",
          7977 => x"05",
          7978 => x"51",
          7979 => x"82",
          7980 => x"55",
          7981 => x"08",
          7982 => x"78",
          7983 => x"08",
          7984 => x"70",
          7985 => x"ae",
          7986 => x"dc",
          7987 => x"bb",
          7988 => x"db",
          7989 => x"fb",
          7990 => x"85",
          7991 => x"06",
          7992 => x"86",
          7993 => x"c7",
          7994 => x"2b",
          7995 => x"24",
          7996 => x"02",
          7997 => x"33",
          7998 => x"58",
          7999 => x"76",
          8000 => x"6b",
          8001 => x"cc",
          8002 => x"bb",
          8003 => x"84",
          8004 => x"06",
          8005 => x"73",
          8006 => x"d4",
          8007 => x"82",
          8008 => x"94",
          8009 => x"81",
          8010 => x"5a",
          8011 => x"08",
          8012 => x"8a",
          8013 => x"54",
          8014 => x"82",
          8015 => x"55",
          8016 => x"08",
          8017 => x"82",
          8018 => x"52",
          8019 => x"e5",
          8020 => x"dc",
          8021 => x"bb",
          8022 => x"38",
          8023 => x"cf",
          8024 => x"dc",
          8025 => x"88",
          8026 => x"dc",
          8027 => x"38",
          8028 => x"c2",
          8029 => x"dc",
          8030 => x"dc",
          8031 => x"82",
          8032 => x"07",
          8033 => x"55",
          8034 => x"2e",
          8035 => x"80",
          8036 => x"80",
          8037 => x"77",
          8038 => x"3f",
          8039 => x"08",
          8040 => x"38",
          8041 => x"ba",
          8042 => x"bb",
          8043 => x"74",
          8044 => x"0c",
          8045 => x"04",
          8046 => x"82",
          8047 => x"c0",
          8048 => x"3d",
          8049 => x"3f",
          8050 => x"08",
          8051 => x"dc",
          8052 => x"38",
          8053 => x"52",
          8054 => x"52",
          8055 => x"3f",
          8056 => x"08",
          8057 => x"dc",
          8058 => x"88",
          8059 => x"39",
          8060 => x"08",
          8061 => x"81",
          8062 => x"38",
          8063 => x"05",
          8064 => x"2a",
          8065 => x"55",
          8066 => x"81",
          8067 => x"5a",
          8068 => x"3d",
          8069 => x"c1",
          8070 => x"bb",
          8071 => x"55",
          8072 => x"dc",
          8073 => x"87",
          8074 => x"dc",
          8075 => x"09",
          8076 => x"38",
          8077 => x"bb",
          8078 => x"2e",
          8079 => x"86",
          8080 => x"81",
          8081 => x"81",
          8082 => x"bb",
          8083 => x"78",
          8084 => x"3f",
          8085 => x"08",
          8086 => x"dc",
          8087 => x"38",
          8088 => x"52",
          8089 => x"ff",
          8090 => x"78",
          8091 => x"b4",
          8092 => x"54",
          8093 => x"15",
          8094 => x"b2",
          8095 => x"ca",
          8096 => x"b6",
          8097 => x"53",
          8098 => x"53",
          8099 => x"3f",
          8100 => x"b4",
          8101 => x"d4",
          8102 => x"b6",
          8103 => x"54",
          8104 => x"d5",
          8105 => x"53",
          8106 => x"11",
          8107 => x"d7",
          8108 => x"81",
          8109 => x"34",
          8110 => x"a4",
          8111 => x"dc",
          8112 => x"bb",
          8113 => x"38",
          8114 => x"0a",
          8115 => x"05",
          8116 => x"d0",
          8117 => x"64",
          8118 => x"c9",
          8119 => x"54",
          8120 => x"15",
          8121 => x"81",
          8122 => x"34",
          8123 => x"b8",
          8124 => x"bb",
          8125 => x"8b",
          8126 => x"75",
          8127 => x"ff",
          8128 => x"73",
          8129 => x"0c",
          8130 => x"04",
          8131 => x"a9",
          8132 => x"51",
          8133 => x"82",
          8134 => x"ff",
          8135 => x"a9",
          8136 => x"ee",
          8137 => x"dc",
          8138 => x"bb",
          8139 => x"d3",
          8140 => x"a9",
          8141 => x"9d",
          8142 => x"58",
          8143 => x"82",
          8144 => x"55",
          8145 => x"08",
          8146 => x"02",
          8147 => x"33",
          8148 => x"54",
          8149 => x"82",
          8150 => x"53",
          8151 => x"52",
          8152 => x"88",
          8153 => x"b4",
          8154 => x"53",
          8155 => x"3d",
          8156 => x"ff",
          8157 => x"aa",
          8158 => x"73",
          8159 => x"3f",
          8160 => x"08",
          8161 => x"dc",
          8162 => x"63",
          8163 => x"81",
          8164 => x"65",
          8165 => x"2e",
          8166 => x"55",
          8167 => x"82",
          8168 => x"84",
          8169 => x"06",
          8170 => x"73",
          8171 => x"3f",
          8172 => x"08",
          8173 => x"dc",
          8174 => x"38",
          8175 => x"53",
          8176 => x"95",
          8177 => x"16",
          8178 => x"87",
          8179 => x"05",
          8180 => x"34",
          8181 => x"70",
          8182 => x"81",
          8183 => x"55",
          8184 => x"74",
          8185 => x"73",
          8186 => x"78",
          8187 => x"83",
          8188 => x"16",
          8189 => x"2a",
          8190 => x"51",
          8191 => x"80",
          8192 => x"38",
          8193 => x"80",
          8194 => x"52",
          8195 => x"be",
          8196 => x"dc",
          8197 => x"51",
          8198 => x"3f",
          8199 => x"bb",
          8200 => x"2e",
          8201 => x"82",
          8202 => x"52",
          8203 => x"b5",
          8204 => x"bb",
          8205 => x"80",
          8206 => x"58",
          8207 => x"dc",
          8208 => x"38",
          8209 => x"54",
          8210 => x"09",
          8211 => x"38",
          8212 => x"52",
          8213 => x"af",
          8214 => x"81",
          8215 => x"34",
          8216 => x"bb",
          8217 => x"38",
          8218 => x"ca",
          8219 => x"dc",
          8220 => x"bb",
          8221 => x"38",
          8222 => x"b5",
          8223 => x"bb",
          8224 => x"74",
          8225 => x"0c",
          8226 => x"04",
          8227 => x"02",
          8228 => x"33",
          8229 => x"80",
          8230 => x"57",
          8231 => x"95",
          8232 => x"52",
          8233 => x"d2",
          8234 => x"bb",
          8235 => x"82",
          8236 => x"80",
          8237 => x"5a",
          8238 => x"3d",
          8239 => x"c9",
          8240 => x"bb",
          8241 => x"82",
          8242 => x"b8",
          8243 => x"cf",
          8244 => x"a0",
          8245 => x"55",
          8246 => x"75",
          8247 => x"71",
          8248 => x"33",
          8249 => x"74",
          8250 => x"57",
          8251 => x"8b",
          8252 => x"54",
          8253 => x"15",
          8254 => x"ff",
          8255 => x"82",
          8256 => x"55",
          8257 => x"dc",
          8258 => x"0d",
          8259 => x"0d",
          8260 => x"53",
          8261 => x"05",
          8262 => x"51",
          8263 => x"82",
          8264 => x"55",
          8265 => x"08",
          8266 => x"76",
          8267 => x"93",
          8268 => x"51",
          8269 => x"82",
          8270 => x"55",
          8271 => x"08",
          8272 => x"80",
          8273 => x"81",
          8274 => x"86",
          8275 => x"38",
          8276 => x"86",
          8277 => x"90",
          8278 => x"54",
          8279 => x"ff",
          8280 => x"76",
          8281 => x"83",
          8282 => x"51",
          8283 => x"3f",
          8284 => x"08",
          8285 => x"bb",
          8286 => x"3d",
          8287 => x"3d",
          8288 => x"5c",
          8289 => x"98",
          8290 => x"52",
          8291 => x"d1",
          8292 => x"bb",
          8293 => x"bb",
          8294 => x"70",
          8295 => x"08",
          8296 => x"51",
          8297 => x"80",
          8298 => x"38",
          8299 => x"06",
          8300 => x"80",
          8301 => x"38",
          8302 => x"5f",
          8303 => x"3d",
          8304 => x"ff",
          8305 => x"82",
          8306 => x"57",
          8307 => x"08",
          8308 => x"74",
          8309 => x"c3",
          8310 => x"bb",
          8311 => x"82",
          8312 => x"bf",
          8313 => x"dc",
          8314 => x"dc",
          8315 => x"59",
          8316 => x"81",
          8317 => x"56",
          8318 => x"33",
          8319 => x"16",
          8320 => x"27",
          8321 => x"56",
          8322 => x"80",
          8323 => x"80",
          8324 => x"ff",
          8325 => x"70",
          8326 => x"56",
          8327 => x"e8",
          8328 => x"76",
          8329 => x"81",
          8330 => x"80",
          8331 => x"57",
          8332 => x"78",
          8333 => x"51",
          8334 => x"2e",
          8335 => x"73",
          8336 => x"38",
          8337 => x"08",
          8338 => x"b1",
          8339 => x"bb",
          8340 => x"82",
          8341 => x"a7",
          8342 => x"33",
          8343 => x"c3",
          8344 => x"2e",
          8345 => x"e4",
          8346 => x"2e",
          8347 => x"56",
          8348 => x"05",
          8349 => x"e3",
          8350 => x"dc",
          8351 => x"76",
          8352 => x"0c",
          8353 => x"04",
          8354 => x"82",
          8355 => x"ff",
          8356 => x"9d",
          8357 => x"fa",
          8358 => x"dc",
          8359 => x"dc",
          8360 => x"82",
          8361 => x"83",
          8362 => x"53",
          8363 => x"3d",
          8364 => x"ff",
          8365 => x"73",
          8366 => x"70",
          8367 => x"52",
          8368 => x"9f",
          8369 => x"bc",
          8370 => x"74",
          8371 => x"6d",
          8372 => x"70",
          8373 => x"af",
          8374 => x"bb",
          8375 => x"2e",
          8376 => x"70",
          8377 => x"57",
          8378 => x"fd",
          8379 => x"dc",
          8380 => x"8d",
          8381 => x"2b",
          8382 => x"81",
          8383 => x"86",
          8384 => x"dc",
          8385 => x"9f",
          8386 => x"ff",
          8387 => x"54",
          8388 => x"8a",
          8389 => x"70",
          8390 => x"06",
          8391 => x"ff",
          8392 => x"38",
          8393 => x"15",
          8394 => x"80",
          8395 => x"74",
          8396 => x"a4",
          8397 => x"89",
          8398 => x"dc",
          8399 => x"81",
          8400 => x"88",
          8401 => x"26",
          8402 => x"39",
          8403 => x"86",
          8404 => x"81",
          8405 => x"ff",
          8406 => x"38",
          8407 => x"54",
          8408 => x"81",
          8409 => x"81",
          8410 => x"78",
          8411 => x"5a",
          8412 => x"6d",
          8413 => x"81",
          8414 => x"57",
          8415 => x"9f",
          8416 => x"38",
          8417 => x"54",
          8418 => x"81",
          8419 => x"b1",
          8420 => x"2e",
          8421 => x"a7",
          8422 => x"15",
          8423 => x"54",
          8424 => x"09",
          8425 => x"38",
          8426 => x"76",
          8427 => x"41",
          8428 => x"52",
          8429 => x"52",
          8430 => x"b3",
          8431 => x"dc",
          8432 => x"bb",
          8433 => x"f7",
          8434 => x"74",
          8435 => x"e5",
          8436 => x"dc",
          8437 => x"bb",
          8438 => x"38",
          8439 => x"38",
          8440 => x"74",
          8441 => x"39",
          8442 => x"08",
          8443 => x"81",
          8444 => x"38",
          8445 => x"74",
          8446 => x"38",
          8447 => x"51",
          8448 => x"3f",
          8449 => x"08",
          8450 => x"dc",
          8451 => x"a0",
          8452 => x"dc",
          8453 => x"51",
          8454 => x"3f",
          8455 => x"0b",
          8456 => x"8b",
          8457 => x"67",
          8458 => x"a7",
          8459 => x"81",
          8460 => x"34",
          8461 => x"ad",
          8462 => x"bb",
          8463 => x"73",
          8464 => x"bb",
          8465 => x"3d",
          8466 => x"3d",
          8467 => x"02",
          8468 => x"cb",
          8469 => x"3d",
          8470 => x"72",
          8471 => x"5a",
          8472 => x"82",
          8473 => x"58",
          8474 => x"08",
          8475 => x"91",
          8476 => x"77",
          8477 => x"7c",
          8478 => x"38",
          8479 => x"59",
          8480 => x"90",
          8481 => x"81",
          8482 => x"06",
          8483 => x"73",
          8484 => x"54",
          8485 => x"82",
          8486 => x"39",
          8487 => x"8b",
          8488 => x"11",
          8489 => x"2b",
          8490 => x"54",
          8491 => x"fe",
          8492 => x"ff",
          8493 => x"70",
          8494 => x"07",
          8495 => x"bb",
          8496 => x"8c",
          8497 => x"40",
          8498 => x"55",
          8499 => x"88",
          8500 => x"08",
          8501 => x"38",
          8502 => x"77",
          8503 => x"56",
          8504 => x"51",
          8505 => x"3f",
          8506 => x"55",
          8507 => x"08",
          8508 => x"38",
          8509 => x"bb",
          8510 => x"2e",
          8511 => x"82",
          8512 => x"ff",
          8513 => x"38",
          8514 => x"08",
          8515 => x"16",
          8516 => x"2e",
          8517 => x"87",
          8518 => x"74",
          8519 => x"74",
          8520 => x"81",
          8521 => x"38",
          8522 => x"ff",
          8523 => x"2e",
          8524 => x"7b",
          8525 => x"80",
          8526 => x"81",
          8527 => x"81",
          8528 => x"06",
          8529 => x"56",
          8530 => x"52",
          8531 => x"af",
          8532 => x"bb",
          8533 => x"82",
          8534 => x"80",
          8535 => x"81",
          8536 => x"56",
          8537 => x"d3",
          8538 => x"ff",
          8539 => x"7c",
          8540 => x"55",
          8541 => x"b3",
          8542 => x"1b",
          8543 => x"1b",
          8544 => x"33",
          8545 => x"54",
          8546 => x"34",
          8547 => x"fe",
          8548 => x"08",
          8549 => x"74",
          8550 => x"75",
          8551 => x"16",
          8552 => x"33",
          8553 => x"73",
          8554 => x"77",
          8555 => x"bb",
          8556 => x"3d",
          8557 => x"3d",
          8558 => x"02",
          8559 => x"eb",
          8560 => x"3d",
          8561 => x"59",
          8562 => x"8b",
          8563 => x"82",
          8564 => x"24",
          8565 => x"82",
          8566 => x"84",
          8567 => x"94",
          8568 => x"51",
          8569 => x"2e",
          8570 => x"75",
          8571 => x"dc",
          8572 => x"06",
          8573 => x"7e",
          8574 => x"d0",
          8575 => x"dc",
          8576 => x"06",
          8577 => x"56",
          8578 => x"74",
          8579 => x"76",
          8580 => x"81",
          8581 => x"8a",
          8582 => x"b2",
          8583 => x"fc",
          8584 => x"52",
          8585 => x"a4",
          8586 => x"bb",
          8587 => x"38",
          8588 => x"80",
          8589 => x"74",
          8590 => x"26",
          8591 => x"15",
          8592 => x"74",
          8593 => x"38",
          8594 => x"80",
          8595 => x"84",
          8596 => x"92",
          8597 => x"80",
          8598 => x"38",
          8599 => x"06",
          8600 => x"2e",
          8601 => x"56",
          8602 => x"78",
          8603 => x"89",
          8604 => x"2b",
          8605 => x"43",
          8606 => x"38",
          8607 => x"30",
          8608 => x"77",
          8609 => x"91",
          8610 => x"c2",
          8611 => x"f8",
          8612 => x"52",
          8613 => x"a4",
          8614 => x"56",
          8615 => x"08",
          8616 => x"77",
          8617 => x"77",
          8618 => x"dc",
          8619 => x"45",
          8620 => x"bf",
          8621 => x"8e",
          8622 => x"26",
          8623 => x"74",
          8624 => x"48",
          8625 => x"75",
          8626 => x"38",
          8627 => x"81",
          8628 => x"fa",
          8629 => x"2a",
          8630 => x"56",
          8631 => x"2e",
          8632 => x"87",
          8633 => x"82",
          8634 => x"38",
          8635 => x"55",
          8636 => x"83",
          8637 => x"81",
          8638 => x"56",
          8639 => x"80",
          8640 => x"38",
          8641 => x"83",
          8642 => x"06",
          8643 => x"78",
          8644 => x"91",
          8645 => x"0b",
          8646 => x"22",
          8647 => x"80",
          8648 => x"74",
          8649 => x"38",
          8650 => x"56",
          8651 => x"17",
          8652 => x"57",
          8653 => x"2e",
          8654 => x"75",
          8655 => x"79",
          8656 => x"fe",
          8657 => x"82",
          8658 => x"84",
          8659 => x"05",
          8660 => x"5e",
          8661 => x"80",
          8662 => x"dc",
          8663 => x"8a",
          8664 => x"fd",
          8665 => x"75",
          8666 => x"38",
          8667 => x"78",
          8668 => x"8c",
          8669 => x"0b",
          8670 => x"22",
          8671 => x"80",
          8672 => x"74",
          8673 => x"38",
          8674 => x"56",
          8675 => x"17",
          8676 => x"57",
          8677 => x"2e",
          8678 => x"75",
          8679 => x"79",
          8680 => x"fe",
          8681 => x"82",
          8682 => x"10",
          8683 => x"82",
          8684 => x"9f",
          8685 => x"38",
          8686 => x"bb",
          8687 => x"82",
          8688 => x"05",
          8689 => x"2a",
          8690 => x"56",
          8691 => x"17",
          8692 => x"81",
          8693 => x"60",
          8694 => x"65",
          8695 => x"12",
          8696 => x"30",
          8697 => x"74",
          8698 => x"59",
          8699 => x"7d",
          8700 => x"81",
          8701 => x"76",
          8702 => x"41",
          8703 => x"76",
          8704 => x"90",
          8705 => x"62",
          8706 => x"51",
          8707 => x"26",
          8708 => x"75",
          8709 => x"31",
          8710 => x"65",
          8711 => x"fe",
          8712 => x"82",
          8713 => x"58",
          8714 => x"09",
          8715 => x"38",
          8716 => x"08",
          8717 => x"26",
          8718 => x"78",
          8719 => x"79",
          8720 => x"78",
          8721 => x"86",
          8722 => x"82",
          8723 => x"06",
          8724 => x"83",
          8725 => x"82",
          8726 => x"27",
          8727 => x"8f",
          8728 => x"55",
          8729 => x"26",
          8730 => x"59",
          8731 => x"62",
          8732 => x"74",
          8733 => x"38",
          8734 => x"88",
          8735 => x"dc",
          8736 => x"26",
          8737 => x"86",
          8738 => x"1a",
          8739 => x"79",
          8740 => x"38",
          8741 => x"80",
          8742 => x"2e",
          8743 => x"83",
          8744 => x"9f",
          8745 => x"8b",
          8746 => x"06",
          8747 => x"74",
          8748 => x"84",
          8749 => x"52",
          8750 => x"a2",
          8751 => x"53",
          8752 => x"52",
          8753 => x"a2",
          8754 => x"80",
          8755 => x"51",
          8756 => x"3f",
          8757 => x"34",
          8758 => x"ff",
          8759 => x"1b",
          8760 => x"a2",
          8761 => x"90",
          8762 => x"83",
          8763 => x"70",
          8764 => x"80",
          8765 => x"55",
          8766 => x"ff",
          8767 => x"66",
          8768 => x"ff",
          8769 => x"38",
          8770 => x"ff",
          8771 => x"1b",
          8772 => x"f2",
          8773 => x"74",
          8774 => x"51",
          8775 => x"3f",
          8776 => x"1c",
          8777 => x"98",
          8778 => x"a0",
          8779 => x"ff",
          8780 => x"51",
          8781 => x"3f",
          8782 => x"1b",
          8783 => x"e4",
          8784 => x"2e",
          8785 => x"80",
          8786 => x"88",
          8787 => x"80",
          8788 => x"ff",
          8789 => x"7c",
          8790 => x"51",
          8791 => x"3f",
          8792 => x"1b",
          8793 => x"bc",
          8794 => x"b0",
          8795 => x"a0",
          8796 => x"52",
          8797 => x"ff",
          8798 => x"ff",
          8799 => x"c0",
          8800 => x"0b",
          8801 => x"34",
          8802 => x"b4",
          8803 => x"c7",
          8804 => x"39",
          8805 => x"0a",
          8806 => x"51",
          8807 => x"3f",
          8808 => x"ff",
          8809 => x"1b",
          8810 => x"da",
          8811 => x"0b",
          8812 => x"a9",
          8813 => x"34",
          8814 => x"b5",
          8815 => x"1b",
          8816 => x"8f",
          8817 => x"d5",
          8818 => x"1b",
          8819 => x"ff",
          8820 => x"81",
          8821 => x"7a",
          8822 => x"ff",
          8823 => x"81",
          8824 => x"dc",
          8825 => x"38",
          8826 => x"09",
          8827 => x"ee",
          8828 => x"60",
          8829 => x"7a",
          8830 => x"ff",
          8831 => x"84",
          8832 => x"52",
          8833 => x"9f",
          8834 => x"8b",
          8835 => x"52",
          8836 => x"9f",
          8837 => x"8a",
          8838 => x"52",
          8839 => x"51",
          8840 => x"3f",
          8841 => x"83",
          8842 => x"ff",
          8843 => x"82",
          8844 => x"1b",
          8845 => x"ec",
          8846 => x"d5",
          8847 => x"ff",
          8848 => x"75",
          8849 => x"05",
          8850 => x"7e",
          8851 => x"e5",
          8852 => x"60",
          8853 => x"52",
          8854 => x"9a",
          8855 => x"53",
          8856 => x"51",
          8857 => x"3f",
          8858 => x"58",
          8859 => x"09",
          8860 => x"38",
          8861 => x"51",
          8862 => x"3f",
          8863 => x"1b",
          8864 => x"a0",
          8865 => x"52",
          8866 => x"91",
          8867 => x"ff",
          8868 => x"81",
          8869 => x"f8",
          8870 => x"7a",
          8871 => x"84",
          8872 => x"61",
          8873 => x"26",
          8874 => x"57",
          8875 => x"53",
          8876 => x"51",
          8877 => x"3f",
          8878 => x"08",
          8879 => x"84",
          8880 => x"bb",
          8881 => x"7a",
          8882 => x"aa",
          8883 => x"75",
          8884 => x"56",
          8885 => x"81",
          8886 => x"80",
          8887 => x"38",
          8888 => x"83",
          8889 => x"63",
          8890 => x"74",
          8891 => x"38",
          8892 => x"54",
          8893 => x"52",
          8894 => x"99",
          8895 => x"bb",
          8896 => x"c1",
          8897 => x"75",
          8898 => x"56",
          8899 => x"8c",
          8900 => x"2e",
          8901 => x"56",
          8902 => x"ff",
          8903 => x"84",
          8904 => x"2e",
          8905 => x"56",
          8906 => x"58",
          8907 => x"38",
          8908 => x"77",
          8909 => x"ff",
          8910 => x"82",
          8911 => x"78",
          8912 => x"c2",
          8913 => x"1b",
          8914 => x"34",
          8915 => x"16",
          8916 => x"82",
          8917 => x"83",
          8918 => x"84",
          8919 => x"67",
          8920 => x"fd",
          8921 => x"51",
          8922 => x"3f",
          8923 => x"16",
          8924 => x"dc",
          8925 => x"bf",
          8926 => x"86",
          8927 => x"bb",
          8928 => x"16",
          8929 => x"83",
          8930 => x"ff",
          8931 => x"66",
          8932 => x"1b",
          8933 => x"8c",
          8934 => x"77",
          8935 => x"7e",
          8936 => x"91",
          8937 => x"82",
          8938 => x"a2",
          8939 => x"80",
          8940 => x"ff",
          8941 => x"81",
          8942 => x"dc",
          8943 => x"89",
          8944 => x"8a",
          8945 => x"86",
          8946 => x"dc",
          8947 => x"82",
          8948 => x"99",
          8949 => x"f5",
          8950 => x"60",
          8951 => x"79",
          8952 => x"5a",
          8953 => x"78",
          8954 => x"8d",
          8955 => x"55",
          8956 => x"fc",
          8957 => x"51",
          8958 => x"7a",
          8959 => x"81",
          8960 => x"8c",
          8961 => x"74",
          8962 => x"38",
          8963 => x"81",
          8964 => x"81",
          8965 => x"8a",
          8966 => x"06",
          8967 => x"76",
          8968 => x"76",
          8969 => x"55",
          8970 => x"dc",
          8971 => x"0d",
          8972 => x"0d",
          8973 => x"05",
          8974 => x"59",
          8975 => x"2e",
          8976 => x"87",
          8977 => x"76",
          8978 => x"84",
          8979 => x"80",
          8980 => x"38",
          8981 => x"77",
          8982 => x"56",
          8983 => x"34",
          8984 => x"bb",
          8985 => x"38",
          8986 => x"05",
          8987 => x"8c",
          8988 => x"08",
          8989 => x"3f",
          8990 => x"70",
          8991 => x"07",
          8992 => x"30",
          8993 => x"56",
          8994 => x"0c",
          8995 => x"18",
          8996 => x"0d",
          8997 => x"0d",
          8998 => x"08",
          8999 => x"75",
          9000 => x"89",
          9001 => x"54",
          9002 => x"16",
          9003 => x"51",
          9004 => x"82",
          9005 => x"91",
          9006 => x"08",
          9007 => x"81",
          9008 => x"88",
          9009 => x"83",
          9010 => x"74",
          9011 => x"0c",
          9012 => x"04",
          9013 => x"75",
          9014 => x"53",
          9015 => x"51",
          9016 => x"3f",
          9017 => x"85",
          9018 => x"ea",
          9019 => x"80",
          9020 => x"6a",
          9021 => x"70",
          9022 => x"d8",
          9023 => x"72",
          9024 => x"3f",
          9025 => x"8d",
          9026 => x"0d",
          9027 => x"ff",
          9028 => x"ff",
          9029 => x"00",
          9030 => x"ff",
          9031 => x"2b",
          9032 => x"2b",
          9033 => x"2b",
          9034 => x"2b",
          9035 => x"2b",
          9036 => x"2b",
          9037 => x"2b",
          9038 => x"2b",
          9039 => x"2b",
          9040 => x"2b",
          9041 => x"2b",
          9042 => x"2b",
          9043 => x"2b",
          9044 => x"2b",
          9045 => x"2b",
          9046 => x"2b",
          9047 => x"2b",
          9048 => x"2b",
          9049 => x"2b",
          9050 => x"2b",
          9051 => x"43",
          9052 => x"43",
          9053 => x"43",
          9054 => x"43",
          9055 => x"43",
          9056 => x"49",
          9057 => x"4a",
          9058 => x"4b",
          9059 => x"4e",
          9060 => x"4a",
          9061 => x"48",
          9062 => x"4c",
          9063 => x"4d",
          9064 => x"4c",
          9065 => x"4d",
          9066 => x"4c",
          9067 => x"4b",
          9068 => x"48",
          9069 => x"4b",
          9070 => x"4b",
          9071 => x"4c",
          9072 => x"48",
          9073 => x"48",
          9074 => x"4c",
          9075 => x"4d",
          9076 => x"4d",
          9077 => x"4e",
          9078 => x"0e",
          9079 => x"17",
          9080 => x"17",
          9081 => x"0e",
          9082 => x"17",
          9083 => x"17",
          9084 => x"17",
          9085 => x"17",
          9086 => x"17",
          9087 => x"17",
          9088 => x"17",
          9089 => x"0e",
          9090 => x"17",
          9091 => x"0e",
          9092 => x"0e",
          9093 => x"17",
          9094 => x"17",
          9095 => x"17",
          9096 => x"17",
          9097 => x"17",
          9098 => x"17",
          9099 => x"17",
          9100 => x"17",
          9101 => x"17",
          9102 => x"17",
          9103 => x"17",
          9104 => x"17",
          9105 => x"17",
          9106 => x"17",
          9107 => x"17",
          9108 => x"17",
          9109 => x"17",
          9110 => x"17",
          9111 => x"17",
          9112 => x"17",
          9113 => x"17",
          9114 => x"17",
          9115 => x"17",
          9116 => x"17",
          9117 => x"17",
          9118 => x"17",
          9119 => x"17",
          9120 => x"17",
          9121 => x"17",
          9122 => x"17",
          9123 => x"17",
          9124 => x"17",
          9125 => x"17",
          9126 => x"17",
          9127 => x"17",
          9128 => x"17",
          9129 => x"0f",
          9130 => x"17",
          9131 => x"17",
          9132 => x"17",
          9133 => x"17",
          9134 => x"11",
          9135 => x"17",
          9136 => x"17",
          9137 => x"17",
          9138 => x"17",
          9139 => x"17",
          9140 => x"17",
          9141 => x"17",
          9142 => x"17",
          9143 => x"17",
          9144 => x"17",
          9145 => x"0e",
          9146 => x"10",
          9147 => x"0e",
          9148 => x"0e",
          9149 => x"0e",
          9150 => x"17",
          9151 => x"10",
          9152 => x"17",
          9153 => x"17",
          9154 => x"0e",
          9155 => x"17",
          9156 => x"17",
          9157 => x"10",
          9158 => x"10",
          9159 => x"17",
          9160 => x"17",
          9161 => x"0f",
          9162 => x"17",
          9163 => x"11",
          9164 => x"17",
          9165 => x"17",
          9166 => x"11",
          9167 => x"6e",
          9168 => x"00",
          9169 => x"6f",
          9170 => x"00",
          9171 => x"6e",
          9172 => x"00",
          9173 => x"6f",
          9174 => x"00",
          9175 => x"78",
          9176 => x"00",
          9177 => x"6c",
          9178 => x"00",
          9179 => x"6f",
          9180 => x"00",
          9181 => x"69",
          9182 => x"00",
          9183 => x"75",
          9184 => x"00",
          9185 => x"62",
          9186 => x"68",
          9187 => x"77",
          9188 => x"64",
          9189 => x"65",
          9190 => x"64",
          9191 => x"65",
          9192 => x"6c",
          9193 => x"00",
          9194 => x"70",
          9195 => x"73",
          9196 => x"74",
          9197 => x"73",
          9198 => x"00",
          9199 => x"66",
          9200 => x"00",
          9201 => x"73",
          9202 => x"00",
          9203 => x"61",
          9204 => x"00",
          9205 => x"61",
          9206 => x"00",
          9207 => x"6c",
          9208 => x"00",
          9209 => x"00",
          9210 => x"73",
          9211 => x"72",
          9212 => x"00",
          9213 => x"74",
          9214 => x"61",
          9215 => x"72",
          9216 => x"2e",
          9217 => x"73",
          9218 => x"6f",
          9219 => x"65",
          9220 => x"2e",
          9221 => x"20",
          9222 => x"65",
          9223 => x"75",
          9224 => x"00",
          9225 => x"20",
          9226 => x"68",
          9227 => x"75",
          9228 => x"00",
          9229 => x"76",
          9230 => x"64",
          9231 => x"6c",
          9232 => x"6d",
          9233 => x"00",
          9234 => x"63",
          9235 => x"20",
          9236 => x"69",
          9237 => x"00",
          9238 => x"6c",
          9239 => x"6c",
          9240 => x"64",
          9241 => x"78",
          9242 => x"73",
          9243 => x"00",
          9244 => x"6c",
          9245 => x"61",
          9246 => x"65",
          9247 => x"76",
          9248 => x"64",
          9249 => x"00",
          9250 => x"20",
          9251 => x"77",
          9252 => x"65",
          9253 => x"6f",
          9254 => x"74",
          9255 => x"00",
          9256 => x"69",
          9257 => x"6e",
          9258 => x"65",
          9259 => x"73",
          9260 => x"76",
          9261 => x"64",
          9262 => x"00",
          9263 => x"73",
          9264 => x"6f",
          9265 => x"6e",
          9266 => x"65",
          9267 => x"00",
          9268 => x"20",
          9269 => x"70",
          9270 => x"62",
          9271 => x"66",
          9272 => x"73",
          9273 => x"65",
          9274 => x"6f",
          9275 => x"20",
          9276 => x"64",
          9277 => x"2e",
          9278 => x"72",
          9279 => x"20",
          9280 => x"72",
          9281 => x"2e",
          9282 => x"6d",
          9283 => x"74",
          9284 => x"70",
          9285 => x"74",
          9286 => x"20",
          9287 => x"63",
          9288 => x"65",
          9289 => x"00",
          9290 => x"6c",
          9291 => x"73",
          9292 => x"63",
          9293 => x"2e",
          9294 => x"73",
          9295 => x"69",
          9296 => x"6e",
          9297 => x"65",
          9298 => x"79",
          9299 => x"00",
          9300 => x"6f",
          9301 => x"6e",
          9302 => x"70",
          9303 => x"66",
          9304 => x"73",
          9305 => x"00",
          9306 => x"72",
          9307 => x"74",
          9308 => x"20",
          9309 => x"6f",
          9310 => x"63",
          9311 => x"00",
          9312 => x"63",
          9313 => x"73",
          9314 => x"00",
          9315 => x"6b",
          9316 => x"6e",
          9317 => x"72",
          9318 => x"00",
          9319 => x"6c",
          9320 => x"79",
          9321 => x"20",
          9322 => x"61",
          9323 => x"6c",
          9324 => x"79",
          9325 => x"2f",
          9326 => x"2e",
          9327 => x"00",
          9328 => x"61",
          9329 => x"00",
          9330 => x"38",
          9331 => x"00",
          9332 => x"20",
          9333 => x"34",
          9334 => x"00",
          9335 => x"20",
          9336 => x"20",
          9337 => x"00",
          9338 => x"32",
          9339 => x"00",
          9340 => x"00",
          9341 => x"00",
          9342 => x"00",
          9343 => x"55",
          9344 => x"00",
          9345 => x"2a",
          9346 => x"20",
          9347 => x"00",
          9348 => x"2f",
          9349 => x"32",
          9350 => x"00",
          9351 => x"2e",
          9352 => x"00",
          9353 => x"50",
          9354 => x"72",
          9355 => x"25",
          9356 => x"29",
          9357 => x"20",
          9358 => x"2a",
          9359 => x"00",
          9360 => x"55",
          9361 => x"49",
          9362 => x"72",
          9363 => x"74",
          9364 => x"6e",
          9365 => x"72",
          9366 => x"6d",
          9367 => x"69",
          9368 => x"72",
          9369 => x"74",
          9370 => x"32",
          9371 => x"74",
          9372 => x"75",
          9373 => x"00",
          9374 => x"43",
          9375 => x"52",
          9376 => x"6e",
          9377 => x"72",
          9378 => x"00",
          9379 => x"43",
          9380 => x"57",
          9381 => x"6e",
          9382 => x"72",
          9383 => x"00",
          9384 => x"52",
          9385 => x"52",
          9386 => x"6e",
          9387 => x"72",
          9388 => x"00",
          9389 => x"52",
          9390 => x"54",
          9391 => x"6e",
          9392 => x"72",
          9393 => x"00",
          9394 => x"52",
          9395 => x"52",
          9396 => x"6e",
          9397 => x"72",
          9398 => x"00",
          9399 => x"52",
          9400 => x"54",
          9401 => x"6e",
          9402 => x"72",
          9403 => x"00",
          9404 => x"74",
          9405 => x"67",
          9406 => x"20",
          9407 => x"65",
          9408 => x"2e",
          9409 => x"61",
          9410 => x"6e",
          9411 => x"69",
          9412 => x"2e",
          9413 => x"00",
          9414 => x"74",
          9415 => x"65",
          9416 => x"61",
          9417 => x"00",
          9418 => x"75",
          9419 => x"68",
          9420 => x"00",
          9421 => x"00",
          9422 => x"69",
          9423 => x"20",
          9424 => x"69",
          9425 => x"69",
          9426 => x"73",
          9427 => x"64",
          9428 => x"72",
          9429 => x"2c",
          9430 => x"65",
          9431 => x"20",
          9432 => x"74",
          9433 => x"6e",
          9434 => x"6c",
          9435 => x"00",
          9436 => x"00",
          9437 => x"64",
          9438 => x"73",
          9439 => x"64",
          9440 => x"00",
          9441 => x"69",
          9442 => x"6c",
          9443 => x"64",
          9444 => x"00",
          9445 => x"69",
          9446 => x"20",
          9447 => x"69",
          9448 => x"69",
          9449 => x"73",
          9450 => x"00",
          9451 => x"3d",
          9452 => x"00",
          9453 => x"3a",
          9454 => x"65",
          9455 => x"6e",
          9456 => x"2e",
          9457 => x"00",
          9458 => x"70",
          9459 => x"67",
          9460 => x"00",
          9461 => x"6d",
          9462 => x"69",
          9463 => x"2e",
          9464 => x"00",
          9465 => x"38",
          9466 => x"25",
          9467 => x"29",
          9468 => x"30",
          9469 => x"28",
          9470 => x"78",
          9471 => x"00",
          9472 => x"6d",
          9473 => x"65",
          9474 => x"79",
          9475 => x"6f",
          9476 => x"65",
          9477 => x"00",
          9478 => x"38",
          9479 => x"25",
          9480 => x"2d",
          9481 => x"3f",
          9482 => x"38",
          9483 => x"25",
          9484 => x"2d",
          9485 => x"38",
          9486 => x"25",
          9487 => x"58",
          9488 => x"00",
          9489 => x"73",
          9490 => x"69",
          9491 => x"69",
          9492 => x"72",
          9493 => x"74",
          9494 => x"00",
          9495 => x"61",
          9496 => x"6e",
          9497 => x"6e",
          9498 => x"72",
          9499 => x"73",
          9500 => x"73",
          9501 => x"65",
          9502 => x"61",
          9503 => x"66",
          9504 => x"00",
          9505 => x"61",
          9506 => x"6e",
          9507 => x"61",
          9508 => x"66",
          9509 => x"00",
          9510 => x"65",
          9511 => x"69",
          9512 => x"63",
          9513 => x"20",
          9514 => x"30",
          9515 => x"20",
          9516 => x"0a",
          9517 => x"6c",
          9518 => x"67",
          9519 => x"64",
          9520 => x"20",
          9521 => x"6c",
          9522 => x"2e",
          9523 => x"00",
          9524 => x"6c",
          9525 => x"65",
          9526 => x"6e",
          9527 => x"63",
          9528 => x"20",
          9529 => x"29",
          9530 => x"00",
          9531 => x"73",
          9532 => x"74",
          9533 => x"20",
          9534 => x"6c",
          9535 => x"74",
          9536 => x"2e",
          9537 => x"00",
          9538 => x"6c",
          9539 => x"65",
          9540 => x"74",
          9541 => x"2e",
          9542 => x"00",
          9543 => x"55",
          9544 => x"6e",
          9545 => x"3a",
          9546 => x"5c",
          9547 => x"25",
          9548 => x"00",
          9549 => x"3a",
          9550 => x"5c",
          9551 => x"00",
          9552 => x"3a",
          9553 => x"00",
          9554 => x"64",
          9555 => x"6d",
          9556 => x"64",
          9557 => x"00",
          9558 => x"6e",
          9559 => x"67",
          9560 => x"00",
          9561 => x"61",
          9562 => x"6e",
          9563 => x"6e",
          9564 => x"72",
          9565 => x"73",
          9566 => x"00",
          9567 => x"2f",
          9568 => x"25",
          9569 => x"64",
          9570 => x"3a",
          9571 => x"25",
          9572 => x"0a",
          9573 => x"43",
          9574 => x"6e",
          9575 => x"75",
          9576 => x"69",
          9577 => x"00",
          9578 => x"66",
          9579 => x"20",
          9580 => x"20",
          9581 => x"66",
          9582 => x"00",
          9583 => x"44",
          9584 => x"63",
          9585 => x"69",
          9586 => x"65",
          9587 => x"74",
          9588 => x"0a",
          9589 => x"20",
          9590 => x"20",
          9591 => x"41",
          9592 => x"28",
          9593 => x"58",
          9594 => x"38",
          9595 => x"0a",
          9596 => x"20",
          9597 => x"52",
          9598 => x"20",
          9599 => x"28",
          9600 => x"58",
          9601 => x"38",
          9602 => x"0a",
          9603 => x"20",
          9604 => x"53",
          9605 => x"52",
          9606 => x"28",
          9607 => x"58",
          9608 => x"38",
          9609 => x"0a",
          9610 => x"20",
          9611 => x"41",
          9612 => x"20",
          9613 => x"28",
          9614 => x"58",
          9615 => x"38",
          9616 => x"0a",
          9617 => x"20",
          9618 => x"4d",
          9619 => x"20",
          9620 => x"28",
          9621 => x"58",
          9622 => x"38",
          9623 => x"0a",
          9624 => x"20",
          9625 => x"20",
          9626 => x"44",
          9627 => x"28",
          9628 => x"69",
          9629 => x"20",
          9630 => x"32",
          9631 => x"0a",
          9632 => x"20",
          9633 => x"4d",
          9634 => x"20",
          9635 => x"28",
          9636 => x"65",
          9637 => x"20",
          9638 => x"32",
          9639 => x"0a",
          9640 => x"20",
          9641 => x"54",
          9642 => x"54",
          9643 => x"28",
          9644 => x"6e",
          9645 => x"73",
          9646 => x"32",
          9647 => x"0a",
          9648 => x"20",
          9649 => x"53",
          9650 => x"4e",
          9651 => x"55",
          9652 => x"00",
          9653 => x"20",
          9654 => x"20",
          9655 => x"0a",
          9656 => x"20",
          9657 => x"43",
          9658 => x"00",
          9659 => x"20",
          9660 => x"32",
          9661 => x"00",
          9662 => x"20",
          9663 => x"49",
          9664 => x"00",
          9665 => x"64",
          9666 => x"73",
          9667 => x"0a",
          9668 => x"20",
          9669 => x"55",
          9670 => x"73",
          9671 => x"56",
          9672 => x"6f",
          9673 => x"64",
          9674 => x"73",
          9675 => x"20",
          9676 => x"58",
          9677 => x"00",
          9678 => x"20",
          9679 => x"55",
          9680 => x"6d",
          9681 => x"20",
          9682 => x"72",
          9683 => x"64",
          9684 => x"73",
          9685 => x"20",
          9686 => x"58",
          9687 => x"00",
          9688 => x"20",
          9689 => x"61",
          9690 => x"53",
          9691 => x"74",
          9692 => x"64",
          9693 => x"73",
          9694 => x"20",
          9695 => x"20",
          9696 => x"58",
          9697 => x"00",
          9698 => x"73",
          9699 => x"00",
          9700 => x"20",
          9701 => x"55",
          9702 => x"20",
          9703 => x"20",
          9704 => x"20",
          9705 => x"20",
          9706 => x"20",
          9707 => x"20",
          9708 => x"58",
          9709 => x"00",
          9710 => x"20",
          9711 => x"73",
          9712 => x"20",
          9713 => x"63",
          9714 => x"72",
          9715 => x"20",
          9716 => x"20",
          9717 => x"20",
          9718 => x"25",
          9719 => x"4d",
          9720 => x"00",
          9721 => x"20",
          9722 => x"52",
          9723 => x"43",
          9724 => x"6b",
          9725 => x"65",
          9726 => x"20",
          9727 => x"20",
          9728 => x"20",
          9729 => x"25",
          9730 => x"4d",
          9731 => x"00",
          9732 => x"20",
          9733 => x"73",
          9734 => x"6e",
          9735 => x"44",
          9736 => x"20",
          9737 => x"63",
          9738 => x"72",
          9739 => x"20",
          9740 => x"25",
          9741 => x"4d",
          9742 => x"00",
          9743 => x"61",
          9744 => x"00",
          9745 => x"64",
          9746 => x"00",
          9747 => x"65",
          9748 => x"00",
          9749 => x"4f",
          9750 => x"4f",
          9751 => x"00",
          9752 => x"6b",
          9753 => x"6e",
          9754 => x"99",
          9755 => x"00",
          9756 => x"00",
          9757 => x"99",
          9758 => x"00",
          9759 => x"00",
          9760 => x"99",
          9761 => x"00",
          9762 => x"00",
          9763 => x"99",
          9764 => x"00",
          9765 => x"00",
          9766 => x"99",
          9767 => x"00",
          9768 => x"00",
          9769 => x"99",
          9770 => x"00",
          9771 => x"00",
          9772 => x"99",
          9773 => x"00",
          9774 => x"00",
          9775 => x"99",
          9776 => x"00",
          9777 => x"00",
          9778 => x"99",
          9779 => x"00",
          9780 => x"00",
          9781 => x"99",
          9782 => x"00",
          9783 => x"00",
          9784 => x"99",
          9785 => x"00",
          9786 => x"00",
          9787 => x"99",
          9788 => x"00",
          9789 => x"00",
          9790 => x"99",
          9791 => x"00",
          9792 => x"00",
          9793 => x"99",
          9794 => x"00",
          9795 => x"00",
          9796 => x"99",
          9797 => x"00",
          9798 => x"00",
          9799 => x"99",
          9800 => x"00",
          9801 => x"00",
          9802 => x"99",
          9803 => x"00",
          9804 => x"00",
          9805 => x"99",
          9806 => x"00",
          9807 => x"00",
          9808 => x"99",
          9809 => x"00",
          9810 => x"00",
          9811 => x"99",
          9812 => x"00",
          9813 => x"00",
          9814 => x"99",
          9815 => x"00",
          9816 => x"00",
          9817 => x"99",
          9818 => x"00",
          9819 => x"00",
          9820 => x"44",
          9821 => x"43",
          9822 => x"42",
          9823 => x"41",
          9824 => x"36",
          9825 => x"35",
          9826 => x"34",
          9827 => x"46",
          9828 => x"33",
          9829 => x"32",
          9830 => x"31",
          9831 => x"00",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"00",
          9836 => x"00",
          9837 => x"00",
          9838 => x"00",
          9839 => x"00",
          9840 => x"00",
          9841 => x"00",
          9842 => x"73",
          9843 => x"79",
          9844 => x"73",
          9845 => x"00",
          9846 => x"00",
          9847 => x"34",
          9848 => x"20",
          9849 => x"00",
          9850 => x"69",
          9851 => x"20",
          9852 => x"72",
          9853 => x"74",
          9854 => x"65",
          9855 => x"73",
          9856 => x"79",
          9857 => x"6c",
          9858 => x"6f",
          9859 => x"46",
          9860 => x"00",
          9861 => x"6e",
          9862 => x"20",
          9863 => x"6e",
          9864 => x"65",
          9865 => x"20",
          9866 => x"74",
          9867 => x"20",
          9868 => x"65",
          9869 => x"69",
          9870 => x"6c",
          9871 => x"2e",
          9872 => x"00",
          9873 => x"2b",
          9874 => x"3c",
          9875 => x"5b",
          9876 => x"00",
          9877 => x"54",
          9878 => x"54",
          9879 => x"00",
          9880 => x"90",
          9881 => x"4f",
          9882 => x"30",
          9883 => x"20",
          9884 => x"45",
          9885 => x"20",
          9886 => x"33",
          9887 => x"20",
          9888 => x"20",
          9889 => x"45",
          9890 => x"20",
          9891 => x"20",
          9892 => x"20",
          9893 => x"9a",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"45",
          9898 => x"8f",
          9899 => x"45",
          9900 => x"8e",
          9901 => x"92",
          9902 => x"55",
          9903 => x"9a",
          9904 => x"9e",
          9905 => x"4f",
          9906 => x"a6",
          9907 => x"aa",
          9908 => x"ae",
          9909 => x"b2",
          9910 => x"b6",
          9911 => x"ba",
          9912 => x"be",
          9913 => x"c2",
          9914 => x"c6",
          9915 => x"ca",
          9916 => x"ce",
          9917 => x"d2",
          9918 => x"d6",
          9919 => x"da",
          9920 => x"de",
          9921 => x"e2",
          9922 => x"e6",
          9923 => x"ea",
          9924 => x"ee",
          9925 => x"f2",
          9926 => x"f6",
          9927 => x"fa",
          9928 => x"fe",
          9929 => x"2c",
          9930 => x"5d",
          9931 => x"2a",
          9932 => x"3f",
          9933 => x"00",
          9934 => x"00",
          9935 => x"00",
          9936 => x"02",
          9937 => x"00",
          9938 => x"00",
          9939 => x"00",
          9940 => x"00",
          9941 => x"00",
          9942 => x"00",
          9943 => x"8f",
          9944 => x"01",
          9945 => x"00",
          9946 => x"00",
          9947 => x"8f",
          9948 => x"01",
          9949 => x"00",
          9950 => x"00",
          9951 => x"8f",
          9952 => x"03",
          9953 => x"00",
          9954 => x"00",
          9955 => x"8f",
          9956 => x"03",
          9957 => x"00",
          9958 => x"00",
          9959 => x"8f",
          9960 => x"03",
          9961 => x"00",
          9962 => x"00",
          9963 => x"8f",
          9964 => x"04",
          9965 => x"00",
          9966 => x"00",
          9967 => x"8f",
          9968 => x"04",
          9969 => x"00",
          9970 => x"00",
          9971 => x"8f",
          9972 => x"04",
          9973 => x"00",
          9974 => x"00",
          9975 => x"8f",
          9976 => x"04",
          9977 => x"00",
          9978 => x"00",
          9979 => x"8f",
          9980 => x"04",
          9981 => x"00",
          9982 => x"00",
          9983 => x"8f",
          9984 => x"04",
          9985 => x"00",
          9986 => x"00",
          9987 => x"8f",
          9988 => x"04",
          9989 => x"00",
          9990 => x"00",
          9991 => x"8f",
          9992 => x"05",
          9993 => x"00",
          9994 => x"00",
          9995 => x"8f",
          9996 => x"05",
          9997 => x"00",
          9998 => x"00",
          9999 => x"8f",
         10000 => x"05",
         10001 => x"00",
         10002 => x"00",
         10003 => x"8f",
         10004 => x"05",
         10005 => x"00",
         10006 => x"00",
         10007 => x"8f",
         10008 => x"07",
         10009 => x"00",
         10010 => x"00",
         10011 => x"8f",
         10012 => x"07",
         10013 => x"00",
         10014 => x"00",
         10015 => x"8f",
         10016 => x"08",
         10017 => x"00",
         10018 => x"00",
         10019 => x"8f",
         10020 => x"08",
         10021 => x"00",
         10022 => x"00",
         10023 => x"8f",
         10024 => x"08",
         10025 => x"00",
         10026 => x"00",
         10027 => x"8f",
         10028 => x"08",
         10029 => x"00",
         10030 => x"00",
         10031 => x"8f",
         10032 => x"09",
         10033 => x"00",
         10034 => x"00",
         10035 => x"8f",
         10036 => x"09",
         10037 => x"00",
         10038 => x"00",
         10039 => x"8f",
         10040 => x"09",
         10041 => x"00",
         10042 => x"00",
         10043 => x"8f",
         10044 => x"09",
         10045 => x"00",
         10046 => x"00",
         10047 => x"00",
         10048 => x"00",
         10049 => x"7f",
         10050 => x"00",
         10051 => x"7f",
         10052 => x"00",
         10053 => x"7f",
         10054 => x"00",
         10055 => x"00",
         10056 => x"00",
         10057 => x"ff",
         10058 => x"00",
         10059 => x"00",
         10060 => x"78",
         10061 => x"00",
         10062 => x"e1",
         10063 => x"e1",
         10064 => x"e1",
         10065 => x"00",
         10066 => x"01",
         10067 => x"01",
         10068 => x"10",
         10069 => x"00",
         10070 => x"00",
         10071 => x"00",
         10072 => x"00",
         10073 => x"00",
         10074 => x"00",
         10075 => x"00",
         10076 => x"00",
         10077 => x"00",
         10078 => x"00",
         10079 => x"00",
         10080 => x"00",
         10081 => x"00",
         10082 => x"00",
         10083 => x"00",
         10084 => x"00",
         10085 => x"00",
         10086 => x"00",
         10087 => x"00",
         10088 => x"00",
         10089 => x"00",
         10090 => x"00",
         10091 => x"00",
         10092 => x"00",
         10093 => x"00",
         10094 => x"99",
         10095 => x"00",
         10096 => x"99",
         10097 => x"00",
         10098 => x"99",
         10099 => x"00",
         10100 => x"00",
         10101 => x"00",
         10102 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"85",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"80",
           387 => x"82",
           388 => x"82",
           389 => x"82",
           390 => x"b3",
           391 => x"bb",
           392 => x"d8",
           393 => x"bb",
           394 => x"e3",
           395 => x"e8",
           396 => x"90",
           397 => x"e8",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"82",
           403 => x"82",
           404 => x"82",
           405 => x"b1",
           406 => x"bb",
           407 => x"d8",
           408 => x"bb",
           409 => x"cf",
           410 => x"bb",
           411 => x"d8",
           412 => x"bb",
           413 => x"c9",
           414 => x"bb",
           415 => x"d8",
           416 => x"bb",
           417 => x"d8",
           418 => x"e8",
           419 => x"90",
           420 => x"e8",
           421 => x"2d",
           422 => x"08",
           423 => x"04",
           424 => x"0c",
           425 => x"82",
           426 => x"82",
           427 => x"82",
           428 => x"80",
           429 => x"82",
           430 => x"82",
           431 => x"82",
           432 => x"80",
           433 => x"82",
           434 => x"82",
           435 => x"82",
           436 => x"80",
           437 => x"82",
           438 => x"82",
           439 => x"82",
           440 => x"80",
           441 => x"82",
           442 => x"82",
           443 => x"82",
           444 => x"80",
           445 => x"82",
           446 => x"82",
           447 => x"82",
           448 => x"81",
           449 => x"82",
           450 => x"82",
           451 => x"82",
           452 => x"81",
           453 => x"82",
           454 => x"82",
           455 => x"82",
           456 => x"81",
           457 => x"82",
           458 => x"82",
           459 => x"82",
           460 => x"81",
           461 => x"82",
           462 => x"82",
           463 => x"82",
           464 => x"81",
           465 => x"82",
           466 => x"82",
           467 => x"82",
           468 => x"81",
           469 => x"82",
           470 => x"82",
           471 => x"82",
           472 => x"81",
           473 => x"82",
           474 => x"82",
           475 => x"82",
           476 => x"81",
           477 => x"82",
           478 => x"82",
           479 => x"82",
           480 => x"81",
           481 => x"82",
           482 => x"82",
           483 => x"82",
           484 => x"81",
           485 => x"82",
           486 => x"82",
           487 => x"82",
           488 => x"81",
           489 => x"82",
           490 => x"82",
           491 => x"82",
           492 => x"81",
           493 => x"82",
           494 => x"82",
           495 => x"82",
           496 => x"81",
           497 => x"82",
           498 => x"82",
           499 => x"82",
           500 => x"81",
           501 => x"82",
           502 => x"82",
           503 => x"82",
           504 => x"82",
           505 => x"82",
           506 => x"82",
           507 => x"82",
           508 => x"82",
           509 => x"82",
           510 => x"82",
           511 => x"82",
           512 => x"81",
           513 => x"82",
           514 => x"82",
           515 => x"82",
           516 => x"81",
           517 => x"82",
           518 => x"82",
           519 => x"82",
           520 => x"81",
           521 => x"82",
           522 => x"82",
           523 => x"82",
           524 => x"81",
           525 => x"82",
           526 => x"82",
           527 => x"82",
           528 => x"82",
           529 => x"82",
           530 => x"82",
           531 => x"82",
           532 => x"82",
           533 => x"82",
           534 => x"82",
           535 => x"82",
           536 => x"82",
           537 => x"82",
           538 => x"82",
           539 => x"82",
           540 => x"81",
           541 => x"82",
           542 => x"82",
           543 => x"82",
           544 => x"82",
           545 => x"82",
           546 => x"82",
           547 => x"82",
           548 => x"82",
           549 => x"82",
           550 => x"82",
           551 => x"82",
           552 => x"82",
           553 => x"82",
           554 => x"82",
           555 => x"82",
           556 => x"81",
           557 => x"82",
           558 => x"82",
           559 => x"82",
           560 => x"81",
           561 => x"82",
           562 => x"82",
           563 => x"82",
           564 => x"81",
           565 => x"82",
           566 => x"82",
           567 => x"82",
           568 => x"80",
           569 => x"82",
           570 => x"82",
           571 => x"82",
           572 => x"80",
           573 => x"82",
           574 => x"82",
           575 => x"82",
           576 => x"80",
           577 => x"82",
           578 => x"82",
           579 => x"82",
           580 => x"80",
           581 => x"82",
           582 => x"82",
           583 => x"82",
           584 => x"81",
           585 => x"82",
           586 => x"82",
           587 => x"82",
           588 => x"81",
           589 => x"82",
           590 => x"82",
           591 => x"82",
           592 => x"81",
           593 => x"82",
           594 => x"82",
           595 => x"82",
           596 => x"81",
           597 => x"82",
           598 => x"82",
           599 => x"3c",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"51",
           609 => x"73",
           610 => x"73",
           611 => x"81",
           612 => x"10",
           613 => x"07",
           614 => x"0c",
           615 => x"72",
           616 => x"81",
           617 => x"09",
           618 => x"71",
           619 => x"0a",
           620 => x"72",
           621 => x"51",
           622 => x"82",
           623 => x"82",
           624 => x"8e",
           625 => x"70",
           626 => x"0c",
           627 => x"93",
           628 => x"81",
           629 => x"95",
           630 => x"bb",
           631 => x"82",
           632 => x"fb",
           633 => x"bb",
           634 => x"05",
           635 => x"e8",
           636 => x"0c",
           637 => x"08",
           638 => x"54",
           639 => x"08",
           640 => x"53",
           641 => x"08",
           642 => x"9a",
           643 => x"dc",
           644 => x"bb",
           645 => x"05",
           646 => x"e8",
           647 => x"08",
           648 => x"dc",
           649 => x"87",
           650 => x"bb",
           651 => x"82",
           652 => x"02",
           653 => x"0c",
           654 => x"82",
           655 => x"90",
           656 => x"11",
           657 => x"32",
           658 => x"51",
           659 => x"71",
           660 => x"0b",
           661 => x"08",
           662 => x"25",
           663 => x"39",
           664 => x"bb",
           665 => x"05",
           666 => x"39",
           667 => x"08",
           668 => x"ff",
           669 => x"e8",
           670 => x"0c",
           671 => x"bb",
           672 => x"05",
           673 => x"e8",
           674 => x"08",
           675 => x"08",
           676 => x"82",
           677 => x"f8",
           678 => x"2e",
           679 => x"80",
           680 => x"e8",
           681 => x"08",
           682 => x"38",
           683 => x"08",
           684 => x"51",
           685 => x"82",
           686 => x"70",
           687 => x"08",
           688 => x"52",
           689 => x"08",
           690 => x"ff",
           691 => x"06",
           692 => x"0b",
           693 => x"08",
           694 => x"80",
           695 => x"bb",
           696 => x"05",
           697 => x"e8",
           698 => x"08",
           699 => x"73",
           700 => x"e8",
           701 => x"08",
           702 => x"bb",
           703 => x"05",
           704 => x"e8",
           705 => x"08",
           706 => x"bb",
           707 => x"05",
           708 => x"39",
           709 => x"08",
           710 => x"52",
           711 => x"82",
           712 => x"88",
           713 => x"82",
           714 => x"f4",
           715 => x"82",
           716 => x"f4",
           717 => x"bb",
           718 => x"3d",
           719 => x"e8",
           720 => x"bb",
           721 => x"82",
           722 => x"f4",
           723 => x"0b",
           724 => x"08",
           725 => x"82",
           726 => x"88",
           727 => x"bb",
           728 => x"05",
           729 => x"0b",
           730 => x"08",
           731 => x"82",
           732 => x"90",
           733 => x"bb",
           734 => x"05",
           735 => x"e8",
           736 => x"08",
           737 => x"e8",
           738 => x"08",
           739 => x"e8",
           740 => x"70",
           741 => x"81",
           742 => x"bb",
           743 => x"82",
           744 => x"dc",
           745 => x"bb",
           746 => x"05",
           747 => x"e8",
           748 => x"08",
           749 => x"80",
           750 => x"bb",
           751 => x"05",
           752 => x"bb",
           753 => x"8e",
           754 => x"bb",
           755 => x"82",
           756 => x"02",
           757 => x"0c",
           758 => x"82",
           759 => x"90",
           760 => x"bb",
           761 => x"05",
           762 => x"e8",
           763 => x"08",
           764 => x"e8",
           765 => x"08",
           766 => x"e8",
           767 => x"08",
           768 => x"3f",
           769 => x"08",
           770 => x"e8",
           771 => x"0c",
           772 => x"08",
           773 => x"70",
           774 => x"0c",
           775 => x"3d",
           776 => x"e8",
           777 => x"bb",
           778 => x"82",
           779 => x"ed",
           780 => x"0b",
           781 => x"08",
           782 => x"82",
           783 => x"88",
           784 => x"80",
           785 => x"0c",
           786 => x"08",
           787 => x"85",
           788 => x"81",
           789 => x"32",
           790 => x"51",
           791 => x"53",
           792 => x"8d",
           793 => x"82",
           794 => x"e0",
           795 => x"ac",
           796 => x"e8",
           797 => x"08",
           798 => x"53",
           799 => x"e8",
           800 => x"34",
           801 => x"06",
           802 => x"2e",
           803 => x"82",
           804 => x"8c",
           805 => x"05",
           806 => x"08",
           807 => x"82",
           808 => x"e4",
           809 => x"81",
           810 => x"72",
           811 => x"8b",
           812 => x"e8",
           813 => x"33",
           814 => x"27",
           815 => x"82",
           816 => x"f8",
           817 => x"72",
           818 => x"ee",
           819 => x"e8",
           820 => x"33",
           821 => x"2e",
           822 => x"80",
           823 => x"bb",
           824 => x"05",
           825 => x"2b",
           826 => x"51",
           827 => x"b2",
           828 => x"e8",
           829 => x"22",
           830 => x"70",
           831 => x"81",
           832 => x"51",
           833 => x"2e",
           834 => x"bb",
           835 => x"05",
           836 => x"80",
           837 => x"72",
           838 => x"08",
           839 => x"fe",
           840 => x"bb",
           841 => x"05",
           842 => x"2b",
           843 => x"70",
           844 => x"72",
           845 => x"51",
           846 => x"51",
           847 => x"82",
           848 => x"e8",
           849 => x"bb",
           850 => x"05",
           851 => x"bb",
           852 => x"05",
           853 => x"d0",
           854 => x"53",
           855 => x"e8",
           856 => x"34",
           857 => x"08",
           858 => x"70",
           859 => x"98",
           860 => x"53",
           861 => x"8b",
           862 => x"0b",
           863 => x"08",
           864 => x"82",
           865 => x"e4",
           866 => x"83",
           867 => x"06",
           868 => x"72",
           869 => x"82",
           870 => x"e8",
           871 => x"88",
           872 => x"2b",
           873 => x"70",
           874 => x"51",
           875 => x"72",
           876 => x"08",
           877 => x"fd",
           878 => x"bb",
           879 => x"05",
           880 => x"2a",
           881 => x"51",
           882 => x"80",
           883 => x"82",
           884 => x"e8",
           885 => x"98",
           886 => x"2c",
           887 => x"72",
           888 => x"0b",
           889 => x"08",
           890 => x"82",
           891 => x"f8",
           892 => x"11",
           893 => x"08",
           894 => x"53",
           895 => x"08",
           896 => x"80",
           897 => x"94",
           898 => x"e8",
           899 => x"08",
           900 => x"82",
           901 => x"70",
           902 => x"51",
           903 => x"82",
           904 => x"e4",
           905 => x"90",
           906 => x"72",
           907 => x"08",
           908 => x"82",
           909 => x"e4",
           910 => x"a0",
           911 => x"72",
           912 => x"08",
           913 => x"fc",
           914 => x"bb",
           915 => x"05",
           916 => x"80",
           917 => x"72",
           918 => x"08",
           919 => x"fc",
           920 => x"bb",
           921 => x"05",
           922 => x"c0",
           923 => x"72",
           924 => x"08",
           925 => x"fb",
           926 => x"bb",
           927 => x"05",
           928 => x"07",
           929 => x"82",
           930 => x"e4",
           931 => x"0b",
           932 => x"08",
           933 => x"fb",
           934 => x"bb",
           935 => x"05",
           936 => x"07",
           937 => x"82",
           938 => x"e4",
           939 => x"c1",
           940 => x"82",
           941 => x"fc",
           942 => x"bb",
           943 => x"05",
           944 => x"51",
           945 => x"bb",
           946 => x"05",
           947 => x"0b",
           948 => x"08",
           949 => x"8d",
           950 => x"bb",
           951 => x"05",
           952 => x"e8",
           953 => x"08",
           954 => x"bb",
           955 => x"05",
           956 => x"51",
           957 => x"bb",
           958 => x"05",
           959 => x"e8",
           960 => x"22",
           961 => x"53",
           962 => x"e8",
           963 => x"23",
           964 => x"82",
           965 => x"90",
           966 => x"bb",
           967 => x"05",
           968 => x"82",
           969 => x"90",
           970 => x"08",
           971 => x"08",
           972 => x"82",
           973 => x"e4",
           974 => x"83",
           975 => x"06",
           976 => x"53",
           977 => x"ab",
           978 => x"e8",
           979 => x"33",
           980 => x"53",
           981 => x"53",
           982 => x"08",
           983 => x"52",
           984 => x"3f",
           985 => x"08",
           986 => x"bb",
           987 => x"05",
           988 => x"82",
           989 => x"fc",
           990 => x"9d",
           991 => x"bb",
           992 => x"72",
           993 => x"08",
           994 => x"82",
           995 => x"ec",
           996 => x"82",
           997 => x"f4",
           998 => x"71",
           999 => x"72",
          1000 => x"08",
          1001 => x"8b",
          1002 => x"bb",
          1003 => x"05",
          1004 => x"e8",
          1005 => x"08",
          1006 => x"bb",
          1007 => x"05",
          1008 => x"82",
          1009 => x"fc",
          1010 => x"bb",
          1011 => x"05",
          1012 => x"2a",
          1013 => x"51",
          1014 => x"72",
          1015 => x"38",
          1016 => x"08",
          1017 => x"70",
          1018 => x"72",
          1019 => x"82",
          1020 => x"fc",
          1021 => x"53",
          1022 => x"82",
          1023 => x"53",
          1024 => x"e8",
          1025 => x"23",
          1026 => x"bb",
          1027 => x"05",
          1028 => x"f3",
          1029 => x"dc",
          1030 => x"82",
          1031 => x"f4",
          1032 => x"bb",
          1033 => x"05",
          1034 => x"bb",
          1035 => x"05",
          1036 => x"31",
          1037 => x"82",
          1038 => x"ec",
          1039 => x"c1",
          1040 => x"e8",
          1041 => x"22",
          1042 => x"70",
          1043 => x"51",
          1044 => x"2e",
          1045 => x"bb",
          1046 => x"05",
          1047 => x"e8",
          1048 => x"08",
          1049 => x"bb",
          1050 => x"05",
          1051 => x"82",
          1052 => x"dc",
          1053 => x"a2",
          1054 => x"e8",
          1055 => x"08",
          1056 => x"08",
          1057 => x"84",
          1058 => x"e8",
          1059 => x"0c",
          1060 => x"bb",
          1061 => x"05",
          1062 => x"bb",
          1063 => x"05",
          1064 => x"e8",
          1065 => x"0c",
          1066 => x"08",
          1067 => x"80",
          1068 => x"82",
          1069 => x"e4",
          1070 => x"82",
          1071 => x"72",
          1072 => x"08",
          1073 => x"82",
          1074 => x"fc",
          1075 => x"82",
          1076 => x"fc",
          1077 => x"bb",
          1078 => x"05",
          1079 => x"bf",
          1080 => x"72",
          1081 => x"08",
          1082 => x"81",
          1083 => x"0b",
          1084 => x"08",
          1085 => x"a9",
          1086 => x"e8",
          1087 => x"22",
          1088 => x"07",
          1089 => x"82",
          1090 => x"e4",
          1091 => x"f8",
          1092 => x"e8",
          1093 => x"34",
          1094 => x"bb",
          1095 => x"05",
          1096 => x"e8",
          1097 => x"22",
          1098 => x"70",
          1099 => x"51",
          1100 => x"2e",
          1101 => x"bb",
          1102 => x"05",
          1103 => x"e8",
          1104 => x"08",
          1105 => x"bb",
          1106 => x"05",
          1107 => x"82",
          1108 => x"d8",
          1109 => x"a2",
          1110 => x"e8",
          1111 => x"08",
          1112 => x"08",
          1113 => x"84",
          1114 => x"e8",
          1115 => x"0c",
          1116 => x"bb",
          1117 => x"05",
          1118 => x"bb",
          1119 => x"05",
          1120 => x"e8",
          1121 => x"0c",
          1122 => x"08",
          1123 => x"70",
          1124 => x"53",
          1125 => x"e8",
          1126 => x"23",
          1127 => x"0b",
          1128 => x"08",
          1129 => x"82",
          1130 => x"f0",
          1131 => x"bb",
          1132 => x"05",
          1133 => x"e8",
          1134 => x"08",
          1135 => x"54",
          1136 => x"a3",
          1137 => x"bb",
          1138 => x"72",
          1139 => x"bb",
          1140 => x"05",
          1141 => x"e8",
          1142 => x"0c",
          1143 => x"08",
          1144 => x"70",
          1145 => x"89",
          1146 => x"38",
          1147 => x"08",
          1148 => x"53",
          1149 => x"82",
          1150 => x"f8",
          1151 => x"15",
          1152 => x"51",
          1153 => x"bb",
          1154 => x"05",
          1155 => x"82",
          1156 => x"f0",
          1157 => x"72",
          1158 => x"51",
          1159 => x"bb",
          1160 => x"05",
          1161 => x"e8",
          1162 => x"08",
          1163 => x"e8",
          1164 => x"33",
          1165 => x"bb",
          1166 => x"05",
          1167 => x"82",
          1168 => x"f0",
          1169 => x"bb",
          1170 => x"05",
          1171 => x"82",
          1172 => x"fc",
          1173 => x"53",
          1174 => x"82",
          1175 => x"70",
          1176 => x"08",
          1177 => x"53",
          1178 => x"08",
          1179 => x"80",
          1180 => x"fe",
          1181 => x"bb",
          1182 => x"05",
          1183 => x"ec",
          1184 => x"54",
          1185 => x"31",
          1186 => x"82",
          1187 => x"fc",
          1188 => x"bb",
          1189 => x"05",
          1190 => x"06",
          1191 => x"80",
          1192 => x"82",
          1193 => x"ec",
          1194 => x"11",
          1195 => x"82",
          1196 => x"ec",
          1197 => x"bb",
          1198 => x"05",
          1199 => x"2a",
          1200 => x"51",
          1201 => x"80",
          1202 => x"38",
          1203 => x"08",
          1204 => x"70",
          1205 => x"bb",
          1206 => x"05",
          1207 => x"e8",
          1208 => x"08",
          1209 => x"bb",
          1210 => x"05",
          1211 => x"e8",
          1212 => x"22",
          1213 => x"90",
          1214 => x"06",
          1215 => x"bb",
          1216 => x"05",
          1217 => x"53",
          1218 => x"e8",
          1219 => x"23",
          1220 => x"bb",
          1221 => x"05",
          1222 => x"53",
          1223 => x"e8",
          1224 => x"23",
          1225 => x"08",
          1226 => x"82",
          1227 => x"ec",
          1228 => x"bb",
          1229 => x"05",
          1230 => x"2a",
          1231 => x"51",
          1232 => x"80",
          1233 => x"38",
          1234 => x"08",
          1235 => x"70",
          1236 => x"98",
          1237 => x"e8",
          1238 => x"33",
          1239 => x"53",
          1240 => x"97",
          1241 => x"e8",
          1242 => x"22",
          1243 => x"51",
          1244 => x"bb",
          1245 => x"05",
          1246 => x"82",
          1247 => x"e8",
          1248 => x"82",
          1249 => x"fc",
          1250 => x"71",
          1251 => x"72",
          1252 => x"08",
          1253 => x"82",
          1254 => x"e4",
          1255 => x"83",
          1256 => x"06",
          1257 => x"72",
          1258 => x"38",
          1259 => x"08",
          1260 => x"70",
          1261 => x"90",
          1262 => x"2c",
          1263 => x"51",
          1264 => x"53",
          1265 => x"bb",
          1266 => x"05",
          1267 => x"31",
          1268 => x"82",
          1269 => x"ec",
          1270 => x"39",
          1271 => x"08",
          1272 => x"70",
          1273 => x"90",
          1274 => x"2c",
          1275 => x"51",
          1276 => x"53",
          1277 => x"bb",
          1278 => x"05",
          1279 => x"31",
          1280 => x"82",
          1281 => x"ec",
          1282 => x"bb",
          1283 => x"05",
          1284 => x"80",
          1285 => x"72",
          1286 => x"bb",
          1287 => x"05",
          1288 => x"54",
          1289 => x"bb",
          1290 => x"05",
          1291 => x"2b",
          1292 => x"51",
          1293 => x"25",
          1294 => x"bb",
          1295 => x"05",
          1296 => x"51",
          1297 => x"d2",
          1298 => x"e8",
          1299 => x"22",
          1300 => x"70",
          1301 => x"51",
          1302 => x"2e",
          1303 => x"bb",
          1304 => x"05",
          1305 => x"51",
          1306 => x"80",
          1307 => x"bb",
          1308 => x"05",
          1309 => x"2a",
          1310 => x"51",
          1311 => x"80",
          1312 => x"82",
          1313 => x"88",
          1314 => x"ab",
          1315 => x"3f",
          1316 => x"bb",
          1317 => x"05",
          1318 => x"2a",
          1319 => x"51",
          1320 => x"80",
          1321 => x"82",
          1322 => x"88",
          1323 => x"a0",
          1324 => x"3f",
          1325 => x"08",
          1326 => x"70",
          1327 => x"81",
          1328 => x"53",
          1329 => x"b1",
          1330 => x"e8",
          1331 => x"08",
          1332 => x"89",
          1333 => x"bb",
          1334 => x"05",
          1335 => x"90",
          1336 => x"06",
          1337 => x"bb",
          1338 => x"05",
          1339 => x"bb",
          1340 => x"05",
          1341 => x"bc",
          1342 => x"e8",
          1343 => x"22",
          1344 => x"70",
          1345 => x"51",
          1346 => x"2e",
          1347 => x"bb",
          1348 => x"05",
          1349 => x"54",
          1350 => x"bb",
          1351 => x"05",
          1352 => x"2b",
          1353 => x"51",
          1354 => x"25",
          1355 => x"bb",
          1356 => x"05",
          1357 => x"51",
          1358 => x"d2",
          1359 => x"e8",
          1360 => x"22",
          1361 => x"70",
          1362 => x"51",
          1363 => x"2e",
          1364 => x"bb",
          1365 => x"05",
          1366 => x"54",
          1367 => x"bb",
          1368 => x"05",
          1369 => x"2b",
          1370 => x"51",
          1371 => x"25",
          1372 => x"bb",
          1373 => x"05",
          1374 => x"51",
          1375 => x"d2",
          1376 => x"e8",
          1377 => x"22",
          1378 => x"70",
          1379 => x"51",
          1380 => x"38",
          1381 => x"08",
          1382 => x"ff",
          1383 => x"72",
          1384 => x"08",
          1385 => x"73",
          1386 => x"90",
          1387 => x"80",
          1388 => x"38",
          1389 => x"08",
          1390 => x"52",
          1391 => x"f4",
          1392 => x"82",
          1393 => x"f8",
          1394 => x"72",
          1395 => x"09",
          1396 => x"38",
          1397 => x"08",
          1398 => x"52",
          1399 => x"08",
          1400 => x"51",
          1401 => x"81",
          1402 => x"bb",
          1403 => x"05",
          1404 => x"80",
          1405 => x"81",
          1406 => x"38",
          1407 => x"08",
          1408 => x"ff",
          1409 => x"72",
          1410 => x"08",
          1411 => x"72",
          1412 => x"06",
          1413 => x"ff",
          1414 => x"bb",
          1415 => x"e8",
          1416 => x"08",
          1417 => x"e8",
          1418 => x"08",
          1419 => x"82",
          1420 => x"fc",
          1421 => x"05",
          1422 => x"08",
          1423 => x"53",
          1424 => x"ff",
          1425 => x"bb",
          1426 => x"05",
          1427 => x"80",
          1428 => x"81",
          1429 => x"38",
          1430 => x"08",
          1431 => x"ff",
          1432 => x"72",
          1433 => x"08",
          1434 => x"72",
          1435 => x"06",
          1436 => x"ff",
          1437 => x"df",
          1438 => x"e8",
          1439 => x"08",
          1440 => x"e8",
          1441 => x"08",
          1442 => x"53",
          1443 => x"82",
          1444 => x"fc",
          1445 => x"05",
          1446 => x"08",
          1447 => x"ff",
          1448 => x"bb",
          1449 => x"05",
          1450 => x"ec",
          1451 => x"82",
          1452 => x"88",
          1453 => x"82",
          1454 => x"f0",
          1455 => x"05",
          1456 => x"08",
          1457 => x"82",
          1458 => x"f0",
          1459 => x"33",
          1460 => x"e0",
          1461 => x"82",
          1462 => x"e4",
          1463 => x"87",
          1464 => x"06",
          1465 => x"72",
          1466 => x"c3",
          1467 => x"e8",
          1468 => x"22",
          1469 => x"54",
          1470 => x"e8",
          1471 => x"23",
          1472 => x"70",
          1473 => x"53",
          1474 => x"a3",
          1475 => x"e8",
          1476 => x"08",
          1477 => x"85",
          1478 => x"39",
          1479 => x"08",
          1480 => x"52",
          1481 => x"08",
          1482 => x"51",
          1483 => x"80",
          1484 => x"e8",
          1485 => x"23",
          1486 => x"82",
          1487 => x"f8",
          1488 => x"72",
          1489 => x"81",
          1490 => x"81",
          1491 => x"e8",
          1492 => x"23",
          1493 => x"bb",
          1494 => x"05",
          1495 => x"82",
          1496 => x"e8",
          1497 => x"0b",
          1498 => x"08",
          1499 => x"ea",
          1500 => x"bb",
          1501 => x"05",
          1502 => x"bb",
          1503 => x"05",
          1504 => x"b0",
          1505 => x"39",
          1506 => x"08",
          1507 => x"8c",
          1508 => x"82",
          1509 => x"e0",
          1510 => x"53",
          1511 => x"08",
          1512 => x"82",
          1513 => x"95",
          1514 => x"bb",
          1515 => x"82",
          1516 => x"02",
          1517 => x"0c",
          1518 => x"82",
          1519 => x"53",
          1520 => x"08",
          1521 => x"52",
          1522 => x"08",
          1523 => x"51",
          1524 => x"82",
          1525 => x"70",
          1526 => x"0c",
          1527 => x"0d",
          1528 => x"0c",
          1529 => x"e8",
          1530 => x"bb",
          1531 => x"3d",
          1532 => x"82",
          1533 => x"f8",
          1534 => x"d3",
          1535 => x"11",
          1536 => x"2a",
          1537 => x"70",
          1538 => x"51",
          1539 => x"72",
          1540 => x"38",
          1541 => x"bb",
          1542 => x"05",
          1543 => x"39",
          1544 => x"08",
          1545 => x"53",
          1546 => x"bb",
          1547 => x"05",
          1548 => x"82",
          1549 => x"88",
          1550 => x"72",
          1551 => x"08",
          1552 => x"72",
          1553 => x"53",
          1554 => x"b0",
          1555 => x"b0",
          1556 => x"b0",
          1557 => x"bb",
          1558 => x"05",
          1559 => x"11",
          1560 => x"72",
          1561 => x"dc",
          1562 => x"80",
          1563 => x"38",
          1564 => x"bb",
          1565 => x"05",
          1566 => x"39",
          1567 => x"08",
          1568 => x"08",
          1569 => x"51",
          1570 => x"53",
          1571 => x"bb",
          1572 => x"72",
          1573 => x"38",
          1574 => x"bb",
          1575 => x"05",
          1576 => x"e8",
          1577 => x"08",
          1578 => x"e8",
          1579 => x"0c",
          1580 => x"e8",
          1581 => x"08",
          1582 => x"0c",
          1583 => x"82",
          1584 => x"04",
          1585 => x"08",
          1586 => x"e8",
          1587 => x"0d",
          1588 => x"bb",
          1589 => x"05",
          1590 => x"e8",
          1591 => x"08",
          1592 => x"70",
          1593 => x"81",
          1594 => x"06",
          1595 => x"51",
          1596 => x"2e",
          1597 => x"0b",
          1598 => x"08",
          1599 => x"80",
          1600 => x"bb",
          1601 => x"05",
          1602 => x"33",
          1603 => x"08",
          1604 => x"81",
          1605 => x"e8",
          1606 => x"0c",
          1607 => x"bb",
          1608 => x"05",
          1609 => x"ff",
          1610 => x"80",
          1611 => x"82",
          1612 => x"8c",
          1613 => x"bb",
          1614 => x"05",
          1615 => x"bb",
          1616 => x"05",
          1617 => x"11",
          1618 => x"72",
          1619 => x"dc",
          1620 => x"80",
          1621 => x"38",
          1622 => x"bb",
          1623 => x"05",
          1624 => x"39",
          1625 => x"08",
          1626 => x"70",
          1627 => x"08",
          1628 => x"53",
          1629 => x"08",
          1630 => x"82",
          1631 => x"87",
          1632 => x"bb",
          1633 => x"82",
          1634 => x"02",
          1635 => x"0c",
          1636 => x"82",
          1637 => x"52",
          1638 => x"08",
          1639 => x"51",
          1640 => x"bb",
          1641 => x"82",
          1642 => x"53",
          1643 => x"82",
          1644 => x"04",
          1645 => x"08",
          1646 => x"e8",
          1647 => x"0d",
          1648 => x"08",
          1649 => x"85",
          1650 => x"81",
          1651 => x"32",
          1652 => x"51",
          1653 => x"53",
          1654 => x"8d",
          1655 => x"82",
          1656 => x"fc",
          1657 => x"cb",
          1658 => x"e8",
          1659 => x"08",
          1660 => x"70",
          1661 => x"81",
          1662 => x"51",
          1663 => x"2e",
          1664 => x"82",
          1665 => x"8c",
          1666 => x"bb",
          1667 => x"05",
          1668 => x"8c",
          1669 => x"14",
          1670 => x"38",
          1671 => x"08",
          1672 => x"70",
          1673 => x"bb",
          1674 => x"05",
          1675 => x"54",
          1676 => x"34",
          1677 => x"05",
          1678 => x"bb",
          1679 => x"05",
          1680 => x"08",
          1681 => x"12",
          1682 => x"e8",
          1683 => x"08",
          1684 => x"e8",
          1685 => x"0c",
          1686 => x"d7",
          1687 => x"e8",
          1688 => x"08",
          1689 => x"08",
          1690 => x"53",
          1691 => x"08",
          1692 => x"70",
          1693 => x"53",
          1694 => x"51",
          1695 => x"2d",
          1696 => x"08",
          1697 => x"38",
          1698 => x"08",
          1699 => x"8c",
          1700 => x"05",
          1701 => x"82",
          1702 => x"88",
          1703 => x"82",
          1704 => x"fc",
          1705 => x"53",
          1706 => x"0b",
          1707 => x"08",
          1708 => x"82",
          1709 => x"fc",
          1710 => x"bb",
          1711 => x"3d",
          1712 => x"e8",
          1713 => x"bb",
          1714 => x"82",
          1715 => x"f9",
          1716 => x"bb",
          1717 => x"05",
          1718 => x"33",
          1719 => x"70",
          1720 => x"51",
          1721 => x"80",
          1722 => x"ff",
          1723 => x"e8",
          1724 => x"0c",
          1725 => x"82",
          1726 => x"88",
          1727 => x"11",
          1728 => x"2a",
          1729 => x"51",
          1730 => x"71",
          1731 => x"c5",
          1732 => x"e8",
          1733 => x"08",
          1734 => x"08",
          1735 => x"53",
          1736 => x"33",
          1737 => x"06",
          1738 => x"85",
          1739 => x"bb",
          1740 => x"05",
          1741 => x"08",
          1742 => x"12",
          1743 => x"e8",
          1744 => x"08",
          1745 => x"70",
          1746 => x"08",
          1747 => x"51",
          1748 => x"b6",
          1749 => x"e8",
          1750 => x"08",
          1751 => x"70",
          1752 => x"81",
          1753 => x"51",
          1754 => x"2e",
          1755 => x"82",
          1756 => x"88",
          1757 => x"08",
          1758 => x"bb",
          1759 => x"05",
          1760 => x"82",
          1761 => x"fc",
          1762 => x"38",
          1763 => x"08",
          1764 => x"82",
          1765 => x"88",
          1766 => x"53",
          1767 => x"70",
          1768 => x"52",
          1769 => x"34",
          1770 => x"bb",
          1771 => x"05",
          1772 => x"39",
          1773 => x"08",
          1774 => x"70",
          1775 => x"71",
          1776 => x"a1",
          1777 => x"e8",
          1778 => x"08",
          1779 => x"08",
          1780 => x"52",
          1781 => x"51",
          1782 => x"82",
          1783 => x"70",
          1784 => x"08",
          1785 => x"52",
          1786 => x"08",
          1787 => x"80",
          1788 => x"38",
          1789 => x"08",
          1790 => x"82",
          1791 => x"f4",
          1792 => x"bb",
          1793 => x"05",
          1794 => x"33",
          1795 => x"08",
          1796 => x"52",
          1797 => x"08",
          1798 => x"ff",
          1799 => x"06",
          1800 => x"bb",
          1801 => x"05",
          1802 => x"52",
          1803 => x"e8",
          1804 => x"34",
          1805 => x"bb",
          1806 => x"05",
          1807 => x"52",
          1808 => x"e8",
          1809 => x"34",
          1810 => x"08",
          1811 => x"52",
          1812 => x"08",
          1813 => x"85",
          1814 => x"0b",
          1815 => x"08",
          1816 => x"a6",
          1817 => x"e8",
          1818 => x"08",
          1819 => x"81",
          1820 => x"0c",
          1821 => x"08",
          1822 => x"70",
          1823 => x"70",
          1824 => x"08",
          1825 => x"51",
          1826 => x"bb",
          1827 => x"05",
          1828 => x"dc",
          1829 => x"0d",
          1830 => x"0c",
          1831 => x"e8",
          1832 => x"bb",
          1833 => x"3d",
          1834 => x"e8",
          1835 => x"08",
          1836 => x"08",
          1837 => x"82",
          1838 => x"8c",
          1839 => x"bb",
          1840 => x"05",
          1841 => x"e8",
          1842 => x"08",
          1843 => x"a2",
          1844 => x"e8",
          1845 => x"08",
          1846 => x"08",
          1847 => x"26",
          1848 => x"82",
          1849 => x"f8",
          1850 => x"bb",
          1851 => x"05",
          1852 => x"82",
          1853 => x"fc",
          1854 => x"27",
          1855 => x"82",
          1856 => x"fc",
          1857 => x"bb",
          1858 => x"05",
          1859 => x"bb",
          1860 => x"05",
          1861 => x"e8",
          1862 => x"08",
          1863 => x"08",
          1864 => x"05",
          1865 => x"08",
          1866 => x"82",
          1867 => x"90",
          1868 => x"05",
          1869 => x"08",
          1870 => x"82",
          1871 => x"90",
          1872 => x"05",
          1873 => x"08",
          1874 => x"82",
          1875 => x"90",
          1876 => x"2e",
          1877 => x"82",
          1878 => x"fc",
          1879 => x"05",
          1880 => x"08",
          1881 => x"82",
          1882 => x"f8",
          1883 => x"05",
          1884 => x"08",
          1885 => x"82",
          1886 => x"fc",
          1887 => x"bb",
          1888 => x"05",
          1889 => x"71",
          1890 => x"ff",
          1891 => x"bb",
          1892 => x"05",
          1893 => x"82",
          1894 => x"90",
          1895 => x"bb",
          1896 => x"05",
          1897 => x"82",
          1898 => x"90",
          1899 => x"bb",
          1900 => x"05",
          1901 => x"ba",
          1902 => x"e8",
          1903 => x"08",
          1904 => x"82",
          1905 => x"f8",
          1906 => x"05",
          1907 => x"08",
          1908 => x"82",
          1909 => x"fc",
          1910 => x"52",
          1911 => x"82",
          1912 => x"fc",
          1913 => x"05",
          1914 => x"08",
          1915 => x"ff",
          1916 => x"bb",
          1917 => x"05",
          1918 => x"bb",
          1919 => x"85",
          1920 => x"bb",
          1921 => x"82",
          1922 => x"02",
          1923 => x"0c",
          1924 => x"82",
          1925 => x"88",
          1926 => x"bb",
          1927 => x"05",
          1928 => x"e8",
          1929 => x"08",
          1930 => x"82",
          1931 => x"fc",
          1932 => x"05",
          1933 => x"08",
          1934 => x"70",
          1935 => x"51",
          1936 => x"2e",
          1937 => x"39",
          1938 => x"08",
          1939 => x"ff",
          1940 => x"e8",
          1941 => x"0c",
          1942 => x"08",
          1943 => x"82",
          1944 => x"88",
          1945 => x"70",
          1946 => x"0c",
          1947 => x"0d",
          1948 => x"0c",
          1949 => x"e8",
          1950 => x"bb",
          1951 => x"3d",
          1952 => x"e8",
          1953 => x"08",
          1954 => x"08",
          1955 => x"82",
          1956 => x"8c",
          1957 => x"71",
          1958 => x"e8",
          1959 => x"08",
          1960 => x"bb",
          1961 => x"05",
          1962 => x"e8",
          1963 => x"08",
          1964 => x"72",
          1965 => x"e8",
          1966 => x"08",
          1967 => x"bb",
          1968 => x"05",
          1969 => x"ff",
          1970 => x"80",
          1971 => x"ff",
          1972 => x"bb",
          1973 => x"05",
          1974 => x"bb",
          1975 => x"84",
          1976 => x"bb",
          1977 => x"82",
          1978 => x"02",
          1979 => x"0c",
          1980 => x"82",
          1981 => x"88",
          1982 => x"bb",
          1983 => x"05",
          1984 => x"e8",
          1985 => x"08",
          1986 => x"08",
          1987 => x"82",
          1988 => x"90",
          1989 => x"2e",
          1990 => x"82",
          1991 => x"90",
          1992 => x"05",
          1993 => x"08",
          1994 => x"82",
          1995 => x"90",
          1996 => x"05",
          1997 => x"08",
          1998 => x"82",
          1999 => x"90",
          2000 => x"2e",
          2001 => x"bb",
          2002 => x"05",
          2003 => x"33",
          2004 => x"08",
          2005 => x"81",
          2006 => x"e8",
          2007 => x"0c",
          2008 => x"08",
          2009 => x"52",
          2010 => x"34",
          2011 => x"08",
          2012 => x"81",
          2013 => x"e8",
          2014 => x"0c",
          2015 => x"82",
          2016 => x"88",
          2017 => x"82",
          2018 => x"51",
          2019 => x"82",
          2020 => x"04",
          2021 => x"08",
          2022 => x"e8",
          2023 => x"0d",
          2024 => x"08",
          2025 => x"80",
          2026 => x"38",
          2027 => x"08",
          2028 => x"52",
          2029 => x"bb",
          2030 => x"05",
          2031 => x"82",
          2032 => x"8c",
          2033 => x"bb",
          2034 => x"05",
          2035 => x"72",
          2036 => x"53",
          2037 => x"71",
          2038 => x"38",
          2039 => x"82",
          2040 => x"88",
          2041 => x"71",
          2042 => x"e8",
          2043 => x"08",
          2044 => x"bb",
          2045 => x"05",
          2046 => x"ff",
          2047 => x"70",
          2048 => x"0b",
          2049 => x"08",
          2050 => x"81",
          2051 => x"bb",
          2052 => x"05",
          2053 => x"82",
          2054 => x"90",
          2055 => x"bb",
          2056 => x"05",
          2057 => x"84",
          2058 => x"39",
          2059 => x"08",
          2060 => x"80",
          2061 => x"38",
          2062 => x"08",
          2063 => x"70",
          2064 => x"70",
          2065 => x"0b",
          2066 => x"08",
          2067 => x"80",
          2068 => x"bb",
          2069 => x"05",
          2070 => x"82",
          2071 => x"8c",
          2072 => x"bb",
          2073 => x"05",
          2074 => x"52",
          2075 => x"38",
          2076 => x"bb",
          2077 => x"05",
          2078 => x"82",
          2079 => x"88",
          2080 => x"33",
          2081 => x"08",
          2082 => x"70",
          2083 => x"31",
          2084 => x"e8",
          2085 => x"0c",
          2086 => x"52",
          2087 => x"80",
          2088 => x"e8",
          2089 => x"0c",
          2090 => x"08",
          2091 => x"82",
          2092 => x"85",
          2093 => x"bb",
          2094 => x"82",
          2095 => x"02",
          2096 => x"0c",
          2097 => x"82",
          2098 => x"88",
          2099 => x"bb",
          2100 => x"05",
          2101 => x"e8",
          2102 => x"08",
          2103 => x"0b",
          2104 => x"08",
          2105 => x"80",
          2106 => x"bb",
          2107 => x"05",
          2108 => x"33",
          2109 => x"08",
          2110 => x"81",
          2111 => x"e8",
          2112 => x"0c",
          2113 => x"06",
          2114 => x"80",
          2115 => x"82",
          2116 => x"8c",
          2117 => x"05",
          2118 => x"08",
          2119 => x"82",
          2120 => x"8c",
          2121 => x"2e",
          2122 => x"be",
          2123 => x"e8",
          2124 => x"08",
          2125 => x"bb",
          2126 => x"05",
          2127 => x"e8",
          2128 => x"08",
          2129 => x"08",
          2130 => x"31",
          2131 => x"e8",
          2132 => x"0c",
          2133 => x"e8",
          2134 => x"08",
          2135 => x"0c",
          2136 => x"82",
          2137 => x"04",
          2138 => x"08",
          2139 => x"e8",
          2140 => x"0d",
          2141 => x"08",
          2142 => x"82",
          2143 => x"fc",
          2144 => x"bb",
          2145 => x"05",
          2146 => x"80",
          2147 => x"bb",
          2148 => x"05",
          2149 => x"82",
          2150 => x"90",
          2151 => x"bb",
          2152 => x"05",
          2153 => x"82",
          2154 => x"90",
          2155 => x"bb",
          2156 => x"05",
          2157 => x"a9",
          2158 => x"e8",
          2159 => x"08",
          2160 => x"bb",
          2161 => x"05",
          2162 => x"71",
          2163 => x"bb",
          2164 => x"05",
          2165 => x"82",
          2166 => x"fc",
          2167 => x"be",
          2168 => x"e8",
          2169 => x"08",
          2170 => x"dc",
          2171 => x"3d",
          2172 => x"e8",
          2173 => x"bb",
          2174 => x"82",
          2175 => x"f9",
          2176 => x"0b",
          2177 => x"08",
          2178 => x"82",
          2179 => x"88",
          2180 => x"25",
          2181 => x"bb",
          2182 => x"05",
          2183 => x"bb",
          2184 => x"05",
          2185 => x"82",
          2186 => x"f4",
          2187 => x"bb",
          2188 => x"05",
          2189 => x"81",
          2190 => x"e8",
          2191 => x"0c",
          2192 => x"08",
          2193 => x"82",
          2194 => x"fc",
          2195 => x"bb",
          2196 => x"05",
          2197 => x"b9",
          2198 => x"e8",
          2199 => x"08",
          2200 => x"e8",
          2201 => x"0c",
          2202 => x"bb",
          2203 => x"05",
          2204 => x"e8",
          2205 => x"08",
          2206 => x"0b",
          2207 => x"08",
          2208 => x"82",
          2209 => x"f0",
          2210 => x"bb",
          2211 => x"05",
          2212 => x"82",
          2213 => x"8c",
          2214 => x"82",
          2215 => x"88",
          2216 => x"82",
          2217 => x"bb",
          2218 => x"82",
          2219 => x"f8",
          2220 => x"82",
          2221 => x"fc",
          2222 => x"2e",
          2223 => x"bb",
          2224 => x"05",
          2225 => x"bb",
          2226 => x"05",
          2227 => x"e8",
          2228 => x"08",
          2229 => x"dc",
          2230 => x"3d",
          2231 => x"e8",
          2232 => x"bb",
          2233 => x"82",
          2234 => x"fb",
          2235 => x"0b",
          2236 => x"08",
          2237 => x"82",
          2238 => x"88",
          2239 => x"25",
          2240 => x"bb",
          2241 => x"05",
          2242 => x"bb",
          2243 => x"05",
          2244 => x"82",
          2245 => x"fc",
          2246 => x"bb",
          2247 => x"05",
          2248 => x"90",
          2249 => x"e8",
          2250 => x"08",
          2251 => x"e8",
          2252 => x"0c",
          2253 => x"bb",
          2254 => x"05",
          2255 => x"bb",
          2256 => x"05",
          2257 => x"a2",
          2258 => x"dc",
          2259 => x"bb",
          2260 => x"05",
          2261 => x"bb",
          2262 => x"05",
          2263 => x"90",
          2264 => x"e8",
          2265 => x"08",
          2266 => x"e8",
          2267 => x"0c",
          2268 => x"08",
          2269 => x"70",
          2270 => x"0c",
          2271 => x"0d",
          2272 => x"0c",
          2273 => x"e8",
          2274 => x"bb",
          2275 => x"3d",
          2276 => x"82",
          2277 => x"8c",
          2278 => x"82",
          2279 => x"88",
          2280 => x"80",
          2281 => x"bb",
          2282 => x"82",
          2283 => x"54",
          2284 => x"82",
          2285 => x"04",
          2286 => x"08",
          2287 => x"e8",
          2288 => x"0d",
          2289 => x"bb",
          2290 => x"05",
          2291 => x"bb",
          2292 => x"05",
          2293 => x"3f",
          2294 => x"08",
          2295 => x"dc",
          2296 => x"3d",
          2297 => x"e8",
          2298 => x"bb",
          2299 => x"82",
          2300 => x"fd",
          2301 => x"0b",
          2302 => x"08",
          2303 => x"80",
          2304 => x"e8",
          2305 => x"0c",
          2306 => x"08",
          2307 => x"82",
          2308 => x"88",
          2309 => x"b9",
          2310 => x"e8",
          2311 => x"08",
          2312 => x"38",
          2313 => x"bb",
          2314 => x"05",
          2315 => x"38",
          2316 => x"08",
          2317 => x"10",
          2318 => x"08",
          2319 => x"82",
          2320 => x"fc",
          2321 => x"82",
          2322 => x"fc",
          2323 => x"b8",
          2324 => x"e8",
          2325 => x"08",
          2326 => x"e1",
          2327 => x"e8",
          2328 => x"08",
          2329 => x"08",
          2330 => x"26",
          2331 => x"bb",
          2332 => x"05",
          2333 => x"e8",
          2334 => x"08",
          2335 => x"e8",
          2336 => x"0c",
          2337 => x"08",
          2338 => x"82",
          2339 => x"fc",
          2340 => x"82",
          2341 => x"f8",
          2342 => x"bb",
          2343 => x"05",
          2344 => x"82",
          2345 => x"fc",
          2346 => x"bb",
          2347 => x"05",
          2348 => x"82",
          2349 => x"8c",
          2350 => x"95",
          2351 => x"e8",
          2352 => x"08",
          2353 => x"38",
          2354 => x"08",
          2355 => x"70",
          2356 => x"08",
          2357 => x"51",
          2358 => x"bb",
          2359 => x"05",
          2360 => x"bb",
          2361 => x"05",
          2362 => x"bb",
          2363 => x"05",
          2364 => x"dc",
          2365 => x"0d",
          2366 => x"0c",
          2367 => x"e8",
          2368 => x"bb",
          2369 => x"3d",
          2370 => x"82",
          2371 => x"f0",
          2372 => x"bb",
          2373 => x"05",
          2374 => x"73",
          2375 => x"e8",
          2376 => x"08",
          2377 => x"53",
          2378 => x"72",
          2379 => x"08",
          2380 => x"72",
          2381 => x"53",
          2382 => x"09",
          2383 => x"38",
          2384 => x"08",
          2385 => x"70",
          2386 => x"71",
          2387 => x"39",
          2388 => x"08",
          2389 => x"53",
          2390 => x"09",
          2391 => x"38",
          2392 => x"bb",
          2393 => x"05",
          2394 => x"e8",
          2395 => x"08",
          2396 => x"05",
          2397 => x"08",
          2398 => x"33",
          2399 => x"08",
          2400 => x"82",
          2401 => x"f8",
          2402 => x"72",
          2403 => x"81",
          2404 => x"38",
          2405 => x"08",
          2406 => x"70",
          2407 => x"71",
          2408 => x"51",
          2409 => x"82",
          2410 => x"f8",
          2411 => x"bb",
          2412 => x"05",
          2413 => x"e8",
          2414 => x"0c",
          2415 => x"08",
          2416 => x"80",
          2417 => x"38",
          2418 => x"08",
          2419 => x"80",
          2420 => x"38",
          2421 => x"90",
          2422 => x"e8",
          2423 => x"34",
          2424 => x"08",
          2425 => x"70",
          2426 => x"71",
          2427 => x"51",
          2428 => x"82",
          2429 => x"f8",
          2430 => x"a4",
          2431 => x"82",
          2432 => x"f4",
          2433 => x"bb",
          2434 => x"05",
          2435 => x"81",
          2436 => x"70",
          2437 => x"72",
          2438 => x"e8",
          2439 => x"34",
          2440 => x"82",
          2441 => x"f8",
          2442 => x"72",
          2443 => x"38",
          2444 => x"bb",
          2445 => x"05",
          2446 => x"39",
          2447 => x"08",
          2448 => x"53",
          2449 => x"90",
          2450 => x"e8",
          2451 => x"33",
          2452 => x"26",
          2453 => x"39",
          2454 => x"bb",
          2455 => x"05",
          2456 => x"39",
          2457 => x"bb",
          2458 => x"05",
          2459 => x"82",
          2460 => x"f8",
          2461 => x"af",
          2462 => x"38",
          2463 => x"08",
          2464 => x"53",
          2465 => x"83",
          2466 => x"80",
          2467 => x"e8",
          2468 => x"0c",
          2469 => x"8a",
          2470 => x"e8",
          2471 => x"34",
          2472 => x"bb",
          2473 => x"05",
          2474 => x"e8",
          2475 => x"33",
          2476 => x"27",
          2477 => x"82",
          2478 => x"f8",
          2479 => x"80",
          2480 => x"94",
          2481 => x"e8",
          2482 => x"33",
          2483 => x"53",
          2484 => x"e8",
          2485 => x"34",
          2486 => x"08",
          2487 => x"d0",
          2488 => x"72",
          2489 => x"08",
          2490 => x"82",
          2491 => x"f8",
          2492 => x"90",
          2493 => x"38",
          2494 => x"08",
          2495 => x"f9",
          2496 => x"72",
          2497 => x"08",
          2498 => x"82",
          2499 => x"f8",
          2500 => x"72",
          2501 => x"38",
          2502 => x"bb",
          2503 => x"05",
          2504 => x"39",
          2505 => x"08",
          2506 => x"82",
          2507 => x"f4",
          2508 => x"54",
          2509 => x"8d",
          2510 => x"82",
          2511 => x"ec",
          2512 => x"f7",
          2513 => x"e8",
          2514 => x"33",
          2515 => x"e8",
          2516 => x"08",
          2517 => x"e8",
          2518 => x"33",
          2519 => x"bb",
          2520 => x"05",
          2521 => x"e8",
          2522 => x"08",
          2523 => x"05",
          2524 => x"08",
          2525 => x"55",
          2526 => x"82",
          2527 => x"f8",
          2528 => x"a5",
          2529 => x"e8",
          2530 => x"33",
          2531 => x"2e",
          2532 => x"bb",
          2533 => x"05",
          2534 => x"bb",
          2535 => x"05",
          2536 => x"e8",
          2537 => x"08",
          2538 => x"08",
          2539 => x"71",
          2540 => x"0b",
          2541 => x"08",
          2542 => x"82",
          2543 => x"ec",
          2544 => x"bb",
          2545 => x"3d",
          2546 => x"e8",
          2547 => x"bb",
          2548 => x"82",
          2549 => x"f7",
          2550 => x"0b",
          2551 => x"08",
          2552 => x"82",
          2553 => x"8c",
          2554 => x"80",
          2555 => x"bb",
          2556 => x"05",
          2557 => x"51",
          2558 => x"53",
          2559 => x"e8",
          2560 => x"34",
          2561 => x"06",
          2562 => x"2e",
          2563 => x"91",
          2564 => x"e8",
          2565 => x"08",
          2566 => x"05",
          2567 => x"ce",
          2568 => x"e8",
          2569 => x"33",
          2570 => x"2e",
          2571 => x"a4",
          2572 => x"82",
          2573 => x"f0",
          2574 => x"bb",
          2575 => x"05",
          2576 => x"81",
          2577 => x"70",
          2578 => x"72",
          2579 => x"e8",
          2580 => x"34",
          2581 => x"08",
          2582 => x"53",
          2583 => x"09",
          2584 => x"dc",
          2585 => x"e8",
          2586 => x"08",
          2587 => x"05",
          2588 => x"08",
          2589 => x"33",
          2590 => x"08",
          2591 => x"82",
          2592 => x"f8",
          2593 => x"bb",
          2594 => x"05",
          2595 => x"e8",
          2596 => x"08",
          2597 => x"b6",
          2598 => x"e8",
          2599 => x"08",
          2600 => x"84",
          2601 => x"39",
          2602 => x"bb",
          2603 => x"05",
          2604 => x"e8",
          2605 => x"08",
          2606 => x"05",
          2607 => x"08",
          2608 => x"33",
          2609 => x"08",
          2610 => x"81",
          2611 => x"0b",
          2612 => x"08",
          2613 => x"82",
          2614 => x"88",
          2615 => x"08",
          2616 => x"0c",
          2617 => x"53",
          2618 => x"bb",
          2619 => x"05",
          2620 => x"39",
          2621 => x"08",
          2622 => x"53",
          2623 => x"8d",
          2624 => x"82",
          2625 => x"ec",
          2626 => x"80",
          2627 => x"e8",
          2628 => x"33",
          2629 => x"27",
          2630 => x"bb",
          2631 => x"05",
          2632 => x"b9",
          2633 => x"8d",
          2634 => x"82",
          2635 => x"ec",
          2636 => x"d8",
          2637 => x"82",
          2638 => x"f4",
          2639 => x"39",
          2640 => x"08",
          2641 => x"53",
          2642 => x"90",
          2643 => x"e8",
          2644 => x"33",
          2645 => x"26",
          2646 => x"39",
          2647 => x"bb",
          2648 => x"05",
          2649 => x"39",
          2650 => x"bb",
          2651 => x"05",
          2652 => x"82",
          2653 => x"fc",
          2654 => x"bb",
          2655 => x"05",
          2656 => x"73",
          2657 => x"38",
          2658 => x"08",
          2659 => x"53",
          2660 => x"27",
          2661 => x"bb",
          2662 => x"05",
          2663 => x"51",
          2664 => x"bb",
          2665 => x"05",
          2666 => x"e8",
          2667 => x"33",
          2668 => x"53",
          2669 => x"e8",
          2670 => x"34",
          2671 => x"08",
          2672 => x"53",
          2673 => x"ad",
          2674 => x"e8",
          2675 => x"33",
          2676 => x"53",
          2677 => x"e8",
          2678 => x"34",
          2679 => x"08",
          2680 => x"53",
          2681 => x"8d",
          2682 => x"82",
          2683 => x"ec",
          2684 => x"98",
          2685 => x"e8",
          2686 => x"33",
          2687 => x"08",
          2688 => x"54",
          2689 => x"26",
          2690 => x"0b",
          2691 => x"08",
          2692 => x"80",
          2693 => x"bb",
          2694 => x"05",
          2695 => x"bb",
          2696 => x"05",
          2697 => x"bb",
          2698 => x"05",
          2699 => x"82",
          2700 => x"fc",
          2701 => x"bb",
          2702 => x"05",
          2703 => x"81",
          2704 => x"70",
          2705 => x"52",
          2706 => x"33",
          2707 => x"08",
          2708 => x"fe",
          2709 => x"bb",
          2710 => x"05",
          2711 => x"80",
          2712 => x"82",
          2713 => x"fc",
          2714 => x"82",
          2715 => x"fc",
          2716 => x"bb",
          2717 => x"05",
          2718 => x"e8",
          2719 => x"08",
          2720 => x"81",
          2721 => x"e8",
          2722 => x"0c",
          2723 => x"08",
          2724 => x"82",
          2725 => x"8b",
          2726 => x"bb",
          2727 => x"f9",
          2728 => x"70",
          2729 => x"56",
          2730 => x"2e",
          2731 => x"95",
          2732 => x"51",
          2733 => x"82",
          2734 => x"15",
          2735 => x"16",
          2736 => x"cd",
          2737 => x"54",
          2738 => x"09",
          2739 => x"38",
          2740 => x"f1",
          2741 => x"76",
          2742 => x"b6",
          2743 => x"08",
          2744 => x"a3",
          2745 => x"dc",
          2746 => x"52",
          2747 => x"e9",
          2748 => x"bb",
          2749 => x"38",
          2750 => x"54",
          2751 => x"ff",
          2752 => x"17",
          2753 => x"06",
          2754 => x"77",
          2755 => x"ff",
          2756 => x"bb",
          2757 => x"3d",
          2758 => x"3d",
          2759 => x"71",
          2760 => x"8e",
          2761 => x"29",
          2762 => x"05",
          2763 => x"04",
          2764 => x"51",
          2765 => x"82",
          2766 => x"80",
          2767 => x"a0",
          2768 => x"f2",
          2769 => x"94",
          2770 => x"39",
          2771 => x"51",
          2772 => x"82",
          2773 => x"80",
          2774 => x"a0",
          2775 => x"d6",
          2776 => x"d8",
          2777 => x"39",
          2778 => x"51",
          2779 => x"82",
          2780 => x"80",
          2781 => x"a1",
          2782 => x"39",
          2783 => x"51",
          2784 => x"a1",
          2785 => x"39",
          2786 => x"51",
          2787 => x"a2",
          2788 => x"39",
          2789 => x"51",
          2790 => x"a2",
          2791 => x"39",
          2792 => x"51",
          2793 => x"a2",
          2794 => x"39",
          2795 => x"51",
          2796 => x"a3",
          2797 => x"ad",
          2798 => x"0d",
          2799 => x"0d",
          2800 => x"56",
          2801 => x"26",
          2802 => x"52",
          2803 => x"29",
          2804 => x"87",
          2805 => x"51",
          2806 => x"82",
          2807 => x"52",
          2808 => x"a1",
          2809 => x"dc",
          2810 => x"53",
          2811 => x"a3",
          2812 => x"bb",
          2813 => x"3d",
          2814 => x"3d",
          2815 => x"84",
          2816 => x"05",
          2817 => x"80",
          2818 => x"70",
          2819 => x"25",
          2820 => x"59",
          2821 => x"87",
          2822 => x"38",
          2823 => x"76",
          2824 => x"ff",
          2825 => x"93",
          2826 => x"82",
          2827 => x"76",
          2828 => x"70",
          2829 => x"84",
          2830 => x"bb",
          2831 => x"82",
          2832 => x"b9",
          2833 => x"dc",
          2834 => x"98",
          2835 => x"bb",
          2836 => x"96",
          2837 => x"54",
          2838 => x"77",
          2839 => x"81",
          2840 => x"82",
          2841 => x"57",
          2842 => x"08",
          2843 => x"55",
          2844 => x"89",
          2845 => x"75",
          2846 => x"d7",
          2847 => x"d8",
          2848 => x"90",
          2849 => x"30",
          2850 => x"80",
          2851 => x"70",
          2852 => x"06",
          2853 => x"56",
          2854 => x"90",
          2855 => x"c0",
          2856 => x"98",
          2857 => x"78",
          2858 => x"3f",
          2859 => x"82",
          2860 => x"96",
          2861 => x"f8",
          2862 => x"02",
          2863 => x"05",
          2864 => x"ff",
          2865 => x"7b",
          2866 => x"fe",
          2867 => x"bb",
          2868 => x"38",
          2869 => x"88",
          2870 => x"2e",
          2871 => x"39",
          2872 => x"56",
          2873 => x"54",
          2874 => x"53",
          2875 => x"51",
          2876 => x"bb",
          2877 => x"83",
          2878 => x"77",
          2879 => x"0c",
          2880 => x"04",
          2881 => x"7f",
          2882 => x"8c",
          2883 => x"05",
          2884 => x"15",
          2885 => x"5c",
          2886 => x"5e",
          2887 => x"a3",
          2888 => x"b9",
          2889 => x"a3",
          2890 => x"b9",
          2891 => x"55",
          2892 => x"81",
          2893 => x"90",
          2894 => x"7b",
          2895 => x"38",
          2896 => x"74",
          2897 => x"7a",
          2898 => x"72",
          2899 => x"a3",
          2900 => x"b9",
          2901 => x"39",
          2902 => x"51",
          2903 => x"3f",
          2904 => x"80",
          2905 => x"18",
          2906 => x"27",
          2907 => x"08",
          2908 => x"c8",
          2909 => x"e2",
          2910 => x"82",
          2911 => x"ff",
          2912 => x"84",
          2913 => x"39",
          2914 => x"72",
          2915 => x"38",
          2916 => x"82",
          2917 => x"ff",
          2918 => x"89",
          2919 => x"f0",
          2920 => x"b6",
          2921 => x"55",
          2922 => x"08",
          2923 => x"d8",
          2924 => x"fc",
          2925 => x"f4",
          2926 => x"9e",
          2927 => x"74",
          2928 => x"c6",
          2929 => x"70",
          2930 => x"80",
          2931 => x"27",
          2932 => x"56",
          2933 => x"74",
          2934 => x"81",
          2935 => x"06",
          2936 => x"06",
          2937 => x"80",
          2938 => x"73",
          2939 => x"8a",
          2940 => x"b0",
          2941 => x"51",
          2942 => x"d3",
          2943 => x"a0",
          2944 => x"3f",
          2945 => x"ff",
          2946 => x"a3",
          2947 => x"d5",
          2948 => x"79",
          2949 => x"a0",
          2950 => x"bb",
          2951 => x"2b",
          2952 => x"51",
          2953 => x"2e",
          2954 => x"aa",
          2955 => x"3f",
          2956 => x"08",
          2957 => x"98",
          2958 => x"32",
          2959 => x"9b",
          2960 => x"70",
          2961 => x"75",
          2962 => x"58",
          2963 => x"51",
          2964 => x"24",
          2965 => x"9b",
          2966 => x"06",
          2967 => x"53",
          2968 => x"1e",
          2969 => x"26",
          2970 => x"ff",
          2971 => x"bb",
          2972 => x"3d",
          2973 => x"3d",
          2974 => x"05",
          2975 => x"fc",
          2976 => x"84",
          2977 => x"b6",
          2978 => x"ba",
          2979 => x"a9",
          2980 => x"a4",
          2981 => x"a4",
          2982 => x"ba",
          2983 => x"82",
          2984 => x"ff",
          2985 => x"74",
          2986 => x"38",
          2987 => x"86",
          2988 => x"fe",
          2989 => x"c0",
          2990 => x"53",
          2991 => x"81",
          2992 => x"3f",
          2993 => x"51",
          2994 => x"80",
          2995 => x"3f",
          2996 => x"70",
          2997 => x"52",
          2998 => x"92",
          2999 => x"9c",
          3000 => x"a4",
          3001 => x"b8",
          3002 => x"9c",
          3003 => x"82",
          3004 => x"06",
          3005 => x"80",
          3006 => x"81",
          3007 => x"3f",
          3008 => x"51",
          3009 => x"80",
          3010 => x"3f",
          3011 => x"70",
          3012 => x"52",
          3013 => x"92",
          3014 => x"9b",
          3015 => x"a4",
          3016 => x"fc",
          3017 => x"9b",
          3018 => x"84",
          3019 => x"06",
          3020 => x"80",
          3021 => x"81",
          3022 => x"3f",
          3023 => x"51",
          3024 => x"80",
          3025 => x"3f",
          3026 => x"70",
          3027 => x"52",
          3028 => x"92",
          3029 => x"9b",
          3030 => x"a5",
          3031 => x"c0",
          3032 => x"9b",
          3033 => x"86",
          3034 => x"06",
          3035 => x"80",
          3036 => x"81",
          3037 => x"3f",
          3038 => x"51",
          3039 => x"80",
          3040 => x"3f",
          3041 => x"70",
          3042 => x"52",
          3043 => x"92",
          3044 => x"9a",
          3045 => x"a5",
          3046 => x"84",
          3047 => x"9a",
          3048 => x"88",
          3049 => x"06",
          3050 => x"80",
          3051 => x"81",
          3052 => x"3f",
          3053 => x"51",
          3054 => x"80",
          3055 => x"3f",
          3056 => x"84",
          3057 => x"fb",
          3058 => x"02",
          3059 => x"05",
          3060 => x"56",
          3061 => x"75",
          3062 => x"3f",
          3063 => x"b6",
          3064 => x"73",
          3065 => x"53",
          3066 => x"52",
          3067 => x"51",
          3068 => x"3f",
          3069 => x"08",
          3070 => x"bb",
          3071 => x"80",
          3072 => x"31",
          3073 => x"73",
          3074 => x"b6",
          3075 => x"0b",
          3076 => x"33",
          3077 => x"2e",
          3078 => x"af",
          3079 => x"dc",
          3080 => x"75",
          3081 => x"b0",
          3082 => x"dc",
          3083 => x"8b",
          3084 => x"dc",
          3085 => x"ad",
          3086 => x"82",
          3087 => x"81",
          3088 => x"82",
          3089 => x"82",
          3090 => x"0b",
          3091 => x"d8",
          3092 => x"82",
          3093 => x"06",
          3094 => x"a6",
          3095 => x"52",
          3096 => x"b2",
          3097 => x"82",
          3098 => x"87",
          3099 => x"ce",
          3100 => x"70",
          3101 => x"d8",
          3102 => x"81",
          3103 => x"80",
          3104 => x"82",
          3105 => x"81",
          3106 => x"78",
          3107 => x"81",
          3108 => x"96",
          3109 => x"53",
          3110 => x"52",
          3111 => x"c7",
          3112 => x"78",
          3113 => x"88",
          3114 => x"e5",
          3115 => x"dc",
          3116 => x"88",
          3117 => x"b8",
          3118 => x"39",
          3119 => x"5d",
          3120 => x"51",
          3121 => x"3f",
          3122 => x"46",
          3123 => x"52",
          3124 => x"f3",
          3125 => x"ff",
          3126 => x"f3",
          3127 => x"bb",
          3128 => x"2b",
          3129 => x"51",
          3130 => x"c1",
          3131 => x"38",
          3132 => x"24",
          3133 => x"78",
          3134 => x"b9",
          3135 => x"24",
          3136 => x"82",
          3137 => x"38",
          3138 => x"8a",
          3139 => x"2e",
          3140 => x"8f",
          3141 => x"84",
          3142 => x"38",
          3143 => x"82",
          3144 => x"f1",
          3145 => x"2e",
          3146 => x"78",
          3147 => x"38",
          3148 => x"83",
          3149 => x"bc",
          3150 => x"38",
          3151 => x"78",
          3152 => x"c4",
          3153 => x"c0",
          3154 => x"38",
          3155 => x"78",
          3156 => x"8d",
          3157 => x"80",
          3158 => x"38",
          3159 => x"2e",
          3160 => x"78",
          3161 => x"92",
          3162 => x"c2",
          3163 => x"38",
          3164 => x"2e",
          3165 => x"8e",
          3166 => x"80",
          3167 => x"ca",
          3168 => x"d4",
          3169 => x"38",
          3170 => x"78",
          3171 => x"8d",
          3172 => x"81",
          3173 => x"38",
          3174 => x"2e",
          3175 => x"78",
          3176 => x"8d",
          3177 => x"ed",
          3178 => x"83",
          3179 => x"38",
          3180 => x"2e",
          3181 => x"8d",
          3182 => x"3d",
          3183 => x"53",
          3184 => x"51",
          3185 => x"82",
          3186 => x"88",
          3187 => x"f4",
          3188 => x"39",
          3189 => x"fc",
          3190 => x"84",
          3191 => x"ee",
          3192 => x"dc",
          3193 => x"88",
          3194 => x"25",
          3195 => x"43",
          3196 => x"05",
          3197 => x"80",
          3198 => x"51",
          3199 => x"3f",
          3200 => x"08",
          3201 => x"59",
          3202 => x"82",
          3203 => x"cb",
          3204 => x"5e",
          3205 => x"82",
          3206 => x"8e",
          3207 => x"3d",
          3208 => x"53",
          3209 => x"51",
          3210 => x"82",
          3211 => x"80",
          3212 => x"38",
          3213 => x"52",
          3214 => x"05",
          3215 => x"cc",
          3216 => x"bb",
          3217 => x"82",
          3218 => x"8c",
          3219 => x"3d",
          3220 => x"53",
          3221 => x"51",
          3222 => x"82",
          3223 => x"80",
          3224 => x"63",
          3225 => x"d8",
          3226 => x"fe",
          3227 => x"ff",
          3228 => x"ea",
          3229 => x"bb",
          3230 => x"38",
          3231 => x"08",
          3232 => x"82",
          3233 => x"79",
          3234 => x"b6",
          3235 => x"cb",
          3236 => x"79",
          3237 => x"b4",
          3238 => x"88",
          3239 => x"f6",
          3240 => x"bb",
          3241 => x"8c",
          3242 => x"84",
          3243 => x"3f",
          3244 => x"8c",
          3245 => x"ff",
          3246 => x"8f",
          3247 => x"bb",
          3248 => x"3d",
          3249 => x"52",
          3250 => x"3f",
          3251 => x"bb",
          3252 => x"7a",
          3253 => x"3f",
          3254 => x"b4",
          3255 => x"05",
          3256 => x"3f",
          3257 => x"08",
          3258 => x"84",
          3259 => x"90",
          3260 => x"bb",
          3261 => x"3d",
          3262 => x"52",
          3263 => x"3f",
          3264 => x"08",
          3265 => x"84",
          3266 => x"90",
          3267 => x"ba",
          3268 => x"bc",
          3269 => x"56",
          3270 => x"bb",
          3271 => x"ff",
          3272 => x"53",
          3273 => x"51",
          3274 => x"82",
          3275 => x"80",
          3276 => x"38",
          3277 => x"08",
          3278 => x"3f",
          3279 => x"b4",
          3280 => x"11",
          3281 => x"05",
          3282 => x"3f",
          3283 => x"08",
          3284 => x"ec",
          3285 => x"fe",
          3286 => x"ff",
          3287 => x"e8",
          3288 => x"bb",
          3289 => x"2e",
          3290 => x"b4",
          3291 => x"11",
          3292 => x"05",
          3293 => x"3f",
          3294 => x"08",
          3295 => x"bb",
          3296 => x"82",
          3297 => x"ff",
          3298 => x"63",
          3299 => x"79",
          3300 => x"ec",
          3301 => x"78",
          3302 => x"05",
          3303 => x"7a",
          3304 => x"81",
          3305 => x"3d",
          3306 => x"53",
          3307 => x"51",
          3308 => x"82",
          3309 => x"80",
          3310 => x"38",
          3311 => x"fc",
          3312 => x"84",
          3313 => x"86",
          3314 => x"dc",
          3315 => x"f9",
          3316 => x"3d",
          3317 => x"53",
          3318 => x"51",
          3319 => x"82",
          3320 => x"80",
          3321 => x"38",
          3322 => x"51",
          3323 => x"3f",
          3324 => x"63",
          3325 => x"38",
          3326 => x"70",
          3327 => x"33",
          3328 => x"81",
          3329 => x"39",
          3330 => x"80",
          3331 => x"84",
          3332 => x"ba",
          3333 => x"dc",
          3334 => x"f9",
          3335 => x"3d",
          3336 => x"53",
          3337 => x"51",
          3338 => x"82",
          3339 => x"80",
          3340 => x"38",
          3341 => x"f8",
          3342 => x"84",
          3343 => x"8e",
          3344 => x"dc",
          3345 => x"f8",
          3346 => x"a7",
          3347 => x"ab",
          3348 => x"5a",
          3349 => x"a8",
          3350 => x"33",
          3351 => x"5a",
          3352 => x"2e",
          3353 => x"55",
          3354 => x"33",
          3355 => x"82",
          3356 => x"ff",
          3357 => x"81",
          3358 => x"05",
          3359 => x"39",
          3360 => x"83",
          3361 => x"39",
          3362 => x"80",
          3363 => x"84",
          3364 => x"ba",
          3365 => x"dc",
          3366 => x"38",
          3367 => x"33",
          3368 => x"2e",
          3369 => x"ba",
          3370 => x"80",
          3371 => x"ba",
          3372 => x"78",
          3373 => x"38",
          3374 => x"08",
          3375 => x"82",
          3376 => x"59",
          3377 => x"88",
          3378 => x"90",
          3379 => x"39",
          3380 => x"33",
          3381 => x"2e",
          3382 => x"ba",
          3383 => x"9a",
          3384 => x"c6",
          3385 => x"80",
          3386 => x"82",
          3387 => x"44",
          3388 => x"ba",
          3389 => x"80",
          3390 => x"3d",
          3391 => x"53",
          3392 => x"51",
          3393 => x"82",
          3394 => x"80",
          3395 => x"ba",
          3396 => x"78",
          3397 => x"38",
          3398 => x"08",
          3399 => x"39",
          3400 => x"33",
          3401 => x"2e",
          3402 => x"ba",
          3403 => x"bb",
          3404 => x"ca",
          3405 => x"80",
          3406 => x"82",
          3407 => x"43",
          3408 => x"ba",
          3409 => x"78",
          3410 => x"38",
          3411 => x"08",
          3412 => x"82",
          3413 => x"59",
          3414 => x"88",
          3415 => x"a4",
          3416 => x"39",
          3417 => x"08",
          3418 => x"b4",
          3419 => x"11",
          3420 => x"05",
          3421 => x"3f",
          3422 => x"08",
          3423 => x"38",
          3424 => x"5c",
          3425 => x"83",
          3426 => x"7a",
          3427 => x"30",
          3428 => x"9f",
          3429 => x"06",
          3430 => x"5a",
          3431 => x"88",
          3432 => x"2e",
          3433 => x"42",
          3434 => x"51",
          3435 => x"a0",
          3436 => x"61",
          3437 => x"63",
          3438 => x"3f",
          3439 => x"51",
          3440 => x"b4",
          3441 => x"11",
          3442 => x"05",
          3443 => x"3f",
          3444 => x"08",
          3445 => x"e8",
          3446 => x"fe",
          3447 => x"ff",
          3448 => x"e3",
          3449 => x"bb",
          3450 => x"2e",
          3451 => x"59",
          3452 => x"05",
          3453 => x"63",
          3454 => x"b4",
          3455 => x"11",
          3456 => x"05",
          3457 => x"3f",
          3458 => x"08",
          3459 => x"b0",
          3460 => x"33",
          3461 => x"a8",
          3462 => x"a7",
          3463 => x"d3",
          3464 => x"80",
          3465 => x"51",
          3466 => x"3f",
          3467 => x"33",
          3468 => x"2e",
          3469 => x"9f",
          3470 => x"38",
          3471 => x"fc",
          3472 => x"84",
          3473 => x"86",
          3474 => x"dc",
          3475 => x"91",
          3476 => x"02",
          3477 => x"33",
          3478 => x"81",
          3479 => x"b1",
          3480 => x"a4",
          3481 => x"3f",
          3482 => x"b4",
          3483 => x"11",
          3484 => x"05",
          3485 => x"3f",
          3486 => x"08",
          3487 => x"c0",
          3488 => x"fe",
          3489 => x"ff",
          3490 => x"dc",
          3491 => x"bb",
          3492 => x"2e",
          3493 => x"59",
          3494 => x"22",
          3495 => x"05",
          3496 => x"41",
          3497 => x"f0",
          3498 => x"84",
          3499 => x"cd",
          3500 => x"dc",
          3501 => x"f4",
          3502 => x"70",
          3503 => x"82",
          3504 => x"ff",
          3505 => x"82",
          3506 => x"53",
          3507 => x"79",
          3508 => x"db",
          3509 => x"79",
          3510 => x"ae",
          3511 => x"38",
          3512 => x"87",
          3513 => x"05",
          3514 => x"b4",
          3515 => x"11",
          3516 => x"05",
          3517 => x"3f",
          3518 => x"08",
          3519 => x"38",
          3520 => x"be",
          3521 => x"70",
          3522 => x"23",
          3523 => x"aa",
          3524 => x"a4",
          3525 => x"3f",
          3526 => x"b4",
          3527 => x"11",
          3528 => x"05",
          3529 => x"3f",
          3530 => x"08",
          3531 => x"90",
          3532 => x"fe",
          3533 => x"ff",
          3534 => x"db",
          3535 => x"bb",
          3536 => x"2e",
          3537 => x"60",
          3538 => x"60",
          3539 => x"b4",
          3540 => x"11",
          3541 => x"05",
          3542 => x"3f",
          3543 => x"08",
          3544 => x"dc",
          3545 => x"08",
          3546 => x"a8",
          3547 => x"a4",
          3548 => x"d3",
          3549 => x"80",
          3550 => x"51",
          3551 => x"3f",
          3552 => x"33",
          3553 => x"2e",
          3554 => x"9f",
          3555 => x"38",
          3556 => x"f0",
          3557 => x"84",
          3558 => x"e1",
          3559 => x"dc",
          3560 => x"8d",
          3561 => x"71",
          3562 => x"84",
          3563 => x"b5",
          3564 => x"a4",
          3565 => x"3f",
          3566 => x"82",
          3567 => x"c0",
          3568 => x"51",
          3569 => x"f1",
          3570 => x"a8",
          3571 => x"95",
          3572 => x"97",
          3573 => x"e8",
          3574 => x"f0",
          3575 => x"3f",
          3576 => x"0b",
          3577 => x"84",
          3578 => x"81",
          3579 => x"94",
          3580 => x"cc",
          3581 => x"84",
          3582 => x"e9",
          3583 => x"83",
          3584 => x"94",
          3585 => x"80",
          3586 => x"c0",
          3587 => x"f1",
          3588 => x"3d",
          3589 => x"53",
          3590 => x"51",
          3591 => x"82",
          3592 => x"80",
          3593 => x"38",
          3594 => x"a9",
          3595 => x"a3",
          3596 => x"59",
          3597 => x"3d",
          3598 => x"53",
          3599 => x"51",
          3600 => x"82",
          3601 => x"80",
          3602 => x"38",
          3603 => x"a9",
          3604 => x"a3",
          3605 => x"59",
          3606 => x"bb",
          3607 => x"2e",
          3608 => x"82",
          3609 => x"52",
          3610 => x"51",
          3611 => x"3f",
          3612 => x"82",
          3613 => x"ff",
          3614 => x"ff",
          3615 => x"f0",
          3616 => x"aa",
          3617 => x"be",
          3618 => x"59",
          3619 => x"91",
          3620 => x"ac",
          3621 => x"79",
          3622 => x"80",
          3623 => x"38",
          3624 => x"59",
          3625 => x"81",
          3626 => x"3d",
          3627 => x"51",
          3628 => x"82",
          3629 => x"5b",
          3630 => x"82",
          3631 => x"7b",
          3632 => x"38",
          3633 => x"8c",
          3634 => x"39",
          3635 => x"ad",
          3636 => x"39",
          3637 => x"56",
          3638 => x"aa",
          3639 => x"53",
          3640 => x"52",
          3641 => x"b0",
          3642 => x"a4",
          3643 => x"39",
          3644 => x"3d",
          3645 => x"51",
          3646 => x"ab",
          3647 => x"82",
          3648 => x"80",
          3649 => x"b4",
          3650 => x"ff",
          3651 => x"ff",
          3652 => x"93",
          3653 => x"80",
          3654 => x"c0",
          3655 => x"ff",
          3656 => x"ff",
          3657 => x"82",
          3658 => x"82",
          3659 => x"80",
          3660 => x"80",
          3661 => x"80",
          3662 => x"80",
          3663 => x"ff",
          3664 => x"e6",
          3665 => x"bb",
          3666 => x"bb",
          3667 => x"70",
          3668 => x"07",
          3669 => x"5b",
          3670 => x"5a",
          3671 => x"83",
          3672 => x"78",
          3673 => x"78",
          3674 => x"38",
          3675 => x"81",
          3676 => x"59",
          3677 => x"38",
          3678 => x"7d",
          3679 => x"59",
          3680 => x"7e",
          3681 => x"81",
          3682 => x"38",
          3683 => x"51",
          3684 => x"3f",
          3685 => x"f5",
          3686 => x"0b",
          3687 => x"34",
          3688 => x"8c",
          3689 => x"55",
          3690 => x"52",
          3691 => x"d5",
          3692 => x"dc",
          3693 => x"75",
          3694 => x"87",
          3695 => x"73",
          3696 => x"3f",
          3697 => x"dc",
          3698 => x"0c",
          3699 => x"9c",
          3700 => x"55",
          3701 => x"52",
          3702 => x"a9",
          3703 => x"dc",
          3704 => x"75",
          3705 => x"87",
          3706 => x"73",
          3707 => x"3f",
          3708 => x"dc",
          3709 => x"0c",
          3710 => x"0b",
          3711 => x"84",
          3712 => x"83",
          3713 => x"94",
          3714 => x"fa",
          3715 => x"fd",
          3716 => x"02",
          3717 => x"05",
          3718 => x"82",
          3719 => x"87",
          3720 => x"13",
          3721 => x"0c",
          3722 => x"0c",
          3723 => x"3f",
          3724 => x"82",
          3725 => x"ff",
          3726 => x"82",
          3727 => x"ff",
          3728 => x"80",
          3729 => x"92",
          3730 => x"51",
          3731 => x"ec",
          3732 => x"04",
          3733 => x"80",
          3734 => x"71",
          3735 => x"87",
          3736 => x"bb",
          3737 => x"ff",
          3738 => x"ff",
          3739 => x"72",
          3740 => x"38",
          3741 => x"dc",
          3742 => x"0d",
          3743 => x"0d",
          3744 => x"54",
          3745 => x"52",
          3746 => x"2e",
          3747 => x"72",
          3748 => x"a0",
          3749 => x"06",
          3750 => x"13",
          3751 => x"72",
          3752 => x"a2",
          3753 => x"06",
          3754 => x"13",
          3755 => x"72",
          3756 => x"2e",
          3757 => x"9f",
          3758 => x"81",
          3759 => x"72",
          3760 => x"70",
          3761 => x"38",
          3762 => x"80",
          3763 => x"73",
          3764 => x"39",
          3765 => x"80",
          3766 => x"54",
          3767 => x"83",
          3768 => x"70",
          3769 => x"38",
          3770 => x"80",
          3771 => x"54",
          3772 => x"09",
          3773 => x"38",
          3774 => x"a2",
          3775 => x"70",
          3776 => x"07",
          3777 => x"70",
          3778 => x"38",
          3779 => x"81",
          3780 => x"71",
          3781 => x"51",
          3782 => x"dc",
          3783 => x"0d",
          3784 => x"0d",
          3785 => x"08",
          3786 => x"38",
          3787 => x"05",
          3788 => x"d3",
          3789 => x"bb",
          3790 => x"38",
          3791 => x"39",
          3792 => x"82",
          3793 => x"86",
          3794 => x"fc",
          3795 => x"82",
          3796 => x"05",
          3797 => x"52",
          3798 => x"81",
          3799 => x"13",
          3800 => x"51",
          3801 => x"9e",
          3802 => x"38",
          3803 => x"51",
          3804 => x"97",
          3805 => x"38",
          3806 => x"51",
          3807 => x"bb",
          3808 => x"38",
          3809 => x"51",
          3810 => x"bb",
          3811 => x"38",
          3812 => x"55",
          3813 => x"87",
          3814 => x"d9",
          3815 => x"22",
          3816 => x"73",
          3817 => x"80",
          3818 => x"0b",
          3819 => x"9c",
          3820 => x"87",
          3821 => x"0c",
          3822 => x"87",
          3823 => x"0c",
          3824 => x"87",
          3825 => x"0c",
          3826 => x"87",
          3827 => x"0c",
          3828 => x"87",
          3829 => x"0c",
          3830 => x"87",
          3831 => x"0c",
          3832 => x"98",
          3833 => x"87",
          3834 => x"0c",
          3835 => x"c0",
          3836 => x"80",
          3837 => x"bb",
          3838 => x"3d",
          3839 => x"3d",
          3840 => x"87",
          3841 => x"5d",
          3842 => x"87",
          3843 => x"08",
          3844 => x"23",
          3845 => x"b8",
          3846 => x"82",
          3847 => x"c0",
          3848 => x"5a",
          3849 => x"34",
          3850 => x"b0",
          3851 => x"84",
          3852 => x"c0",
          3853 => x"5a",
          3854 => x"34",
          3855 => x"a8",
          3856 => x"86",
          3857 => x"c0",
          3858 => x"5c",
          3859 => x"23",
          3860 => x"a0",
          3861 => x"8a",
          3862 => x"7d",
          3863 => x"ff",
          3864 => x"7b",
          3865 => x"06",
          3866 => x"33",
          3867 => x"33",
          3868 => x"33",
          3869 => x"33",
          3870 => x"33",
          3871 => x"ff",
          3872 => x"82",
          3873 => x"ff",
          3874 => x"8f",
          3875 => x"fb",
          3876 => x"9f",
          3877 => x"b9",
          3878 => x"81",
          3879 => x"55",
          3880 => x"94",
          3881 => x"80",
          3882 => x"87",
          3883 => x"51",
          3884 => x"96",
          3885 => x"06",
          3886 => x"70",
          3887 => x"38",
          3888 => x"70",
          3889 => x"51",
          3890 => x"72",
          3891 => x"81",
          3892 => x"70",
          3893 => x"38",
          3894 => x"70",
          3895 => x"51",
          3896 => x"38",
          3897 => x"06",
          3898 => x"94",
          3899 => x"80",
          3900 => x"87",
          3901 => x"52",
          3902 => x"74",
          3903 => x"0c",
          3904 => x"04",
          3905 => x"02",
          3906 => x"70",
          3907 => x"2a",
          3908 => x"70",
          3909 => x"34",
          3910 => x"04",
          3911 => x"02",
          3912 => x"58",
          3913 => x"09",
          3914 => x"38",
          3915 => x"51",
          3916 => x"b9",
          3917 => x"81",
          3918 => x"56",
          3919 => x"84",
          3920 => x"2e",
          3921 => x"c0",
          3922 => x"72",
          3923 => x"2a",
          3924 => x"55",
          3925 => x"80",
          3926 => x"73",
          3927 => x"81",
          3928 => x"72",
          3929 => x"81",
          3930 => x"06",
          3931 => x"80",
          3932 => x"73",
          3933 => x"81",
          3934 => x"72",
          3935 => x"75",
          3936 => x"53",
          3937 => x"80",
          3938 => x"2e",
          3939 => x"c0",
          3940 => x"77",
          3941 => x"0b",
          3942 => x"0c",
          3943 => x"04",
          3944 => x"79",
          3945 => x"33",
          3946 => x"06",
          3947 => x"70",
          3948 => x"fc",
          3949 => x"ff",
          3950 => x"82",
          3951 => x"70",
          3952 => x"59",
          3953 => x"87",
          3954 => x"51",
          3955 => x"86",
          3956 => x"94",
          3957 => x"08",
          3958 => x"70",
          3959 => x"54",
          3960 => x"2e",
          3961 => x"91",
          3962 => x"06",
          3963 => x"d7",
          3964 => x"32",
          3965 => x"51",
          3966 => x"2e",
          3967 => x"93",
          3968 => x"06",
          3969 => x"ff",
          3970 => x"81",
          3971 => x"87",
          3972 => x"52",
          3973 => x"86",
          3974 => x"94",
          3975 => x"72",
          3976 => x"74",
          3977 => x"ff",
          3978 => x"57",
          3979 => x"38",
          3980 => x"dc",
          3981 => x"0d",
          3982 => x"0d",
          3983 => x"33",
          3984 => x"06",
          3985 => x"c0",
          3986 => x"72",
          3987 => x"38",
          3988 => x"94",
          3989 => x"70",
          3990 => x"81",
          3991 => x"51",
          3992 => x"e2",
          3993 => x"ff",
          3994 => x"c0",
          3995 => x"70",
          3996 => x"38",
          3997 => x"90",
          3998 => x"70",
          3999 => x"82",
          4000 => x"51",
          4001 => x"04",
          4002 => x"82",
          4003 => x"81",
          4004 => x"bb",
          4005 => x"fe",
          4006 => x"b9",
          4007 => x"81",
          4008 => x"53",
          4009 => x"84",
          4010 => x"2e",
          4011 => x"c0",
          4012 => x"71",
          4013 => x"2a",
          4014 => x"51",
          4015 => x"52",
          4016 => x"a0",
          4017 => x"ff",
          4018 => x"c0",
          4019 => x"70",
          4020 => x"38",
          4021 => x"90",
          4022 => x"70",
          4023 => x"98",
          4024 => x"51",
          4025 => x"dc",
          4026 => x"0d",
          4027 => x"0d",
          4028 => x"80",
          4029 => x"2a",
          4030 => x"51",
          4031 => x"84",
          4032 => x"c0",
          4033 => x"82",
          4034 => x"87",
          4035 => x"08",
          4036 => x"0c",
          4037 => x"94",
          4038 => x"88",
          4039 => x"9e",
          4040 => x"ba",
          4041 => x"c0",
          4042 => x"82",
          4043 => x"87",
          4044 => x"08",
          4045 => x"0c",
          4046 => x"ac",
          4047 => x"98",
          4048 => x"9e",
          4049 => x"ba",
          4050 => x"c0",
          4051 => x"82",
          4052 => x"87",
          4053 => x"08",
          4054 => x"0c",
          4055 => x"bc",
          4056 => x"a8",
          4057 => x"9e",
          4058 => x"ba",
          4059 => x"c0",
          4060 => x"82",
          4061 => x"87",
          4062 => x"08",
          4063 => x"ba",
          4064 => x"c0",
          4065 => x"82",
          4066 => x"87",
          4067 => x"08",
          4068 => x"0c",
          4069 => x"8c",
          4070 => x"c0",
          4071 => x"82",
          4072 => x"80",
          4073 => x"9e",
          4074 => x"84",
          4075 => x"51",
          4076 => x"80",
          4077 => x"81",
          4078 => x"ba",
          4079 => x"0b",
          4080 => x"90",
          4081 => x"80",
          4082 => x"52",
          4083 => x"2e",
          4084 => x"52",
          4085 => x"c6",
          4086 => x"87",
          4087 => x"08",
          4088 => x"0a",
          4089 => x"52",
          4090 => x"83",
          4091 => x"71",
          4092 => x"34",
          4093 => x"c0",
          4094 => x"70",
          4095 => x"06",
          4096 => x"70",
          4097 => x"38",
          4098 => x"82",
          4099 => x"80",
          4100 => x"9e",
          4101 => x"a0",
          4102 => x"51",
          4103 => x"80",
          4104 => x"81",
          4105 => x"ba",
          4106 => x"0b",
          4107 => x"90",
          4108 => x"80",
          4109 => x"52",
          4110 => x"2e",
          4111 => x"52",
          4112 => x"ca",
          4113 => x"87",
          4114 => x"08",
          4115 => x"80",
          4116 => x"52",
          4117 => x"83",
          4118 => x"71",
          4119 => x"34",
          4120 => x"c0",
          4121 => x"70",
          4122 => x"06",
          4123 => x"70",
          4124 => x"38",
          4125 => x"82",
          4126 => x"80",
          4127 => x"9e",
          4128 => x"81",
          4129 => x"51",
          4130 => x"80",
          4131 => x"81",
          4132 => x"ba",
          4133 => x"0b",
          4134 => x"90",
          4135 => x"c0",
          4136 => x"52",
          4137 => x"2e",
          4138 => x"52",
          4139 => x"ce",
          4140 => x"87",
          4141 => x"08",
          4142 => x"06",
          4143 => x"70",
          4144 => x"38",
          4145 => x"82",
          4146 => x"87",
          4147 => x"08",
          4148 => x"06",
          4149 => x"51",
          4150 => x"82",
          4151 => x"80",
          4152 => x"9e",
          4153 => x"84",
          4154 => x"52",
          4155 => x"2e",
          4156 => x"52",
          4157 => x"d1",
          4158 => x"9e",
          4159 => x"83",
          4160 => x"84",
          4161 => x"51",
          4162 => x"d2",
          4163 => x"87",
          4164 => x"08",
          4165 => x"51",
          4166 => x"80",
          4167 => x"81",
          4168 => x"ba",
          4169 => x"c0",
          4170 => x"70",
          4171 => x"51",
          4172 => x"d4",
          4173 => x"0d",
          4174 => x"0d",
          4175 => x"51",
          4176 => x"3f",
          4177 => x"33",
          4178 => x"2e",
          4179 => x"ab",
          4180 => x"ad",
          4181 => x"ab",
          4182 => x"ad",
          4183 => x"ba",
          4184 => x"73",
          4185 => x"38",
          4186 => x"08",
          4187 => x"08",
          4188 => x"82",
          4189 => x"ff",
          4190 => x"82",
          4191 => x"54",
          4192 => x"94",
          4193 => x"98",
          4194 => x"9c",
          4195 => x"52",
          4196 => x"51",
          4197 => x"3f",
          4198 => x"33",
          4199 => x"2e",
          4200 => x"ba",
          4201 => x"ba",
          4202 => x"54",
          4203 => x"8c",
          4204 => x"a6",
          4205 => x"c9",
          4206 => x"80",
          4207 => x"82",
          4208 => x"82",
          4209 => x"11",
          4210 => x"ac",
          4211 => x"90",
          4212 => x"ba",
          4213 => x"73",
          4214 => x"38",
          4215 => x"08",
          4216 => x"08",
          4217 => x"82",
          4218 => x"ff",
          4219 => x"82",
          4220 => x"54",
          4221 => x"8e",
          4222 => x"d0",
          4223 => x"ac",
          4224 => x"8f",
          4225 => x"ba",
          4226 => x"73",
          4227 => x"38",
          4228 => x"33",
          4229 => x"80",
          4230 => x"be",
          4231 => x"d1",
          4232 => x"80",
          4233 => x"82",
          4234 => x"52",
          4235 => x"51",
          4236 => x"3f",
          4237 => x"33",
          4238 => x"2e",
          4239 => x"ad",
          4240 => x"ab",
          4241 => x"ba",
          4242 => x"73",
          4243 => x"38",
          4244 => x"51",
          4245 => x"3f",
          4246 => x"33",
          4247 => x"2e",
          4248 => x"ad",
          4249 => x"aa",
          4250 => x"ba",
          4251 => x"73",
          4252 => x"38",
          4253 => x"51",
          4254 => x"3f",
          4255 => x"33",
          4256 => x"2e",
          4257 => x"ad",
          4258 => x"aa",
          4259 => x"ae",
          4260 => x"aa",
          4261 => x"ba",
          4262 => x"82",
          4263 => x"ff",
          4264 => x"82",
          4265 => x"52",
          4266 => x"51",
          4267 => x"3f",
          4268 => x"08",
          4269 => x"e0",
          4270 => x"9e",
          4271 => x"88",
          4272 => x"a1",
          4273 => x"b4",
          4274 => x"af",
          4275 => x"8e",
          4276 => x"ba",
          4277 => x"bd",
          4278 => x"75",
          4279 => x"3f",
          4280 => x"08",
          4281 => x"29",
          4282 => x"54",
          4283 => x"dc",
          4284 => x"af",
          4285 => x"8d",
          4286 => x"ba",
          4287 => x"73",
          4288 => x"38",
          4289 => x"08",
          4290 => x"c0",
          4291 => x"c0",
          4292 => x"bb",
          4293 => x"84",
          4294 => x"71",
          4295 => x"82",
          4296 => x"52",
          4297 => x"51",
          4298 => x"3f",
          4299 => x"33",
          4300 => x"2e",
          4301 => x"ba",
          4302 => x"bd",
          4303 => x"75",
          4304 => x"3f",
          4305 => x"08",
          4306 => x"29",
          4307 => x"54",
          4308 => x"dc",
          4309 => x"b0",
          4310 => x"8c",
          4311 => x"a7",
          4312 => x"a9",
          4313 => x"3d",
          4314 => x"3d",
          4315 => x"05",
          4316 => x"52",
          4317 => x"aa",
          4318 => x"29",
          4319 => x"05",
          4320 => x"04",
          4321 => x"51",
          4322 => x"b0",
          4323 => x"39",
          4324 => x"51",
          4325 => x"b0",
          4326 => x"39",
          4327 => x"51",
          4328 => x"b0",
          4329 => x"a8",
          4330 => x"3d",
          4331 => x"88",
          4332 => x"ff",
          4333 => x"c0",
          4334 => x"08",
          4335 => x"72",
          4336 => x"07",
          4337 => x"d8",
          4338 => x"83",
          4339 => x"ff",
          4340 => x"c0",
          4341 => x"08",
          4342 => x"0c",
          4343 => x"0c",
          4344 => x"82",
          4345 => x"06",
          4346 => x"d8",
          4347 => x"51",
          4348 => x"04",
          4349 => x"c0",
          4350 => x"04",
          4351 => x"08",
          4352 => x"84",
          4353 => x"3d",
          4354 => x"2b",
          4355 => x"79",
          4356 => x"98",
          4357 => x"13",
          4358 => x"51",
          4359 => x"51",
          4360 => x"82",
          4361 => x"33",
          4362 => x"74",
          4363 => x"82",
          4364 => x"08",
          4365 => x"05",
          4366 => x"71",
          4367 => x"52",
          4368 => x"09",
          4369 => x"38",
          4370 => x"82",
          4371 => x"85",
          4372 => x"fb",
          4373 => x"02",
          4374 => x"05",
          4375 => x"55",
          4376 => x"80",
          4377 => x"82",
          4378 => x"52",
          4379 => x"aa",
          4380 => x"d3",
          4381 => x"a0",
          4382 => x"b8",
          4383 => x"b0",
          4384 => x"51",
          4385 => x"3f",
          4386 => x"05",
          4387 => x"34",
          4388 => x"06",
          4389 => x"77",
          4390 => x"be",
          4391 => x"34",
          4392 => x"04",
          4393 => x"7c",
          4394 => x"b7",
          4395 => x"88",
          4396 => x"33",
          4397 => x"33",
          4398 => x"82",
          4399 => x"70",
          4400 => x"59",
          4401 => x"74",
          4402 => x"38",
          4403 => x"fa",
          4404 => x"b4",
          4405 => x"29",
          4406 => x"05",
          4407 => x"54",
          4408 => x"9d",
          4409 => x"bb",
          4410 => x"0c",
          4411 => x"33",
          4412 => x"82",
          4413 => x"70",
          4414 => x"5a",
          4415 => x"a7",
          4416 => x"78",
          4417 => x"ff",
          4418 => x"82",
          4419 => x"81",
          4420 => x"82",
          4421 => x"74",
          4422 => x"55",
          4423 => x"87",
          4424 => x"82",
          4425 => x"77",
          4426 => x"38",
          4427 => x"08",
          4428 => x"2e",
          4429 => x"bb",
          4430 => x"74",
          4431 => x"3d",
          4432 => x"76",
          4433 => x"75",
          4434 => x"88",
          4435 => x"b0",
          4436 => x"51",
          4437 => x"3f",
          4438 => x"08",
          4439 => x"e5",
          4440 => x"0d",
          4441 => x"0d",
          4442 => x"53",
          4443 => x"08",
          4444 => x"2e",
          4445 => x"51",
          4446 => x"80",
          4447 => x"14",
          4448 => x"54",
          4449 => x"e6",
          4450 => x"82",
          4451 => x"82",
          4452 => x"52",
          4453 => x"95",
          4454 => x"80",
          4455 => x"82",
          4456 => x"51",
          4457 => x"80",
          4458 => x"b0",
          4459 => x"0d",
          4460 => x"0d",
          4461 => x"52",
          4462 => x"08",
          4463 => x"b2",
          4464 => x"dc",
          4465 => x"38",
          4466 => x"08",
          4467 => x"52",
          4468 => x"52",
          4469 => x"80",
          4470 => x"dc",
          4471 => x"ba",
          4472 => x"ff",
          4473 => x"82",
          4474 => x"55",
          4475 => x"bb",
          4476 => x"9d",
          4477 => x"dc",
          4478 => x"70",
          4479 => x"80",
          4480 => x"53",
          4481 => x"17",
          4482 => x"52",
          4483 => x"ca",
          4484 => x"2e",
          4485 => x"ff",
          4486 => x"3d",
          4487 => x"3d",
          4488 => x"08",
          4489 => x"5a",
          4490 => x"58",
          4491 => x"82",
          4492 => x"51",
          4493 => x"3f",
          4494 => x"08",
          4495 => x"ff",
          4496 => x"b0",
          4497 => x"80",
          4498 => x"3d",
          4499 => x"81",
          4500 => x"82",
          4501 => x"80",
          4502 => x"75",
          4503 => x"a7",
          4504 => x"dc",
          4505 => x"58",
          4506 => x"82",
          4507 => x"25",
          4508 => x"bb",
          4509 => x"05",
          4510 => x"55",
          4511 => x"74",
          4512 => x"70",
          4513 => x"2a",
          4514 => x"78",
          4515 => x"38",
          4516 => x"38",
          4517 => x"08",
          4518 => x"53",
          4519 => x"d2",
          4520 => x"dc",
          4521 => x"89",
          4522 => x"e8",
          4523 => x"aa",
          4524 => x"2e",
          4525 => x"9b",
          4526 => x"79",
          4527 => x"b5",
          4528 => x"ff",
          4529 => x"ab",
          4530 => x"82",
          4531 => x"74",
          4532 => x"77",
          4533 => x"0c",
          4534 => x"04",
          4535 => x"7c",
          4536 => x"71",
          4537 => x"59",
          4538 => x"a0",
          4539 => x"06",
          4540 => x"33",
          4541 => x"77",
          4542 => x"38",
          4543 => x"5b",
          4544 => x"56",
          4545 => x"a0",
          4546 => x"06",
          4547 => x"75",
          4548 => x"80",
          4549 => x"29",
          4550 => x"05",
          4551 => x"55",
          4552 => x"3f",
          4553 => x"08",
          4554 => x"74",
          4555 => x"b0",
          4556 => x"bb",
          4557 => x"c5",
          4558 => x"33",
          4559 => x"2e",
          4560 => x"82",
          4561 => x"b5",
          4562 => x"3f",
          4563 => x"1a",
          4564 => x"fc",
          4565 => x"05",
          4566 => x"3f",
          4567 => x"08",
          4568 => x"38",
          4569 => x"78",
          4570 => x"fd",
          4571 => x"bb",
          4572 => x"ff",
          4573 => x"85",
          4574 => x"91",
          4575 => x"70",
          4576 => x"51",
          4577 => x"27",
          4578 => x"80",
          4579 => x"bb",
          4580 => x"3d",
          4581 => x"3d",
          4582 => x"08",
          4583 => x"b4",
          4584 => x"5f",
          4585 => x"af",
          4586 => x"bb",
          4587 => x"bb",
          4588 => x"5b",
          4589 => x"38",
          4590 => x"ac",
          4591 => x"73",
          4592 => x"55",
          4593 => x"81",
          4594 => x"70",
          4595 => x"56",
          4596 => x"81",
          4597 => x"51",
          4598 => x"82",
          4599 => x"82",
          4600 => x"82",
          4601 => x"80",
          4602 => x"38",
          4603 => x"52",
          4604 => x"08",
          4605 => x"fa",
          4606 => x"dc",
          4607 => x"8c",
          4608 => x"94",
          4609 => x"dd",
          4610 => x"39",
          4611 => x"08",
          4612 => x"b0",
          4613 => x"f8",
          4614 => x"70",
          4615 => x"87",
          4616 => x"bb",
          4617 => x"82",
          4618 => x"74",
          4619 => x"06",
          4620 => x"82",
          4621 => x"51",
          4622 => x"3f",
          4623 => x"08",
          4624 => x"82",
          4625 => x"25",
          4626 => x"bb",
          4627 => x"05",
          4628 => x"55",
          4629 => x"80",
          4630 => x"ff",
          4631 => x"51",
          4632 => x"81",
          4633 => x"ff",
          4634 => x"93",
          4635 => x"38",
          4636 => x"ff",
          4637 => x"06",
          4638 => x"86",
          4639 => x"bb",
          4640 => x"8c",
          4641 => x"b0",
          4642 => x"84",
          4643 => x"3f",
          4644 => x"ec",
          4645 => x"bb",
          4646 => x"2b",
          4647 => x"51",
          4648 => x"2e",
          4649 => x"81",
          4650 => x"d3",
          4651 => x"98",
          4652 => x"2c",
          4653 => x"33",
          4654 => x"70",
          4655 => x"98",
          4656 => x"84",
          4657 => x"e8",
          4658 => x"15",
          4659 => x"51",
          4660 => x"59",
          4661 => x"58",
          4662 => x"78",
          4663 => x"38",
          4664 => x"b4",
          4665 => x"80",
          4666 => x"ff",
          4667 => x"98",
          4668 => x"80",
          4669 => x"ce",
          4670 => x"74",
          4671 => x"f6",
          4672 => x"bb",
          4673 => x"ff",
          4674 => x"80",
          4675 => x"74",
          4676 => x"34",
          4677 => x"39",
          4678 => x"0a",
          4679 => x"0a",
          4680 => x"2c",
          4681 => x"06",
          4682 => x"73",
          4683 => x"38",
          4684 => x"52",
          4685 => x"ce",
          4686 => x"dc",
          4687 => x"06",
          4688 => x"38",
          4689 => x"56",
          4690 => x"80",
          4691 => x"1c",
          4692 => x"d3",
          4693 => x"98",
          4694 => x"2c",
          4695 => x"33",
          4696 => x"70",
          4697 => x"10",
          4698 => x"2b",
          4699 => x"11",
          4700 => x"51",
          4701 => x"51",
          4702 => x"2e",
          4703 => x"fe",
          4704 => x"b0",
          4705 => x"7d",
          4706 => x"82",
          4707 => x"80",
          4708 => x"84",
          4709 => x"75",
          4710 => x"34",
          4711 => x"84",
          4712 => x"3d",
          4713 => x"0c",
          4714 => x"95",
          4715 => x"38",
          4716 => x"82",
          4717 => x"54",
          4718 => x"82",
          4719 => x"54",
          4720 => x"fd",
          4721 => x"d3",
          4722 => x"73",
          4723 => x"38",
          4724 => x"70",
          4725 => x"55",
          4726 => x"9e",
          4727 => x"54",
          4728 => x"15",
          4729 => x"80",
          4730 => x"ff",
          4731 => x"98",
          4732 => x"90",
          4733 => x"55",
          4734 => x"d3",
          4735 => x"11",
          4736 => x"82",
          4737 => x"73",
          4738 => x"3d",
          4739 => x"82",
          4740 => x"54",
          4741 => x"89",
          4742 => x"54",
          4743 => x"8c",
          4744 => x"90",
          4745 => x"80",
          4746 => x"ff",
          4747 => x"98",
          4748 => x"8c",
          4749 => x"56",
          4750 => x"25",
          4751 => x"d3",
          4752 => x"74",
          4753 => x"52",
          4754 => x"e8",
          4755 => x"80",
          4756 => x"80",
          4757 => x"98",
          4758 => x"8c",
          4759 => x"55",
          4760 => x"da",
          4761 => x"90",
          4762 => x"2b",
          4763 => x"82",
          4764 => x"5a",
          4765 => x"74",
          4766 => x"94",
          4767 => x"b0",
          4768 => x"51",
          4769 => x"3f",
          4770 => x"0a",
          4771 => x"0a",
          4772 => x"2c",
          4773 => x"33",
          4774 => x"73",
          4775 => x"38",
          4776 => x"83",
          4777 => x"0b",
          4778 => x"82",
          4779 => x"80",
          4780 => x"bc",
          4781 => x"3f",
          4782 => x"82",
          4783 => x"70",
          4784 => x"55",
          4785 => x"2e",
          4786 => x"82",
          4787 => x"ff",
          4788 => x"82",
          4789 => x"ff",
          4790 => x"82",
          4791 => x"82",
          4792 => x"52",
          4793 => x"9d",
          4794 => x"d3",
          4795 => x"98",
          4796 => x"2c",
          4797 => x"33",
          4798 => x"57",
          4799 => x"ad",
          4800 => x"54",
          4801 => x"74",
          4802 => x"b0",
          4803 => x"33",
          4804 => x"a0",
          4805 => x"80",
          4806 => x"80",
          4807 => x"98",
          4808 => x"8c",
          4809 => x"55",
          4810 => x"d5",
          4811 => x"b0",
          4812 => x"51",
          4813 => x"3f",
          4814 => x"33",
          4815 => x"70",
          4816 => x"d3",
          4817 => x"51",
          4818 => x"74",
          4819 => x"38",
          4820 => x"08",
          4821 => x"ff",
          4822 => x"74",
          4823 => x"29",
          4824 => x"05",
          4825 => x"82",
          4826 => x"58",
          4827 => x"75",
          4828 => x"fa",
          4829 => x"d3",
          4830 => x"05",
          4831 => x"34",
          4832 => x"08",
          4833 => x"ff",
          4834 => x"82",
          4835 => x"79",
          4836 => x"3f",
          4837 => x"08",
          4838 => x"54",
          4839 => x"82",
          4840 => x"54",
          4841 => x"8f",
          4842 => x"73",
          4843 => x"f1",
          4844 => x"39",
          4845 => x"80",
          4846 => x"90",
          4847 => x"82",
          4848 => x"79",
          4849 => x"0c",
          4850 => x"04",
          4851 => x"33",
          4852 => x"2e",
          4853 => x"82",
          4854 => x"52",
          4855 => x"9b",
          4856 => x"d3",
          4857 => x"05",
          4858 => x"d3",
          4859 => x"81",
          4860 => x"dd",
          4861 => x"90",
          4862 => x"8c",
          4863 => x"73",
          4864 => x"8c",
          4865 => x"54",
          4866 => x"8c",
          4867 => x"2b",
          4868 => x"75",
          4869 => x"56",
          4870 => x"74",
          4871 => x"74",
          4872 => x"14",
          4873 => x"82",
          4874 => x"52",
          4875 => x"ff",
          4876 => x"74",
          4877 => x"29",
          4878 => x"05",
          4879 => x"82",
          4880 => x"58",
          4881 => x"75",
          4882 => x"82",
          4883 => x"52",
          4884 => x"9a",
          4885 => x"d3",
          4886 => x"98",
          4887 => x"2c",
          4888 => x"33",
          4889 => x"57",
          4890 => x"f8",
          4891 => x"d3",
          4892 => x"88",
          4893 => x"bc",
          4894 => x"80",
          4895 => x"80",
          4896 => x"98",
          4897 => x"8c",
          4898 => x"55",
          4899 => x"de",
          4900 => x"39",
          4901 => x"33",
          4902 => x"06",
          4903 => x"33",
          4904 => x"74",
          4905 => x"e8",
          4906 => x"b0",
          4907 => x"14",
          4908 => x"d3",
          4909 => x"1a",
          4910 => x"54",
          4911 => x"3f",
          4912 => x"33",
          4913 => x"06",
          4914 => x"33",
          4915 => x"75",
          4916 => x"38",
          4917 => x"82",
          4918 => x"80",
          4919 => x"bc",
          4920 => x"3f",
          4921 => x"d3",
          4922 => x"0b",
          4923 => x"34",
          4924 => x"7a",
          4925 => x"bb",
          4926 => x"74",
          4927 => x"38",
          4928 => x"a2",
          4929 => x"bb",
          4930 => x"d3",
          4931 => x"bb",
          4932 => x"ff",
          4933 => x"53",
          4934 => x"51",
          4935 => x"3f",
          4936 => x"c0",
          4937 => x"29",
          4938 => x"05",
          4939 => x"56",
          4940 => x"2e",
          4941 => x"51",
          4942 => x"3f",
          4943 => x"08",
          4944 => x"34",
          4945 => x"08",
          4946 => x"81",
          4947 => x"52",
          4948 => x"a3",
          4949 => x"1b",
          4950 => x"39",
          4951 => x"74",
          4952 => x"ac",
          4953 => x"ff",
          4954 => x"99",
          4955 => x"2e",
          4956 => x"ae",
          4957 => x"dc",
          4958 => x"80",
          4959 => x"74",
          4960 => x"83",
          4961 => x"dc",
          4962 => x"8c",
          4963 => x"dc",
          4964 => x"06",
          4965 => x"74",
          4966 => x"ff",
          4967 => x"80",
          4968 => x"84",
          4969 => x"e0",
          4970 => x"56",
          4971 => x"2e",
          4972 => x"51",
          4973 => x"3f",
          4974 => x"08",
          4975 => x"34",
          4976 => x"08",
          4977 => x"81",
          4978 => x"52",
          4979 => x"a2",
          4980 => x"1b",
          4981 => x"ff",
          4982 => x"39",
          4983 => x"8c",
          4984 => x"34",
          4985 => x"53",
          4986 => x"33",
          4987 => x"ec",
          4988 => x"9c",
          4989 => x"90",
          4990 => x"ff",
          4991 => x"8c",
          4992 => x"54",
          4993 => x"f5",
          4994 => x"d3",
          4995 => x"81",
          4996 => x"82",
          4997 => x"74",
          4998 => x"52",
          4999 => x"94",
          5000 => x"39",
          5001 => x"33",
          5002 => x"2e",
          5003 => x"82",
          5004 => x"52",
          5005 => x"96",
          5006 => x"d3",
          5007 => x"05",
          5008 => x"d3",
          5009 => x"c8",
          5010 => x"0d",
          5011 => x"0b",
          5012 => x"0c",
          5013 => x"82",
          5014 => x"a0",
          5015 => x"52",
          5016 => x"51",
          5017 => x"3f",
          5018 => x"08",
          5019 => x"77",
          5020 => x"57",
          5021 => x"34",
          5022 => x"08",
          5023 => x"15",
          5024 => x"15",
          5025 => x"d4",
          5026 => x"86",
          5027 => x"87",
          5028 => x"bb",
          5029 => x"bb",
          5030 => x"05",
          5031 => x"07",
          5032 => x"ff",
          5033 => x"2a",
          5034 => x"56",
          5035 => x"34",
          5036 => x"34",
          5037 => x"22",
          5038 => x"82",
          5039 => x"05",
          5040 => x"55",
          5041 => x"15",
          5042 => x"15",
          5043 => x"0d",
          5044 => x"0d",
          5045 => x"51",
          5046 => x"8f",
          5047 => x"83",
          5048 => x"70",
          5049 => x"06",
          5050 => x"70",
          5051 => x"0c",
          5052 => x"04",
          5053 => x"02",
          5054 => x"02",
          5055 => x"05",
          5056 => x"82",
          5057 => x"71",
          5058 => x"11",
          5059 => x"73",
          5060 => x"81",
          5061 => x"88",
          5062 => x"a4",
          5063 => x"22",
          5064 => x"ff",
          5065 => x"88",
          5066 => x"52",
          5067 => x"5b",
          5068 => x"55",
          5069 => x"70",
          5070 => x"82",
          5071 => x"14",
          5072 => x"52",
          5073 => x"15",
          5074 => x"15",
          5075 => x"d4",
          5076 => x"70",
          5077 => x"33",
          5078 => x"07",
          5079 => x"8f",
          5080 => x"51",
          5081 => x"71",
          5082 => x"ff",
          5083 => x"88",
          5084 => x"51",
          5085 => x"34",
          5086 => x"06",
          5087 => x"12",
          5088 => x"d4",
          5089 => x"71",
          5090 => x"81",
          5091 => x"3d",
          5092 => x"3d",
          5093 => x"d4",
          5094 => x"05",
          5095 => x"70",
          5096 => x"11",
          5097 => x"87",
          5098 => x"8b",
          5099 => x"2b",
          5100 => x"59",
          5101 => x"72",
          5102 => x"33",
          5103 => x"71",
          5104 => x"70",
          5105 => x"56",
          5106 => x"84",
          5107 => x"85",
          5108 => x"bb",
          5109 => x"14",
          5110 => x"85",
          5111 => x"8b",
          5112 => x"2b",
          5113 => x"57",
          5114 => x"86",
          5115 => x"13",
          5116 => x"2b",
          5117 => x"2a",
          5118 => x"52",
          5119 => x"34",
          5120 => x"34",
          5121 => x"08",
          5122 => x"81",
          5123 => x"88",
          5124 => x"81",
          5125 => x"70",
          5126 => x"51",
          5127 => x"71",
          5128 => x"81",
          5129 => x"3d",
          5130 => x"3d",
          5131 => x"05",
          5132 => x"d4",
          5133 => x"2b",
          5134 => x"33",
          5135 => x"71",
          5136 => x"70",
          5137 => x"70",
          5138 => x"33",
          5139 => x"71",
          5140 => x"53",
          5141 => x"52",
          5142 => x"53",
          5143 => x"25",
          5144 => x"72",
          5145 => x"3f",
          5146 => x"08",
          5147 => x"33",
          5148 => x"71",
          5149 => x"83",
          5150 => x"11",
          5151 => x"12",
          5152 => x"2b",
          5153 => x"2b",
          5154 => x"06",
          5155 => x"51",
          5156 => x"53",
          5157 => x"88",
          5158 => x"72",
          5159 => x"73",
          5160 => x"82",
          5161 => x"70",
          5162 => x"81",
          5163 => x"8b",
          5164 => x"2b",
          5165 => x"57",
          5166 => x"70",
          5167 => x"33",
          5168 => x"07",
          5169 => x"ff",
          5170 => x"2a",
          5171 => x"58",
          5172 => x"34",
          5173 => x"34",
          5174 => x"04",
          5175 => x"82",
          5176 => x"02",
          5177 => x"05",
          5178 => x"2b",
          5179 => x"11",
          5180 => x"33",
          5181 => x"71",
          5182 => x"59",
          5183 => x"56",
          5184 => x"71",
          5185 => x"33",
          5186 => x"07",
          5187 => x"a2",
          5188 => x"07",
          5189 => x"53",
          5190 => x"53",
          5191 => x"70",
          5192 => x"82",
          5193 => x"70",
          5194 => x"81",
          5195 => x"8b",
          5196 => x"2b",
          5197 => x"57",
          5198 => x"82",
          5199 => x"13",
          5200 => x"2b",
          5201 => x"2a",
          5202 => x"52",
          5203 => x"34",
          5204 => x"34",
          5205 => x"08",
          5206 => x"33",
          5207 => x"71",
          5208 => x"82",
          5209 => x"52",
          5210 => x"0d",
          5211 => x"0d",
          5212 => x"d4",
          5213 => x"2a",
          5214 => x"ff",
          5215 => x"57",
          5216 => x"3f",
          5217 => x"08",
          5218 => x"71",
          5219 => x"33",
          5220 => x"71",
          5221 => x"83",
          5222 => x"11",
          5223 => x"12",
          5224 => x"2b",
          5225 => x"07",
          5226 => x"51",
          5227 => x"55",
          5228 => x"80",
          5229 => x"82",
          5230 => x"75",
          5231 => x"3f",
          5232 => x"84",
          5233 => x"15",
          5234 => x"2b",
          5235 => x"07",
          5236 => x"88",
          5237 => x"55",
          5238 => x"86",
          5239 => x"81",
          5240 => x"75",
          5241 => x"82",
          5242 => x"70",
          5243 => x"33",
          5244 => x"71",
          5245 => x"70",
          5246 => x"57",
          5247 => x"72",
          5248 => x"73",
          5249 => x"82",
          5250 => x"18",
          5251 => x"86",
          5252 => x"0b",
          5253 => x"82",
          5254 => x"53",
          5255 => x"34",
          5256 => x"34",
          5257 => x"08",
          5258 => x"81",
          5259 => x"88",
          5260 => x"82",
          5261 => x"70",
          5262 => x"51",
          5263 => x"74",
          5264 => x"81",
          5265 => x"3d",
          5266 => x"3d",
          5267 => x"82",
          5268 => x"84",
          5269 => x"3f",
          5270 => x"86",
          5271 => x"fe",
          5272 => x"3d",
          5273 => x"3d",
          5274 => x"52",
          5275 => x"3f",
          5276 => x"08",
          5277 => x"06",
          5278 => x"08",
          5279 => x"85",
          5280 => x"88",
          5281 => x"5f",
          5282 => x"5a",
          5283 => x"59",
          5284 => x"80",
          5285 => x"88",
          5286 => x"33",
          5287 => x"71",
          5288 => x"70",
          5289 => x"06",
          5290 => x"83",
          5291 => x"70",
          5292 => x"53",
          5293 => x"55",
          5294 => x"8a",
          5295 => x"2e",
          5296 => x"78",
          5297 => x"15",
          5298 => x"33",
          5299 => x"07",
          5300 => x"c2",
          5301 => x"ff",
          5302 => x"38",
          5303 => x"56",
          5304 => x"2b",
          5305 => x"08",
          5306 => x"81",
          5307 => x"88",
          5308 => x"81",
          5309 => x"51",
          5310 => x"5c",
          5311 => x"2e",
          5312 => x"55",
          5313 => x"78",
          5314 => x"38",
          5315 => x"80",
          5316 => x"38",
          5317 => x"09",
          5318 => x"38",
          5319 => x"f2",
          5320 => x"39",
          5321 => x"53",
          5322 => x"51",
          5323 => x"82",
          5324 => x"70",
          5325 => x"33",
          5326 => x"71",
          5327 => x"83",
          5328 => x"5a",
          5329 => x"05",
          5330 => x"83",
          5331 => x"70",
          5332 => x"59",
          5333 => x"84",
          5334 => x"81",
          5335 => x"76",
          5336 => x"82",
          5337 => x"75",
          5338 => x"11",
          5339 => x"11",
          5340 => x"33",
          5341 => x"07",
          5342 => x"53",
          5343 => x"5a",
          5344 => x"86",
          5345 => x"87",
          5346 => x"bb",
          5347 => x"1c",
          5348 => x"85",
          5349 => x"8b",
          5350 => x"2b",
          5351 => x"5a",
          5352 => x"54",
          5353 => x"34",
          5354 => x"34",
          5355 => x"08",
          5356 => x"1d",
          5357 => x"85",
          5358 => x"88",
          5359 => x"88",
          5360 => x"5f",
          5361 => x"73",
          5362 => x"75",
          5363 => x"82",
          5364 => x"1b",
          5365 => x"73",
          5366 => x"0c",
          5367 => x"04",
          5368 => x"74",
          5369 => x"d4",
          5370 => x"f4",
          5371 => x"53",
          5372 => x"8b",
          5373 => x"fc",
          5374 => x"bb",
          5375 => x"72",
          5376 => x"0c",
          5377 => x"04",
          5378 => x"64",
          5379 => x"80",
          5380 => x"82",
          5381 => x"60",
          5382 => x"06",
          5383 => x"a9",
          5384 => x"38",
          5385 => x"b8",
          5386 => x"dc",
          5387 => x"c7",
          5388 => x"38",
          5389 => x"92",
          5390 => x"83",
          5391 => x"51",
          5392 => x"82",
          5393 => x"83",
          5394 => x"82",
          5395 => x"7d",
          5396 => x"2a",
          5397 => x"ff",
          5398 => x"2b",
          5399 => x"33",
          5400 => x"71",
          5401 => x"70",
          5402 => x"83",
          5403 => x"70",
          5404 => x"05",
          5405 => x"1a",
          5406 => x"12",
          5407 => x"2b",
          5408 => x"2b",
          5409 => x"53",
          5410 => x"5c",
          5411 => x"5c",
          5412 => x"73",
          5413 => x"38",
          5414 => x"ff",
          5415 => x"70",
          5416 => x"06",
          5417 => x"16",
          5418 => x"33",
          5419 => x"07",
          5420 => x"1c",
          5421 => x"12",
          5422 => x"2b",
          5423 => x"07",
          5424 => x"52",
          5425 => x"80",
          5426 => x"78",
          5427 => x"83",
          5428 => x"41",
          5429 => x"27",
          5430 => x"60",
          5431 => x"7b",
          5432 => x"06",
          5433 => x"51",
          5434 => x"7a",
          5435 => x"06",
          5436 => x"39",
          5437 => x"7a",
          5438 => x"38",
          5439 => x"aa",
          5440 => x"39",
          5441 => x"7a",
          5442 => x"c8",
          5443 => x"82",
          5444 => x"12",
          5445 => x"2b",
          5446 => x"54",
          5447 => x"80",
          5448 => x"f7",
          5449 => x"bb",
          5450 => x"ff",
          5451 => x"54",
          5452 => x"83",
          5453 => x"d4",
          5454 => x"05",
          5455 => x"ff",
          5456 => x"82",
          5457 => x"14",
          5458 => x"83",
          5459 => x"59",
          5460 => x"39",
          5461 => x"7a",
          5462 => x"d4",
          5463 => x"f5",
          5464 => x"bb",
          5465 => x"82",
          5466 => x"12",
          5467 => x"2b",
          5468 => x"54",
          5469 => x"80",
          5470 => x"f6",
          5471 => x"bb",
          5472 => x"ff",
          5473 => x"54",
          5474 => x"83",
          5475 => x"d4",
          5476 => x"05",
          5477 => x"ff",
          5478 => x"82",
          5479 => x"14",
          5480 => x"62",
          5481 => x"5c",
          5482 => x"ff",
          5483 => x"39",
          5484 => x"54",
          5485 => x"82",
          5486 => x"5c",
          5487 => x"08",
          5488 => x"38",
          5489 => x"52",
          5490 => x"08",
          5491 => x"97",
          5492 => x"f7",
          5493 => x"58",
          5494 => x"99",
          5495 => x"7a",
          5496 => x"f2",
          5497 => x"19",
          5498 => x"bb",
          5499 => x"84",
          5500 => x"f9",
          5501 => x"73",
          5502 => x"0c",
          5503 => x"04",
          5504 => x"77",
          5505 => x"52",
          5506 => x"3f",
          5507 => x"08",
          5508 => x"dc",
          5509 => x"8e",
          5510 => x"80",
          5511 => x"dc",
          5512 => x"96",
          5513 => x"82",
          5514 => x"86",
          5515 => x"ff",
          5516 => x"8f",
          5517 => x"81",
          5518 => x"26",
          5519 => x"bb",
          5520 => x"52",
          5521 => x"dc",
          5522 => x"0d",
          5523 => x"0d",
          5524 => x"33",
          5525 => x"9f",
          5526 => x"53",
          5527 => x"81",
          5528 => x"38",
          5529 => x"87",
          5530 => x"11",
          5531 => x"54",
          5532 => x"84",
          5533 => x"54",
          5534 => x"87",
          5535 => x"11",
          5536 => x"0c",
          5537 => x"c0",
          5538 => x"70",
          5539 => x"70",
          5540 => x"51",
          5541 => x"8a",
          5542 => x"98",
          5543 => x"70",
          5544 => x"08",
          5545 => x"06",
          5546 => x"38",
          5547 => x"8c",
          5548 => x"80",
          5549 => x"71",
          5550 => x"14",
          5551 => x"d8",
          5552 => x"70",
          5553 => x"0c",
          5554 => x"04",
          5555 => x"60",
          5556 => x"8c",
          5557 => x"33",
          5558 => x"5b",
          5559 => x"5a",
          5560 => x"82",
          5561 => x"81",
          5562 => x"52",
          5563 => x"38",
          5564 => x"84",
          5565 => x"92",
          5566 => x"c0",
          5567 => x"87",
          5568 => x"13",
          5569 => x"57",
          5570 => x"0b",
          5571 => x"8c",
          5572 => x"0c",
          5573 => x"75",
          5574 => x"2a",
          5575 => x"51",
          5576 => x"80",
          5577 => x"7b",
          5578 => x"7b",
          5579 => x"5d",
          5580 => x"59",
          5581 => x"06",
          5582 => x"73",
          5583 => x"81",
          5584 => x"ff",
          5585 => x"72",
          5586 => x"38",
          5587 => x"8c",
          5588 => x"c3",
          5589 => x"98",
          5590 => x"71",
          5591 => x"38",
          5592 => x"2e",
          5593 => x"76",
          5594 => x"92",
          5595 => x"72",
          5596 => x"06",
          5597 => x"f7",
          5598 => x"5a",
          5599 => x"80",
          5600 => x"70",
          5601 => x"5a",
          5602 => x"80",
          5603 => x"73",
          5604 => x"06",
          5605 => x"38",
          5606 => x"fe",
          5607 => x"fc",
          5608 => x"52",
          5609 => x"83",
          5610 => x"71",
          5611 => x"bb",
          5612 => x"3d",
          5613 => x"3d",
          5614 => x"64",
          5615 => x"bf",
          5616 => x"40",
          5617 => x"59",
          5618 => x"58",
          5619 => x"82",
          5620 => x"81",
          5621 => x"52",
          5622 => x"09",
          5623 => x"b1",
          5624 => x"84",
          5625 => x"92",
          5626 => x"c0",
          5627 => x"87",
          5628 => x"13",
          5629 => x"56",
          5630 => x"87",
          5631 => x"0c",
          5632 => x"82",
          5633 => x"58",
          5634 => x"84",
          5635 => x"06",
          5636 => x"71",
          5637 => x"38",
          5638 => x"05",
          5639 => x"0c",
          5640 => x"73",
          5641 => x"81",
          5642 => x"71",
          5643 => x"38",
          5644 => x"8c",
          5645 => x"d0",
          5646 => x"98",
          5647 => x"71",
          5648 => x"38",
          5649 => x"2e",
          5650 => x"76",
          5651 => x"92",
          5652 => x"72",
          5653 => x"06",
          5654 => x"f7",
          5655 => x"59",
          5656 => x"1a",
          5657 => x"06",
          5658 => x"59",
          5659 => x"80",
          5660 => x"73",
          5661 => x"06",
          5662 => x"38",
          5663 => x"fe",
          5664 => x"fc",
          5665 => x"52",
          5666 => x"83",
          5667 => x"71",
          5668 => x"bb",
          5669 => x"3d",
          5670 => x"3d",
          5671 => x"84",
          5672 => x"33",
          5673 => x"a7",
          5674 => x"54",
          5675 => x"fa",
          5676 => x"bb",
          5677 => x"06",
          5678 => x"72",
          5679 => x"85",
          5680 => x"98",
          5681 => x"56",
          5682 => x"80",
          5683 => x"76",
          5684 => x"74",
          5685 => x"c0",
          5686 => x"54",
          5687 => x"2e",
          5688 => x"d4",
          5689 => x"2e",
          5690 => x"80",
          5691 => x"08",
          5692 => x"70",
          5693 => x"51",
          5694 => x"2e",
          5695 => x"c0",
          5696 => x"52",
          5697 => x"87",
          5698 => x"08",
          5699 => x"38",
          5700 => x"87",
          5701 => x"14",
          5702 => x"70",
          5703 => x"52",
          5704 => x"96",
          5705 => x"92",
          5706 => x"0a",
          5707 => x"39",
          5708 => x"0c",
          5709 => x"39",
          5710 => x"54",
          5711 => x"dc",
          5712 => x"0d",
          5713 => x"0d",
          5714 => x"33",
          5715 => x"88",
          5716 => x"bb",
          5717 => x"51",
          5718 => x"04",
          5719 => x"75",
          5720 => x"82",
          5721 => x"90",
          5722 => x"2b",
          5723 => x"33",
          5724 => x"88",
          5725 => x"71",
          5726 => x"dc",
          5727 => x"54",
          5728 => x"85",
          5729 => x"ff",
          5730 => x"02",
          5731 => x"05",
          5732 => x"70",
          5733 => x"05",
          5734 => x"88",
          5735 => x"72",
          5736 => x"0d",
          5737 => x"0d",
          5738 => x"52",
          5739 => x"81",
          5740 => x"70",
          5741 => x"70",
          5742 => x"05",
          5743 => x"88",
          5744 => x"72",
          5745 => x"54",
          5746 => x"2a",
          5747 => x"34",
          5748 => x"04",
          5749 => x"76",
          5750 => x"54",
          5751 => x"2e",
          5752 => x"70",
          5753 => x"33",
          5754 => x"05",
          5755 => x"11",
          5756 => x"84",
          5757 => x"fe",
          5758 => x"77",
          5759 => x"53",
          5760 => x"81",
          5761 => x"ff",
          5762 => x"f4",
          5763 => x"0d",
          5764 => x"0d",
          5765 => x"56",
          5766 => x"70",
          5767 => x"33",
          5768 => x"05",
          5769 => x"71",
          5770 => x"56",
          5771 => x"72",
          5772 => x"38",
          5773 => x"e2",
          5774 => x"bb",
          5775 => x"3d",
          5776 => x"3d",
          5777 => x"54",
          5778 => x"71",
          5779 => x"38",
          5780 => x"70",
          5781 => x"f3",
          5782 => x"82",
          5783 => x"84",
          5784 => x"80",
          5785 => x"dc",
          5786 => x"0b",
          5787 => x"0c",
          5788 => x"0d",
          5789 => x"0b",
          5790 => x"56",
          5791 => x"2e",
          5792 => x"81",
          5793 => x"08",
          5794 => x"70",
          5795 => x"33",
          5796 => x"a2",
          5797 => x"dc",
          5798 => x"09",
          5799 => x"38",
          5800 => x"08",
          5801 => x"b0",
          5802 => x"a4",
          5803 => x"9c",
          5804 => x"56",
          5805 => x"27",
          5806 => x"16",
          5807 => x"82",
          5808 => x"06",
          5809 => x"54",
          5810 => x"78",
          5811 => x"33",
          5812 => x"3f",
          5813 => x"5a",
          5814 => x"dc",
          5815 => x"0d",
          5816 => x"0d",
          5817 => x"56",
          5818 => x"b0",
          5819 => x"af",
          5820 => x"fe",
          5821 => x"bb",
          5822 => x"82",
          5823 => x"9f",
          5824 => x"74",
          5825 => x"52",
          5826 => x"51",
          5827 => x"82",
          5828 => x"80",
          5829 => x"ff",
          5830 => x"74",
          5831 => x"76",
          5832 => x"0c",
          5833 => x"04",
          5834 => x"7a",
          5835 => x"fe",
          5836 => x"bb",
          5837 => x"82",
          5838 => x"81",
          5839 => x"33",
          5840 => x"2e",
          5841 => x"80",
          5842 => x"17",
          5843 => x"81",
          5844 => x"06",
          5845 => x"84",
          5846 => x"bb",
          5847 => x"b4",
          5848 => x"56",
          5849 => x"82",
          5850 => x"84",
          5851 => x"fc",
          5852 => x"8b",
          5853 => x"52",
          5854 => x"a9",
          5855 => x"85",
          5856 => x"84",
          5857 => x"fc",
          5858 => x"17",
          5859 => x"9c",
          5860 => x"91",
          5861 => x"08",
          5862 => x"17",
          5863 => x"3f",
          5864 => x"81",
          5865 => x"19",
          5866 => x"53",
          5867 => x"17",
          5868 => x"82",
          5869 => x"18",
          5870 => x"80",
          5871 => x"33",
          5872 => x"3f",
          5873 => x"08",
          5874 => x"38",
          5875 => x"82",
          5876 => x"8a",
          5877 => x"fb",
          5878 => x"fe",
          5879 => x"08",
          5880 => x"56",
          5881 => x"74",
          5882 => x"38",
          5883 => x"75",
          5884 => x"16",
          5885 => x"53",
          5886 => x"dc",
          5887 => x"0d",
          5888 => x"0d",
          5889 => x"08",
          5890 => x"81",
          5891 => x"df",
          5892 => x"15",
          5893 => x"d7",
          5894 => x"33",
          5895 => x"82",
          5896 => x"38",
          5897 => x"89",
          5898 => x"2e",
          5899 => x"bf",
          5900 => x"2e",
          5901 => x"81",
          5902 => x"81",
          5903 => x"89",
          5904 => x"08",
          5905 => x"52",
          5906 => x"3f",
          5907 => x"08",
          5908 => x"74",
          5909 => x"14",
          5910 => x"81",
          5911 => x"2a",
          5912 => x"05",
          5913 => x"57",
          5914 => x"f5",
          5915 => x"dc",
          5916 => x"38",
          5917 => x"06",
          5918 => x"33",
          5919 => x"78",
          5920 => x"06",
          5921 => x"5c",
          5922 => x"53",
          5923 => x"38",
          5924 => x"06",
          5925 => x"39",
          5926 => x"a4",
          5927 => x"52",
          5928 => x"bd",
          5929 => x"dc",
          5930 => x"38",
          5931 => x"fe",
          5932 => x"b4",
          5933 => x"8d",
          5934 => x"dc",
          5935 => x"ff",
          5936 => x"39",
          5937 => x"a4",
          5938 => x"52",
          5939 => x"91",
          5940 => x"dc",
          5941 => x"76",
          5942 => x"fc",
          5943 => x"b4",
          5944 => x"f8",
          5945 => x"dc",
          5946 => x"06",
          5947 => x"81",
          5948 => x"bb",
          5949 => x"3d",
          5950 => x"3d",
          5951 => x"7e",
          5952 => x"82",
          5953 => x"27",
          5954 => x"76",
          5955 => x"27",
          5956 => x"75",
          5957 => x"79",
          5958 => x"38",
          5959 => x"89",
          5960 => x"2e",
          5961 => x"80",
          5962 => x"2e",
          5963 => x"81",
          5964 => x"81",
          5965 => x"89",
          5966 => x"08",
          5967 => x"52",
          5968 => x"3f",
          5969 => x"08",
          5970 => x"dc",
          5971 => x"38",
          5972 => x"06",
          5973 => x"81",
          5974 => x"06",
          5975 => x"77",
          5976 => x"2e",
          5977 => x"84",
          5978 => x"06",
          5979 => x"06",
          5980 => x"53",
          5981 => x"81",
          5982 => x"34",
          5983 => x"a4",
          5984 => x"52",
          5985 => x"d9",
          5986 => x"dc",
          5987 => x"bb",
          5988 => x"94",
          5989 => x"ff",
          5990 => x"05",
          5991 => x"54",
          5992 => x"38",
          5993 => x"74",
          5994 => x"06",
          5995 => x"07",
          5996 => x"74",
          5997 => x"39",
          5998 => x"a4",
          5999 => x"52",
          6000 => x"9d",
          6001 => x"dc",
          6002 => x"bb",
          6003 => x"d8",
          6004 => x"ff",
          6005 => x"76",
          6006 => x"06",
          6007 => x"05",
          6008 => x"3f",
          6009 => x"87",
          6010 => x"08",
          6011 => x"51",
          6012 => x"82",
          6013 => x"59",
          6014 => x"08",
          6015 => x"f0",
          6016 => x"82",
          6017 => x"06",
          6018 => x"05",
          6019 => x"54",
          6020 => x"3f",
          6021 => x"08",
          6022 => x"74",
          6023 => x"51",
          6024 => x"81",
          6025 => x"34",
          6026 => x"dc",
          6027 => x"0d",
          6028 => x"0d",
          6029 => x"72",
          6030 => x"56",
          6031 => x"27",
          6032 => x"98",
          6033 => x"9d",
          6034 => x"2e",
          6035 => x"53",
          6036 => x"51",
          6037 => x"82",
          6038 => x"54",
          6039 => x"08",
          6040 => x"93",
          6041 => x"80",
          6042 => x"54",
          6043 => x"82",
          6044 => x"54",
          6045 => x"74",
          6046 => x"fb",
          6047 => x"bb",
          6048 => x"82",
          6049 => x"80",
          6050 => x"38",
          6051 => x"08",
          6052 => x"38",
          6053 => x"08",
          6054 => x"38",
          6055 => x"52",
          6056 => x"d6",
          6057 => x"dc",
          6058 => x"98",
          6059 => x"11",
          6060 => x"57",
          6061 => x"74",
          6062 => x"81",
          6063 => x"0c",
          6064 => x"81",
          6065 => x"84",
          6066 => x"55",
          6067 => x"ff",
          6068 => x"54",
          6069 => x"dc",
          6070 => x"0d",
          6071 => x"0d",
          6072 => x"08",
          6073 => x"79",
          6074 => x"17",
          6075 => x"80",
          6076 => x"98",
          6077 => x"26",
          6078 => x"58",
          6079 => x"52",
          6080 => x"fd",
          6081 => x"74",
          6082 => x"08",
          6083 => x"38",
          6084 => x"08",
          6085 => x"dc",
          6086 => x"82",
          6087 => x"17",
          6088 => x"dc",
          6089 => x"c7",
          6090 => x"90",
          6091 => x"56",
          6092 => x"2e",
          6093 => x"77",
          6094 => x"81",
          6095 => x"38",
          6096 => x"98",
          6097 => x"26",
          6098 => x"56",
          6099 => x"51",
          6100 => x"80",
          6101 => x"dc",
          6102 => x"09",
          6103 => x"38",
          6104 => x"08",
          6105 => x"dc",
          6106 => x"30",
          6107 => x"80",
          6108 => x"07",
          6109 => x"08",
          6110 => x"55",
          6111 => x"ef",
          6112 => x"dc",
          6113 => x"95",
          6114 => x"08",
          6115 => x"27",
          6116 => x"98",
          6117 => x"89",
          6118 => x"85",
          6119 => x"db",
          6120 => x"81",
          6121 => x"17",
          6122 => x"89",
          6123 => x"75",
          6124 => x"ac",
          6125 => x"7a",
          6126 => x"3f",
          6127 => x"08",
          6128 => x"38",
          6129 => x"bb",
          6130 => x"2e",
          6131 => x"86",
          6132 => x"dc",
          6133 => x"bb",
          6134 => x"70",
          6135 => x"07",
          6136 => x"7c",
          6137 => x"55",
          6138 => x"f8",
          6139 => x"2e",
          6140 => x"ff",
          6141 => x"55",
          6142 => x"ff",
          6143 => x"76",
          6144 => x"3f",
          6145 => x"08",
          6146 => x"08",
          6147 => x"bb",
          6148 => x"80",
          6149 => x"55",
          6150 => x"94",
          6151 => x"2e",
          6152 => x"53",
          6153 => x"51",
          6154 => x"82",
          6155 => x"55",
          6156 => x"75",
          6157 => x"98",
          6158 => x"05",
          6159 => x"56",
          6160 => x"26",
          6161 => x"15",
          6162 => x"84",
          6163 => x"07",
          6164 => x"18",
          6165 => x"ff",
          6166 => x"2e",
          6167 => x"39",
          6168 => x"39",
          6169 => x"08",
          6170 => x"81",
          6171 => x"74",
          6172 => x"0c",
          6173 => x"04",
          6174 => x"7a",
          6175 => x"f3",
          6176 => x"bb",
          6177 => x"81",
          6178 => x"dc",
          6179 => x"38",
          6180 => x"51",
          6181 => x"82",
          6182 => x"82",
          6183 => x"b0",
          6184 => x"84",
          6185 => x"52",
          6186 => x"52",
          6187 => x"3f",
          6188 => x"39",
          6189 => x"8a",
          6190 => x"75",
          6191 => x"38",
          6192 => x"19",
          6193 => x"81",
          6194 => x"ed",
          6195 => x"bb",
          6196 => x"2e",
          6197 => x"15",
          6198 => x"70",
          6199 => x"07",
          6200 => x"53",
          6201 => x"75",
          6202 => x"0c",
          6203 => x"04",
          6204 => x"7a",
          6205 => x"58",
          6206 => x"f0",
          6207 => x"80",
          6208 => x"9f",
          6209 => x"80",
          6210 => x"90",
          6211 => x"17",
          6212 => x"aa",
          6213 => x"53",
          6214 => x"88",
          6215 => x"08",
          6216 => x"38",
          6217 => x"53",
          6218 => x"17",
          6219 => x"72",
          6220 => x"fe",
          6221 => x"08",
          6222 => x"80",
          6223 => x"16",
          6224 => x"2b",
          6225 => x"75",
          6226 => x"73",
          6227 => x"f5",
          6228 => x"bb",
          6229 => x"82",
          6230 => x"ff",
          6231 => x"81",
          6232 => x"dc",
          6233 => x"38",
          6234 => x"82",
          6235 => x"26",
          6236 => x"58",
          6237 => x"73",
          6238 => x"39",
          6239 => x"51",
          6240 => x"82",
          6241 => x"98",
          6242 => x"94",
          6243 => x"17",
          6244 => x"58",
          6245 => x"9a",
          6246 => x"81",
          6247 => x"74",
          6248 => x"98",
          6249 => x"83",
          6250 => x"b4",
          6251 => x"0c",
          6252 => x"82",
          6253 => x"8a",
          6254 => x"f8",
          6255 => x"70",
          6256 => x"08",
          6257 => x"57",
          6258 => x"0a",
          6259 => x"38",
          6260 => x"15",
          6261 => x"08",
          6262 => x"72",
          6263 => x"cb",
          6264 => x"ff",
          6265 => x"81",
          6266 => x"13",
          6267 => x"94",
          6268 => x"74",
          6269 => x"85",
          6270 => x"22",
          6271 => x"73",
          6272 => x"38",
          6273 => x"8a",
          6274 => x"05",
          6275 => x"06",
          6276 => x"8a",
          6277 => x"73",
          6278 => x"3f",
          6279 => x"08",
          6280 => x"81",
          6281 => x"dc",
          6282 => x"ff",
          6283 => x"82",
          6284 => x"ff",
          6285 => x"38",
          6286 => x"82",
          6287 => x"26",
          6288 => x"7b",
          6289 => x"98",
          6290 => x"55",
          6291 => x"94",
          6292 => x"73",
          6293 => x"3f",
          6294 => x"08",
          6295 => x"82",
          6296 => x"80",
          6297 => x"38",
          6298 => x"bb",
          6299 => x"2e",
          6300 => x"55",
          6301 => x"08",
          6302 => x"38",
          6303 => x"08",
          6304 => x"fb",
          6305 => x"bb",
          6306 => x"38",
          6307 => x"0c",
          6308 => x"51",
          6309 => x"82",
          6310 => x"98",
          6311 => x"90",
          6312 => x"16",
          6313 => x"15",
          6314 => x"74",
          6315 => x"0c",
          6316 => x"04",
          6317 => x"7b",
          6318 => x"5b",
          6319 => x"52",
          6320 => x"ac",
          6321 => x"dc",
          6322 => x"bb",
          6323 => x"ec",
          6324 => x"dc",
          6325 => x"17",
          6326 => x"51",
          6327 => x"82",
          6328 => x"54",
          6329 => x"08",
          6330 => x"82",
          6331 => x"9c",
          6332 => x"33",
          6333 => x"72",
          6334 => x"09",
          6335 => x"38",
          6336 => x"bb",
          6337 => x"72",
          6338 => x"55",
          6339 => x"53",
          6340 => x"8e",
          6341 => x"56",
          6342 => x"09",
          6343 => x"38",
          6344 => x"bb",
          6345 => x"81",
          6346 => x"fd",
          6347 => x"bb",
          6348 => x"82",
          6349 => x"80",
          6350 => x"38",
          6351 => x"09",
          6352 => x"38",
          6353 => x"82",
          6354 => x"8b",
          6355 => x"fd",
          6356 => x"9a",
          6357 => x"eb",
          6358 => x"bb",
          6359 => x"ff",
          6360 => x"70",
          6361 => x"53",
          6362 => x"09",
          6363 => x"38",
          6364 => x"eb",
          6365 => x"bb",
          6366 => x"2b",
          6367 => x"72",
          6368 => x"0c",
          6369 => x"04",
          6370 => x"77",
          6371 => x"ff",
          6372 => x"9a",
          6373 => x"55",
          6374 => x"76",
          6375 => x"53",
          6376 => x"09",
          6377 => x"38",
          6378 => x"52",
          6379 => x"eb",
          6380 => x"3d",
          6381 => x"3d",
          6382 => x"5b",
          6383 => x"08",
          6384 => x"15",
          6385 => x"81",
          6386 => x"15",
          6387 => x"51",
          6388 => x"82",
          6389 => x"58",
          6390 => x"08",
          6391 => x"9c",
          6392 => x"33",
          6393 => x"86",
          6394 => x"80",
          6395 => x"13",
          6396 => x"06",
          6397 => x"06",
          6398 => x"72",
          6399 => x"82",
          6400 => x"53",
          6401 => x"2e",
          6402 => x"53",
          6403 => x"a9",
          6404 => x"74",
          6405 => x"72",
          6406 => x"38",
          6407 => x"99",
          6408 => x"dc",
          6409 => x"06",
          6410 => x"88",
          6411 => x"06",
          6412 => x"54",
          6413 => x"a0",
          6414 => x"74",
          6415 => x"3f",
          6416 => x"08",
          6417 => x"dc",
          6418 => x"98",
          6419 => x"fa",
          6420 => x"80",
          6421 => x"0c",
          6422 => x"dc",
          6423 => x"0d",
          6424 => x"0d",
          6425 => x"57",
          6426 => x"73",
          6427 => x"3f",
          6428 => x"08",
          6429 => x"dc",
          6430 => x"98",
          6431 => x"75",
          6432 => x"3f",
          6433 => x"08",
          6434 => x"dc",
          6435 => x"a0",
          6436 => x"dc",
          6437 => x"14",
          6438 => x"db",
          6439 => x"a0",
          6440 => x"14",
          6441 => x"ac",
          6442 => x"83",
          6443 => x"82",
          6444 => x"87",
          6445 => x"fd",
          6446 => x"70",
          6447 => x"08",
          6448 => x"55",
          6449 => x"3f",
          6450 => x"08",
          6451 => x"13",
          6452 => x"73",
          6453 => x"83",
          6454 => x"3d",
          6455 => x"3d",
          6456 => x"57",
          6457 => x"89",
          6458 => x"17",
          6459 => x"81",
          6460 => x"70",
          6461 => x"55",
          6462 => x"08",
          6463 => x"81",
          6464 => x"52",
          6465 => x"a8",
          6466 => x"2e",
          6467 => x"84",
          6468 => x"52",
          6469 => x"09",
          6470 => x"38",
          6471 => x"81",
          6472 => x"81",
          6473 => x"73",
          6474 => x"55",
          6475 => x"55",
          6476 => x"c5",
          6477 => x"88",
          6478 => x"0b",
          6479 => x"9c",
          6480 => x"8b",
          6481 => x"17",
          6482 => x"08",
          6483 => x"52",
          6484 => x"82",
          6485 => x"76",
          6486 => x"51",
          6487 => x"82",
          6488 => x"86",
          6489 => x"12",
          6490 => x"3f",
          6491 => x"08",
          6492 => x"88",
          6493 => x"f3",
          6494 => x"70",
          6495 => x"80",
          6496 => x"51",
          6497 => x"af",
          6498 => x"81",
          6499 => x"dc",
          6500 => x"74",
          6501 => x"38",
          6502 => x"88",
          6503 => x"39",
          6504 => x"80",
          6505 => x"56",
          6506 => x"af",
          6507 => x"06",
          6508 => x"56",
          6509 => x"32",
          6510 => x"80",
          6511 => x"51",
          6512 => x"dc",
          6513 => x"1c",
          6514 => x"33",
          6515 => x"9f",
          6516 => x"ff",
          6517 => x"1c",
          6518 => x"7a",
          6519 => x"3f",
          6520 => x"08",
          6521 => x"39",
          6522 => x"a0",
          6523 => x"5e",
          6524 => x"52",
          6525 => x"ff",
          6526 => x"59",
          6527 => x"33",
          6528 => x"ae",
          6529 => x"06",
          6530 => x"78",
          6531 => x"81",
          6532 => x"32",
          6533 => x"9f",
          6534 => x"26",
          6535 => x"53",
          6536 => x"73",
          6537 => x"17",
          6538 => x"34",
          6539 => x"db",
          6540 => x"32",
          6541 => x"9f",
          6542 => x"54",
          6543 => x"2e",
          6544 => x"80",
          6545 => x"75",
          6546 => x"bd",
          6547 => x"7e",
          6548 => x"a0",
          6549 => x"bd",
          6550 => x"82",
          6551 => x"18",
          6552 => x"1a",
          6553 => x"a0",
          6554 => x"fc",
          6555 => x"32",
          6556 => x"80",
          6557 => x"30",
          6558 => x"71",
          6559 => x"51",
          6560 => x"55",
          6561 => x"ac",
          6562 => x"81",
          6563 => x"78",
          6564 => x"51",
          6565 => x"af",
          6566 => x"06",
          6567 => x"55",
          6568 => x"32",
          6569 => x"80",
          6570 => x"51",
          6571 => x"db",
          6572 => x"39",
          6573 => x"09",
          6574 => x"38",
          6575 => x"7c",
          6576 => x"54",
          6577 => x"a2",
          6578 => x"32",
          6579 => x"ae",
          6580 => x"72",
          6581 => x"9f",
          6582 => x"51",
          6583 => x"74",
          6584 => x"88",
          6585 => x"fe",
          6586 => x"98",
          6587 => x"80",
          6588 => x"75",
          6589 => x"82",
          6590 => x"33",
          6591 => x"51",
          6592 => x"82",
          6593 => x"80",
          6594 => x"78",
          6595 => x"81",
          6596 => x"5a",
          6597 => x"d2",
          6598 => x"dc",
          6599 => x"80",
          6600 => x"1c",
          6601 => x"27",
          6602 => x"79",
          6603 => x"74",
          6604 => x"7a",
          6605 => x"74",
          6606 => x"39",
          6607 => x"b4",
          6608 => x"fe",
          6609 => x"dc",
          6610 => x"ff",
          6611 => x"73",
          6612 => x"38",
          6613 => x"81",
          6614 => x"54",
          6615 => x"75",
          6616 => x"17",
          6617 => x"39",
          6618 => x"0c",
          6619 => x"99",
          6620 => x"54",
          6621 => x"2e",
          6622 => x"84",
          6623 => x"34",
          6624 => x"76",
          6625 => x"8b",
          6626 => x"81",
          6627 => x"56",
          6628 => x"80",
          6629 => x"1b",
          6630 => x"08",
          6631 => x"51",
          6632 => x"82",
          6633 => x"56",
          6634 => x"08",
          6635 => x"98",
          6636 => x"76",
          6637 => x"3f",
          6638 => x"08",
          6639 => x"dc",
          6640 => x"38",
          6641 => x"70",
          6642 => x"73",
          6643 => x"be",
          6644 => x"33",
          6645 => x"73",
          6646 => x"8b",
          6647 => x"83",
          6648 => x"06",
          6649 => x"73",
          6650 => x"53",
          6651 => x"51",
          6652 => x"82",
          6653 => x"80",
          6654 => x"75",
          6655 => x"f3",
          6656 => x"9f",
          6657 => x"1c",
          6658 => x"74",
          6659 => x"38",
          6660 => x"09",
          6661 => x"e7",
          6662 => x"2a",
          6663 => x"77",
          6664 => x"51",
          6665 => x"2e",
          6666 => x"81",
          6667 => x"80",
          6668 => x"38",
          6669 => x"ab",
          6670 => x"55",
          6671 => x"75",
          6672 => x"73",
          6673 => x"55",
          6674 => x"82",
          6675 => x"06",
          6676 => x"ab",
          6677 => x"33",
          6678 => x"70",
          6679 => x"55",
          6680 => x"2e",
          6681 => x"1b",
          6682 => x"06",
          6683 => x"52",
          6684 => x"db",
          6685 => x"dc",
          6686 => x"0c",
          6687 => x"74",
          6688 => x"0c",
          6689 => x"04",
          6690 => x"7c",
          6691 => x"08",
          6692 => x"55",
          6693 => x"59",
          6694 => x"81",
          6695 => x"70",
          6696 => x"33",
          6697 => x"52",
          6698 => x"2e",
          6699 => x"ee",
          6700 => x"2e",
          6701 => x"81",
          6702 => x"33",
          6703 => x"81",
          6704 => x"52",
          6705 => x"26",
          6706 => x"14",
          6707 => x"06",
          6708 => x"52",
          6709 => x"80",
          6710 => x"0b",
          6711 => x"59",
          6712 => x"7a",
          6713 => x"70",
          6714 => x"33",
          6715 => x"05",
          6716 => x"9f",
          6717 => x"53",
          6718 => x"89",
          6719 => x"70",
          6720 => x"54",
          6721 => x"12",
          6722 => x"26",
          6723 => x"12",
          6724 => x"06",
          6725 => x"30",
          6726 => x"51",
          6727 => x"2e",
          6728 => x"85",
          6729 => x"be",
          6730 => x"74",
          6731 => x"30",
          6732 => x"9f",
          6733 => x"2a",
          6734 => x"54",
          6735 => x"2e",
          6736 => x"15",
          6737 => x"55",
          6738 => x"ff",
          6739 => x"39",
          6740 => x"86",
          6741 => x"7c",
          6742 => x"51",
          6743 => x"d3",
          6744 => x"70",
          6745 => x"0c",
          6746 => x"04",
          6747 => x"78",
          6748 => x"83",
          6749 => x"0b",
          6750 => x"79",
          6751 => x"e2",
          6752 => x"55",
          6753 => x"08",
          6754 => x"84",
          6755 => x"df",
          6756 => x"bb",
          6757 => x"ff",
          6758 => x"83",
          6759 => x"d4",
          6760 => x"81",
          6761 => x"38",
          6762 => x"17",
          6763 => x"74",
          6764 => x"09",
          6765 => x"38",
          6766 => x"81",
          6767 => x"30",
          6768 => x"79",
          6769 => x"54",
          6770 => x"74",
          6771 => x"09",
          6772 => x"38",
          6773 => x"b4",
          6774 => x"ea",
          6775 => x"b1",
          6776 => x"dc",
          6777 => x"bb",
          6778 => x"2e",
          6779 => x"53",
          6780 => x"52",
          6781 => x"51",
          6782 => x"82",
          6783 => x"55",
          6784 => x"08",
          6785 => x"38",
          6786 => x"82",
          6787 => x"88",
          6788 => x"f2",
          6789 => x"02",
          6790 => x"cb",
          6791 => x"55",
          6792 => x"60",
          6793 => x"3f",
          6794 => x"08",
          6795 => x"80",
          6796 => x"dc",
          6797 => x"fc",
          6798 => x"dc",
          6799 => x"82",
          6800 => x"70",
          6801 => x"8c",
          6802 => x"2e",
          6803 => x"73",
          6804 => x"81",
          6805 => x"33",
          6806 => x"80",
          6807 => x"81",
          6808 => x"d7",
          6809 => x"bb",
          6810 => x"ff",
          6811 => x"06",
          6812 => x"98",
          6813 => x"2e",
          6814 => x"74",
          6815 => x"81",
          6816 => x"8a",
          6817 => x"ac",
          6818 => x"39",
          6819 => x"77",
          6820 => x"81",
          6821 => x"33",
          6822 => x"3f",
          6823 => x"08",
          6824 => x"70",
          6825 => x"55",
          6826 => x"86",
          6827 => x"80",
          6828 => x"74",
          6829 => x"81",
          6830 => x"8a",
          6831 => x"f4",
          6832 => x"53",
          6833 => x"fd",
          6834 => x"bb",
          6835 => x"ff",
          6836 => x"82",
          6837 => x"06",
          6838 => x"8c",
          6839 => x"58",
          6840 => x"f6",
          6841 => x"58",
          6842 => x"2e",
          6843 => x"fa",
          6844 => x"e8",
          6845 => x"dc",
          6846 => x"78",
          6847 => x"5a",
          6848 => x"90",
          6849 => x"75",
          6850 => x"38",
          6851 => x"3d",
          6852 => x"70",
          6853 => x"08",
          6854 => x"7a",
          6855 => x"38",
          6856 => x"51",
          6857 => x"82",
          6858 => x"81",
          6859 => x"81",
          6860 => x"38",
          6861 => x"83",
          6862 => x"38",
          6863 => x"84",
          6864 => x"38",
          6865 => x"81",
          6866 => x"38",
          6867 => x"db",
          6868 => x"bb",
          6869 => x"ff",
          6870 => x"72",
          6871 => x"09",
          6872 => x"d0",
          6873 => x"14",
          6874 => x"3f",
          6875 => x"08",
          6876 => x"06",
          6877 => x"38",
          6878 => x"51",
          6879 => x"82",
          6880 => x"58",
          6881 => x"0c",
          6882 => x"33",
          6883 => x"80",
          6884 => x"ff",
          6885 => x"ff",
          6886 => x"55",
          6887 => x"81",
          6888 => x"38",
          6889 => x"06",
          6890 => x"80",
          6891 => x"52",
          6892 => x"8a",
          6893 => x"80",
          6894 => x"ff",
          6895 => x"53",
          6896 => x"86",
          6897 => x"83",
          6898 => x"c5",
          6899 => x"f5",
          6900 => x"dc",
          6901 => x"bb",
          6902 => x"15",
          6903 => x"06",
          6904 => x"76",
          6905 => x"80",
          6906 => x"da",
          6907 => x"bb",
          6908 => x"ff",
          6909 => x"74",
          6910 => x"d4",
          6911 => x"dc",
          6912 => x"dc",
          6913 => x"c2",
          6914 => x"b9",
          6915 => x"dc",
          6916 => x"ff",
          6917 => x"56",
          6918 => x"83",
          6919 => x"14",
          6920 => x"71",
          6921 => x"5a",
          6922 => x"26",
          6923 => x"8a",
          6924 => x"74",
          6925 => x"fe",
          6926 => x"82",
          6927 => x"55",
          6928 => x"08",
          6929 => x"ec",
          6930 => x"dc",
          6931 => x"ff",
          6932 => x"83",
          6933 => x"74",
          6934 => x"26",
          6935 => x"57",
          6936 => x"26",
          6937 => x"57",
          6938 => x"56",
          6939 => x"82",
          6940 => x"15",
          6941 => x"0c",
          6942 => x"0c",
          6943 => x"a4",
          6944 => x"1d",
          6945 => x"54",
          6946 => x"2e",
          6947 => x"af",
          6948 => x"14",
          6949 => x"3f",
          6950 => x"08",
          6951 => x"06",
          6952 => x"72",
          6953 => x"79",
          6954 => x"80",
          6955 => x"d9",
          6956 => x"bb",
          6957 => x"15",
          6958 => x"2b",
          6959 => x"8d",
          6960 => x"2e",
          6961 => x"77",
          6962 => x"0c",
          6963 => x"76",
          6964 => x"38",
          6965 => x"70",
          6966 => x"81",
          6967 => x"53",
          6968 => x"89",
          6969 => x"56",
          6970 => x"08",
          6971 => x"38",
          6972 => x"15",
          6973 => x"8c",
          6974 => x"80",
          6975 => x"34",
          6976 => x"09",
          6977 => x"92",
          6978 => x"14",
          6979 => x"3f",
          6980 => x"08",
          6981 => x"06",
          6982 => x"2e",
          6983 => x"80",
          6984 => x"1b",
          6985 => x"db",
          6986 => x"bb",
          6987 => x"ea",
          6988 => x"dc",
          6989 => x"34",
          6990 => x"51",
          6991 => x"82",
          6992 => x"83",
          6993 => x"53",
          6994 => x"d5",
          6995 => x"06",
          6996 => x"b4",
          6997 => x"84",
          6998 => x"dc",
          6999 => x"85",
          7000 => x"09",
          7001 => x"38",
          7002 => x"51",
          7003 => x"82",
          7004 => x"86",
          7005 => x"f2",
          7006 => x"06",
          7007 => x"9c",
          7008 => x"d8",
          7009 => x"dc",
          7010 => x"0c",
          7011 => x"51",
          7012 => x"82",
          7013 => x"8c",
          7014 => x"74",
          7015 => x"a4",
          7016 => x"53",
          7017 => x"a4",
          7018 => x"15",
          7019 => x"94",
          7020 => x"56",
          7021 => x"dc",
          7022 => x"0d",
          7023 => x"0d",
          7024 => x"55",
          7025 => x"b9",
          7026 => x"53",
          7027 => x"b1",
          7028 => x"52",
          7029 => x"a9",
          7030 => x"22",
          7031 => x"57",
          7032 => x"2e",
          7033 => x"99",
          7034 => x"33",
          7035 => x"3f",
          7036 => x"08",
          7037 => x"71",
          7038 => x"74",
          7039 => x"83",
          7040 => x"78",
          7041 => x"52",
          7042 => x"dc",
          7043 => x"0d",
          7044 => x"0d",
          7045 => x"33",
          7046 => x"3d",
          7047 => x"56",
          7048 => x"8b",
          7049 => x"82",
          7050 => x"24",
          7051 => x"bb",
          7052 => x"29",
          7053 => x"05",
          7054 => x"55",
          7055 => x"84",
          7056 => x"34",
          7057 => x"80",
          7058 => x"80",
          7059 => x"75",
          7060 => x"75",
          7061 => x"38",
          7062 => x"3d",
          7063 => x"05",
          7064 => x"3f",
          7065 => x"08",
          7066 => x"bb",
          7067 => x"3d",
          7068 => x"3d",
          7069 => x"84",
          7070 => x"05",
          7071 => x"89",
          7072 => x"2e",
          7073 => x"77",
          7074 => x"54",
          7075 => x"05",
          7076 => x"84",
          7077 => x"f6",
          7078 => x"bb",
          7079 => x"82",
          7080 => x"84",
          7081 => x"5c",
          7082 => x"3d",
          7083 => x"ed",
          7084 => x"bb",
          7085 => x"82",
          7086 => x"92",
          7087 => x"d7",
          7088 => x"98",
          7089 => x"73",
          7090 => x"38",
          7091 => x"9c",
          7092 => x"80",
          7093 => x"38",
          7094 => x"95",
          7095 => x"2e",
          7096 => x"aa",
          7097 => x"ea",
          7098 => x"bb",
          7099 => x"9e",
          7100 => x"05",
          7101 => x"54",
          7102 => x"38",
          7103 => x"70",
          7104 => x"54",
          7105 => x"8e",
          7106 => x"83",
          7107 => x"88",
          7108 => x"83",
          7109 => x"83",
          7110 => x"06",
          7111 => x"80",
          7112 => x"38",
          7113 => x"51",
          7114 => x"82",
          7115 => x"56",
          7116 => x"0a",
          7117 => x"05",
          7118 => x"3f",
          7119 => x"0b",
          7120 => x"80",
          7121 => x"7a",
          7122 => x"3f",
          7123 => x"9c",
          7124 => x"d1",
          7125 => x"81",
          7126 => x"34",
          7127 => x"80",
          7128 => x"b0",
          7129 => x"54",
          7130 => x"52",
          7131 => x"05",
          7132 => x"3f",
          7133 => x"08",
          7134 => x"dc",
          7135 => x"38",
          7136 => x"82",
          7137 => x"b2",
          7138 => x"84",
          7139 => x"06",
          7140 => x"73",
          7141 => x"38",
          7142 => x"ad",
          7143 => x"2a",
          7144 => x"51",
          7145 => x"2e",
          7146 => x"81",
          7147 => x"80",
          7148 => x"87",
          7149 => x"39",
          7150 => x"51",
          7151 => x"82",
          7152 => x"7b",
          7153 => x"12",
          7154 => x"82",
          7155 => x"81",
          7156 => x"83",
          7157 => x"06",
          7158 => x"80",
          7159 => x"77",
          7160 => x"58",
          7161 => x"08",
          7162 => x"63",
          7163 => x"63",
          7164 => x"57",
          7165 => x"82",
          7166 => x"82",
          7167 => x"88",
          7168 => x"9c",
          7169 => x"d2",
          7170 => x"bb",
          7171 => x"bb",
          7172 => x"1b",
          7173 => x"0c",
          7174 => x"22",
          7175 => x"77",
          7176 => x"80",
          7177 => x"34",
          7178 => x"1a",
          7179 => x"94",
          7180 => x"85",
          7181 => x"06",
          7182 => x"80",
          7183 => x"38",
          7184 => x"08",
          7185 => x"84",
          7186 => x"dc",
          7187 => x"0c",
          7188 => x"70",
          7189 => x"52",
          7190 => x"39",
          7191 => x"51",
          7192 => x"82",
          7193 => x"57",
          7194 => x"08",
          7195 => x"38",
          7196 => x"bb",
          7197 => x"2e",
          7198 => x"83",
          7199 => x"75",
          7200 => x"74",
          7201 => x"07",
          7202 => x"54",
          7203 => x"8a",
          7204 => x"75",
          7205 => x"73",
          7206 => x"98",
          7207 => x"a9",
          7208 => x"ff",
          7209 => x"80",
          7210 => x"76",
          7211 => x"d6",
          7212 => x"bb",
          7213 => x"38",
          7214 => x"39",
          7215 => x"82",
          7216 => x"05",
          7217 => x"84",
          7218 => x"0c",
          7219 => x"82",
          7220 => x"97",
          7221 => x"f2",
          7222 => x"63",
          7223 => x"40",
          7224 => x"7e",
          7225 => x"fc",
          7226 => x"51",
          7227 => x"82",
          7228 => x"55",
          7229 => x"08",
          7230 => x"19",
          7231 => x"80",
          7232 => x"74",
          7233 => x"39",
          7234 => x"81",
          7235 => x"56",
          7236 => x"82",
          7237 => x"39",
          7238 => x"1a",
          7239 => x"82",
          7240 => x"0b",
          7241 => x"81",
          7242 => x"39",
          7243 => x"94",
          7244 => x"55",
          7245 => x"83",
          7246 => x"7b",
          7247 => x"89",
          7248 => x"08",
          7249 => x"06",
          7250 => x"81",
          7251 => x"8a",
          7252 => x"05",
          7253 => x"06",
          7254 => x"a8",
          7255 => x"38",
          7256 => x"55",
          7257 => x"19",
          7258 => x"51",
          7259 => x"82",
          7260 => x"55",
          7261 => x"ff",
          7262 => x"ff",
          7263 => x"38",
          7264 => x"0c",
          7265 => x"52",
          7266 => x"cb",
          7267 => x"dc",
          7268 => x"ff",
          7269 => x"bb",
          7270 => x"7c",
          7271 => x"57",
          7272 => x"80",
          7273 => x"1a",
          7274 => x"22",
          7275 => x"75",
          7276 => x"38",
          7277 => x"58",
          7278 => x"53",
          7279 => x"1b",
          7280 => x"88",
          7281 => x"dc",
          7282 => x"38",
          7283 => x"33",
          7284 => x"80",
          7285 => x"b0",
          7286 => x"31",
          7287 => x"27",
          7288 => x"80",
          7289 => x"52",
          7290 => x"77",
          7291 => x"7d",
          7292 => x"e0",
          7293 => x"2b",
          7294 => x"76",
          7295 => x"94",
          7296 => x"ff",
          7297 => x"71",
          7298 => x"7b",
          7299 => x"38",
          7300 => x"19",
          7301 => x"51",
          7302 => x"82",
          7303 => x"fe",
          7304 => x"53",
          7305 => x"83",
          7306 => x"b4",
          7307 => x"51",
          7308 => x"7b",
          7309 => x"08",
          7310 => x"76",
          7311 => x"08",
          7312 => x"0c",
          7313 => x"f3",
          7314 => x"75",
          7315 => x"0c",
          7316 => x"04",
          7317 => x"60",
          7318 => x"40",
          7319 => x"80",
          7320 => x"3d",
          7321 => x"77",
          7322 => x"3f",
          7323 => x"08",
          7324 => x"dc",
          7325 => x"91",
          7326 => x"74",
          7327 => x"38",
          7328 => x"b8",
          7329 => x"33",
          7330 => x"70",
          7331 => x"56",
          7332 => x"74",
          7333 => x"a4",
          7334 => x"82",
          7335 => x"34",
          7336 => x"98",
          7337 => x"91",
          7338 => x"56",
          7339 => x"94",
          7340 => x"11",
          7341 => x"76",
          7342 => x"75",
          7343 => x"80",
          7344 => x"38",
          7345 => x"70",
          7346 => x"56",
          7347 => x"fd",
          7348 => x"11",
          7349 => x"77",
          7350 => x"5c",
          7351 => x"38",
          7352 => x"88",
          7353 => x"74",
          7354 => x"52",
          7355 => x"18",
          7356 => x"51",
          7357 => x"82",
          7358 => x"55",
          7359 => x"08",
          7360 => x"ab",
          7361 => x"2e",
          7362 => x"74",
          7363 => x"95",
          7364 => x"19",
          7365 => x"08",
          7366 => x"88",
          7367 => x"55",
          7368 => x"9c",
          7369 => x"09",
          7370 => x"38",
          7371 => x"c1",
          7372 => x"dc",
          7373 => x"38",
          7374 => x"52",
          7375 => x"97",
          7376 => x"dc",
          7377 => x"fe",
          7378 => x"bb",
          7379 => x"7c",
          7380 => x"57",
          7381 => x"80",
          7382 => x"1b",
          7383 => x"22",
          7384 => x"75",
          7385 => x"38",
          7386 => x"59",
          7387 => x"53",
          7388 => x"1a",
          7389 => x"be",
          7390 => x"dc",
          7391 => x"38",
          7392 => x"08",
          7393 => x"56",
          7394 => x"9b",
          7395 => x"53",
          7396 => x"77",
          7397 => x"7d",
          7398 => x"16",
          7399 => x"3f",
          7400 => x"0b",
          7401 => x"78",
          7402 => x"80",
          7403 => x"18",
          7404 => x"08",
          7405 => x"7e",
          7406 => x"3f",
          7407 => x"08",
          7408 => x"7e",
          7409 => x"0c",
          7410 => x"19",
          7411 => x"08",
          7412 => x"84",
          7413 => x"57",
          7414 => x"27",
          7415 => x"56",
          7416 => x"52",
          7417 => x"f9",
          7418 => x"dc",
          7419 => x"38",
          7420 => x"52",
          7421 => x"83",
          7422 => x"b4",
          7423 => x"d4",
          7424 => x"81",
          7425 => x"34",
          7426 => x"7e",
          7427 => x"0c",
          7428 => x"1a",
          7429 => x"94",
          7430 => x"1b",
          7431 => x"5e",
          7432 => x"27",
          7433 => x"55",
          7434 => x"0c",
          7435 => x"90",
          7436 => x"c0",
          7437 => x"90",
          7438 => x"56",
          7439 => x"dc",
          7440 => x"0d",
          7441 => x"0d",
          7442 => x"fc",
          7443 => x"52",
          7444 => x"3f",
          7445 => x"08",
          7446 => x"dc",
          7447 => x"38",
          7448 => x"70",
          7449 => x"81",
          7450 => x"55",
          7451 => x"80",
          7452 => x"16",
          7453 => x"51",
          7454 => x"82",
          7455 => x"57",
          7456 => x"08",
          7457 => x"a4",
          7458 => x"11",
          7459 => x"55",
          7460 => x"16",
          7461 => x"08",
          7462 => x"75",
          7463 => x"e8",
          7464 => x"08",
          7465 => x"51",
          7466 => x"82",
          7467 => x"52",
          7468 => x"c9",
          7469 => x"52",
          7470 => x"c9",
          7471 => x"54",
          7472 => x"15",
          7473 => x"cc",
          7474 => x"bb",
          7475 => x"17",
          7476 => x"06",
          7477 => x"90",
          7478 => x"82",
          7479 => x"8a",
          7480 => x"fc",
          7481 => x"70",
          7482 => x"d9",
          7483 => x"dc",
          7484 => x"bb",
          7485 => x"38",
          7486 => x"05",
          7487 => x"f1",
          7488 => x"bb",
          7489 => x"82",
          7490 => x"87",
          7491 => x"dc",
          7492 => x"72",
          7493 => x"0c",
          7494 => x"04",
          7495 => x"84",
          7496 => x"e4",
          7497 => x"80",
          7498 => x"dc",
          7499 => x"38",
          7500 => x"08",
          7501 => x"34",
          7502 => x"82",
          7503 => x"83",
          7504 => x"ef",
          7505 => x"53",
          7506 => x"05",
          7507 => x"51",
          7508 => x"82",
          7509 => x"55",
          7510 => x"08",
          7511 => x"76",
          7512 => x"93",
          7513 => x"51",
          7514 => x"82",
          7515 => x"55",
          7516 => x"08",
          7517 => x"80",
          7518 => x"70",
          7519 => x"56",
          7520 => x"89",
          7521 => x"94",
          7522 => x"b2",
          7523 => x"05",
          7524 => x"2a",
          7525 => x"51",
          7526 => x"80",
          7527 => x"76",
          7528 => x"52",
          7529 => x"3f",
          7530 => x"08",
          7531 => x"8e",
          7532 => x"dc",
          7533 => x"09",
          7534 => x"38",
          7535 => x"82",
          7536 => x"93",
          7537 => x"e4",
          7538 => x"6f",
          7539 => x"7a",
          7540 => x"9e",
          7541 => x"05",
          7542 => x"51",
          7543 => x"82",
          7544 => x"57",
          7545 => x"08",
          7546 => x"7b",
          7547 => x"94",
          7548 => x"55",
          7549 => x"73",
          7550 => x"ed",
          7551 => x"93",
          7552 => x"55",
          7553 => x"82",
          7554 => x"57",
          7555 => x"08",
          7556 => x"68",
          7557 => x"c9",
          7558 => x"bb",
          7559 => x"82",
          7560 => x"82",
          7561 => x"52",
          7562 => x"a3",
          7563 => x"dc",
          7564 => x"52",
          7565 => x"b8",
          7566 => x"dc",
          7567 => x"bb",
          7568 => x"a2",
          7569 => x"74",
          7570 => x"3f",
          7571 => x"08",
          7572 => x"dc",
          7573 => x"69",
          7574 => x"d9",
          7575 => x"82",
          7576 => x"2e",
          7577 => x"52",
          7578 => x"cf",
          7579 => x"dc",
          7580 => x"bb",
          7581 => x"2e",
          7582 => x"84",
          7583 => x"06",
          7584 => x"57",
          7585 => x"76",
          7586 => x"9e",
          7587 => x"05",
          7588 => x"dc",
          7589 => x"90",
          7590 => x"81",
          7591 => x"56",
          7592 => x"80",
          7593 => x"02",
          7594 => x"81",
          7595 => x"70",
          7596 => x"56",
          7597 => x"81",
          7598 => x"78",
          7599 => x"38",
          7600 => x"99",
          7601 => x"81",
          7602 => x"18",
          7603 => x"18",
          7604 => x"58",
          7605 => x"33",
          7606 => x"ee",
          7607 => x"6f",
          7608 => x"af",
          7609 => x"8d",
          7610 => x"2e",
          7611 => x"8a",
          7612 => x"6f",
          7613 => x"af",
          7614 => x"0b",
          7615 => x"33",
          7616 => x"82",
          7617 => x"70",
          7618 => x"52",
          7619 => x"56",
          7620 => x"8d",
          7621 => x"70",
          7622 => x"51",
          7623 => x"f5",
          7624 => x"54",
          7625 => x"a7",
          7626 => x"74",
          7627 => x"38",
          7628 => x"73",
          7629 => x"81",
          7630 => x"81",
          7631 => x"39",
          7632 => x"81",
          7633 => x"74",
          7634 => x"81",
          7635 => x"91",
          7636 => x"6e",
          7637 => x"59",
          7638 => x"7a",
          7639 => x"5c",
          7640 => x"26",
          7641 => x"7a",
          7642 => x"bb",
          7643 => x"3d",
          7644 => x"3d",
          7645 => x"8d",
          7646 => x"54",
          7647 => x"55",
          7648 => x"82",
          7649 => x"53",
          7650 => x"08",
          7651 => x"91",
          7652 => x"72",
          7653 => x"8c",
          7654 => x"73",
          7655 => x"38",
          7656 => x"70",
          7657 => x"81",
          7658 => x"57",
          7659 => x"73",
          7660 => x"08",
          7661 => x"94",
          7662 => x"75",
          7663 => x"97",
          7664 => x"11",
          7665 => x"2b",
          7666 => x"73",
          7667 => x"38",
          7668 => x"16",
          7669 => x"ad",
          7670 => x"dc",
          7671 => x"78",
          7672 => x"55",
          7673 => x"9d",
          7674 => x"dc",
          7675 => x"96",
          7676 => x"70",
          7677 => x"94",
          7678 => x"71",
          7679 => x"08",
          7680 => x"53",
          7681 => x"15",
          7682 => x"a6",
          7683 => x"74",
          7684 => x"3f",
          7685 => x"08",
          7686 => x"dc",
          7687 => x"81",
          7688 => x"bb",
          7689 => x"2e",
          7690 => x"82",
          7691 => x"88",
          7692 => x"98",
          7693 => x"80",
          7694 => x"38",
          7695 => x"80",
          7696 => x"77",
          7697 => x"08",
          7698 => x"0c",
          7699 => x"70",
          7700 => x"81",
          7701 => x"5a",
          7702 => x"2e",
          7703 => x"52",
          7704 => x"f9",
          7705 => x"dc",
          7706 => x"bb",
          7707 => x"38",
          7708 => x"08",
          7709 => x"73",
          7710 => x"c7",
          7711 => x"bb",
          7712 => x"73",
          7713 => x"38",
          7714 => x"af",
          7715 => x"73",
          7716 => x"27",
          7717 => x"98",
          7718 => x"a0",
          7719 => x"08",
          7720 => x"0c",
          7721 => x"06",
          7722 => x"2e",
          7723 => x"52",
          7724 => x"a3",
          7725 => x"dc",
          7726 => x"82",
          7727 => x"34",
          7728 => x"c4",
          7729 => x"91",
          7730 => x"53",
          7731 => x"89",
          7732 => x"dc",
          7733 => x"94",
          7734 => x"8c",
          7735 => x"27",
          7736 => x"8c",
          7737 => x"15",
          7738 => x"07",
          7739 => x"16",
          7740 => x"ff",
          7741 => x"80",
          7742 => x"77",
          7743 => x"2e",
          7744 => x"9c",
          7745 => x"53",
          7746 => x"dc",
          7747 => x"0d",
          7748 => x"0d",
          7749 => x"54",
          7750 => x"81",
          7751 => x"53",
          7752 => x"05",
          7753 => x"84",
          7754 => x"e7",
          7755 => x"dc",
          7756 => x"bb",
          7757 => x"ea",
          7758 => x"0c",
          7759 => x"51",
          7760 => x"82",
          7761 => x"55",
          7762 => x"08",
          7763 => x"ab",
          7764 => x"98",
          7765 => x"80",
          7766 => x"38",
          7767 => x"70",
          7768 => x"81",
          7769 => x"57",
          7770 => x"ad",
          7771 => x"08",
          7772 => x"d3",
          7773 => x"bb",
          7774 => x"17",
          7775 => x"86",
          7776 => x"17",
          7777 => x"75",
          7778 => x"3f",
          7779 => x"08",
          7780 => x"2e",
          7781 => x"85",
          7782 => x"86",
          7783 => x"2e",
          7784 => x"76",
          7785 => x"73",
          7786 => x"0c",
          7787 => x"04",
          7788 => x"76",
          7789 => x"05",
          7790 => x"53",
          7791 => x"82",
          7792 => x"87",
          7793 => x"dc",
          7794 => x"86",
          7795 => x"fb",
          7796 => x"79",
          7797 => x"05",
          7798 => x"56",
          7799 => x"3f",
          7800 => x"08",
          7801 => x"dc",
          7802 => x"38",
          7803 => x"82",
          7804 => x"52",
          7805 => x"f8",
          7806 => x"dc",
          7807 => x"ca",
          7808 => x"dc",
          7809 => x"51",
          7810 => x"82",
          7811 => x"53",
          7812 => x"08",
          7813 => x"81",
          7814 => x"80",
          7815 => x"82",
          7816 => x"a6",
          7817 => x"73",
          7818 => x"3f",
          7819 => x"51",
          7820 => x"82",
          7821 => x"84",
          7822 => x"70",
          7823 => x"2c",
          7824 => x"dc",
          7825 => x"51",
          7826 => x"82",
          7827 => x"87",
          7828 => x"ee",
          7829 => x"57",
          7830 => x"3d",
          7831 => x"3d",
          7832 => x"af",
          7833 => x"dc",
          7834 => x"bb",
          7835 => x"38",
          7836 => x"51",
          7837 => x"82",
          7838 => x"55",
          7839 => x"08",
          7840 => x"80",
          7841 => x"70",
          7842 => x"58",
          7843 => x"85",
          7844 => x"8d",
          7845 => x"2e",
          7846 => x"52",
          7847 => x"be",
          7848 => x"bb",
          7849 => x"3d",
          7850 => x"3d",
          7851 => x"55",
          7852 => x"92",
          7853 => x"52",
          7854 => x"de",
          7855 => x"bb",
          7856 => x"82",
          7857 => x"82",
          7858 => x"74",
          7859 => x"98",
          7860 => x"11",
          7861 => x"59",
          7862 => x"75",
          7863 => x"38",
          7864 => x"81",
          7865 => x"5b",
          7866 => x"82",
          7867 => x"39",
          7868 => x"08",
          7869 => x"59",
          7870 => x"09",
          7871 => x"38",
          7872 => x"57",
          7873 => x"3d",
          7874 => x"c1",
          7875 => x"bb",
          7876 => x"2e",
          7877 => x"bb",
          7878 => x"2e",
          7879 => x"bb",
          7880 => x"70",
          7881 => x"08",
          7882 => x"7a",
          7883 => x"7f",
          7884 => x"54",
          7885 => x"77",
          7886 => x"80",
          7887 => x"15",
          7888 => x"dc",
          7889 => x"75",
          7890 => x"52",
          7891 => x"52",
          7892 => x"8d",
          7893 => x"dc",
          7894 => x"bb",
          7895 => x"d6",
          7896 => x"33",
          7897 => x"1a",
          7898 => x"54",
          7899 => x"09",
          7900 => x"38",
          7901 => x"ff",
          7902 => x"82",
          7903 => x"83",
          7904 => x"70",
          7905 => x"25",
          7906 => x"59",
          7907 => x"9b",
          7908 => x"51",
          7909 => x"3f",
          7910 => x"08",
          7911 => x"70",
          7912 => x"25",
          7913 => x"59",
          7914 => x"75",
          7915 => x"7a",
          7916 => x"ff",
          7917 => x"7c",
          7918 => x"90",
          7919 => x"11",
          7920 => x"56",
          7921 => x"15",
          7922 => x"bb",
          7923 => x"3d",
          7924 => x"3d",
          7925 => x"3d",
          7926 => x"70",
          7927 => x"dd",
          7928 => x"dc",
          7929 => x"bb",
          7930 => x"a8",
          7931 => x"33",
          7932 => x"a0",
          7933 => x"33",
          7934 => x"70",
          7935 => x"55",
          7936 => x"73",
          7937 => x"8e",
          7938 => x"08",
          7939 => x"18",
          7940 => x"80",
          7941 => x"38",
          7942 => x"08",
          7943 => x"08",
          7944 => x"c4",
          7945 => x"bb",
          7946 => x"88",
          7947 => x"80",
          7948 => x"17",
          7949 => x"51",
          7950 => x"3f",
          7951 => x"08",
          7952 => x"81",
          7953 => x"81",
          7954 => x"dc",
          7955 => x"09",
          7956 => x"38",
          7957 => x"39",
          7958 => x"77",
          7959 => x"dc",
          7960 => x"08",
          7961 => x"98",
          7962 => x"82",
          7963 => x"52",
          7964 => x"bd",
          7965 => x"dc",
          7966 => x"17",
          7967 => x"0c",
          7968 => x"80",
          7969 => x"73",
          7970 => x"75",
          7971 => x"38",
          7972 => x"34",
          7973 => x"82",
          7974 => x"89",
          7975 => x"e2",
          7976 => x"53",
          7977 => x"a4",
          7978 => x"3d",
          7979 => x"3f",
          7980 => x"08",
          7981 => x"dc",
          7982 => x"38",
          7983 => x"3d",
          7984 => x"3d",
          7985 => x"d1",
          7986 => x"bb",
          7987 => x"82",
          7988 => x"81",
          7989 => x"80",
          7990 => x"70",
          7991 => x"81",
          7992 => x"56",
          7993 => x"81",
          7994 => x"98",
          7995 => x"74",
          7996 => x"38",
          7997 => x"05",
          7998 => x"06",
          7999 => x"55",
          8000 => x"38",
          8001 => x"51",
          8002 => x"82",
          8003 => x"74",
          8004 => x"81",
          8005 => x"56",
          8006 => x"80",
          8007 => x"54",
          8008 => x"08",
          8009 => x"2e",
          8010 => x"73",
          8011 => x"dc",
          8012 => x"52",
          8013 => x"52",
          8014 => x"3f",
          8015 => x"08",
          8016 => x"dc",
          8017 => x"38",
          8018 => x"08",
          8019 => x"cc",
          8020 => x"bb",
          8021 => x"82",
          8022 => x"86",
          8023 => x"80",
          8024 => x"bb",
          8025 => x"2e",
          8026 => x"bb",
          8027 => x"c0",
          8028 => x"ce",
          8029 => x"bb",
          8030 => x"bb",
          8031 => x"70",
          8032 => x"08",
          8033 => x"51",
          8034 => x"80",
          8035 => x"73",
          8036 => x"38",
          8037 => x"52",
          8038 => x"95",
          8039 => x"dc",
          8040 => x"8c",
          8041 => x"ff",
          8042 => x"82",
          8043 => x"55",
          8044 => x"dc",
          8045 => x"0d",
          8046 => x"0d",
          8047 => x"3d",
          8048 => x"9a",
          8049 => x"cb",
          8050 => x"dc",
          8051 => x"bb",
          8052 => x"b0",
          8053 => x"69",
          8054 => x"70",
          8055 => x"97",
          8056 => x"dc",
          8057 => x"bb",
          8058 => x"38",
          8059 => x"94",
          8060 => x"dc",
          8061 => x"09",
          8062 => x"88",
          8063 => x"df",
          8064 => x"85",
          8065 => x"51",
          8066 => x"74",
          8067 => x"78",
          8068 => x"8a",
          8069 => x"57",
          8070 => x"82",
          8071 => x"75",
          8072 => x"bb",
          8073 => x"38",
          8074 => x"bb",
          8075 => x"2e",
          8076 => x"83",
          8077 => x"82",
          8078 => x"ff",
          8079 => x"06",
          8080 => x"54",
          8081 => x"73",
          8082 => x"82",
          8083 => x"52",
          8084 => x"a4",
          8085 => x"dc",
          8086 => x"bb",
          8087 => x"9a",
          8088 => x"a0",
          8089 => x"51",
          8090 => x"3f",
          8091 => x"0b",
          8092 => x"78",
          8093 => x"bf",
          8094 => x"88",
          8095 => x"80",
          8096 => x"ff",
          8097 => x"75",
          8098 => x"11",
          8099 => x"f8",
          8100 => x"78",
          8101 => x"80",
          8102 => x"ff",
          8103 => x"78",
          8104 => x"80",
          8105 => x"7f",
          8106 => x"d4",
          8107 => x"c9",
          8108 => x"54",
          8109 => x"15",
          8110 => x"cb",
          8111 => x"bb",
          8112 => x"82",
          8113 => x"b2",
          8114 => x"b2",
          8115 => x"96",
          8116 => x"b5",
          8117 => x"53",
          8118 => x"51",
          8119 => x"64",
          8120 => x"8b",
          8121 => x"54",
          8122 => x"15",
          8123 => x"ff",
          8124 => x"82",
          8125 => x"54",
          8126 => x"53",
          8127 => x"51",
          8128 => x"3f",
          8129 => x"dc",
          8130 => x"0d",
          8131 => x"0d",
          8132 => x"05",
          8133 => x"3f",
          8134 => x"3d",
          8135 => x"52",
          8136 => x"d5",
          8137 => x"bb",
          8138 => x"82",
          8139 => x"82",
          8140 => x"4d",
          8141 => x"52",
          8142 => x"52",
          8143 => x"3f",
          8144 => x"08",
          8145 => x"dc",
          8146 => x"38",
          8147 => x"05",
          8148 => x"06",
          8149 => x"73",
          8150 => x"a0",
          8151 => x"08",
          8152 => x"ff",
          8153 => x"ff",
          8154 => x"ac",
          8155 => x"92",
          8156 => x"54",
          8157 => x"3f",
          8158 => x"52",
          8159 => x"f7",
          8160 => x"dc",
          8161 => x"bb",
          8162 => x"38",
          8163 => x"09",
          8164 => x"38",
          8165 => x"08",
          8166 => x"88",
          8167 => x"39",
          8168 => x"08",
          8169 => x"81",
          8170 => x"38",
          8171 => x"b1",
          8172 => x"dc",
          8173 => x"bb",
          8174 => x"c8",
          8175 => x"93",
          8176 => x"ff",
          8177 => x"8d",
          8178 => x"b4",
          8179 => x"af",
          8180 => x"17",
          8181 => x"33",
          8182 => x"70",
          8183 => x"55",
          8184 => x"38",
          8185 => x"54",
          8186 => x"34",
          8187 => x"0b",
          8188 => x"8b",
          8189 => x"84",
          8190 => x"06",
          8191 => x"73",
          8192 => x"e5",
          8193 => x"2e",
          8194 => x"75",
          8195 => x"c6",
          8196 => x"bb",
          8197 => x"78",
          8198 => x"bb",
          8199 => x"82",
          8200 => x"80",
          8201 => x"38",
          8202 => x"08",
          8203 => x"ff",
          8204 => x"82",
          8205 => x"79",
          8206 => x"58",
          8207 => x"bb",
          8208 => x"c0",
          8209 => x"33",
          8210 => x"2e",
          8211 => x"99",
          8212 => x"75",
          8213 => x"c6",
          8214 => x"54",
          8215 => x"15",
          8216 => x"82",
          8217 => x"9c",
          8218 => x"c8",
          8219 => x"bb",
          8220 => x"82",
          8221 => x"8c",
          8222 => x"ff",
          8223 => x"82",
          8224 => x"55",
          8225 => x"dc",
          8226 => x"0d",
          8227 => x"0d",
          8228 => x"05",
          8229 => x"05",
          8230 => x"33",
          8231 => x"53",
          8232 => x"05",
          8233 => x"51",
          8234 => x"82",
          8235 => x"55",
          8236 => x"08",
          8237 => x"78",
          8238 => x"95",
          8239 => x"51",
          8240 => x"82",
          8241 => x"55",
          8242 => x"08",
          8243 => x"80",
          8244 => x"81",
          8245 => x"86",
          8246 => x"38",
          8247 => x"61",
          8248 => x"12",
          8249 => x"7a",
          8250 => x"51",
          8251 => x"74",
          8252 => x"78",
          8253 => x"83",
          8254 => x"51",
          8255 => x"3f",
          8256 => x"08",
          8257 => x"bb",
          8258 => x"3d",
          8259 => x"3d",
          8260 => x"82",
          8261 => x"d0",
          8262 => x"3d",
          8263 => x"3f",
          8264 => x"08",
          8265 => x"dc",
          8266 => x"38",
          8267 => x"52",
          8268 => x"05",
          8269 => x"3f",
          8270 => x"08",
          8271 => x"dc",
          8272 => x"02",
          8273 => x"33",
          8274 => x"54",
          8275 => x"a6",
          8276 => x"22",
          8277 => x"71",
          8278 => x"53",
          8279 => x"51",
          8280 => x"3f",
          8281 => x"0b",
          8282 => x"76",
          8283 => x"b8",
          8284 => x"dc",
          8285 => x"82",
          8286 => x"93",
          8287 => x"ea",
          8288 => x"6b",
          8289 => x"53",
          8290 => x"05",
          8291 => x"51",
          8292 => x"82",
          8293 => x"82",
          8294 => x"30",
          8295 => x"dc",
          8296 => x"25",
          8297 => x"79",
          8298 => x"85",
          8299 => x"75",
          8300 => x"73",
          8301 => x"f9",
          8302 => x"80",
          8303 => x"8d",
          8304 => x"54",
          8305 => x"3f",
          8306 => x"08",
          8307 => x"dc",
          8308 => x"38",
          8309 => x"51",
          8310 => x"82",
          8311 => x"57",
          8312 => x"08",
          8313 => x"bb",
          8314 => x"bb",
          8315 => x"5b",
          8316 => x"18",
          8317 => x"18",
          8318 => x"74",
          8319 => x"81",
          8320 => x"78",
          8321 => x"8b",
          8322 => x"54",
          8323 => x"75",
          8324 => x"38",
          8325 => x"1b",
          8326 => x"55",
          8327 => x"2e",
          8328 => x"39",
          8329 => x"09",
          8330 => x"38",
          8331 => x"80",
          8332 => x"70",
          8333 => x"25",
          8334 => x"80",
          8335 => x"38",
          8336 => x"bc",
          8337 => x"11",
          8338 => x"ff",
          8339 => x"82",
          8340 => x"57",
          8341 => x"08",
          8342 => x"70",
          8343 => x"80",
          8344 => x"83",
          8345 => x"80",
          8346 => x"84",
          8347 => x"a7",
          8348 => x"b4",
          8349 => x"ad",
          8350 => x"bb",
          8351 => x"0c",
          8352 => x"dc",
          8353 => x"0d",
          8354 => x"0d",
          8355 => x"3d",
          8356 => x"52",
          8357 => x"ce",
          8358 => x"bb",
          8359 => x"bb",
          8360 => x"54",
          8361 => x"08",
          8362 => x"8b",
          8363 => x"8b",
          8364 => x"59",
          8365 => x"3f",
          8366 => x"33",
          8367 => x"06",
          8368 => x"57",
          8369 => x"81",
          8370 => x"58",
          8371 => x"06",
          8372 => x"4e",
          8373 => x"ff",
          8374 => x"82",
          8375 => x"80",
          8376 => x"6c",
          8377 => x"53",
          8378 => x"ae",
          8379 => x"bb",
          8380 => x"2e",
          8381 => x"88",
          8382 => x"6d",
          8383 => x"55",
          8384 => x"bb",
          8385 => x"ff",
          8386 => x"83",
          8387 => x"51",
          8388 => x"26",
          8389 => x"15",
          8390 => x"ff",
          8391 => x"80",
          8392 => x"87",
          8393 => x"a4",
          8394 => x"74",
          8395 => x"38",
          8396 => x"b6",
          8397 => x"ae",
          8398 => x"bb",
          8399 => x"38",
          8400 => x"27",
          8401 => x"89",
          8402 => x"8b",
          8403 => x"27",
          8404 => x"55",
          8405 => x"81",
          8406 => x"8f",
          8407 => x"2a",
          8408 => x"70",
          8409 => x"34",
          8410 => x"74",
          8411 => x"05",
          8412 => x"17",
          8413 => x"70",
          8414 => x"52",
          8415 => x"73",
          8416 => x"c8",
          8417 => x"33",
          8418 => x"73",
          8419 => x"81",
          8420 => x"80",
          8421 => x"02",
          8422 => x"76",
          8423 => x"51",
          8424 => x"2e",
          8425 => x"87",
          8426 => x"57",
          8427 => x"79",
          8428 => x"80",
          8429 => x"70",
          8430 => x"ba",
          8431 => x"bb",
          8432 => x"82",
          8433 => x"80",
          8434 => x"52",
          8435 => x"bf",
          8436 => x"bb",
          8437 => x"82",
          8438 => x"8d",
          8439 => x"c4",
          8440 => x"e5",
          8441 => x"c6",
          8442 => x"dc",
          8443 => x"09",
          8444 => x"cc",
          8445 => x"76",
          8446 => x"c4",
          8447 => x"74",
          8448 => x"b0",
          8449 => x"dc",
          8450 => x"bb",
          8451 => x"38",
          8452 => x"bb",
          8453 => x"67",
          8454 => x"db",
          8455 => x"88",
          8456 => x"34",
          8457 => x"52",
          8458 => x"ab",
          8459 => x"54",
          8460 => x"15",
          8461 => x"ff",
          8462 => x"82",
          8463 => x"54",
          8464 => x"82",
          8465 => x"9c",
          8466 => x"f2",
          8467 => x"62",
          8468 => x"80",
          8469 => x"93",
          8470 => x"55",
          8471 => x"5e",
          8472 => x"3f",
          8473 => x"08",
          8474 => x"dc",
          8475 => x"38",
          8476 => x"58",
          8477 => x"38",
          8478 => x"97",
          8479 => x"08",
          8480 => x"38",
          8481 => x"70",
          8482 => x"81",
          8483 => x"55",
          8484 => x"87",
          8485 => x"39",
          8486 => x"90",
          8487 => x"82",
          8488 => x"8a",
          8489 => x"89",
          8490 => x"7f",
          8491 => x"56",
          8492 => x"3f",
          8493 => x"06",
          8494 => x"72",
          8495 => x"82",
          8496 => x"05",
          8497 => x"7c",
          8498 => x"55",
          8499 => x"27",
          8500 => x"16",
          8501 => x"83",
          8502 => x"76",
          8503 => x"80",
          8504 => x"79",
          8505 => x"99",
          8506 => x"7f",
          8507 => x"14",
          8508 => x"83",
          8509 => x"82",
          8510 => x"81",
          8511 => x"38",
          8512 => x"08",
          8513 => x"95",
          8514 => x"dc",
          8515 => x"81",
          8516 => x"7b",
          8517 => x"06",
          8518 => x"39",
          8519 => x"56",
          8520 => x"09",
          8521 => x"b9",
          8522 => x"80",
          8523 => x"80",
          8524 => x"78",
          8525 => x"7a",
          8526 => x"38",
          8527 => x"73",
          8528 => x"81",
          8529 => x"ff",
          8530 => x"74",
          8531 => x"ff",
          8532 => x"82",
          8533 => x"58",
          8534 => x"08",
          8535 => x"74",
          8536 => x"16",
          8537 => x"73",
          8538 => x"39",
          8539 => x"7e",
          8540 => x"0c",
          8541 => x"2e",
          8542 => x"88",
          8543 => x"8c",
          8544 => x"1a",
          8545 => x"07",
          8546 => x"1b",
          8547 => x"08",
          8548 => x"16",
          8549 => x"75",
          8550 => x"38",
          8551 => x"90",
          8552 => x"15",
          8553 => x"54",
          8554 => x"34",
          8555 => x"82",
          8556 => x"90",
          8557 => x"e9",
          8558 => x"6d",
          8559 => x"80",
          8560 => x"9d",
          8561 => x"5c",
          8562 => x"3f",
          8563 => x"0b",
          8564 => x"08",
          8565 => x"38",
          8566 => x"08",
          8567 => x"d3",
          8568 => x"08",
          8569 => x"80",
          8570 => x"80",
          8571 => x"bb",
          8572 => x"ff",
          8573 => x"52",
          8574 => x"a0",
          8575 => x"bb",
          8576 => x"ff",
          8577 => x"06",
          8578 => x"56",
          8579 => x"38",
          8580 => x"70",
          8581 => x"55",
          8582 => x"8b",
          8583 => x"3d",
          8584 => x"83",
          8585 => x"ff",
          8586 => x"82",
          8587 => x"99",
          8588 => x"74",
          8589 => x"38",
          8590 => x"80",
          8591 => x"ff",
          8592 => x"55",
          8593 => x"83",
          8594 => x"78",
          8595 => x"38",
          8596 => x"26",
          8597 => x"81",
          8598 => x"8b",
          8599 => x"79",
          8600 => x"80",
          8601 => x"93",
          8602 => x"39",
          8603 => x"6e",
          8604 => x"89",
          8605 => x"48",
          8606 => x"83",
          8607 => x"61",
          8608 => x"25",
          8609 => x"55",
          8610 => x"8a",
          8611 => x"3d",
          8612 => x"81",
          8613 => x"ff",
          8614 => x"81",
          8615 => x"dc",
          8616 => x"38",
          8617 => x"70",
          8618 => x"bb",
          8619 => x"56",
          8620 => x"38",
          8621 => x"55",
          8622 => x"75",
          8623 => x"38",
          8624 => x"70",
          8625 => x"ff",
          8626 => x"83",
          8627 => x"78",
          8628 => x"89",
          8629 => x"81",
          8630 => x"06",
          8631 => x"80",
          8632 => x"77",
          8633 => x"74",
          8634 => x"8d",
          8635 => x"06",
          8636 => x"2e",
          8637 => x"77",
          8638 => x"93",
          8639 => x"74",
          8640 => x"cb",
          8641 => x"7d",
          8642 => x"81",
          8643 => x"38",
          8644 => x"66",
          8645 => x"81",
          8646 => x"c8",
          8647 => x"74",
          8648 => x"38",
          8649 => x"98",
          8650 => x"c8",
          8651 => x"82",
          8652 => x"57",
          8653 => x"80",
          8654 => x"76",
          8655 => x"38",
          8656 => x"51",
          8657 => x"3f",
          8658 => x"08",
          8659 => x"87",
          8660 => x"2a",
          8661 => x"5c",
          8662 => x"bb",
          8663 => x"80",
          8664 => x"44",
          8665 => x"0a",
          8666 => x"ec",
          8667 => x"39",
          8668 => x"66",
          8669 => x"81",
          8670 => x"b8",
          8671 => x"74",
          8672 => x"38",
          8673 => x"98",
          8674 => x"b8",
          8675 => x"82",
          8676 => x"57",
          8677 => x"80",
          8678 => x"76",
          8679 => x"38",
          8680 => x"51",
          8681 => x"3f",
          8682 => x"08",
          8683 => x"57",
          8684 => x"08",
          8685 => x"96",
          8686 => x"82",
          8687 => x"10",
          8688 => x"08",
          8689 => x"72",
          8690 => x"59",
          8691 => x"ff",
          8692 => x"5d",
          8693 => x"44",
          8694 => x"11",
          8695 => x"70",
          8696 => x"71",
          8697 => x"06",
          8698 => x"52",
          8699 => x"40",
          8700 => x"09",
          8701 => x"38",
          8702 => x"18",
          8703 => x"39",
          8704 => x"79",
          8705 => x"70",
          8706 => x"58",
          8707 => x"76",
          8708 => x"38",
          8709 => x"7d",
          8710 => x"70",
          8711 => x"55",
          8712 => x"3f",
          8713 => x"08",
          8714 => x"2e",
          8715 => x"9b",
          8716 => x"dc",
          8717 => x"f5",
          8718 => x"38",
          8719 => x"38",
          8720 => x"59",
          8721 => x"38",
          8722 => x"7d",
          8723 => x"81",
          8724 => x"38",
          8725 => x"0b",
          8726 => x"08",
          8727 => x"78",
          8728 => x"1a",
          8729 => x"c0",
          8730 => x"74",
          8731 => x"39",
          8732 => x"55",
          8733 => x"8f",
          8734 => x"fd",
          8735 => x"bb",
          8736 => x"f5",
          8737 => x"78",
          8738 => x"79",
          8739 => x"80",
          8740 => x"f1",
          8741 => x"39",
          8742 => x"81",
          8743 => x"06",
          8744 => x"55",
          8745 => x"27",
          8746 => x"81",
          8747 => x"56",
          8748 => x"38",
          8749 => x"80",
          8750 => x"ff",
          8751 => x"8b",
          8752 => x"e0",
          8753 => x"ff",
          8754 => x"84",
          8755 => x"1b",
          8756 => x"b3",
          8757 => x"1c",
          8758 => x"ff",
          8759 => x"8e",
          8760 => x"a1",
          8761 => x"0b",
          8762 => x"7d",
          8763 => x"30",
          8764 => x"84",
          8765 => x"51",
          8766 => x"51",
          8767 => x"3f",
          8768 => x"83",
          8769 => x"90",
          8770 => x"ff",
          8771 => x"93",
          8772 => x"a0",
          8773 => x"39",
          8774 => x"1b",
          8775 => x"85",
          8776 => x"95",
          8777 => x"52",
          8778 => x"ff",
          8779 => x"81",
          8780 => x"1b",
          8781 => x"cf",
          8782 => x"9c",
          8783 => x"a0",
          8784 => x"83",
          8785 => x"06",
          8786 => x"82",
          8787 => x"52",
          8788 => x"51",
          8789 => x"3f",
          8790 => x"1b",
          8791 => x"c5",
          8792 => x"ac",
          8793 => x"a0",
          8794 => x"52",
          8795 => x"ff",
          8796 => x"86",
          8797 => x"51",
          8798 => x"3f",
          8799 => x"80",
          8800 => x"a9",
          8801 => x"1c",
          8802 => x"82",
          8803 => x"80",
          8804 => x"ae",
          8805 => x"b2",
          8806 => x"1b",
          8807 => x"85",
          8808 => x"ff",
          8809 => x"96",
          8810 => x"9f",
          8811 => x"80",
          8812 => x"34",
          8813 => x"1c",
          8814 => x"82",
          8815 => x"ab",
          8816 => x"a0",
          8817 => x"d4",
          8818 => x"fe",
          8819 => x"59",
          8820 => x"3f",
          8821 => x"53",
          8822 => x"51",
          8823 => x"3f",
          8824 => x"bb",
          8825 => x"e7",
          8826 => x"2e",
          8827 => x"80",
          8828 => x"54",
          8829 => x"53",
          8830 => x"51",
          8831 => x"3f",
          8832 => x"80",
          8833 => x"ff",
          8834 => x"84",
          8835 => x"d2",
          8836 => x"ff",
          8837 => x"86",
          8838 => x"f2",
          8839 => x"1b",
          8840 => x"81",
          8841 => x"52",
          8842 => x"51",
          8843 => x"3f",
          8844 => x"ec",
          8845 => x"9e",
          8846 => x"d4",
          8847 => x"51",
          8848 => x"3f",
          8849 => x"87",
          8850 => x"52",
          8851 => x"9a",
          8852 => x"54",
          8853 => x"7a",
          8854 => x"ff",
          8855 => x"65",
          8856 => x"7a",
          8857 => x"8f",
          8858 => x"80",
          8859 => x"2e",
          8860 => x"9a",
          8861 => x"7a",
          8862 => x"a9",
          8863 => x"84",
          8864 => x"9e",
          8865 => x"0a",
          8866 => x"51",
          8867 => x"ff",
          8868 => x"7d",
          8869 => x"38",
          8870 => x"52",
          8871 => x"9e",
          8872 => x"55",
          8873 => x"62",
          8874 => x"74",
          8875 => x"75",
          8876 => x"7e",
          8877 => x"fe",
          8878 => x"dc",
          8879 => x"38",
          8880 => x"82",
          8881 => x"52",
          8882 => x"9e",
          8883 => x"16",
          8884 => x"56",
          8885 => x"38",
          8886 => x"77",
          8887 => x"8d",
          8888 => x"7d",
          8889 => x"38",
          8890 => x"57",
          8891 => x"83",
          8892 => x"76",
          8893 => x"7a",
          8894 => x"ff",
          8895 => x"82",
          8896 => x"81",
          8897 => x"16",
          8898 => x"56",
          8899 => x"38",
          8900 => x"83",
          8901 => x"86",
          8902 => x"ff",
          8903 => x"38",
          8904 => x"82",
          8905 => x"81",
          8906 => x"06",
          8907 => x"fe",
          8908 => x"53",
          8909 => x"51",
          8910 => x"3f",
          8911 => x"52",
          8912 => x"9c",
          8913 => x"be",
          8914 => x"75",
          8915 => x"81",
          8916 => x"0b",
          8917 => x"77",
          8918 => x"75",
          8919 => x"60",
          8920 => x"80",
          8921 => x"75",
          8922 => x"99",
          8923 => x"85",
          8924 => x"bb",
          8925 => x"2a",
          8926 => x"75",
          8927 => x"82",
          8928 => x"87",
          8929 => x"52",
          8930 => x"51",
          8931 => x"3f",
          8932 => x"ca",
          8933 => x"9c",
          8934 => x"54",
          8935 => x"52",
          8936 => x"98",
          8937 => x"56",
          8938 => x"08",
          8939 => x"53",
          8940 => x"51",
          8941 => x"3f",
          8942 => x"bb",
          8943 => x"38",
          8944 => x"56",
          8945 => x"56",
          8946 => x"bb",
          8947 => x"75",
          8948 => x"0c",
          8949 => x"04",
          8950 => x"7d",
          8951 => x"80",
          8952 => x"05",
          8953 => x"76",
          8954 => x"38",
          8955 => x"11",
          8956 => x"53",
          8957 => x"79",
          8958 => x"3f",
          8959 => x"09",
          8960 => x"38",
          8961 => x"55",
          8962 => x"db",
          8963 => x"70",
          8964 => x"34",
          8965 => x"74",
          8966 => x"81",
          8967 => x"80",
          8968 => x"55",
          8969 => x"76",
          8970 => x"bb",
          8971 => x"3d",
          8972 => x"3d",
          8973 => x"84",
          8974 => x"33",
          8975 => x"8a",
          8976 => x"06",
          8977 => x"52",
          8978 => x"3f",
          8979 => x"56",
          8980 => x"be",
          8981 => x"08",
          8982 => x"05",
          8983 => x"75",
          8984 => x"56",
          8985 => x"a1",
          8986 => x"fc",
          8987 => x"53",
          8988 => x"76",
          8989 => x"dc",
          8990 => x"32",
          8991 => x"72",
          8992 => x"70",
          8993 => x"56",
          8994 => x"18",
          8995 => x"88",
          8996 => x"3d",
          8997 => x"3d",
          8998 => x"11",
          8999 => x"80",
          9000 => x"38",
          9001 => x"05",
          9002 => x"8c",
          9003 => x"08",
          9004 => x"3f",
          9005 => x"08",
          9006 => x"16",
          9007 => x"09",
          9008 => x"38",
          9009 => x"55",
          9010 => x"55",
          9011 => x"dc",
          9012 => x"0d",
          9013 => x"0d",
          9014 => x"cc",
          9015 => x"73",
          9016 => x"93",
          9017 => x"0c",
          9018 => x"04",
          9019 => x"02",
          9020 => x"33",
          9021 => x"3d",
          9022 => x"54",
          9023 => x"52",
          9024 => x"ae",
          9025 => x"ff",
          9026 => x"3d",
          9027 => x"ff",
          9028 => x"00",
          9029 => x"ff",
          9030 => x"ff",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"00",
          9136 => x"00",
          9137 => x"00",
          9138 => x"00",
          9139 => x"00",
          9140 => x"00",
          9141 => x"00",
          9142 => x"00",
          9143 => x"00",
          9144 => x"00",
          9145 => x"00",
          9146 => x"00",
          9147 => x"00",
          9148 => x"00",
          9149 => x"00",
          9150 => x"00",
          9151 => x"00",
          9152 => x"00",
          9153 => x"00",
          9154 => x"00",
          9155 => x"00",
          9156 => x"00",
          9157 => x"00",
          9158 => x"00",
          9159 => x"00",
          9160 => x"00",
          9161 => x"00",
          9162 => x"00",
          9163 => x"00",
          9164 => x"00",
          9165 => x"00",
          9166 => x"00",
          9167 => x"69",
          9168 => x"00",
          9169 => x"69",
          9170 => x"6c",
          9171 => x"69",
          9172 => x"00",
          9173 => x"6c",
          9174 => x"00",
          9175 => x"65",
          9176 => x"00",
          9177 => x"63",
          9178 => x"72",
          9179 => x"63",
          9180 => x"00",
          9181 => x"64",
          9182 => x"00",
          9183 => x"64",
          9184 => x"00",
          9185 => x"65",
          9186 => x"65",
          9187 => x"65",
          9188 => x"69",
          9189 => x"69",
          9190 => x"66",
          9191 => x"66",
          9192 => x"61",
          9193 => x"00",
          9194 => x"6d",
          9195 => x"65",
          9196 => x"72",
          9197 => x"65",
          9198 => x"00",
          9199 => x"6e",
          9200 => x"00",
          9201 => x"65",
          9202 => x"00",
          9203 => x"62",
          9204 => x"63",
          9205 => x"62",
          9206 => x"63",
          9207 => x"69",
          9208 => x"00",
          9209 => x"64",
          9210 => x"69",
          9211 => x"45",
          9212 => x"72",
          9213 => x"6e",
          9214 => x"6e",
          9215 => x"65",
          9216 => x"72",
          9217 => x"69",
          9218 => x"6e",
          9219 => x"72",
          9220 => x"79",
          9221 => x"6f",
          9222 => x"6c",
          9223 => x"6f",
          9224 => x"2e",
          9225 => x"6f",
          9226 => x"74",
          9227 => x"6f",
          9228 => x"2e",
          9229 => x"6e",
          9230 => x"69",
          9231 => x"69",
          9232 => x"61",
          9233 => x"00",
          9234 => x"63",
          9235 => x"73",
          9236 => x"6e",
          9237 => x"2e",
          9238 => x"69",
          9239 => x"61",
          9240 => x"61",
          9241 => x"65",
          9242 => x"74",
          9243 => x"00",
          9244 => x"69",
          9245 => x"68",
          9246 => x"6c",
          9247 => x"6e",
          9248 => x"69",
          9249 => x"00",
          9250 => x"44",
          9251 => x"20",
          9252 => x"74",
          9253 => x"72",
          9254 => x"63",
          9255 => x"2e",
          9256 => x"72",
          9257 => x"20",
          9258 => x"62",
          9259 => x"69",
          9260 => x"6e",
          9261 => x"69",
          9262 => x"00",
          9263 => x"69",
          9264 => x"6e",
          9265 => x"65",
          9266 => x"6c",
          9267 => x"00",
          9268 => x"6f",
          9269 => x"6d",
          9270 => x"69",
          9271 => x"20",
          9272 => x"65",
          9273 => x"74",
          9274 => x"66",
          9275 => x"64",
          9276 => x"20",
          9277 => x"6b",
          9278 => x"6f",
          9279 => x"74",
          9280 => x"6f",
          9281 => x"64",
          9282 => x"69",
          9283 => x"75",
          9284 => x"6f",
          9285 => x"61",
          9286 => x"6e",
          9287 => x"6e",
          9288 => x"6c",
          9289 => x"00",
          9290 => x"69",
          9291 => x"69",
          9292 => x"6f",
          9293 => x"64",
          9294 => x"6e",
          9295 => x"66",
          9296 => x"65",
          9297 => x"6d",
          9298 => x"72",
          9299 => x"00",
          9300 => x"6f",
          9301 => x"61",
          9302 => x"6f",
          9303 => x"20",
          9304 => x"65",
          9305 => x"00",
          9306 => x"61",
          9307 => x"65",
          9308 => x"73",
          9309 => x"63",
          9310 => x"65",
          9311 => x"00",
          9312 => x"75",
          9313 => x"73",
          9314 => x"00",
          9315 => x"6e",
          9316 => x"77",
          9317 => x"72",
          9318 => x"2e",
          9319 => x"25",
          9320 => x"62",
          9321 => x"73",
          9322 => x"20",
          9323 => x"25",
          9324 => x"62",
          9325 => x"73",
          9326 => x"63",
          9327 => x"00",
          9328 => x"65",
          9329 => x"00",
          9330 => x"30",
          9331 => x"00",
          9332 => x"20",
          9333 => x"30",
          9334 => x"00",
          9335 => x"20",
          9336 => x"20",
          9337 => x"00",
          9338 => x"30",
          9339 => x"00",
          9340 => x"20",
          9341 => x"7c",
          9342 => x"00",
          9343 => x"50",
          9344 => x"00",
          9345 => x"2a",
          9346 => x"73",
          9347 => x"00",
          9348 => x"32",
          9349 => x"2f",
          9350 => x"30",
          9351 => x"31",
          9352 => x"00",
          9353 => x"5a",
          9354 => x"20",
          9355 => x"20",
          9356 => x"78",
          9357 => x"73",
          9358 => x"20",
          9359 => x"0a",
          9360 => x"50",
          9361 => x"20",
          9362 => x"65",
          9363 => x"70",
          9364 => x"61",
          9365 => x"65",
          9366 => x"69",
          9367 => x"20",
          9368 => x"65",
          9369 => x"70",
          9370 => x"53",
          9371 => x"6e",
          9372 => x"72",
          9373 => x"00",
          9374 => x"4f",
          9375 => x"20",
          9376 => x"69",
          9377 => x"72",
          9378 => x"74",
          9379 => x"4f",
          9380 => x"20",
          9381 => x"69",
          9382 => x"72",
          9383 => x"74",
          9384 => x"41",
          9385 => x"20",
          9386 => x"69",
          9387 => x"72",
          9388 => x"74",
          9389 => x"41",
          9390 => x"20",
          9391 => x"69",
          9392 => x"72",
          9393 => x"74",
          9394 => x"41",
          9395 => x"20",
          9396 => x"69",
          9397 => x"72",
          9398 => x"74",
          9399 => x"41",
          9400 => x"20",
          9401 => x"69",
          9402 => x"72",
          9403 => x"74",
          9404 => x"65",
          9405 => x"6e",
          9406 => x"70",
          9407 => x"6d",
          9408 => x"2e",
          9409 => x"6e",
          9410 => x"69",
          9411 => x"74",
          9412 => x"72",
          9413 => x"00",
          9414 => x"75",
          9415 => x"78",
          9416 => x"62",
          9417 => x"00",
          9418 => x"70",
          9419 => x"2e",
          9420 => x"00",
          9421 => x"3a",
          9422 => x"61",
          9423 => x"64",
          9424 => x"20",
          9425 => x"74",
          9426 => x"69",
          9427 => x"73",
          9428 => x"61",
          9429 => x"30",
          9430 => x"6c",
          9431 => x"65",
          9432 => x"69",
          9433 => x"61",
          9434 => x"6c",
          9435 => x"00",
          9436 => x"20",
          9437 => x"61",
          9438 => x"69",
          9439 => x"69",
          9440 => x"00",
          9441 => x"6e",
          9442 => x"61",
          9443 => x"65",
          9444 => x"00",
          9445 => x"61",
          9446 => x"64",
          9447 => x"20",
          9448 => x"74",
          9449 => x"69",
          9450 => x"00",
          9451 => x"63",
          9452 => x"0a",
          9453 => x"75",
          9454 => x"6c",
          9455 => x"69",
          9456 => x"2e",
          9457 => x"00",
          9458 => x"6f",
          9459 => x"6e",
          9460 => x"2e",
          9461 => x"6f",
          9462 => x"72",
          9463 => x"2e",
          9464 => x"00",
          9465 => x"30",
          9466 => x"28",
          9467 => x"78",
          9468 => x"25",
          9469 => x"78",
          9470 => x"38",
          9471 => x"00",
          9472 => x"75",
          9473 => x"4d",
          9474 => x"72",
          9475 => x"43",
          9476 => x"6c",
          9477 => x"2e",
          9478 => x"30",
          9479 => x"20",
          9480 => x"58",
          9481 => x"3f",
          9482 => x"30",
          9483 => x"20",
          9484 => x"58",
          9485 => x"30",
          9486 => x"20",
          9487 => x"6c",
          9488 => x"00",
          9489 => x"69",
          9490 => x"6c",
          9491 => x"20",
          9492 => x"65",
          9493 => x"70",
          9494 => x"00",
          9495 => x"6e",
          9496 => x"69",
          9497 => x"69",
          9498 => x"72",
          9499 => x"74",
          9500 => x"69",
          9501 => x"6c",
          9502 => x"75",
          9503 => x"20",
          9504 => x"6f",
          9505 => x"6e",
          9506 => x"69",
          9507 => x"75",
          9508 => x"20",
          9509 => x"6f",
          9510 => x"78",
          9511 => x"74",
          9512 => x"20",
          9513 => x"65",
          9514 => x"25",
          9515 => x"78",
          9516 => x"2e",
          9517 => x"61",
          9518 => x"6e",
          9519 => x"6f",
          9520 => x"40",
          9521 => x"38",
          9522 => x"2e",
          9523 => x"00",
          9524 => x"61",
          9525 => x"72",
          9526 => x"72",
          9527 => x"20",
          9528 => x"65",
          9529 => x"64",
          9530 => x"00",
          9531 => x"65",
          9532 => x"72",
          9533 => x"67",
          9534 => x"70",
          9535 => x"61",
          9536 => x"6e",
          9537 => x"00",
          9538 => x"6f",
          9539 => x"72",
          9540 => x"6f",
          9541 => x"67",
          9542 => x"00",
          9543 => x"50",
          9544 => x"69",
          9545 => x"64",
          9546 => x"73",
          9547 => x"2e",
          9548 => x"00",
          9549 => x"64",
          9550 => x"73",
          9551 => x"00",
          9552 => x"64",
          9553 => x"73",
          9554 => x"61",
          9555 => x"6f",
          9556 => x"6e",
          9557 => x"00",
          9558 => x"75",
          9559 => x"6e",
          9560 => x"2e",
          9561 => x"6e",
          9562 => x"69",
          9563 => x"69",
          9564 => x"72",
          9565 => x"74",
          9566 => x"2e",
          9567 => x"64",
          9568 => x"2f",
          9569 => x"25",
          9570 => x"64",
          9571 => x"2e",
          9572 => x"64",
          9573 => x"6f",
          9574 => x"6f",
          9575 => x"67",
          9576 => x"74",
          9577 => x"00",
          9578 => x"28",
          9579 => x"6d",
          9580 => x"43",
          9581 => x"6e",
          9582 => x"29",
          9583 => x"0a",
          9584 => x"69",
          9585 => x"20",
          9586 => x"6c",
          9587 => x"6e",
          9588 => x"3a",
          9589 => x"20",
          9590 => x"42",
          9591 => x"52",
          9592 => x"20",
          9593 => x"38",
          9594 => x"30",
          9595 => x"2e",
          9596 => x"20",
          9597 => x"44",
          9598 => x"20",
          9599 => x"20",
          9600 => x"38",
          9601 => x"30",
          9602 => x"2e",
          9603 => x"20",
          9604 => x"4e",
          9605 => x"42",
          9606 => x"20",
          9607 => x"38",
          9608 => x"30",
          9609 => x"2e",
          9610 => x"20",
          9611 => x"52",
          9612 => x"20",
          9613 => x"20",
          9614 => x"38",
          9615 => x"30",
          9616 => x"2e",
          9617 => x"20",
          9618 => x"41",
          9619 => x"20",
          9620 => x"20",
          9621 => x"38",
          9622 => x"30",
          9623 => x"2e",
          9624 => x"20",
          9625 => x"44",
          9626 => x"52",
          9627 => x"20",
          9628 => x"76",
          9629 => x"73",
          9630 => x"30",
          9631 => x"2e",
          9632 => x"20",
          9633 => x"49",
          9634 => x"31",
          9635 => x"20",
          9636 => x"6d",
          9637 => x"20",
          9638 => x"30",
          9639 => x"2e",
          9640 => x"20",
          9641 => x"4e",
          9642 => x"43",
          9643 => x"20",
          9644 => x"61",
          9645 => x"6c",
          9646 => x"30",
          9647 => x"2e",
          9648 => x"20",
          9649 => x"49",
          9650 => x"4f",
          9651 => x"42",
          9652 => x"00",
          9653 => x"20",
          9654 => x"42",
          9655 => x"43",
          9656 => x"20",
          9657 => x"4f",
          9658 => x"0a",
          9659 => x"20",
          9660 => x"53",
          9661 => x"00",
          9662 => x"20",
          9663 => x"50",
          9664 => x"00",
          9665 => x"64",
          9666 => x"73",
          9667 => x"3a",
          9668 => x"20",
          9669 => x"50",
          9670 => x"65",
          9671 => x"20",
          9672 => x"74",
          9673 => x"41",
          9674 => x"65",
          9675 => x"3d",
          9676 => x"38",
          9677 => x"00",
          9678 => x"20",
          9679 => x"50",
          9680 => x"65",
          9681 => x"79",
          9682 => x"61",
          9683 => x"41",
          9684 => x"65",
          9685 => x"3d",
          9686 => x"38",
          9687 => x"00",
          9688 => x"20",
          9689 => x"74",
          9690 => x"20",
          9691 => x"72",
          9692 => x"64",
          9693 => x"73",
          9694 => x"20",
          9695 => x"3d",
          9696 => x"38",
          9697 => x"00",
          9698 => x"69",
          9699 => x"0a",
          9700 => x"20",
          9701 => x"50",
          9702 => x"64",
          9703 => x"20",
          9704 => x"20",
          9705 => x"20",
          9706 => x"20",
          9707 => x"3d",
          9708 => x"34",
          9709 => x"00",
          9710 => x"20",
          9711 => x"79",
          9712 => x"6d",
          9713 => x"6f",
          9714 => x"46",
          9715 => x"20",
          9716 => x"20",
          9717 => x"3d",
          9718 => x"2e",
          9719 => x"64",
          9720 => x"0a",
          9721 => x"20",
          9722 => x"44",
          9723 => x"20",
          9724 => x"63",
          9725 => x"72",
          9726 => x"20",
          9727 => x"20",
          9728 => x"3d",
          9729 => x"2e",
          9730 => x"64",
          9731 => x"0a",
          9732 => x"20",
          9733 => x"69",
          9734 => x"6f",
          9735 => x"53",
          9736 => x"4d",
          9737 => x"6f",
          9738 => x"46",
          9739 => x"3d",
          9740 => x"2e",
          9741 => x"64",
          9742 => x"0a",
          9743 => x"6d",
          9744 => x"00",
          9745 => x"65",
          9746 => x"6d",
          9747 => x"6c",
          9748 => x"00",
          9749 => x"56",
          9750 => x"56",
          9751 => x"6e",
          9752 => x"6e",
          9753 => x"77",
          9754 => x"00",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"00",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"00",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"00",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"00",
          9788 => x"00",
          9789 => x"00",
          9790 => x"00",
          9791 => x"00",
          9792 => x"00",
          9793 => x"00",
          9794 => x"00",
          9795 => x"00",
          9796 => x"00",
          9797 => x"00",
          9798 => x"00",
          9799 => x"00",
          9800 => x"00",
          9801 => x"00",
          9802 => x"00",
          9803 => x"00",
          9804 => x"00",
          9805 => x"00",
          9806 => x"00",
          9807 => x"00",
          9808 => x"00",
          9809 => x"00",
          9810 => x"00",
          9811 => x"00",
          9812 => x"00",
          9813 => x"00",
          9814 => x"00",
          9815 => x"00",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"00",
          9820 => x"5b",
          9821 => x"5b",
          9822 => x"5b",
          9823 => x"5b",
          9824 => x"5b",
          9825 => x"5b",
          9826 => x"5b",
          9827 => x"30",
          9828 => x"5b",
          9829 => x"5b",
          9830 => x"5b",
          9831 => x"00",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"00",
          9836 => x"00",
          9837 => x"00",
          9838 => x"00",
          9839 => x"00",
          9840 => x"00",
          9841 => x"00",
          9842 => x"69",
          9843 => x"72",
          9844 => x"69",
          9845 => x"00",
          9846 => x"00",
          9847 => x"30",
          9848 => x"20",
          9849 => x"0a",
          9850 => x"61",
          9851 => x"64",
          9852 => x"20",
          9853 => x"65",
          9854 => x"68",
          9855 => x"69",
          9856 => x"72",
          9857 => x"69",
          9858 => x"74",
          9859 => x"4f",
          9860 => x"00",
          9861 => x"61",
          9862 => x"74",
          9863 => x"65",
          9864 => x"72",
          9865 => x"65",
          9866 => x"73",
          9867 => x"79",
          9868 => x"6c",
          9869 => x"64",
          9870 => x"62",
          9871 => x"67",
          9872 => x"44",
          9873 => x"2a",
          9874 => x"3b",
          9875 => x"3f",
          9876 => x"7f",
          9877 => x"41",
          9878 => x"41",
          9879 => x"00",
          9880 => x"fe",
          9881 => x"44",
          9882 => x"2e",
          9883 => x"4f",
          9884 => x"4d",
          9885 => x"20",
          9886 => x"54",
          9887 => x"20",
          9888 => x"4f",
          9889 => x"4d",
          9890 => x"20",
          9891 => x"54",
          9892 => x"20",
          9893 => x"00",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"9a",
          9898 => x"41",
          9899 => x"45",
          9900 => x"49",
          9901 => x"92",
          9902 => x"4f",
          9903 => x"99",
          9904 => x"9d",
          9905 => x"49",
          9906 => x"a5",
          9907 => x"a9",
          9908 => x"ad",
          9909 => x"b1",
          9910 => x"b5",
          9911 => x"b9",
          9912 => x"bd",
          9913 => x"c1",
          9914 => x"c5",
          9915 => x"c9",
          9916 => x"cd",
          9917 => x"d1",
          9918 => x"d5",
          9919 => x"d9",
          9920 => x"dd",
          9921 => x"e1",
          9922 => x"e5",
          9923 => x"e9",
          9924 => x"ed",
          9925 => x"f1",
          9926 => x"f5",
          9927 => x"f9",
          9928 => x"fd",
          9929 => x"2e",
          9930 => x"5b",
          9931 => x"22",
          9932 => x"3e",
          9933 => x"00",
          9934 => x"01",
          9935 => x"10",
          9936 => x"00",
          9937 => x"00",
          9938 => x"01",
          9939 => x"04",
          9940 => x"10",
          9941 => x"00",
          9942 => x"00",
          9943 => x"00",
          9944 => x"02",
          9945 => x"00",
          9946 => x"00",
          9947 => x"00",
          9948 => x"04",
          9949 => x"00",
          9950 => x"00",
          9951 => x"00",
          9952 => x"14",
          9953 => x"00",
          9954 => x"00",
          9955 => x"00",
          9956 => x"2b",
          9957 => x"00",
          9958 => x"00",
          9959 => x"00",
          9960 => x"30",
          9961 => x"00",
          9962 => x"00",
          9963 => x"00",
          9964 => x"3c",
          9965 => x"00",
          9966 => x"00",
          9967 => x"00",
          9968 => x"3d",
          9969 => x"00",
          9970 => x"00",
          9971 => x"00",
          9972 => x"3f",
          9973 => x"00",
          9974 => x"00",
          9975 => x"00",
          9976 => x"40",
          9977 => x"00",
          9978 => x"00",
          9979 => x"00",
          9980 => x"41",
          9981 => x"00",
          9982 => x"00",
          9983 => x"00",
          9984 => x"42",
          9985 => x"00",
          9986 => x"00",
          9987 => x"00",
          9988 => x"43",
          9989 => x"00",
          9990 => x"00",
          9991 => x"00",
          9992 => x"50",
          9993 => x"00",
          9994 => x"00",
          9995 => x"00",
          9996 => x"51",
          9997 => x"00",
          9998 => x"00",
          9999 => x"00",
         10000 => x"54",
         10001 => x"00",
         10002 => x"00",
         10003 => x"00",
         10004 => x"55",
         10005 => x"00",
         10006 => x"00",
         10007 => x"00",
         10008 => x"79",
         10009 => x"00",
         10010 => x"00",
         10011 => x"00",
         10012 => x"78",
         10013 => x"00",
         10014 => x"00",
         10015 => x"00",
         10016 => x"82",
         10017 => x"00",
         10018 => x"00",
         10019 => x"00",
         10020 => x"83",
         10021 => x"00",
         10022 => x"00",
         10023 => x"00",
         10024 => x"85",
         10025 => x"00",
         10026 => x"00",
         10027 => x"00",
         10028 => x"87",
         10029 => x"00",
         10030 => x"00",
         10031 => x"00",
         10032 => x"8c",
         10033 => x"00",
         10034 => x"00",
         10035 => x"00",
         10036 => x"8d",
         10037 => x"00",
         10038 => x"00",
         10039 => x"00",
         10040 => x"8e",
         10041 => x"00",
         10042 => x"00",
         10043 => x"00",
         10044 => x"8f",
         10045 => x"00",
         10046 => x"00",
         10047 => x"00",
         10048 => x"00",
         10049 => x"00",
         10050 => x"00",
         10051 => x"00",
         10052 => x"01",
         10053 => x"00",
         10054 => x"01",
         10055 => x"81",
         10056 => x"00",
         10057 => x"7f",
         10058 => x"00",
         10059 => x"00",
         10060 => x"00",
         10061 => x"00",
         10062 => x"f5",
         10063 => x"f5",
         10064 => x"f5",
         10065 => x"00",
         10066 => x"01",
         10067 => x"01",
         10068 => x"01",
         10069 => x"00",
         10070 => x"00",
         10071 => x"00",
         10072 => x"00",
         10073 => x"00",
         10074 => x"00",
         10075 => x"00",
         10076 => x"00",
         10077 => x"00",
         10078 => x"00",
         10079 => x"00",
         10080 => x"00",
         10081 => x"00",
         10082 => x"00",
         10083 => x"00",
         10084 => x"00",
         10085 => x"00",
         10086 => x"00",
         10087 => x"00",
         10088 => x"00",
         10089 => x"00",
         10090 => x"00",
         10091 => x"00",
         10092 => x"00",
         10093 => x"00",
         10094 => x"00",
         10095 => x"00",
         10096 => x"00",
         10097 => x"00",
         10098 => x"00",
         10099 => x"00",
         10100 => x"00",
         10101 => x"00",
         10102 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"9d",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"8c",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"f4",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"e0",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"95",
           269 => x"0b",
           270 => x"0b",
           271 => x"b3",
           272 => x"0b",
           273 => x"0b",
           274 => x"d1",
           275 => x"0b",
           276 => x"0b",
           277 => x"f0",
           278 => x"0b",
           279 => x"0b",
           280 => x"8f",
           281 => x"0b",
           282 => x"0b",
           283 => x"ad",
           284 => x"0b",
           285 => x"0b",
           286 => x"cd",
           287 => x"0b",
           288 => x"0b",
           289 => x"ed",
           290 => x"0b",
           291 => x"0b",
           292 => x"8d",
           293 => x"0b",
           294 => x"0b",
           295 => x"ad",
           296 => x"0b",
           297 => x"0b",
           298 => x"cd",
           299 => x"0b",
           300 => x"0b",
           301 => x"ed",
           302 => x"0b",
           303 => x"0b",
           304 => x"8d",
           305 => x"0b",
           306 => x"0b",
           307 => x"ad",
           308 => x"0b",
           309 => x"0b",
           310 => x"cd",
           311 => x"0b",
           312 => x"0b",
           313 => x"ed",
           314 => x"0b",
           315 => x"0b",
           316 => x"8d",
           317 => x"0b",
           318 => x"0b",
           319 => x"ad",
           320 => x"0b",
           321 => x"0b",
           322 => x"cd",
           323 => x"0b",
           324 => x"0b",
           325 => x"ed",
           326 => x"0b",
           327 => x"0b",
           328 => x"8d",
           329 => x"0b",
           330 => x"0b",
           331 => x"ad",
           332 => x"0b",
           333 => x"0b",
           334 => x"cd",
           335 => x"0b",
           336 => x"0b",
           337 => x"ed",
           338 => x"0b",
           339 => x"0b",
           340 => x"8d",
           341 => x"0b",
           342 => x"0b",
           343 => x"ad",
           344 => x"0b",
           345 => x"0b",
           346 => x"cd",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"04",
           390 => x"0c",
           391 => x"82",
           392 => x"82",
           393 => x"82",
           394 => x"af",
           395 => x"bb",
           396 => x"d8",
           397 => x"bb",
           398 => x"ad",
           399 => x"e8",
           400 => x"90",
           401 => x"e8",
           402 => x"2d",
           403 => x"08",
           404 => x"04",
           405 => x"0c",
           406 => x"82",
           407 => x"82",
           408 => x"82",
           409 => x"80",
           410 => x"82",
           411 => x"82",
           412 => x"82",
           413 => x"80",
           414 => x"82",
           415 => x"82",
           416 => x"82",
           417 => x"93",
           418 => x"bb",
           419 => x"d8",
           420 => x"bb",
           421 => x"c0",
           422 => x"e8",
           423 => x"90",
           424 => x"e8",
           425 => x"2d",
           426 => x"08",
           427 => x"04",
           428 => x"0c",
           429 => x"2d",
           430 => x"08",
           431 => x"04",
           432 => x"0c",
           433 => x"2d",
           434 => x"08",
           435 => x"04",
           436 => x"0c",
           437 => x"2d",
           438 => x"08",
           439 => x"04",
           440 => x"0c",
           441 => x"2d",
           442 => x"08",
           443 => x"04",
           444 => x"0c",
           445 => x"2d",
           446 => x"08",
           447 => x"04",
           448 => x"0c",
           449 => x"2d",
           450 => x"08",
           451 => x"04",
           452 => x"0c",
           453 => x"2d",
           454 => x"08",
           455 => x"04",
           456 => x"0c",
           457 => x"2d",
           458 => x"08",
           459 => x"04",
           460 => x"0c",
           461 => x"2d",
           462 => x"08",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"04",
           468 => x"0c",
           469 => x"2d",
           470 => x"08",
           471 => x"04",
           472 => x"0c",
           473 => x"2d",
           474 => x"08",
           475 => x"04",
           476 => x"0c",
           477 => x"2d",
           478 => x"08",
           479 => x"04",
           480 => x"0c",
           481 => x"2d",
           482 => x"08",
           483 => x"04",
           484 => x"0c",
           485 => x"2d",
           486 => x"08",
           487 => x"04",
           488 => x"0c",
           489 => x"2d",
           490 => x"08",
           491 => x"04",
           492 => x"0c",
           493 => x"2d",
           494 => x"08",
           495 => x"04",
           496 => x"0c",
           497 => x"2d",
           498 => x"08",
           499 => x"04",
           500 => x"0c",
           501 => x"2d",
           502 => x"08",
           503 => x"04",
           504 => x"0c",
           505 => x"2d",
           506 => x"08",
           507 => x"04",
           508 => x"0c",
           509 => x"2d",
           510 => x"08",
           511 => x"04",
           512 => x"0c",
           513 => x"2d",
           514 => x"08",
           515 => x"04",
           516 => x"0c",
           517 => x"2d",
           518 => x"08",
           519 => x"04",
           520 => x"0c",
           521 => x"2d",
           522 => x"08",
           523 => x"04",
           524 => x"0c",
           525 => x"2d",
           526 => x"08",
           527 => x"04",
           528 => x"0c",
           529 => x"2d",
           530 => x"08",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"04",
           536 => x"0c",
           537 => x"2d",
           538 => x"08",
           539 => x"04",
           540 => x"0c",
           541 => x"2d",
           542 => x"08",
           543 => x"04",
           544 => x"0c",
           545 => x"2d",
           546 => x"08",
           547 => x"04",
           548 => x"0c",
           549 => x"2d",
           550 => x"08",
           551 => x"04",
           552 => x"0c",
           553 => x"2d",
           554 => x"08",
           555 => x"04",
           556 => x"0c",
           557 => x"2d",
           558 => x"08",
           559 => x"04",
           560 => x"0c",
           561 => x"2d",
           562 => x"08",
           563 => x"04",
           564 => x"0c",
           565 => x"2d",
           566 => x"08",
           567 => x"04",
           568 => x"0c",
           569 => x"2d",
           570 => x"08",
           571 => x"04",
           572 => x"0c",
           573 => x"2d",
           574 => x"08",
           575 => x"04",
           576 => x"0c",
           577 => x"2d",
           578 => x"08",
           579 => x"04",
           580 => x"0c",
           581 => x"2d",
           582 => x"08",
           583 => x"04",
           584 => x"0c",
           585 => x"2d",
           586 => x"08",
           587 => x"04",
           588 => x"0c",
           589 => x"2d",
           590 => x"08",
           591 => x"04",
           592 => x"0c",
           593 => x"2d",
           594 => x"08",
           595 => x"04",
           596 => x"0c",
           597 => x"2d",
           598 => x"08",
           599 => x"04",
           600 => x"00",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"53",
           609 => x"00",
           610 => x"06",
           611 => x"09",
           612 => x"05",
           613 => x"2b",
           614 => x"06",
           615 => x"04",
           616 => x"72",
           617 => x"05",
           618 => x"05",
           619 => x"72",
           620 => x"53",
           621 => x"51",
           622 => x"04",
           623 => x"70",
           624 => x"27",
           625 => x"71",
           626 => x"53",
           627 => x"0b",
           628 => x"8c",
           629 => x"f3",
           630 => x"82",
           631 => x"02",
           632 => x"0c",
           633 => x"82",
           634 => x"8c",
           635 => x"bb",
           636 => x"05",
           637 => x"e8",
           638 => x"08",
           639 => x"e8",
           640 => x"08",
           641 => x"b0",
           642 => x"84",
           643 => x"bb",
           644 => x"82",
           645 => x"f8",
           646 => x"bb",
           647 => x"05",
           648 => x"bb",
           649 => x"54",
           650 => x"82",
           651 => x"04",
           652 => x"08",
           653 => x"e8",
           654 => x"0d",
           655 => x"08",
           656 => x"85",
           657 => x"81",
           658 => x"06",
           659 => x"52",
           660 => x"80",
           661 => x"e8",
           662 => x"08",
           663 => x"8d",
           664 => x"82",
           665 => x"f4",
           666 => x"c4",
           667 => x"e8",
           668 => x"08",
           669 => x"bb",
           670 => x"05",
           671 => x"82",
           672 => x"f8",
           673 => x"bb",
           674 => x"05",
           675 => x"e8",
           676 => x"0c",
           677 => x"08",
           678 => x"8a",
           679 => x"38",
           680 => x"bb",
           681 => x"05",
           682 => x"e9",
           683 => x"e8",
           684 => x"08",
           685 => x"3f",
           686 => x"08",
           687 => x"e8",
           688 => x"0c",
           689 => x"e8",
           690 => x"08",
           691 => x"81",
           692 => x"80",
           693 => x"e8",
           694 => x"0c",
           695 => x"82",
           696 => x"fc",
           697 => x"bb",
           698 => x"05",
           699 => x"71",
           700 => x"bb",
           701 => x"05",
           702 => x"82",
           703 => x"8c",
           704 => x"bb",
           705 => x"05",
           706 => x"82",
           707 => x"fc",
           708 => x"80",
           709 => x"e8",
           710 => x"08",
           711 => x"34",
           712 => x"08",
           713 => x"70",
           714 => x"08",
           715 => x"52",
           716 => x"08",
           717 => x"82",
           718 => x"87",
           719 => x"bb",
           720 => x"82",
           721 => x"02",
           722 => x"0c",
           723 => x"86",
           724 => x"e8",
           725 => x"34",
           726 => x"08",
           727 => x"82",
           728 => x"e0",
           729 => x"0a",
           730 => x"e8",
           731 => x"0c",
           732 => x"08",
           733 => x"82",
           734 => x"fc",
           735 => x"bb",
           736 => x"05",
           737 => x"bb",
           738 => x"05",
           739 => x"bb",
           740 => x"05",
           741 => x"54",
           742 => x"82",
           743 => x"70",
           744 => x"08",
           745 => x"82",
           746 => x"ec",
           747 => x"bb",
           748 => x"05",
           749 => x"54",
           750 => x"82",
           751 => x"dc",
           752 => x"82",
           753 => x"54",
           754 => x"82",
           755 => x"04",
           756 => x"08",
           757 => x"e8",
           758 => x"0d",
           759 => x"08",
           760 => x"82",
           761 => x"fc",
           762 => x"bb",
           763 => x"05",
           764 => x"bb",
           765 => x"05",
           766 => x"bb",
           767 => x"05",
           768 => x"a3",
           769 => x"dc",
           770 => x"bb",
           771 => x"05",
           772 => x"e8",
           773 => x"08",
           774 => x"dc",
           775 => x"87",
           776 => x"bb",
           777 => x"82",
           778 => x"02",
           779 => x"0c",
           780 => x"80",
           781 => x"e8",
           782 => x"23",
           783 => x"08",
           784 => x"53",
           785 => x"14",
           786 => x"e8",
           787 => x"08",
           788 => x"70",
           789 => x"81",
           790 => x"06",
           791 => x"51",
           792 => x"2e",
           793 => x"0b",
           794 => x"08",
           795 => x"96",
           796 => x"bb",
           797 => x"05",
           798 => x"33",
           799 => x"bb",
           800 => x"05",
           801 => x"ff",
           802 => x"80",
           803 => x"38",
           804 => x"08",
           805 => x"81",
           806 => x"e8",
           807 => x"0c",
           808 => x"08",
           809 => x"70",
           810 => x"53",
           811 => x"95",
           812 => x"bb",
           813 => x"05",
           814 => x"73",
           815 => x"38",
           816 => x"08",
           817 => x"53",
           818 => x"81",
           819 => x"bb",
           820 => x"05",
           821 => x"b0",
           822 => x"06",
           823 => x"82",
           824 => x"e8",
           825 => x"98",
           826 => x"2c",
           827 => x"72",
           828 => x"bb",
           829 => x"05",
           830 => x"2a",
           831 => x"70",
           832 => x"51",
           833 => x"80",
           834 => x"82",
           835 => x"e4",
           836 => x"82",
           837 => x"53",
           838 => x"e8",
           839 => x"23",
           840 => x"82",
           841 => x"e8",
           842 => x"98",
           843 => x"2c",
           844 => x"2b",
           845 => x"11",
           846 => x"53",
           847 => x"72",
           848 => x"08",
           849 => x"82",
           850 => x"e8",
           851 => x"82",
           852 => x"f8",
           853 => x"15",
           854 => x"51",
           855 => x"bb",
           856 => x"05",
           857 => x"e8",
           858 => x"33",
           859 => x"70",
           860 => x"51",
           861 => x"25",
           862 => x"ff",
           863 => x"e8",
           864 => x"34",
           865 => x"08",
           866 => x"70",
           867 => x"81",
           868 => x"53",
           869 => x"38",
           870 => x"08",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"53",
           876 => x"e8",
           877 => x"23",
           878 => x"82",
           879 => x"e4",
           880 => x"83",
           881 => x"06",
           882 => x"72",
           883 => x"38",
           884 => x"08",
           885 => x"70",
           886 => x"98",
           887 => x"53",
           888 => x"81",
           889 => x"e8",
           890 => x"34",
           891 => x"08",
           892 => x"e0",
           893 => x"e8",
           894 => x"0c",
           895 => x"e8",
           896 => x"08",
           897 => x"92",
           898 => x"bb",
           899 => x"05",
           900 => x"2b",
           901 => x"11",
           902 => x"51",
           903 => x"04",
           904 => x"08",
           905 => x"70",
           906 => x"53",
           907 => x"e8",
           908 => x"23",
           909 => x"08",
           910 => x"70",
           911 => x"53",
           912 => x"e8",
           913 => x"23",
           914 => x"82",
           915 => x"e4",
           916 => x"81",
           917 => x"53",
           918 => x"e8",
           919 => x"23",
           920 => x"82",
           921 => x"e4",
           922 => x"80",
           923 => x"53",
           924 => x"e8",
           925 => x"23",
           926 => x"82",
           927 => x"e4",
           928 => x"88",
           929 => x"72",
           930 => x"08",
           931 => x"80",
           932 => x"e8",
           933 => x"34",
           934 => x"82",
           935 => x"e4",
           936 => x"84",
           937 => x"72",
           938 => x"08",
           939 => x"fb",
           940 => x"0b",
           941 => x"08",
           942 => x"82",
           943 => x"ec",
           944 => x"11",
           945 => x"82",
           946 => x"ec",
           947 => x"e3",
           948 => x"e8",
           949 => x"34",
           950 => x"82",
           951 => x"90",
           952 => x"bb",
           953 => x"05",
           954 => x"82",
           955 => x"90",
           956 => x"08",
           957 => x"82",
           958 => x"fc",
           959 => x"bb",
           960 => x"05",
           961 => x"51",
           962 => x"bb",
           963 => x"05",
           964 => x"39",
           965 => x"08",
           966 => x"82",
           967 => x"90",
           968 => x"05",
           969 => x"08",
           970 => x"70",
           971 => x"e8",
           972 => x"0c",
           973 => x"08",
           974 => x"70",
           975 => x"81",
           976 => x"51",
           977 => x"2e",
           978 => x"bb",
           979 => x"05",
           980 => x"2b",
           981 => x"2c",
           982 => x"e8",
           983 => x"08",
           984 => x"d8",
           985 => x"dc",
           986 => x"82",
           987 => x"f4",
           988 => x"39",
           989 => x"08",
           990 => x"51",
           991 => x"82",
           992 => x"53",
           993 => x"e8",
           994 => x"23",
           995 => x"08",
           996 => x"53",
           997 => x"08",
           998 => x"73",
           999 => x"54",
          1000 => x"e8",
          1001 => x"23",
          1002 => x"82",
          1003 => x"90",
          1004 => x"bb",
          1005 => x"05",
          1006 => x"82",
          1007 => x"90",
          1008 => x"08",
          1009 => x"08",
          1010 => x"82",
          1011 => x"e4",
          1012 => x"83",
          1013 => x"06",
          1014 => x"53",
          1015 => x"ab",
          1016 => x"e8",
          1017 => x"33",
          1018 => x"53",
          1019 => x"53",
          1020 => x"08",
          1021 => x"52",
          1022 => x"3f",
          1023 => x"08",
          1024 => x"bb",
          1025 => x"05",
          1026 => x"82",
          1027 => x"fc",
          1028 => x"9b",
          1029 => x"bb",
          1030 => x"72",
          1031 => x"08",
          1032 => x"82",
          1033 => x"ec",
          1034 => x"82",
          1035 => x"f4",
          1036 => x"71",
          1037 => x"72",
          1038 => x"08",
          1039 => x"8a",
          1040 => x"bb",
          1041 => x"05",
          1042 => x"2a",
          1043 => x"51",
          1044 => x"80",
          1045 => x"82",
          1046 => x"90",
          1047 => x"bb",
          1048 => x"05",
          1049 => x"82",
          1050 => x"90",
          1051 => x"08",
          1052 => x"08",
          1053 => x"53",
          1054 => x"bb",
          1055 => x"05",
          1056 => x"e8",
          1057 => x"08",
          1058 => x"bb",
          1059 => x"05",
          1060 => x"82",
          1061 => x"dc",
          1062 => x"82",
          1063 => x"dc",
          1064 => x"bb",
          1065 => x"05",
          1066 => x"e8",
          1067 => x"08",
          1068 => x"38",
          1069 => x"08",
          1070 => x"70",
          1071 => x"53",
          1072 => x"e8",
          1073 => x"23",
          1074 => x"08",
          1075 => x"30",
          1076 => x"08",
          1077 => x"82",
          1078 => x"e4",
          1079 => x"ff",
          1080 => x"53",
          1081 => x"e8",
          1082 => x"23",
          1083 => x"88",
          1084 => x"e8",
          1085 => x"23",
          1086 => x"bb",
          1087 => x"05",
          1088 => x"c0",
          1089 => x"72",
          1090 => x"08",
          1091 => x"80",
          1092 => x"bb",
          1093 => x"05",
          1094 => x"82",
          1095 => x"f4",
          1096 => x"bb",
          1097 => x"05",
          1098 => x"2a",
          1099 => x"51",
          1100 => x"80",
          1101 => x"82",
          1102 => x"90",
          1103 => x"bb",
          1104 => x"05",
          1105 => x"82",
          1106 => x"90",
          1107 => x"08",
          1108 => x"08",
          1109 => x"53",
          1110 => x"bb",
          1111 => x"05",
          1112 => x"e8",
          1113 => x"08",
          1114 => x"bb",
          1115 => x"05",
          1116 => x"82",
          1117 => x"d8",
          1118 => x"82",
          1119 => x"d8",
          1120 => x"bb",
          1121 => x"05",
          1122 => x"e8",
          1123 => x"22",
          1124 => x"51",
          1125 => x"bb",
          1126 => x"05",
          1127 => x"ec",
          1128 => x"e8",
          1129 => x"0c",
          1130 => x"08",
          1131 => x"82",
          1132 => x"f4",
          1133 => x"bb",
          1134 => x"05",
          1135 => x"70",
          1136 => x"55",
          1137 => x"82",
          1138 => x"53",
          1139 => x"82",
          1140 => x"f0",
          1141 => x"bb",
          1142 => x"05",
          1143 => x"e8",
          1144 => x"08",
          1145 => x"53",
          1146 => x"a4",
          1147 => x"e8",
          1148 => x"08",
          1149 => x"54",
          1150 => x"08",
          1151 => x"70",
          1152 => x"51",
          1153 => x"82",
          1154 => x"d0",
          1155 => x"39",
          1156 => x"08",
          1157 => x"53",
          1158 => x"11",
          1159 => x"82",
          1160 => x"d0",
          1161 => x"bb",
          1162 => x"05",
          1163 => x"bb",
          1164 => x"05",
          1165 => x"82",
          1166 => x"f0",
          1167 => x"05",
          1168 => x"08",
          1169 => x"82",
          1170 => x"f4",
          1171 => x"53",
          1172 => x"08",
          1173 => x"52",
          1174 => x"3f",
          1175 => x"08",
          1176 => x"e8",
          1177 => x"0c",
          1178 => x"e8",
          1179 => x"08",
          1180 => x"38",
          1181 => x"82",
          1182 => x"f0",
          1183 => x"bb",
          1184 => x"72",
          1185 => x"75",
          1186 => x"72",
          1187 => x"08",
          1188 => x"82",
          1189 => x"e4",
          1190 => x"b2",
          1191 => x"72",
          1192 => x"38",
          1193 => x"08",
          1194 => x"ff",
          1195 => x"72",
          1196 => x"08",
          1197 => x"82",
          1198 => x"e4",
          1199 => x"86",
          1200 => x"06",
          1201 => x"72",
          1202 => x"e7",
          1203 => x"e8",
          1204 => x"22",
          1205 => x"82",
          1206 => x"cc",
          1207 => x"bb",
          1208 => x"05",
          1209 => x"82",
          1210 => x"cc",
          1211 => x"bb",
          1212 => x"05",
          1213 => x"72",
          1214 => x"81",
          1215 => x"82",
          1216 => x"cc",
          1217 => x"05",
          1218 => x"bb",
          1219 => x"05",
          1220 => x"82",
          1221 => x"cc",
          1222 => x"05",
          1223 => x"bb",
          1224 => x"05",
          1225 => x"e8",
          1226 => x"22",
          1227 => x"08",
          1228 => x"82",
          1229 => x"e4",
          1230 => x"83",
          1231 => x"06",
          1232 => x"72",
          1233 => x"d0",
          1234 => x"e8",
          1235 => x"33",
          1236 => x"70",
          1237 => x"bb",
          1238 => x"05",
          1239 => x"51",
          1240 => x"24",
          1241 => x"bb",
          1242 => x"05",
          1243 => x"06",
          1244 => x"82",
          1245 => x"e4",
          1246 => x"39",
          1247 => x"08",
          1248 => x"53",
          1249 => x"08",
          1250 => x"73",
          1251 => x"54",
          1252 => x"e8",
          1253 => x"34",
          1254 => x"08",
          1255 => x"70",
          1256 => x"81",
          1257 => x"53",
          1258 => x"b1",
          1259 => x"e8",
          1260 => x"33",
          1261 => x"70",
          1262 => x"90",
          1263 => x"2c",
          1264 => x"51",
          1265 => x"82",
          1266 => x"ec",
          1267 => x"75",
          1268 => x"72",
          1269 => x"08",
          1270 => x"af",
          1271 => x"e8",
          1272 => x"33",
          1273 => x"70",
          1274 => x"90",
          1275 => x"2c",
          1276 => x"51",
          1277 => x"82",
          1278 => x"ec",
          1279 => x"75",
          1280 => x"72",
          1281 => x"08",
          1282 => x"82",
          1283 => x"e4",
          1284 => x"83",
          1285 => x"53",
          1286 => x"82",
          1287 => x"ec",
          1288 => x"11",
          1289 => x"82",
          1290 => x"ec",
          1291 => x"90",
          1292 => x"2c",
          1293 => x"73",
          1294 => x"82",
          1295 => x"88",
          1296 => x"a0",
          1297 => x"3f",
          1298 => x"bb",
          1299 => x"05",
          1300 => x"2a",
          1301 => x"51",
          1302 => x"80",
          1303 => x"82",
          1304 => x"88",
          1305 => x"ad",
          1306 => x"3f",
          1307 => x"82",
          1308 => x"e4",
          1309 => x"84",
          1310 => x"06",
          1311 => x"72",
          1312 => x"38",
          1313 => x"08",
          1314 => x"52",
          1315 => x"a5",
          1316 => x"82",
          1317 => x"e4",
          1318 => x"85",
          1319 => x"06",
          1320 => x"72",
          1321 => x"38",
          1322 => x"08",
          1323 => x"52",
          1324 => x"81",
          1325 => x"e8",
          1326 => x"22",
          1327 => x"70",
          1328 => x"51",
          1329 => x"2e",
          1330 => x"bb",
          1331 => x"05",
          1332 => x"51",
          1333 => x"82",
          1334 => x"f4",
          1335 => x"72",
          1336 => x"81",
          1337 => x"82",
          1338 => x"88",
          1339 => x"82",
          1340 => x"f8",
          1341 => x"89",
          1342 => x"bb",
          1343 => x"05",
          1344 => x"2a",
          1345 => x"51",
          1346 => x"80",
          1347 => x"82",
          1348 => x"ec",
          1349 => x"11",
          1350 => x"82",
          1351 => x"ec",
          1352 => x"90",
          1353 => x"2c",
          1354 => x"73",
          1355 => x"82",
          1356 => x"88",
          1357 => x"b0",
          1358 => x"3f",
          1359 => x"bb",
          1360 => x"05",
          1361 => x"2a",
          1362 => x"51",
          1363 => x"80",
          1364 => x"82",
          1365 => x"e8",
          1366 => x"11",
          1367 => x"82",
          1368 => x"e8",
          1369 => x"98",
          1370 => x"2c",
          1371 => x"73",
          1372 => x"82",
          1373 => x"88",
          1374 => x"b0",
          1375 => x"3f",
          1376 => x"bb",
          1377 => x"05",
          1378 => x"2a",
          1379 => x"51",
          1380 => x"b0",
          1381 => x"e8",
          1382 => x"22",
          1383 => x"54",
          1384 => x"e8",
          1385 => x"23",
          1386 => x"70",
          1387 => x"53",
          1388 => x"90",
          1389 => x"e8",
          1390 => x"08",
          1391 => x"87",
          1392 => x"39",
          1393 => x"08",
          1394 => x"53",
          1395 => x"2e",
          1396 => x"97",
          1397 => x"e8",
          1398 => x"08",
          1399 => x"e8",
          1400 => x"33",
          1401 => x"3f",
          1402 => x"82",
          1403 => x"f8",
          1404 => x"72",
          1405 => x"09",
          1406 => x"cb",
          1407 => x"e8",
          1408 => x"22",
          1409 => x"53",
          1410 => x"e8",
          1411 => x"23",
          1412 => x"ff",
          1413 => x"83",
          1414 => x"81",
          1415 => x"bb",
          1416 => x"05",
          1417 => x"bb",
          1418 => x"05",
          1419 => x"52",
          1420 => x"08",
          1421 => x"81",
          1422 => x"e8",
          1423 => x"0c",
          1424 => x"3f",
          1425 => x"82",
          1426 => x"f8",
          1427 => x"72",
          1428 => x"09",
          1429 => x"cb",
          1430 => x"e8",
          1431 => x"22",
          1432 => x"53",
          1433 => x"e8",
          1434 => x"23",
          1435 => x"ff",
          1436 => x"83",
          1437 => x"80",
          1438 => x"bb",
          1439 => x"05",
          1440 => x"bb",
          1441 => x"05",
          1442 => x"52",
          1443 => x"3f",
          1444 => x"08",
          1445 => x"81",
          1446 => x"e8",
          1447 => x"0c",
          1448 => x"82",
          1449 => x"f0",
          1450 => x"bb",
          1451 => x"38",
          1452 => x"08",
          1453 => x"52",
          1454 => x"08",
          1455 => x"ff",
          1456 => x"e8",
          1457 => x"0c",
          1458 => x"08",
          1459 => x"70",
          1460 => x"85",
          1461 => x"39",
          1462 => x"08",
          1463 => x"70",
          1464 => x"81",
          1465 => x"53",
          1466 => x"80",
          1467 => x"bb",
          1468 => x"05",
          1469 => x"54",
          1470 => x"bb",
          1471 => x"05",
          1472 => x"2b",
          1473 => x"51",
          1474 => x"25",
          1475 => x"bb",
          1476 => x"05",
          1477 => x"51",
          1478 => x"d2",
          1479 => x"e8",
          1480 => x"08",
          1481 => x"e8",
          1482 => x"33",
          1483 => x"3f",
          1484 => x"bb",
          1485 => x"05",
          1486 => x"39",
          1487 => x"08",
          1488 => x"53",
          1489 => x"09",
          1490 => x"38",
          1491 => x"bb",
          1492 => x"05",
          1493 => x"82",
          1494 => x"ec",
          1495 => x"0b",
          1496 => x"08",
          1497 => x"8a",
          1498 => x"e8",
          1499 => x"23",
          1500 => x"82",
          1501 => x"88",
          1502 => x"82",
          1503 => x"f8",
          1504 => x"84",
          1505 => x"ea",
          1506 => x"e8",
          1507 => x"08",
          1508 => x"70",
          1509 => x"08",
          1510 => x"51",
          1511 => x"e8",
          1512 => x"08",
          1513 => x"0c",
          1514 => x"82",
          1515 => x"04",
          1516 => x"08",
          1517 => x"e8",
          1518 => x"0d",
          1519 => x"08",
          1520 => x"e8",
          1521 => x"08",
          1522 => x"e8",
          1523 => x"08",
          1524 => x"3f",
          1525 => x"08",
          1526 => x"dc",
          1527 => x"3d",
          1528 => x"e8",
          1529 => x"bb",
          1530 => x"82",
          1531 => x"fb",
          1532 => x"0b",
          1533 => x"08",
          1534 => x"82",
          1535 => x"85",
          1536 => x"81",
          1537 => x"32",
          1538 => x"51",
          1539 => x"53",
          1540 => x"8d",
          1541 => x"82",
          1542 => x"f4",
          1543 => x"92",
          1544 => x"e8",
          1545 => x"08",
          1546 => x"82",
          1547 => x"88",
          1548 => x"05",
          1549 => x"08",
          1550 => x"53",
          1551 => x"e8",
          1552 => x"34",
          1553 => x"06",
          1554 => x"2e",
          1555 => x"d3",
          1556 => x"d3",
          1557 => x"82",
          1558 => x"fc",
          1559 => x"90",
          1560 => x"53",
          1561 => x"bb",
          1562 => x"72",
          1563 => x"b1",
          1564 => x"82",
          1565 => x"f8",
          1566 => x"a5",
          1567 => x"b0",
          1568 => x"b0",
          1569 => x"8a",
          1570 => x"08",
          1571 => x"82",
          1572 => x"53",
          1573 => x"8a",
          1574 => x"82",
          1575 => x"f8",
          1576 => x"bb",
          1577 => x"05",
          1578 => x"bb",
          1579 => x"05",
          1580 => x"bb",
          1581 => x"05",
          1582 => x"dc",
          1583 => x"0d",
          1584 => x"0c",
          1585 => x"e8",
          1586 => x"bb",
          1587 => x"3d",
          1588 => x"82",
          1589 => x"f8",
          1590 => x"bb",
          1591 => x"05",
          1592 => x"33",
          1593 => x"70",
          1594 => x"81",
          1595 => x"51",
          1596 => x"80",
          1597 => x"ff",
          1598 => x"e8",
          1599 => x"0c",
          1600 => x"82",
          1601 => x"88",
          1602 => x"72",
          1603 => x"e8",
          1604 => x"08",
          1605 => x"bb",
          1606 => x"05",
          1607 => x"82",
          1608 => x"fc",
          1609 => x"81",
          1610 => x"72",
          1611 => x"38",
          1612 => x"08",
          1613 => x"82",
          1614 => x"8c",
          1615 => x"82",
          1616 => x"fc",
          1617 => x"90",
          1618 => x"53",
          1619 => x"bb",
          1620 => x"72",
          1621 => x"ab",
          1622 => x"82",
          1623 => x"f8",
          1624 => x"9f",
          1625 => x"e8",
          1626 => x"08",
          1627 => x"e8",
          1628 => x"0c",
          1629 => x"e8",
          1630 => x"08",
          1631 => x"0c",
          1632 => x"82",
          1633 => x"04",
          1634 => x"08",
          1635 => x"e8",
          1636 => x"0d",
          1637 => x"08",
          1638 => x"e8",
          1639 => x"08",
          1640 => x"82",
          1641 => x"70",
          1642 => x"0c",
          1643 => x"0d",
          1644 => x"0c",
          1645 => x"e8",
          1646 => x"bb",
          1647 => x"3d",
          1648 => x"e8",
          1649 => x"08",
          1650 => x"70",
          1651 => x"81",
          1652 => x"06",
          1653 => x"51",
          1654 => x"2e",
          1655 => x"0b",
          1656 => x"08",
          1657 => x"81",
          1658 => x"bb",
          1659 => x"05",
          1660 => x"33",
          1661 => x"70",
          1662 => x"51",
          1663 => x"80",
          1664 => x"38",
          1665 => x"08",
          1666 => x"82",
          1667 => x"8c",
          1668 => x"54",
          1669 => x"88",
          1670 => x"9f",
          1671 => x"e8",
          1672 => x"08",
          1673 => x"82",
          1674 => x"88",
          1675 => x"57",
          1676 => x"75",
          1677 => x"81",
          1678 => x"82",
          1679 => x"8c",
          1680 => x"11",
          1681 => x"8c",
          1682 => x"bb",
          1683 => x"05",
          1684 => x"bb",
          1685 => x"05",
          1686 => x"80",
          1687 => x"bb",
          1688 => x"05",
          1689 => x"e8",
          1690 => x"08",
          1691 => x"e8",
          1692 => x"08",
          1693 => x"06",
          1694 => x"08",
          1695 => x"72",
          1696 => x"dc",
          1697 => x"a3",
          1698 => x"e8",
          1699 => x"08",
          1700 => x"81",
          1701 => x"0c",
          1702 => x"08",
          1703 => x"70",
          1704 => x"08",
          1705 => x"51",
          1706 => x"ff",
          1707 => x"e8",
          1708 => x"0c",
          1709 => x"08",
          1710 => x"82",
          1711 => x"87",
          1712 => x"bb",
          1713 => x"82",
          1714 => x"02",
          1715 => x"0c",
          1716 => x"82",
          1717 => x"88",
          1718 => x"11",
          1719 => x"32",
          1720 => x"51",
          1721 => x"71",
          1722 => x"38",
          1723 => x"bb",
          1724 => x"05",
          1725 => x"39",
          1726 => x"08",
          1727 => x"85",
          1728 => x"86",
          1729 => x"06",
          1730 => x"52",
          1731 => x"80",
          1732 => x"bb",
          1733 => x"05",
          1734 => x"e8",
          1735 => x"08",
          1736 => x"12",
          1737 => x"bf",
          1738 => x"71",
          1739 => x"82",
          1740 => x"88",
          1741 => x"11",
          1742 => x"8c",
          1743 => x"bb",
          1744 => x"05",
          1745 => x"33",
          1746 => x"e8",
          1747 => x"0c",
          1748 => x"82",
          1749 => x"bb",
          1750 => x"05",
          1751 => x"33",
          1752 => x"70",
          1753 => x"51",
          1754 => x"80",
          1755 => x"38",
          1756 => x"08",
          1757 => x"70",
          1758 => x"82",
          1759 => x"fc",
          1760 => x"52",
          1761 => x"08",
          1762 => x"a9",
          1763 => x"e8",
          1764 => x"08",
          1765 => x"08",
          1766 => x"53",
          1767 => x"33",
          1768 => x"51",
          1769 => x"14",
          1770 => x"82",
          1771 => x"f8",
          1772 => x"d7",
          1773 => x"e8",
          1774 => x"08",
          1775 => x"05",
          1776 => x"81",
          1777 => x"bb",
          1778 => x"05",
          1779 => x"e8",
          1780 => x"08",
          1781 => x"08",
          1782 => x"2d",
          1783 => x"08",
          1784 => x"e8",
          1785 => x"0c",
          1786 => x"e8",
          1787 => x"08",
          1788 => x"f2",
          1789 => x"e8",
          1790 => x"08",
          1791 => x"08",
          1792 => x"82",
          1793 => x"88",
          1794 => x"11",
          1795 => x"e8",
          1796 => x"0c",
          1797 => x"e8",
          1798 => x"08",
          1799 => x"81",
          1800 => x"82",
          1801 => x"f0",
          1802 => x"07",
          1803 => x"bb",
          1804 => x"05",
          1805 => x"82",
          1806 => x"f0",
          1807 => x"07",
          1808 => x"bb",
          1809 => x"05",
          1810 => x"e8",
          1811 => x"08",
          1812 => x"e8",
          1813 => x"33",
          1814 => x"ff",
          1815 => x"e8",
          1816 => x"0c",
          1817 => x"bb",
          1818 => x"05",
          1819 => x"08",
          1820 => x"12",
          1821 => x"e8",
          1822 => x"08",
          1823 => x"06",
          1824 => x"e8",
          1825 => x"0c",
          1826 => x"82",
          1827 => x"f8",
          1828 => x"bb",
          1829 => x"3d",
          1830 => x"e8",
          1831 => x"bb",
          1832 => x"82",
          1833 => x"fd",
          1834 => x"bb",
          1835 => x"05",
          1836 => x"e8",
          1837 => x"0c",
          1838 => x"08",
          1839 => x"82",
          1840 => x"f8",
          1841 => x"bb",
          1842 => x"05",
          1843 => x"82",
          1844 => x"bb",
          1845 => x"05",
          1846 => x"e8",
          1847 => x"08",
          1848 => x"38",
          1849 => x"08",
          1850 => x"82",
          1851 => x"90",
          1852 => x"51",
          1853 => x"08",
          1854 => x"71",
          1855 => x"38",
          1856 => x"08",
          1857 => x"82",
          1858 => x"90",
          1859 => x"82",
          1860 => x"fc",
          1861 => x"bb",
          1862 => x"05",
          1863 => x"e8",
          1864 => x"08",
          1865 => x"e8",
          1866 => x"0c",
          1867 => x"08",
          1868 => x"81",
          1869 => x"e8",
          1870 => x"0c",
          1871 => x"08",
          1872 => x"ff",
          1873 => x"e8",
          1874 => x"0c",
          1875 => x"08",
          1876 => x"80",
          1877 => x"38",
          1878 => x"08",
          1879 => x"ff",
          1880 => x"e8",
          1881 => x"0c",
          1882 => x"08",
          1883 => x"ff",
          1884 => x"e8",
          1885 => x"0c",
          1886 => x"08",
          1887 => x"82",
          1888 => x"f8",
          1889 => x"51",
          1890 => x"34",
          1891 => x"82",
          1892 => x"90",
          1893 => x"05",
          1894 => x"08",
          1895 => x"82",
          1896 => x"90",
          1897 => x"05",
          1898 => x"08",
          1899 => x"82",
          1900 => x"90",
          1901 => x"2e",
          1902 => x"bb",
          1903 => x"05",
          1904 => x"33",
          1905 => x"08",
          1906 => x"81",
          1907 => x"e8",
          1908 => x"0c",
          1909 => x"08",
          1910 => x"52",
          1911 => x"34",
          1912 => x"08",
          1913 => x"81",
          1914 => x"e8",
          1915 => x"0c",
          1916 => x"82",
          1917 => x"88",
          1918 => x"82",
          1919 => x"51",
          1920 => x"82",
          1921 => x"04",
          1922 => x"08",
          1923 => x"e8",
          1924 => x"0d",
          1925 => x"08",
          1926 => x"82",
          1927 => x"fc",
          1928 => x"bb",
          1929 => x"05",
          1930 => x"33",
          1931 => x"08",
          1932 => x"81",
          1933 => x"e8",
          1934 => x"0c",
          1935 => x"06",
          1936 => x"80",
          1937 => x"da",
          1938 => x"e8",
          1939 => x"08",
          1940 => x"bb",
          1941 => x"05",
          1942 => x"e8",
          1943 => x"08",
          1944 => x"08",
          1945 => x"31",
          1946 => x"dc",
          1947 => x"3d",
          1948 => x"e8",
          1949 => x"bb",
          1950 => x"82",
          1951 => x"fe",
          1952 => x"bb",
          1953 => x"05",
          1954 => x"e8",
          1955 => x"0c",
          1956 => x"08",
          1957 => x"52",
          1958 => x"bb",
          1959 => x"05",
          1960 => x"82",
          1961 => x"8c",
          1962 => x"bb",
          1963 => x"05",
          1964 => x"70",
          1965 => x"bb",
          1966 => x"05",
          1967 => x"82",
          1968 => x"fc",
          1969 => x"81",
          1970 => x"70",
          1971 => x"38",
          1972 => x"82",
          1973 => x"88",
          1974 => x"82",
          1975 => x"51",
          1976 => x"82",
          1977 => x"04",
          1978 => x"08",
          1979 => x"e8",
          1980 => x"0d",
          1981 => x"08",
          1982 => x"82",
          1983 => x"fc",
          1984 => x"bb",
          1985 => x"05",
          1986 => x"e8",
          1987 => x"0c",
          1988 => x"08",
          1989 => x"80",
          1990 => x"38",
          1991 => x"08",
          1992 => x"81",
          1993 => x"e8",
          1994 => x"0c",
          1995 => x"08",
          1996 => x"ff",
          1997 => x"e8",
          1998 => x"0c",
          1999 => x"08",
          2000 => x"80",
          2001 => x"82",
          2002 => x"f8",
          2003 => x"70",
          2004 => x"e8",
          2005 => x"08",
          2006 => x"bb",
          2007 => x"05",
          2008 => x"e8",
          2009 => x"08",
          2010 => x"71",
          2011 => x"e8",
          2012 => x"08",
          2013 => x"bb",
          2014 => x"05",
          2015 => x"39",
          2016 => x"08",
          2017 => x"70",
          2018 => x"0c",
          2019 => x"0d",
          2020 => x"0c",
          2021 => x"e8",
          2022 => x"bb",
          2023 => x"3d",
          2024 => x"e8",
          2025 => x"08",
          2026 => x"f4",
          2027 => x"e8",
          2028 => x"08",
          2029 => x"82",
          2030 => x"8c",
          2031 => x"05",
          2032 => x"08",
          2033 => x"82",
          2034 => x"88",
          2035 => x"33",
          2036 => x"06",
          2037 => x"51",
          2038 => x"84",
          2039 => x"39",
          2040 => x"08",
          2041 => x"52",
          2042 => x"bb",
          2043 => x"05",
          2044 => x"82",
          2045 => x"88",
          2046 => x"81",
          2047 => x"51",
          2048 => x"80",
          2049 => x"e8",
          2050 => x"0c",
          2051 => x"82",
          2052 => x"90",
          2053 => x"05",
          2054 => x"08",
          2055 => x"82",
          2056 => x"90",
          2057 => x"2e",
          2058 => x"81",
          2059 => x"e8",
          2060 => x"08",
          2061 => x"e8",
          2062 => x"e8",
          2063 => x"08",
          2064 => x"53",
          2065 => x"ff",
          2066 => x"e8",
          2067 => x"0c",
          2068 => x"82",
          2069 => x"8c",
          2070 => x"05",
          2071 => x"08",
          2072 => x"82",
          2073 => x"8c",
          2074 => x"33",
          2075 => x"8c",
          2076 => x"82",
          2077 => x"fc",
          2078 => x"39",
          2079 => x"08",
          2080 => x"70",
          2081 => x"e8",
          2082 => x"08",
          2083 => x"71",
          2084 => x"bb",
          2085 => x"05",
          2086 => x"52",
          2087 => x"39",
          2088 => x"bb",
          2089 => x"05",
          2090 => x"e8",
          2091 => x"08",
          2092 => x"0c",
          2093 => x"82",
          2094 => x"04",
          2095 => x"08",
          2096 => x"e8",
          2097 => x"0d",
          2098 => x"08",
          2099 => x"82",
          2100 => x"f8",
          2101 => x"bb",
          2102 => x"05",
          2103 => x"80",
          2104 => x"e8",
          2105 => x"0c",
          2106 => x"82",
          2107 => x"f8",
          2108 => x"71",
          2109 => x"e8",
          2110 => x"08",
          2111 => x"bb",
          2112 => x"05",
          2113 => x"ff",
          2114 => x"70",
          2115 => x"38",
          2116 => x"08",
          2117 => x"ff",
          2118 => x"e8",
          2119 => x"0c",
          2120 => x"08",
          2121 => x"ff",
          2122 => x"ff",
          2123 => x"bb",
          2124 => x"05",
          2125 => x"82",
          2126 => x"f8",
          2127 => x"bb",
          2128 => x"05",
          2129 => x"e8",
          2130 => x"08",
          2131 => x"bb",
          2132 => x"05",
          2133 => x"bb",
          2134 => x"05",
          2135 => x"dc",
          2136 => x"0d",
          2137 => x"0c",
          2138 => x"e8",
          2139 => x"bb",
          2140 => x"3d",
          2141 => x"e8",
          2142 => x"08",
          2143 => x"08",
          2144 => x"82",
          2145 => x"90",
          2146 => x"2e",
          2147 => x"82",
          2148 => x"90",
          2149 => x"05",
          2150 => x"08",
          2151 => x"82",
          2152 => x"90",
          2153 => x"05",
          2154 => x"08",
          2155 => x"82",
          2156 => x"90",
          2157 => x"2e",
          2158 => x"bb",
          2159 => x"05",
          2160 => x"82",
          2161 => x"fc",
          2162 => x"52",
          2163 => x"82",
          2164 => x"fc",
          2165 => x"05",
          2166 => x"08",
          2167 => x"ff",
          2168 => x"bb",
          2169 => x"05",
          2170 => x"bb",
          2171 => x"84",
          2172 => x"bb",
          2173 => x"82",
          2174 => x"02",
          2175 => x"0c",
          2176 => x"80",
          2177 => x"e8",
          2178 => x"0c",
          2179 => x"08",
          2180 => x"80",
          2181 => x"82",
          2182 => x"88",
          2183 => x"82",
          2184 => x"88",
          2185 => x"0b",
          2186 => x"08",
          2187 => x"82",
          2188 => x"fc",
          2189 => x"38",
          2190 => x"bb",
          2191 => x"05",
          2192 => x"e8",
          2193 => x"08",
          2194 => x"08",
          2195 => x"82",
          2196 => x"8c",
          2197 => x"25",
          2198 => x"bb",
          2199 => x"05",
          2200 => x"bb",
          2201 => x"05",
          2202 => x"82",
          2203 => x"f0",
          2204 => x"bb",
          2205 => x"05",
          2206 => x"81",
          2207 => x"e8",
          2208 => x"0c",
          2209 => x"08",
          2210 => x"82",
          2211 => x"fc",
          2212 => x"53",
          2213 => x"08",
          2214 => x"52",
          2215 => x"08",
          2216 => x"51",
          2217 => x"82",
          2218 => x"70",
          2219 => x"08",
          2220 => x"54",
          2221 => x"08",
          2222 => x"80",
          2223 => x"82",
          2224 => x"f8",
          2225 => x"82",
          2226 => x"f8",
          2227 => x"bb",
          2228 => x"05",
          2229 => x"bb",
          2230 => x"89",
          2231 => x"bb",
          2232 => x"82",
          2233 => x"02",
          2234 => x"0c",
          2235 => x"80",
          2236 => x"e8",
          2237 => x"0c",
          2238 => x"08",
          2239 => x"80",
          2240 => x"82",
          2241 => x"88",
          2242 => x"82",
          2243 => x"88",
          2244 => x"0b",
          2245 => x"08",
          2246 => x"82",
          2247 => x"8c",
          2248 => x"25",
          2249 => x"bb",
          2250 => x"05",
          2251 => x"bb",
          2252 => x"05",
          2253 => x"82",
          2254 => x"8c",
          2255 => x"82",
          2256 => x"88",
          2257 => x"81",
          2258 => x"bb",
          2259 => x"82",
          2260 => x"f8",
          2261 => x"82",
          2262 => x"fc",
          2263 => x"2e",
          2264 => x"bb",
          2265 => x"05",
          2266 => x"bb",
          2267 => x"05",
          2268 => x"e8",
          2269 => x"08",
          2270 => x"dc",
          2271 => x"3d",
          2272 => x"e8",
          2273 => x"bb",
          2274 => x"82",
          2275 => x"fd",
          2276 => x"53",
          2277 => x"08",
          2278 => x"52",
          2279 => x"08",
          2280 => x"51",
          2281 => x"82",
          2282 => x"70",
          2283 => x"0c",
          2284 => x"0d",
          2285 => x"0c",
          2286 => x"e8",
          2287 => x"bb",
          2288 => x"3d",
          2289 => x"82",
          2290 => x"8c",
          2291 => x"82",
          2292 => x"88",
          2293 => x"93",
          2294 => x"dc",
          2295 => x"bb",
          2296 => x"85",
          2297 => x"bb",
          2298 => x"82",
          2299 => x"02",
          2300 => x"0c",
          2301 => x"81",
          2302 => x"e8",
          2303 => x"0c",
          2304 => x"bb",
          2305 => x"05",
          2306 => x"e8",
          2307 => x"08",
          2308 => x"08",
          2309 => x"27",
          2310 => x"bb",
          2311 => x"05",
          2312 => x"ae",
          2313 => x"82",
          2314 => x"8c",
          2315 => x"a2",
          2316 => x"e8",
          2317 => x"08",
          2318 => x"e8",
          2319 => x"0c",
          2320 => x"08",
          2321 => x"10",
          2322 => x"08",
          2323 => x"ff",
          2324 => x"bb",
          2325 => x"05",
          2326 => x"80",
          2327 => x"bb",
          2328 => x"05",
          2329 => x"e8",
          2330 => x"08",
          2331 => x"82",
          2332 => x"88",
          2333 => x"bb",
          2334 => x"05",
          2335 => x"bb",
          2336 => x"05",
          2337 => x"e8",
          2338 => x"08",
          2339 => x"08",
          2340 => x"07",
          2341 => x"08",
          2342 => x"82",
          2343 => x"fc",
          2344 => x"2a",
          2345 => x"08",
          2346 => x"82",
          2347 => x"8c",
          2348 => x"2a",
          2349 => x"08",
          2350 => x"ff",
          2351 => x"bb",
          2352 => x"05",
          2353 => x"93",
          2354 => x"e8",
          2355 => x"08",
          2356 => x"e8",
          2357 => x"0c",
          2358 => x"82",
          2359 => x"f8",
          2360 => x"82",
          2361 => x"f4",
          2362 => x"82",
          2363 => x"f4",
          2364 => x"bb",
          2365 => x"3d",
          2366 => x"e8",
          2367 => x"bb",
          2368 => x"82",
          2369 => x"f7",
          2370 => x"0b",
          2371 => x"08",
          2372 => x"82",
          2373 => x"8c",
          2374 => x"80",
          2375 => x"bb",
          2376 => x"05",
          2377 => x"51",
          2378 => x"53",
          2379 => x"e8",
          2380 => x"34",
          2381 => x"06",
          2382 => x"2e",
          2383 => x"91",
          2384 => x"e8",
          2385 => x"08",
          2386 => x"05",
          2387 => x"ce",
          2388 => x"e8",
          2389 => x"33",
          2390 => x"2e",
          2391 => x"a4",
          2392 => x"82",
          2393 => x"f0",
          2394 => x"bb",
          2395 => x"05",
          2396 => x"81",
          2397 => x"70",
          2398 => x"72",
          2399 => x"e8",
          2400 => x"34",
          2401 => x"08",
          2402 => x"53",
          2403 => x"09",
          2404 => x"dc",
          2405 => x"e8",
          2406 => x"08",
          2407 => x"05",
          2408 => x"08",
          2409 => x"33",
          2410 => x"08",
          2411 => x"82",
          2412 => x"f8",
          2413 => x"bb",
          2414 => x"05",
          2415 => x"e8",
          2416 => x"08",
          2417 => x"b6",
          2418 => x"e8",
          2419 => x"08",
          2420 => x"84",
          2421 => x"39",
          2422 => x"bb",
          2423 => x"05",
          2424 => x"e8",
          2425 => x"08",
          2426 => x"05",
          2427 => x"08",
          2428 => x"33",
          2429 => x"08",
          2430 => x"81",
          2431 => x"0b",
          2432 => x"08",
          2433 => x"82",
          2434 => x"88",
          2435 => x"08",
          2436 => x"0c",
          2437 => x"53",
          2438 => x"bb",
          2439 => x"05",
          2440 => x"39",
          2441 => x"08",
          2442 => x"53",
          2443 => x"8d",
          2444 => x"82",
          2445 => x"ec",
          2446 => x"80",
          2447 => x"e8",
          2448 => x"33",
          2449 => x"27",
          2450 => x"bb",
          2451 => x"05",
          2452 => x"b9",
          2453 => x"8d",
          2454 => x"82",
          2455 => x"ec",
          2456 => x"d8",
          2457 => x"82",
          2458 => x"f4",
          2459 => x"39",
          2460 => x"08",
          2461 => x"53",
          2462 => x"90",
          2463 => x"e8",
          2464 => x"33",
          2465 => x"26",
          2466 => x"39",
          2467 => x"bb",
          2468 => x"05",
          2469 => x"39",
          2470 => x"bb",
          2471 => x"05",
          2472 => x"82",
          2473 => x"fc",
          2474 => x"bb",
          2475 => x"05",
          2476 => x"73",
          2477 => x"38",
          2478 => x"08",
          2479 => x"53",
          2480 => x"27",
          2481 => x"bb",
          2482 => x"05",
          2483 => x"51",
          2484 => x"bb",
          2485 => x"05",
          2486 => x"e8",
          2487 => x"33",
          2488 => x"53",
          2489 => x"e8",
          2490 => x"34",
          2491 => x"08",
          2492 => x"53",
          2493 => x"ad",
          2494 => x"e8",
          2495 => x"33",
          2496 => x"53",
          2497 => x"e8",
          2498 => x"34",
          2499 => x"08",
          2500 => x"53",
          2501 => x"8d",
          2502 => x"82",
          2503 => x"ec",
          2504 => x"98",
          2505 => x"e8",
          2506 => x"33",
          2507 => x"08",
          2508 => x"54",
          2509 => x"26",
          2510 => x"0b",
          2511 => x"08",
          2512 => x"80",
          2513 => x"bb",
          2514 => x"05",
          2515 => x"bb",
          2516 => x"05",
          2517 => x"bb",
          2518 => x"05",
          2519 => x"82",
          2520 => x"fc",
          2521 => x"bb",
          2522 => x"05",
          2523 => x"81",
          2524 => x"70",
          2525 => x"52",
          2526 => x"33",
          2527 => x"08",
          2528 => x"fe",
          2529 => x"bb",
          2530 => x"05",
          2531 => x"80",
          2532 => x"82",
          2533 => x"fc",
          2534 => x"82",
          2535 => x"fc",
          2536 => x"bb",
          2537 => x"05",
          2538 => x"e8",
          2539 => x"08",
          2540 => x"81",
          2541 => x"e8",
          2542 => x"0c",
          2543 => x"08",
          2544 => x"82",
          2545 => x"8b",
          2546 => x"bb",
          2547 => x"82",
          2548 => x"02",
          2549 => x"0c",
          2550 => x"80",
          2551 => x"e8",
          2552 => x"34",
          2553 => x"08",
          2554 => x"53",
          2555 => x"82",
          2556 => x"88",
          2557 => x"08",
          2558 => x"33",
          2559 => x"bb",
          2560 => x"05",
          2561 => x"ff",
          2562 => x"a0",
          2563 => x"06",
          2564 => x"bb",
          2565 => x"05",
          2566 => x"81",
          2567 => x"53",
          2568 => x"bb",
          2569 => x"05",
          2570 => x"ad",
          2571 => x"06",
          2572 => x"0b",
          2573 => x"08",
          2574 => x"82",
          2575 => x"88",
          2576 => x"08",
          2577 => x"0c",
          2578 => x"53",
          2579 => x"bb",
          2580 => x"05",
          2581 => x"e8",
          2582 => x"33",
          2583 => x"2e",
          2584 => x"81",
          2585 => x"bb",
          2586 => x"05",
          2587 => x"81",
          2588 => x"70",
          2589 => x"72",
          2590 => x"e8",
          2591 => x"34",
          2592 => x"08",
          2593 => x"82",
          2594 => x"e8",
          2595 => x"bb",
          2596 => x"05",
          2597 => x"2e",
          2598 => x"bb",
          2599 => x"05",
          2600 => x"2e",
          2601 => x"cd",
          2602 => x"82",
          2603 => x"f4",
          2604 => x"bb",
          2605 => x"05",
          2606 => x"81",
          2607 => x"70",
          2608 => x"72",
          2609 => x"e8",
          2610 => x"34",
          2611 => x"82",
          2612 => x"e8",
          2613 => x"34",
          2614 => x"08",
          2615 => x"70",
          2616 => x"71",
          2617 => x"51",
          2618 => x"82",
          2619 => x"f8",
          2620 => x"fe",
          2621 => x"e8",
          2622 => x"33",
          2623 => x"26",
          2624 => x"0b",
          2625 => x"08",
          2626 => x"83",
          2627 => x"bb",
          2628 => x"05",
          2629 => x"73",
          2630 => x"82",
          2631 => x"f8",
          2632 => x"72",
          2633 => x"38",
          2634 => x"0b",
          2635 => x"08",
          2636 => x"82",
          2637 => x"0b",
          2638 => x"08",
          2639 => x"b2",
          2640 => x"e8",
          2641 => x"33",
          2642 => x"27",
          2643 => x"bb",
          2644 => x"05",
          2645 => x"b9",
          2646 => x"8d",
          2647 => x"82",
          2648 => x"ec",
          2649 => x"a5",
          2650 => x"82",
          2651 => x"f4",
          2652 => x"0b",
          2653 => x"08",
          2654 => x"82",
          2655 => x"f8",
          2656 => x"a0",
          2657 => x"cf",
          2658 => x"e8",
          2659 => x"33",
          2660 => x"73",
          2661 => x"82",
          2662 => x"f8",
          2663 => x"11",
          2664 => x"82",
          2665 => x"f8",
          2666 => x"bb",
          2667 => x"05",
          2668 => x"51",
          2669 => x"bb",
          2670 => x"05",
          2671 => x"e8",
          2672 => x"33",
          2673 => x"27",
          2674 => x"bb",
          2675 => x"05",
          2676 => x"51",
          2677 => x"bb",
          2678 => x"05",
          2679 => x"e8",
          2680 => x"33",
          2681 => x"26",
          2682 => x"0b",
          2683 => x"08",
          2684 => x"81",
          2685 => x"bb",
          2686 => x"05",
          2687 => x"e8",
          2688 => x"33",
          2689 => x"74",
          2690 => x"80",
          2691 => x"e8",
          2692 => x"0c",
          2693 => x"82",
          2694 => x"f4",
          2695 => x"82",
          2696 => x"fc",
          2697 => x"82",
          2698 => x"f8",
          2699 => x"12",
          2700 => x"08",
          2701 => x"82",
          2702 => x"88",
          2703 => x"08",
          2704 => x"0c",
          2705 => x"51",
          2706 => x"72",
          2707 => x"e8",
          2708 => x"34",
          2709 => x"82",
          2710 => x"f0",
          2711 => x"72",
          2712 => x"38",
          2713 => x"08",
          2714 => x"30",
          2715 => x"08",
          2716 => x"82",
          2717 => x"8c",
          2718 => x"bb",
          2719 => x"05",
          2720 => x"53",
          2721 => x"bb",
          2722 => x"05",
          2723 => x"e8",
          2724 => x"08",
          2725 => x"0c",
          2726 => x"82",
          2727 => x"04",
          2728 => x"79",
          2729 => x"56",
          2730 => x"80",
          2731 => x"38",
          2732 => x"08",
          2733 => x"3f",
          2734 => x"08",
          2735 => x"85",
          2736 => x"80",
          2737 => x"33",
          2738 => x"2e",
          2739 => x"86",
          2740 => x"55",
          2741 => x"57",
          2742 => x"82",
          2743 => x"70",
          2744 => x"e6",
          2745 => x"bb",
          2746 => x"74",
          2747 => x"51",
          2748 => x"82",
          2749 => x"8b",
          2750 => x"33",
          2751 => x"2e",
          2752 => x"81",
          2753 => x"ff",
          2754 => x"99",
          2755 => x"38",
          2756 => x"82",
          2757 => x"89",
          2758 => x"ff",
          2759 => x"52",
          2760 => x"81",
          2761 => x"84",
          2762 => x"9c",
          2763 => x"08",
          2764 => x"e8",
          2765 => x"39",
          2766 => x"51",
          2767 => x"82",
          2768 => x"80",
          2769 => x"a0",
          2770 => x"eb",
          2771 => x"a4",
          2772 => x"39",
          2773 => x"51",
          2774 => x"82",
          2775 => x"80",
          2776 => x"a0",
          2777 => x"cf",
          2778 => x"f0",
          2779 => x"39",
          2780 => x"51",
          2781 => x"82",
          2782 => x"bb",
          2783 => x"bc",
          2784 => x"82",
          2785 => x"af",
          2786 => x"f8",
          2787 => x"82",
          2788 => x"a3",
          2789 => x"a8",
          2790 => x"82",
          2791 => x"97",
          2792 => x"d0",
          2793 => x"82",
          2794 => x"8b",
          2795 => x"80",
          2796 => x"82",
          2797 => x"d8",
          2798 => x"3d",
          2799 => x"3d",
          2800 => x"56",
          2801 => x"e7",
          2802 => x"74",
          2803 => x"e8",
          2804 => x"39",
          2805 => x"74",
          2806 => x"3f",
          2807 => x"08",
          2808 => x"ef",
          2809 => x"bb",
          2810 => x"79",
          2811 => x"82",
          2812 => x"ff",
          2813 => x"87",
          2814 => x"ec",
          2815 => x"02",
          2816 => x"e3",
          2817 => x"57",
          2818 => x"30",
          2819 => x"73",
          2820 => x"59",
          2821 => x"77",
          2822 => x"83",
          2823 => x"74",
          2824 => x"81",
          2825 => x"55",
          2826 => x"81",
          2827 => x"53",
          2828 => x"3d",
          2829 => x"81",
          2830 => x"82",
          2831 => x"57",
          2832 => x"08",
          2833 => x"bb",
          2834 => x"c0",
          2835 => x"82",
          2836 => x"59",
          2837 => x"05",
          2838 => x"53",
          2839 => x"51",
          2840 => x"3f",
          2841 => x"08",
          2842 => x"dc",
          2843 => x"7a",
          2844 => x"2e",
          2845 => x"19",
          2846 => x"59",
          2847 => x"3d",
          2848 => x"81",
          2849 => x"76",
          2850 => x"07",
          2851 => x"30",
          2852 => x"72",
          2853 => x"51",
          2854 => x"2e",
          2855 => x"a3",
          2856 => x"c0",
          2857 => x"52",
          2858 => x"92",
          2859 => x"75",
          2860 => x"0c",
          2861 => x"04",
          2862 => x"7c",
          2863 => x"b7",
          2864 => x"59",
          2865 => x"53",
          2866 => x"51",
          2867 => x"82",
          2868 => x"a8",
          2869 => x"2e",
          2870 => x"81",
          2871 => x"9c",
          2872 => x"ac",
          2873 => x"60",
          2874 => x"dc",
          2875 => x"7e",
          2876 => x"82",
          2877 => x"58",
          2878 => x"04",
          2879 => x"dc",
          2880 => x"0d",
          2881 => x"0d",
          2882 => x"02",
          2883 => x"cf",
          2884 => x"73",
          2885 => x"5f",
          2886 => x"5e",
          2887 => x"82",
          2888 => x"ff",
          2889 => x"82",
          2890 => x"ff",
          2891 => x"80",
          2892 => x"27",
          2893 => x"7b",
          2894 => x"38",
          2895 => x"a7",
          2896 => x"39",
          2897 => x"72",
          2898 => x"38",
          2899 => x"82",
          2900 => x"ff",
          2901 => x"89",
          2902 => x"e0",
          2903 => x"fb",
          2904 => x"55",
          2905 => x"74",
          2906 => x"7a",
          2907 => x"72",
          2908 => x"a3",
          2909 => x"b8",
          2910 => x"39",
          2911 => x"51",
          2912 => x"3f",
          2913 => x"a1",
          2914 => x"53",
          2915 => x"8e",
          2916 => x"52",
          2917 => x"51",
          2918 => x"3f",
          2919 => x"a3",
          2920 => x"b8",
          2921 => x"15",
          2922 => x"b0",
          2923 => x"51",
          2924 => x"fe",
          2925 => x"a3",
          2926 => x"b8",
          2927 => x"55",
          2928 => x"80",
          2929 => x"18",
          2930 => x"53",
          2931 => x"7a",
          2932 => x"81",
          2933 => x"9f",
          2934 => x"38",
          2935 => x"73",
          2936 => x"ff",
          2937 => x"72",
          2938 => x"38",
          2939 => x"26",
          2940 => x"d3",
          2941 => x"73",
          2942 => x"82",
          2943 => x"52",
          2944 => x"b1",
          2945 => x"55",
          2946 => x"82",
          2947 => x"d3",
          2948 => x"18",
          2949 => x"58",
          2950 => x"82",
          2951 => x"98",
          2952 => x"2c",
          2953 => x"a0",
          2954 => x"06",
          2955 => x"e8",
          2956 => x"dc",
          2957 => x"70",
          2958 => x"a0",
          2959 => x"72",
          2960 => x"30",
          2961 => x"73",
          2962 => x"51",
          2963 => x"57",
          2964 => x"73",
          2965 => x"76",
          2966 => x"81",
          2967 => x"80",
          2968 => x"7c",
          2969 => x"78",
          2970 => x"38",
          2971 => x"82",
          2972 => x"8f",
          2973 => x"fc",
          2974 => x"9b",
          2975 => x"a3",
          2976 => x"a4",
          2977 => x"ff",
          2978 => x"82",
          2979 => x"51",
          2980 => x"82",
          2981 => x"82",
          2982 => x"82",
          2983 => x"52",
          2984 => x"51",
          2985 => x"3f",
          2986 => x"84",
          2987 => x"3f",
          2988 => x"04",
          2989 => x"87",
          2990 => x"08",
          2991 => x"3f",
          2992 => x"c1",
          2993 => x"c0",
          2994 => x"3f",
          2995 => x"b5",
          2996 => x"2a",
          2997 => x"51",
          2998 => x"2e",
          2999 => x"51",
          3000 => x"82",
          3001 => x"9d",
          3002 => x"51",
          3003 => x"72",
          3004 => x"81",
          3005 => x"71",
          3006 => x"38",
          3007 => x"85",
          3008 => x"e8",
          3009 => x"3f",
          3010 => x"f9",
          3011 => x"2a",
          3012 => x"51",
          3013 => x"2e",
          3014 => x"51",
          3015 => x"82",
          3016 => x"9c",
          3017 => x"51",
          3018 => x"72",
          3019 => x"81",
          3020 => x"71",
          3021 => x"38",
          3022 => x"c9",
          3023 => x"8c",
          3024 => x"3f",
          3025 => x"bd",
          3026 => x"2a",
          3027 => x"51",
          3028 => x"2e",
          3029 => x"51",
          3030 => x"82",
          3031 => x"9c",
          3032 => x"51",
          3033 => x"72",
          3034 => x"81",
          3035 => x"71",
          3036 => x"38",
          3037 => x"8d",
          3038 => x"b4",
          3039 => x"3f",
          3040 => x"81",
          3041 => x"2a",
          3042 => x"51",
          3043 => x"2e",
          3044 => x"51",
          3045 => x"82",
          3046 => x"9c",
          3047 => x"51",
          3048 => x"72",
          3049 => x"81",
          3050 => x"71",
          3051 => x"38",
          3052 => x"d1",
          3053 => x"dc",
          3054 => x"3f",
          3055 => x"c5",
          3056 => x"3f",
          3057 => x"04",
          3058 => x"77",
          3059 => x"a3",
          3060 => x"55",
          3061 => x"52",
          3062 => x"8d",
          3063 => x"82",
          3064 => x"54",
          3065 => x"81",
          3066 => x"98",
          3067 => x"dc",
          3068 => x"ff",
          3069 => x"dc",
          3070 => x"82",
          3071 => x"07",
          3072 => x"71",
          3073 => x"54",
          3074 => x"82",
          3075 => x"0b",
          3076 => x"d8",
          3077 => x"81",
          3078 => x"06",
          3079 => x"d2",
          3080 => x"52",
          3081 => x"b7",
          3082 => x"bb",
          3083 => x"2e",
          3084 => x"bb",
          3085 => x"cf",
          3086 => x"39",
          3087 => x"51",
          3088 => x"3f",
          3089 => x"0b",
          3090 => x"34",
          3091 => x"b6",
          3092 => x"73",
          3093 => x"81",
          3094 => x"82",
          3095 => x"74",
          3096 => x"ae",
          3097 => x"0b",
          3098 => x"0c",
          3099 => x"04",
          3100 => x"80",
          3101 => x"d2",
          3102 => x"5d",
          3103 => x"51",
          3104 => x"3f",
          3105 => x"08",
          3106 => x"59",
          3107 => x"09",
          3108 => x"38",
          3109 => x"83",
          3110 => x"b4",
          3111 => x"dc",
          3112 => x"53",
          3113 => x"bd",
          3114 => x"fa",
          3115 => x"bb",
          3116 => x"2e",
          3117 => x"a6",
          3118 => x"d5",
          3119 => x"5f",
          3120 => x"f0",
          3121 => x"93",
          3122 => x"70",
          3123 => x"f8",
          3124 => x"fd",
          3125 => x"3d",
          3126 => x"51",
          3127 => x"82",
          3128 => x"90",
          3129 => x"2c",
          3130 => x"80",
          3131 => x"d4",
          3132 => x"c1",
          3133 => x"38",
          3134 => x"83",
          3135 => x"ab",
          3136 => x"78",
          3137 => x"b3",
          3138 => x"24",
          3139 => x"80",
          3140 => x"38",
          3141 => x"78",
          3142 => x"83",
          3143 => x"2e",
          3144 => x"8e",
          3145 => x"bd",
          3146 => x"38",
          3147 => x"90",
          3148 => x"2e",
          3149 => x"78",
          3150 => x"84",
          3151 => x"39",
          3152 => x"85",
          3153 => x"80",
          3154 => x"bd",
          3155 => x"39",
          3156 => x"2e",
          3157 => x"78",
          3158 => x"b0",
          3159 => x"d0",
          3160 => x"38",
          3161 => x"24",
          3162 => x"80",
          3163 => x"fc",
          3164 => x"c3",
          3165 => x"38",
          3166 => x"78",
          3167 => x"8c",
          3168 => x"80",
          3169 => x"d2",
          3170 => x"39",
          3171 => x"2e",
          3172 => x"78",
          3173 => x"92",
          3174 => x"f8",
          3175 => x"38",
          3176 => x"2e",
          3177 => x"8d",
          3178 => x"81",
          3179 => x"d3",
          3180 => x"85",
          3181 => x"38",
          3182 => x"b4",
          3183 => x"11",
          3184 => x"05",
          3185 => x"3f",
          3186 => x"08",
          3187 => x"a6",
          3188 => x"bd",
          3189 => x"fe",
          3190 => x"ff",
          3191 => x"eb",
          3192 => x"bb",
          3193 => x"2e",
          3194 => x"63",
          3195 => x"80",
          3196 => x"cb",
          3197 => x"02",
          3198 => x"33",
          3199 => x"ce",
          3200 => x"dc",
          3201 => x"06",
          3202 => x"38",
          3203 => x"51",
          3204 => x"81",
          3205 => x"39",
          3206 => x"51",
          3207 => x"b4",
          3208 => x"11",
          3209 => x"05",
          3210 => x"3f",
          3211 => x"08",
          3212 => x"8d",
          3213 => x"80",
          3214 => x"cf",
          3215 => x"80",
          3216 => x"82",
          3217 => x"52",
          3218 => x"51",
          3219 => x"b4",
          3220 => x"11",
          3221 => x"05",
          3222 => x"3f",
          3223 => x"08",
          3224 => x"38",
          3225 => x"fc",
          3226 => x"3d",
          3227 => x"53",
          3228 => x"51",
          3229 => x"82",
          3230 => x"86",
          3231 => x"dc",
          3232 => x"53",
          3233 => x"52",
          3234 => x"b1",
          3235 => x"80",
          3236 => x"53",
          3237 => x"84",
          3238 => x"bd",
          3239 => x"80",
          3240 => x"82",
          3241 => x"81",
          3242 => x"a7",
          3243 => x"b6",
          3244 => x"fc",
          3245 => x"3d",
          3246 => x"51",
          3247 => x"82",
          3248 => x"b5",
          3249 => x"05",
          3250 => x"d6",
          3251 => x"82",
          3252 => x"52",
          3253 => x"a3",
          3254 => x"39",
          3255 => x"84",
          3256 => x"9a",
          3257 => x"dc",
          3258 => x"ff",
          3259 => x"5b",
          3260 => x"82",
          3261 => x"b5",
          3262 => x"05",
          3263 => x"a2",
          3264 => x"dc",
          3265 => x"ff",
          3266 => x"59",
          3267 => x"82",
          3268 => x"82",
          3269 => x"80",
          3270 => x"82",
          3271 => x"81",
          3272 => x"78",
          3273 => x"7a",
          3274 => x"3f",
          3275 => x"08",
          3276 => x"8d",
          3277 => x"dc",
          3278 => x"df",
          3279 => x"39",
          3280 => x"80",
          3281 => x"84",
          3282 => x"83",
          3283 => x"dc",
          3284 => x"fa",
          3285 => x"3d",
          3286 => x"53",
          3287 => x"51",
          3288 => x"82",
          3289 => x"80",
          3290 => x"38",
          3291 => x"f8",
          3292 => x"84",
          3293 => x"d7",
          3294 => x"dc",
          3295 => x"82",
          3296 => x"42",
          3297 => x"51",
          3298 => x"3f",
          3299 => x"5a",
          3300 => x"81",
          3301 => x"59",
          3302 => x"84",
          3303 => x"7a",
          3304 => x"38",
          3305 => x"b4",
          3306 => x"11",
          3307 => x"05",
          3308 => x"3f",
          3309 => x"08",
          3310 => x"85",
          3311 => x"fe",
          3312 => x"ff",
          3313 => x"e8",
          3314 => x"bb",
          3315 => x"2e",
          3316 => x"b4",
          3317 => x"11",
          3318 => x"05",
          3319 => x"3f",
          3320 => x"08",
          3321 => x"d9",
          3322 => x"c8",
          3323 => x"eb",
          3324 => x"79",
          3325 => x"89",
          3326 => x"79",
          3327 => x"5b",
          3328 => x"61",
          3329 => x"eb",
          3330 => x"ff",
          3331 => x"ff",
          3332 => x"e7",
          3333 => x"bb",
          3334 => x"2e",
          3335 => x"b4",
          3336 => x"11",
          3337 => x"05",
          3338 => x"3f",
          3339 => x"08",
          3340 => x"8d",
          3341 => x"fe",
          3342 => x"ff",
          3343 => x"e7",
          3344 => x"bb",
          3345 => x"2e",
          3346 => x"82",
          3347 => x"ff",
          3348 => x"63",
          3349 => x"27",
          3350 => x"70",
          3351 => x"5e",
          3352 => x"7c",
          3353 => x"78",
          3354 => x"79",
          3355 => x"52",
          3356 => x"51",
          3357 => x"3f",
          3358 => x"81",
          3359 => x"d5",
          3360 => x"ca",
          3361 => x"b9",
          3362 => x"ff",
          3363 => x"ff",
          3364 => x"e6",
          3365 => x"bb",
          3366 => x"df",
          3367 => x"c8",
          3368 => x"80",
          3369 => x"82",
          3370 => x"44",
          3371 => x"82",
          3372 => x"59",
          3373 => x"88",
          3374 => x"88",
          3375 => x"39",
          3376 => x"33",
          3377 => x"2e",
          3378 => x"ba",
          3379 => x"ab",
          3380 => x"cb",
          3381 => x"80",
          3382 => x"82",
          3383 => x"44",
          3384 => x"ba",
          3385 => x"78",
          3386 => x"38",
          3387 => x"08",
          3388 => x"82",
          3389 => x"fc",
          3390 => x"b4",
          3391 => x"11",
          3392 => x"05",
          3393 => x"3f",
          3394 => x"08",
          3395 => x"82",
          3396 => x"59",
          3397 => x"89",
          3398 => x"84",
          3399 => x"cc",
          3400 => x"c9",
          3401 => x"80",
          3402 => x"82",
          3403 => x"43",
          3404 => x"ba",
          3405 => x"78",
          3406 => x"38",
          3407 => x"08",
          3408 => x"82",
          3409 => x"59",
          3410 => x"88",
          3411 => x"9c",
          3412 => x"39",
          3413 => x"33",
          3414 => x"2e",
          3415 => x"ba",
          3416 => x"88",
          3417 => x"b0",
          3418 => x"43",
          3419 => x"f8",
          3420 => x"84",
          3421 => x"d7",
          3422 => x"dc",
          3423 => x"a7",
          3424 => x"5c",
          3425 => x"2e",
          3426 => x"5c",
          3427 => x"70",
          3428 => x"07",
          3429 => x"7f",
          3430 => x"5a",
          3431 => x"2e",
          3432 => x"a0",
          3433 => x"88",
          3434 => x"80",
          3435 => x"3f",
          3436 => x"54",
          3437 => x"52",
          3438 => x"c9",
          3439 => x"8c",
          3440 => x"39",
          3441 => x"80",
          3442 => x"84",
          3443 => x"ff",
          3444 => x"dc",
          3445 => x"f5",
          3446 => x"3d",
          3447 => x"53",
          3448 => x"51",
          3449 => x"82",
          3450 => x"80",
          3451 => x"63",
          3452 => x"cb",
          3453 => x"34",
          3454 => x"44",
          3455 => x"fc",
          3456 => x"84",
          3457 => x"c7",
          3458 => x"dc",
          3459 => x"f5",
          3460 => x"70",
          3461 => x"82",
          3462 => x"ff",
          3463 => x"82",
          3464 => x"53",
          3465 => x"79",
          3466 => x"84",
          3467 => x"79",
          3468 => x"ae",
          3469 => x"38",
          3470 => x"9f",
          3471 => x"fe",
          3472 => x"ff",
          3473 => x"e3",
          3474 => x"bb",
          3475 => x"2e",
          3476 => x"59",
          3477 => x"05",
          3478 => x"63",
          3479 => x"ff",
          3480 => x"a8",
          3481 => x"fe",
          3482 => x"39",
          3483 => x"f4",
          3484 => x"84",
          3485 => x"86",
          3486 => x"dc",
          3487 => x"f4",
          3488 => x"3d",
          3489 => x"53",
          3490 => x"51",
          3491 => x"82",
          3492 => x"80",
          3493 => x"60",
          3494 => x"05",
          3495 => x"82",
          3496 => x"78",
          3497 => x"fe",
          3498 => x"ff",
          3499 => x"dc",
          3500 => x"bb",
          3501 => x"38",
          3502 => x"60",
          3503 => x"52",
          3504 => x"51",
          3505 => x"3f",
          3506 => x"08",
          3507 => x"52",
          3508 => x"a6",
          3509 => x"45",
          3510 => x"78",
          3511 => x"e1",
          3512 => x"26",
          3513 => x"82",
          3514 => x"39",
          3515 => x"f0",
          3516 => x"84",
          3517 => x"86",
          3518 => x"dc",
          3519 => x"92",
          3520 => x"02",
          3521 => x"79",
          3522 => x"5b",
          3523 => x"ff",
          3524 => x"a8",
          3525 => x"ce",
          3526 => x"39",
          3527 => x"f4",
          3528 => x"84",
          3529 => x"d6",
          3530 => x"dc",
          3531 => x"f3",
          3532 => x"3d",
          3533 => x"53",
          3534 => x"51",
          3535 => x"82",
          3536 => x"80",
          3537 => x"60",
          3538 => x"59",
          3539 => x"41",
          3540 => x"f0",
          3541 => x"84",
          3542 => x"a2",
          3543 => x"dc",
          3544 => x"f2",
          3545 => x"70",
          3546 => x"82",
          3547 => x"ff",
          3548 => x"82",
          3549 => x"53",
          3550 => x"79",
          3551 => x"b0",
          3552 => x"79",
          3553 => x"ae",
          3554 => x"38",
          3555 => x"9b",
          3556 => x"fe",
          3557 => x"ff",
          3558 => x"da",
          3559 => x"bb",
          3560 => x"2e",
          3561 => x"60",
          3562 => x"60",
          3563 => x"ff",
          3564 => x"a8",
          3565 => x"ae",
          3566 => x"39",
          3567 => x"51",
          3568 => x"82",
          3569 => x"3f",
          3570 => x"82",
          3571 => x"c0",
          3572 => x"51",
          3573 => x"f1",
          3574 => x"a8",
          3575 => x"86",
          3576 => x"81",
          3577 => x"94",
          3578 => x"80",
          3579 => x"c0",
          3580 => x"f1",
          3581 => x"a9",
          3582 => x"bf",
          3583 => x"80",
          3584 => x"c0",
          3585 => x"8c",
          3586 => x"87",
          3587 => x"0c",
          3588 => x"b4",
          3589 => x"11",
          3590 => x"05",
          3591 => x"3f",
          3592 => x"08",
          3593 => x"99",
          3594 => x"82",
          3595 => x"ff",
          3596 => x"63",
          3597 => x"b4",
          3598 => x"11",
          3599 => x"05",
          3600 => x"3f",
          3601 => x"08",
          3602 => x"f5",
          3603 => x"82",
          3604 => x"ff",
          3605 => x"63",
          3606 => x"82",
          3607 => x"80",
          3608 => x"38",
          3609 => x"08",
          3610 => x"d0",
          3611 => x"eb",
          3612 => x"39",
          3613 => x"51",
          3614 => x"3f",
          3615 => x"3f",
          3616 => x"82",
          3617 => x"ff",
          3618 => x"80",
          3619 => x"39",
          3620 => x"f0",
          3621 => x"45",
          3622 => x"78",
          3623 => x"a1",
          3624 => x"06",
          3625 => x"2e",
          3626 => x"b4",
          3627 => x"05",
          3628 => x"3f",
          3629 => x"08",
          3630 => x"7b",
          3631 => x"38",
          3632 => x"89",
          3633 => x"2e",
          3634 => x"ca",
          3635 => x"2e",
          3636 => x"c2",
          3637 => x"9c",
          3638 => x"82",
          3639 => x"80",
          3640 => x"a4",
          3641 => x"ff",
          3642 => x"ff",
          3643 => x"b8",
          3644 => x"b4",
          3645 => x"05",
          3646 => x"3f",
          3647 => x"55",
          3648 => x"54",
          3649 => x"aa",
          3650 => x"3d",
          3651 => x"51",
          3652 => x"3f",
          3653 => x"54",
          3654 => x"aa",
          3655 => x"3d",
          3656 => x"51",
          3657 => x"3f",
          3658 => x"58",
          3659 => x"57",
          3660 => x"55",
          3661 => x"d8",
          3662 => x"d8",
          3663 => x"3d",
          3664 => x"51",
          3665 => x"82",
          3666 => x"82",
          3667 => x"09",
          3668 => x"72",
          3669 => x"51",
          3670 => x"80",
          3671 => x"26",
          3672 => x"5a",
          3673 => x"59",
          3674 => x"8d",
          3675 => x"70",
          3676 => x"5d",
          3677 => x"c3",
          3678 => x"32",
          3679 => x"07",
          3680 => x"38",
          3681 => x"09",
          3682 => x"b5",
          3683 => x"c8",
          3684 => x"d2",
          3685 => x"39",
          3686 => x"80",
          3687 => x"8c",
          3688 => x"94",
          3689 => x"54",
          3690 => x"80",
          3691 => x"d3",
          3692 => x"bb",
          3693 => x"2b",
          3694 => x"53",
          3695 => x"52",
          3696 => x"c2",
          3697 => x"bb",
          3698 => x"75",
          3699 => x"94",
          3700 => x"54",
          3701 => x"80",
          3702 => x"d3",
          3703 => x"bb",
          3704 => x"2b",
          3705 => x"53",
          3706 => x"52",
          3707 => x"96",
          3708 => x"bb",
          3709 => x"75",
          3710 => x"83",
          3711 => x"94",
          3712 => x"80",
          3713 => x"c0",
          3714 => x"80",
          3715 => x"80",
          3716 => x"83",
          3717 => x"99",
          3718 => x"5c",
          3719 => x"0b",
          3720 => x"88",
          3721 => x"72",
          3722 => x"b0",
          3723 => x"be",
          3724 => x"3f",
          3725 => x"51",
          3726 => x"3f",
          3727 => x"51",
          3728 => x"3f",
          3729 => x"51",
          3730 => x"81",
          3731 => x"3f",
          3732 => x"80",
          3733 => x"0d",
          3734 => x"53",
          3735 => x"52",
          3736 => x"82",
          3737 => x"81",
          3738 => x"07",
          3739 => x"52",
          3740 => x"e8",
          3741 => x"bb",
          3742 => x"3d",
          3743 => x"3d",
          3744 => x"08",
          3745 => x"73",
          3746 => x"74",
          3747 => x"38",
          3748 => x"70",
          3749 => x"81",
          3750 => x"81",
          3751 => x"39",
          3752 => x"70",
          3753 => x"81",
          3754 => x"81",
          3755 => x"54",
          3756 => x"81",
          3757 => x"06",
          3758 => x"39",
          3759 => x"80",
          3760 => x"54",
          3761 => x"83",
          3762 => x"70",
          3763 => x"38",
          3764 => x"98",
          3765 => x"52",
          3766 => x"52",
          3767 => x"2e",
          3768 => x"54",
          3769 => x"84",
          3770 => x"38",
          3771 => x"52",
          3772 => x"2e",
          3773 => x"83",
          3774 => x"70",
          3775 => x"30",
          3776 => x"76",
          3777 => x"51",
          3778 => x"88",
          3779 => x"70",
          3780 => x"34",
          3781 => x"72",
          3782 => x"bb",
          3783 => x"3d",
          3784 => x"3d",
          3785 => x"72",
          3786 => x"91",
          3787 => x"fc",
          3788 => x"51",
          3789 => x"82",
          3790 => x"85",
          3791 => x"83",
          3792 => x"72",
          3793 => x"0c",
          3794 => x"04",
          3795 => x"76",
          3796 => x"ff",
          3797 => x"81",
          3798 => x"26",
          3799 => x"83",
          3800 => x"05",
          3801 => x"70",
          3802 => x"8a",
          3803 => x"33",
          3804 => x"70",
          3805 => x"fe",
          3806 => x"33",
          3807 => x"70",
          3808 => x"f2",
          3809 => x"33",
          3810 => x"70",
          3811 => x"e6",
          3812 => x"22",
          3813 => x"74",
          3814 => x"80",
          3815 => x"13",
          3816 => x"52",
          3817 => x"26",
          3818 => x"81",
          3819 => x"98",
          3820 => x"22",
          3821 => x"bc",
          3822 => x"33",
          3823 => x"b8",
          3824 => x"33",
          3825 => x"b4",
          3826 => x"33",
          3827 => x"b0",
          3828 => x"33",
          3829 => x"ac",
          3830 => x"33",
          3831 => x"a8",
          3832 => x"c0",
          3833 => x"73",
          3834 => x"a0",
          3835 => x"87",
          3836 => x"0c",
          3837 => x"82",
          3838 => x"86",
          3839 => x"f3",
          3840 => x"5b",
          3841 => x"9c",
          3842 => x"0c",
          3843 => x"bc",
          3844 => x"7b",
          3845 => x"98",
          3846 => x"79",
          3847 => x"87",
          3848 => x"08",
          3849 => x"1c",
          3850 => x"98",
          3851 => x"79",
          3852 => x"87",
          3853 => x"08",
          3854 => x"1c",
          3855 => x"98",
          3856 => x"79",
          3857 => x"87",
          3858 => x"08",
          3859 => x"1c",
          3860 => x"98",
          3861 => x"79",
          3862 => x"80",
          3863 => x"83",
          3864 => x"59",
          3865 => x"ff",
          3866 => x"1b",
          3867 => x"1b",
          3868 => x"1b",
          3869 => x"1b",
          3870 => x"1b",
          3871 => x"83",
          3872 => x"52",
          3873 => x"51",
          3874 => x"3f",
          3875 => x"04",
          3876 => x"02",
          3877 => x"82",
          3878 => x"70",
          3879 => x"58",
          3880 => x"c0",
          3881 => x"75",
          3882 => x"38",
          3883 => x"94",
          3884 => x"70",
          3885 => x"81",
          3886 => x"52",
          3887 => x"8c",
          3888 => x"2a",
          3889 => x"51",
          3890 => x"38",
          3891 => x"70",
          3892 => x"51",
          3893 => x"8d",
          3894 => x"2a",
          3895 => x"51",
          3896 => x"be",
          3897 => x"ff",
          3898 => x"c0",
          3899 => x"70",
          3900 => x"38",
          3901 => x"90",
          3902 => x"0c",
          3903 => x"dc",
          3904 => x"0d",
          3905 => x"0d",
          3906 => x"33",
          3907 => x"9f",
          3908 => x"52",
          3909 => x"fc",
          3910 => x"0d",
          3911 => x"0d",
          3912 => x"33",
          3913 => x"2e",
          3914 => x"87",
          3915 => x"8d",
          3916 => x"82",
          3917 => x"70",
          3918 => x"58",
          3919 => x"94",
          3920 => x"80",
          3921 => x"87",
          3922 => x"53",
          3923 => x"96",
          3924 => x"06",
          3925 => x"72",
          3926 => x"38",
          3927 => x"70",
          3928 => x"53",
          3929 => x"74",
          3930 => x"81",
          3931 => x"72",
          3932 => x"38",
          3933 => x"70",
          3934 => x"53",
          3935 => x"38",
          3936 => x"06",
          3937 => x"94",
          3938 => x"80",
          3939 => x"87",
          3940 => x"54",
          3941 => x"80",
          3942 => x"dc",
          3943 => x"0d",
          3944 => x"0d",
          3945 => x"74",
          3946 => x"ff",
          3947 => x"57",
          3948 => x"80",
          3949 => x"81",
          3950 => x"15",
          3951 => x"33",
          3952 => x"06",
          3953 => x"58",
          3954 => x"84",
          3955 => x"2e",
          3956 => x"c0",
          3957 => x"70",
          3958 => x"2a",
          3959 => x"53",
          3960 => x"80",
          3961 => x"71",
          3962 => x"81",
          3963 => x"70",
          3964 => x"81",
          3965 => x"06",
          3966 => x"80",
          3967 => x"71",
          3968 => x"81",
          3969 => x"70",
          3970 => x"74",
          3971 => x"51",
          3972 => x"80",
          3973 => x"2e",
          3974 => x"c0",
          3975 => x"77",
          3976 => x"17",
          3977 => x"81",
          3978 => x"53",
          3979 => x"86",
          3980 => x"bb",
          3981 => x"3d",
          3982 => x"3d",
          3983 => x"fc",
          3984 => x"ff",
          3985 => x"87",
          3986 => x"51",
          3987 => x"86",
          3988 => x"94",
          3989 => x"08",
          3990 => x"70",
          3991 => x"51",
          3992 => x"2e",
          3993 => x"81",
          3994 => x"87",
          3995 => x"52",
          3996 => x"86",
          3997 => x"94",
          3998 => x"08",
          3999 => x"06",
          4000 => x"0c",
          4001 => x"0d",
          4002 => x"3f",
          4003 => x"08",
          4004 => x"82",
          4005 => x"04",
          4006 => x"82",
          4007 => x"70",
          4008 => x"52",
          4009 => x"94",
          4010 => x"80",
          4011 => x"87",
          4012 => x"52",
          4013 => x"82",
          4014 => x"06",
          4015 => x"ff",
          4016 => x"2e",
          4017 => x"81",
          4018 => x"87",
          4019 => x"52",
          4020 => x"86",
          4021 => x"94",
          4022 => x"08",
          4023 => x"70",
          4024 => x"53",
          4025 => x"bb",
          4026 => x"3d",
          4027 => x"3d",
          4028 => x"9e",
          4029 => x"9c",
          4030 => x"51",
          4031 => x"2e",
          4032 => x"87",
          4033 => x"08",
          4034 => x"0c",
          4035 => x"a8",
          4036 => x"84",
          4037 => x"9e",
          4038 => x"ba",
          4039 => x"c0",
          4040 => x"82",
          4041 => x"87",
          4042 => x"08",
          4043 => x"0c",
          4044 => x"a0",
          4045 => x"94",
          4046 => x"9e",
          4047 => x"ba",
          4048 => x"c0",
          4049 => x"82",
          4050 => x"87",
          4051 => x"08",
          4052 => x"0c",
          4053 => x"b8",
          4054 => x"a4",
          4055 => x"9e",
          4056 => x"ba",
          4057 => x"c0",
          4058 => x"82",
          4059 => x"87",
          4060 => x"08",
          4061 => x"0c",
          4062 => x"80",
          4063 => x"82",
          4064 => x"87",
          4065 => x"08",
          4066 => x"0c",
          4067 => x"88",
          4068 => x"bc",
          4069 => x"9e",
          4070 => x"ba",
          4071 => x"0b",
          4072 => x"34",
          4073 => x"c0",
          4074 => x"70",
          4075 => x"06",
          4076 => x"70",
          4077 => x"38",
          4078 => x"82",
          4079 => x"80",
          4080 => x"9e",
          4081 => x"88",
          4082 => x"51",
          4083 => x"80",
          4084 => x"81",
          4085 => x"ba",
          4086 => x"0b",
          4087 => x"90",
          4088 => x"80",
          4089 => x"52",
          4090 => x"2e",
          4091 => x"52",
          4092 => x"c7",
          4093 => x"87",
          4094 => x"08",
          4095 => x"80",
          4096 => x"52",
          4097 => x"83",
          4098 => x"71",
          4099 => x"34",
          4100 => x"c0",
          4101 => x"70",
          4102 => x"06",
          4103 => x"70",
          4104 => x"38",
          4105 => x"82",
          4106 => x"80",
          4107 => x"9e",
          4108 => x"90",
          4109 => x"51",
          4110 => x"80",
          4111 => x"81",
          4112 => x"ba",
          4113 => x"0b",
          4114 => x"90",
          4115 => x"80",
          4116 => x"52",
          4117 => x"2e",
          4118 => x"52",
          4119 => x"cb",
          4120 => x"87",
          4121 => x"08",
          4122 => x"80",
          4123 => x"52",
          4124 => x"83",
          4125 => x"71",
          4126 => x"34",
          4127 => x"c0",
          4128 => x"70",
          4129 => x"06",
          4130 => x"70",
          4131 => x"38",
          4132 => x"82",
          4133 => x"80",
          4134 => x"9e",
          4135 => x"80",
          4136 => x"51",
          4137 => x"80",
          4138 => x"81",
          4139 => x"ba",
          4140 => x"0b",
          4141 => x"90",
          4142 => x"80",
          4143 => x"52",
          4144 => x"83",
          4145 => x"71",
          4146 => x"34",
          4147 => x"90",
          4148 => x"80",
          4149 => x"2a",
          4150 => x"70",
          4151 => x"34",
          4152 => x"c0",
          4153 => x"70",
          4154 => x"51",
          4155 => x"80",
          4156 => x"81",
          4157 => x"ba",
          4158 => x"c0",
          4159 => x"70",
          4160 => x"70",
          4161 => x"51",
          4162 => x"ba",
          4163 => x"0b",
          4164 => x"90",
          4165 => x"06",
          4166 => x"70",
          4167 => x"38",
          4168 => x"82",
          4169 => x"87",
          4170 => x"08",
          4171 => x"51",
          4172 => x"ba",
          4173 => x"3d",
          4174 => x"3d",
          4175 => x"94",
          4176 => x"a2",
          4177 => x"c4",
          4178 => x"80",
          4179 => x"82",
          4180 => x"ff",
          4181 => x"82",
          4182 => x"ff",
          4183 => x"82",
          4184 => x"54",
          4185 => x"94",
          4186 => x"a0",
          4187 => x"a4",
          4188 => x"52",
          4189 => x"51",
          4190 => x"3f",
          4191 => x"33",
          4192 => x"2e",
          4193 => x"ba",
          4194 => x"ba",
          4195 => x"54",
          4196 => x"f0",
          4197 => x"c3",
          4198 => x"c8",
          4199 => x"80",
          4200 => x"82",
          4201 => x"82",
          4202 => x"11",
          4203 => x"ac",
          4204 => x"90",
          4205 => x"ba",
          4206 => x"73",
          4207 => x"38",
          4208 => x"08",
          4209 => x"08",
          4210 => x"82",
          4211 => x"ff",
          4212 => x"82",
          4213 => x"54",
          4214 => x"94",
          4215 => x"90",
          4216 => x"94",
          4217 => x"52",
          4218 => x"51",
          4219 => x"3f",
          4220 => x"33",
          4221 => x"2e",
          4222 => x"ba",
          4223 => x"82",
          4224 => x"ff",
          4225 => x"82",
          4226 => x"54",
          4227 => x"8e",
          4228 => x"d4",
          4229 => x"ad",
          4230 => x"8f",
          4231 => x"ba",
          4232 => x"73",
          4233 => x"38",
          4234 => x"33",
          4235 => x"a0",
          4236 => x"a7",
          4237 => x"c5",
          4238 => x"80",
          4239 => x"82",
          4240 => x"ff",
          4241 => x"82",
          4242 => x"54",
          4243 => x"89",
          4244 => x"d4",
          4245 => x"8e",
          4246 => x"cc",
          4247 => x"80",
          4248 => x"82",
          4249 => x"ff",
          4250 => x"82",
          4251 => x"54",
          4252 => x"89",
          4253 => x"ec",
          4254 => x"ea",
          4255 => x"ce",
          4256 => x"80",
          4257 => x"82",
          4258 => x"ff",
          4259 => x"82",
          4260 => x"ff",
          4261 => x"82",
          4262 => x"52",
          4263 => x"51",
          4264 => x"3f",
          4265 => x"08",
          4266 => x"b8",
          4267 => x"ab",
          4268 => x"b0",
          4269 => x"ae",
          4270 => x"8e",
          4271 => x"af",
          4272 => x"aa",
          4273 => x"ba",
          4274 => x"82",
          4275 => x"ff",
          4276 => x"82",
          4277 => x"56",
          4278 => x"52",
          4279 => x"a6",
          4280 => x"dc",
          4281 => x"c0",
          4282 => x"31",
          4283 => x"bb",
          4284 => x"82",
          4285 => x"ff",
          4286 => x"82",
          4287 => x"54",
          4288 => x"a9",
          4289 => x"bc",
          4290 => x"84",
          4291 => x"51",
          4292 => x"82",
          4293 => x"bd",
          4294 => x"76",
          4295 => x"54",
          4296 => x"08",
          4297 => x"e4",
          4298 => x"af",
          4299 => x"c6",
          4300 => x"80",
          4301 => x"82",
          4302 => x"56",
          4303 => x"52",
          4304 => x"c2",
          4305 => x"dc",
          4306 => x"c0",
          4307 => x"31",
          4308 => x"bb",
          4309 => x"82",
          4310 => x"ff",
          4311 => x"82",
          4312 => x"ff",
          4313 => x"87",
          4314 => x"fe",
          4315 => x"92",
          4316 => x"05",
          4317 => x"26",
          4318 => x"84",
          4319 => x"ec",
          4320 => x"08",
          4321 => x"bc",
          4322 => x"82",
          4323 => x"97",
          4324 => x"cc",
          4325 => x"82",
          4326 => x"8b",
          4327 => x"d8",
          4328 => x"82",
          4329 => x"ff",
          4330 => x"84",
          4331 => x"71",
          4332 => x"04",
          4333 => x"87",
          4334 => x"70",
          4335 => x"80",
          4336 => x"74",
          4337 => x"ba",
          4338 => x"0c",
          4339 => x"04",
          4340 => x"87",
          4341 => x"70",
          4342 => x"d8",
          4343 => x"72",
          4344 => x"70",
          4345 => x"08",
          4346 => x"ba",
          4347 => x"0c",
          4348 => x"0d",
          4349 => x"87",
          4350 => x"0c",
          4351 => x"d8",
          4352 => x"96",
          4353 => x"fd",
          4354 => x"98",
          4355 => x"2c",
          4356 => x"70",
          4357 => x"10",
          4358 => x"2b",
          4359 => x"54",
          4360 => x"0b",
          4361 => x"12",
          4362 => x"71",
          4363 => x"38",
          4364 => x"11",
          4365 => x"84",
          4366 => x"33",
          4367 => x"52",
          4368 => x"2e",
          4369 => x"83",
          4370 => x"72",
          4371 => x"0c",
          4372 => x"04",
          4373 => x"79",
          4374 => x"a3",
          4375 => x"33",
          4376 => x"72",
          4377 => x"38",
          4378 => x"08",
          4379 => x"ff",
          4380 => x"82",
          4381 => x"52",
          4382 => x"aa",
          4383 => x"d3",
          4384 => x"88",
          4385 => x"ad",
          4386 => x"ff",
          4387 => x"74",
          4388 => x"ff",
          4389 => x"39",
          4390 => x"8a",
          4391 => x"74",
          4392 => x"0d",
          4393 => x"0d",
          4394 => x"05",
          4395 => x"02",
          4396 => x"05",
          4397 => x"b4",
          4398 => x"29",
          4399 => x"05",
          4400 => x"59",
          4401 => x"59",
          4402 => x"86",
          4403 => x"9a",
          4404 => x"bb",
          4405 => x"84",
          4406 => x"dc",
          4407 => x"70",
          4408 => x"5a",
          4409 => x"82",
          4410 => x"75",
          4411 => x"b4",
          4412 => x"29",
          4413 => x"05",
          4414 => x"56",
          4415 => x"2e",
          4416 => x"53",
          4417 => x"51",
          4418 => x"3f",
          4419 => x"33",
          4420 => x"74",
          4421 => x"34",
          4422 => x"06",
          4423 => x"27",
          4424 => x"0b",
          4425 => x"34",
          4426 => x"b6",
          4427 => x"b0",
          4428 => x"80",
          4429 => x"82",
          4430 => x"55",
          4431 => x"8c",
          4432 => x"54",
          4433 => x"52",
          4434 => x"da",
          4435 => x"bb",
          4436 => x"8a",
          4437 => x"95",
          4438 => x"b0",
          4439 => x"dd",
          4440 => x"3d",
          4441 => x"3d",
          4442 => x"dc",
          4443 => x"72",
          4444 => x"80",
          4445 => x"71",
          4446 => x"3f",
          4447 => x"ff",
          4448 => x"54",
          4449 => x"25",
          4450 => x"0b",
          4451 => x"34",
          4452 => x"08",
          4453 => x"2e",
          4454 => x"51",
          4455 => x"3f",
          4456 => x"08",
          4457 => x"3f",
          4458 => x"bb",
          4459 => x"3d",
          4460 => x"3d",
          4461 => x"80",
          4462 => x"b0",
          4463 => x"e3",
          4464 => x"bb",
          4465 => x"d3",
          4466 => x"b0",
          4467 => x"f8",
          4468 => x"70",
          4469 => x"8c",
          4470 => x"bb",
          4471 => x"2e",
          4472 => x"51",
          4473 => x"3f",
          4474 => x"08",
          4475 => x"82",
          4476 => x"25",
          4477 => x"bb",
          4478 => x"05",
          4479 => x"55",
          4480 => x"75",
          4481 => x"81",
          4482 => x"dc",
          4483 => x"87",
          4484 => x"ff",
          4485 => x"06",
          4486 => x"a6",
          4487 => x"d9",
          4488 => x"3d",
          4489 => x"08",
          4490 => x"70",
          4491 => x"52",
          4492 => x"08",
          4493 => x"bb",
          4494 => x"dc",
          4495 => x"38",
          4496 => x"bb",
          4497 => x"55",
          4498 => x"8b",
          4499 => x"56",
          4500 => x"3f",
          4501 => x"08",
          4502 => x"38",
          4503 => x"af",
          4504 => x"bb",
          4505 => x"18",
          4506 => x"0b",
          4507 => x"08",
          4508 => x"82",
          4509 => x"ff",
          4510 => x"55",
          4511 => x"34",
          4512 => x"30",
          4513 => x"9f",
          4514 => x"55",
          4515 => x"85",
          4516 => x"ac",
          4517 => x"b0",
          4518 => x"08",
          4519 => x"e1",
          4520 => x"bb",
          4521 => x"2e",
          4522 => x"b3",
          4523 => x"86",
          4524 => x"77",
          4525 => x"06",
          4526 => x"52",
          4527 => x"af",
          4528 => x"51",
          4529 => x"3f",
          4530 => x"54",
          4531 => x"08",
          4532 => x"58",
          4533 => x"dc",
          4534 => x"0d",
          4535 => x"0d",
          4536 => x"5c",
          4537 => x"57",
          4538 => x"73",
          4539 => x"81",
          4540 => x"78",
          4541 => x"56",
          4542 => x"98",
          4543 => x"70",
          4544 => x"33",
          4545 => x"73",
          4546 => x"81",
          4547 => x"75",
          4548 => x"38",
          4549 => x"88",
          4550 => x"b8",
          4551 => x"52",
          4552 => x"e4",
          4553 => x"dc",
          4554 => x"52",
          4555 => x"ff",
          4556 => x"82",
          4557 => x"80",
          4558 => x"15",
          4559 => x"81",
          4560 => x"74",
          4561 => x"38",
          4562 => x"e6",
          4563 => x"81",
          4564 => x"3d",
          4565 => x"f8",
          4566 => x"f3",
          4567 => x"dc",
          4568 => x"9a",
          4569 => x"53",
          4570 => x"51",
          4571 => x"82",
          4572 => x"81",
          4573 => x"74",
          4574 => x"54",
          4575 => x"14",
          4576 => x"06",
          4577 => x"74",
          4578 => x"38",
          4579 => x"82",
          4580 => x"8c",
          4581 => x"d3",
          4582 => x"3d",
          4583 => x"08",
          4584 => x"59",
          4585 => x"0b",
          4586 => x"82",
          4587 => x"82",
          4588 => x"55",
          4589 => x"cb",
          4590 => x"bb",
          4591 => x"55",
          4592 => x"81",
          4593 => x"2e",
          4594 => x"81",
          4595 => x"55",
          4596 => x"2e",
          4597 => x"a8",
          4598 => x"3f",
          4599 => x"08",
          4600 => x"0c",
          4601 => x"08",
          4602 => x"92",
          4603 => x"76",
          4604 => x"dc",
          4605 => x"cc",
          4606 => x"bb",
          4607 => x"2e",
          4608 => x"b4",
          4609 => x"9f",
          4610 => x"f7",
          4611 => x"dc",
          4612 => x"bb",
          4613 => x"80",
          4614 => x"3d",
          4615 => x"81",
          4616 => x"82",
          4617 => x"56",
          4618 => x"08",
          4619 => x"81",
          4620 => x"38",
          4621 => x"08",
          4622 => x"cc",
          4623 => x"dc",
          4624 => x"0b",
          4625 => x"08",
          4626 => x"82",
          4627 => x"ff",
          4628 => x"55",
          4629 => x"34",
          4630 => x"81",
          4631 => x"75",
          4632 => x"3f",
          4633 => x"81",
          4634 => x"54",
          4635 => x"83",
          4636 => x"74",
          4637 => x"81",
          4638 => x"38",
          4639 => x"82",
          4640 => x"76",
          4641 => x"bb",
          4642 => x"2e",
          4643 => x"d6",
          4644 => x"5d",
          4645 => x"82",
          4646 => x"98",
          4647 => x"2c",
          4648 => x"ff",
          4649 => x"78",
          4650 => x"82",
          4651 => x"70",
          4652 => x"98",
          4653 => x"84",
          4654 => x"2b",
          4655 => x"71",
          4656 => x"70",
          4657 => x"b0",
          4658 => x"08",
          4659 => x"51",
          4660 => x"59",
          4661 => x"5d",
          4662 => x"73",
          4663 => x"e9",
          4664 => x"27",
          4665 => x"81",
          4666 => x"81",
          4667 => x"70",
          4668 => x"55",
          4669 => x"80",
          4670 => x"53",
          4671 => x"51",
          4672 => x"82",
          4673 => x"81",
          4674 => x"73",
          4675 => x"38",
          4676 => x"84",
          4677 => x"b1",
          4678 => x"80",
          4679 => x"80",
          4680 => x"98",
          4681 => x"ff",
          4682 => x"55",
          4683 => x"97",
          4684 => x"74",
          4685 => x"f5",
          4686 => x"bb",
          4687 => x"ff",
          4688 => x"cc",
          4689 => x"80",
          4690 => x"2e",
          4691 => x"81",
          4692 => x"82",
          4693 => x"74",
          4694 => x"98",
          4695 => x"84",
          4696 => x"2b",
          4697 => x"70",
          4698 => x"82",
          4699 => x"ec",
          4700 => x"51",
          4701 => x"58",
          4702 => x"77",
          4703 => x"06",
          4704 => x"82",
          4705 => x"08",
          4706 => x"0b",
          4707 => x"34",
          4708 => x"d3",
          4709 => x"39",
          4710 => x"88",
          4711 => x"d3",
          4712 => x"af",
          4713 => x"7d",
          4714 => x"73",
          4715 => x"e1",
          4716 => x"29",
          4717 => x"05",
          4718 => x"04",
          4719 => x"33",
          4720 => x"2e",
          4721 => x"82",
          4722 => x"55",
          4723 => x"ab",
          4724 => x"2b",
          4725 => x"51",
          4726 => x"24",
          4727 => x"1a",
          4728 => x"81",
          4729 => x"81",
          4730 => x"81",
          4731 => x"70",
          4732 => x"d3",
          4733 => x"51",
          4734 => x"82",
          4735 => x"81",
          4736 => x"74",
          4737 => x"34",
          4738 => x"ae",
          4739 => x"34",
          4740 => x"33",
          4741 => x"25",
          4742 => x"14",
          4743 => x"d3",
          4744 => x"d3",
          4745 => x"81",
          4746 => x"81",
          4747 => x"70",
          4748 => x"d3",
          4749 => x"51",
          4750 => x"77",
          4751 => x"82",
          4752 => x"52",
          4753 => x"33",
          4754 => x"9e",
          4755 => x"81",
          4756 => x"81",
          4757 => x"70",
          4758 => x"d3",
          4759 => x"51",
          4760 => x"24",
          4761 => x"d3",
          4762 => x"98",
          4763 => x"2c",
          4764 => x"33",
          4765 => x"56",
          4766 => x"fc",
          4767 => x"d3",
          4768 => x"88",
          4769 => x"ad",
          4770 => x"80",
          4771 => x"80",
          4772 => x"98",
          4773 => x"8c",
          4774 => x"55",
          4775 => x"de",
          4776 => x"39",
          4777 => x"80",
          4778 => x"34",
          4779 => x"53",
          4780 => x"a3",
          4781 => x"9c",
          4782 => x"39",
          4783 => x"33",
          4784 => x"06",
          4785 => x"80",
          4786 => x"38",
          4787 => x"33",
          4788 => x"73",
          4789 => x"34",
          4790 => x"73",
          4791 => x"34",
          4792 => x"08",
          4793 => x"ff",
          4794 => x"82",
          4795 => x"70",
          4796 => x"98",
          4797 => x"8c",
          4798 => x"56",
          4799 => x"25",
          4800 => x"1a",
          4801 => x"33",
          4802 => x"d3",
          4803 => x"73",
          4804 => x"9d",
          4805 => x"81",
          4806 => x"81",
          4807 => x"70",
          4808 => x"d3",
          4809 => x"51",
          4810 => x"24",
          4811 => x"d3",
          4812 => x"a0",
          4813 => x"fd",
          4814 => x"90",
          4815 => x"2b",
          4816 => x"82",
          4817 => x"57",
          4818 => x"74",
          4819 => x"c1",
          4820 => x"b0",
          4821 => x"51",
          4822 => x"3f",
          4823 => x"0a",
          4824 => x"0a",
          4825 => x"2c",
          4826 => x"33",
          4827 => x"75",
          4828 => x"38",
          4829 => x"82",
          4830 => x"7a",
          4831 => x"74",
          4832 => x"b0",
          4833 => x"51",
          4834 => x"3f",
          4835 => x"52",
          4836 => x"c9",
          4837 => x"dc",
          4838 => x"06",
          4839 => x"38",
          4840 => x"33",
          4841 => x"2e",
          4842 => x"53",
          4843 => x"51",
          4844 => x"84",
          4845 => x"34",
          4846 => x"d3",
          4847 => x"0b",
          4848 => x"34",
          4849 => x"dc",
          4850 => x"0d",
          4851 => x"90",
          4852 => x"80",
          4853 => x"38",
          4854 => x"08",
          4855 => x"ff",
          4856 => x"82",
          4857 => x"ff",
          4858 => x"82",
          4859 => x"73",
          4860 => x"54",
          4861 => x"d3",
          4862 => x"d3",
          4863 => x"55",
          4864 => x"f9",
          4865 => x"14",
          4866 => x"d3",
          4867 => x"98",
          4868 => x"2c",
          4869 => x"06",
          4870 => x"74",
          4871 => x"38",
          4872 => x"81",
          4873 => x"34",
          4874 => x"08",
          4875 => x"51",
          4876 => x"3f",
          4877 => x"0a",
          4878 => x"0a",
          4879 => x"2c",
          4880 => x"33",
          4881 => x"75",
          4882 => x"38",
          4883 => x"08",
          4884 => x"ff",
          4885 => x"82",
          4886 => x"70",
          4887 => x"98",
          4888 => x"8c",
          4889 => x"56",
          4890 => x"24",
          4891 => x"82",
          4892 => x"52",
          4893 => x"9a",
          4894 => x"81",
          4895 => x"81",
          4896 => x"70",
          4897 => x"d3",
          4898 => x"51",
          4899 => x"25",
          4900 => x"fd",
          4901 => x"90",
          4902 => x"ff",
          4903 => x"8c",
          4904 => x"54",
          4905 => x"f7",
          4906 => x"d3",
          4907 => x"81",
          4908 => x"82",
          4909 => x"74",
          4910 => x"52",
          4911 => x"f5",
          4912 => x"90",
          4913 => x"ff",
          4914 => x"8c",
          4915 => x"54",
          4916 => x"d6",
          4917 => x"39",
          4918 => x"53",
          4919 => x"a3",
          4920 => x"f0",
          4921 => x"82",
          4922 => x"80",
          4923 => x"8c",
          4924 => x"39",
          4925 => x"82",
          4926 => x"55",
          4927 => x"a6",
          4928 => x"ff",
          4929 => x"82",
          4930 => x"82",
          4931 => x"82",
          4932 => x"81",
          4933 => x"05",
          4934 => x"79",
          4935 => x"c8",
          4936 => x"81",
          4937 => x"84",
          4938 => x"dc",
          4939 => x"08",
          4940 => x"80",
          4941 => x"74",
          4942 => x"cc",
          4943 => x"dc",
          4944 => x"8c",
          4945 => x"dc",
          4946 => x"06",
          4947 => x"74",
          4948 => x"ff",
          4949 => x"ff",
          4950 => x"fa",
          4951 => x"55",
          4952 => x"f6",
          4953 => x"51",
          4954 => x"3f",
          4955 => x"93",
          4956 => x"06",
          4957 => x"ba",
          4958 => x"74",
          4959 => x"38",
          4960 => x"a1",
          4961 => x"bb",
          4962 => x"d3",
          4963 => x"bb",
          4964 => x"ff",
          4965 => x"53",
          4966 => x"51",
          4967 => x"3f",
          4968 => x"7a",
          4969 => x"ba",
          4970 => x"08",
          4971 => x"80",
          4972 => x"74",
          4973 => x"d0",
          4974 => x"dc",
          4975 => x"8c",
          4976 => x"dc",
          4977 => x"06",
          4978 => x"74",
          4979 => x"ff",
          4980 => x"81",
          4981 => x"81",
          4982 => x"89",
          4983 => x"d3",
          4984 => x"7a",
          4985 => x"90",
          4986 => x"8c",
          4987 => x"51",
          4988 => x"f5",
          4989 => x"d3",
          4990 => x"81",
          4991 => x"d3",
          4992 => x"56",
          4993 => x"27",
          4994 => x"82",
          4995 => x"52",
          4996 => x"73",
          4997 => x"34",
          4998 => x"33",
          4999 => x"97",
          5000 => x"ed",
          5001 => x"90",
          5002 => x"80",
          5003 => x"38",
          5004 => x"08",
          5005 => x"ff",
          5006 => x"82",
          5007 => x"ff",
          5008 => x"82",
          5009 => x"f4",
          5010 => x"3d",
          5011 => x"80",
          5012 => x"d4",
          5013 => x"0b",
          5014 => x"23",
          5015 => x"80",
          5016 => x"80",
          5017 => x"81",
          5018 => x"d4",
          5019 => x"58",
          5020 => x"81",
          5021 => x"15",
          5022 => x"d4",
          5023 => x"84",
          5024 => x"85",
          5025 => x"bb",
          5026 => x"77",
          5027 => x"76",
          5028 => x"82",
          5029 => x"82",
          5030 => x"ff",
          5031 => x"80",
          5032 => x"ff",
          5033 => x"88",
          5034 => x"55",
          5035 => x"17",
          5036 => x"17",
          5037 => x"d0",
          5038 => x"29",
          5039 => x"08",
          5040 => x"51",
          5041 => x"82",
          5042 => x"83",
          5043 => x"3d",
          5044 => x"3d",
          5045 => x"81",
          5046 => x"27",
          5047 => x"12",
          5048 => x"11",
          5049 => x"ff",
          5050 => x"51",
          5051 => x"dc",
          5052 => x"0d",
          5053 => x"0d",
          5054 => x"22",
          5055 => x"aa",
          5056 => x"05",
          5057 => x"08",
          5058 => x"71",
          5059 => x"2b",
          5060 => x"33",
          5061 => x"71",
          5062 => x"02",
          5063 => x"05",
          5064 => x"ff",
          5065 => x"70",
          5066 => x"51",
          5067 => x"5b",
          5068 => x"54",
          5069 => x"34",
          5070 => x"34",
          5071 => x"08",
          5072 => x"2a",
          5073 => x"82",
          5074 => x"83",
          5075 => x"bb",
          5076 => x"17",
          5077 => x"12",
          5078 => x"2b",
          5079 => x"2b",
          5080 => x"06",
          5081 => x"52",
          5082 => x"83",
          5083 => x"70",
          5084 => x"54",
          5085 => x"12",
          5086 => x"ff",
          5087 => x"83",
          5088 => x"bb",
          5089 => x"56",
          5090 => x"72",
          5091 => x"89",
          5092 => x"fb",
          5093 => x"bb",
          5094 => x"84",
          5095 => x"22",
          5096 => x"72",
          5097 => x"33",
          5098 => x"71",
          5099 => x"83",
          5100 => x"5b",
          5101 => x"52",
          5102 => x"12",
          5103 => x"33",
          5104 => x"07",
          5105 => x"54",
          5106 => x"70",
          5107 => x"73",
          5108 => x"82",
          5109 => x"70",
          5110 => x"33",
          5111 => x"71",
          5112 => x"83",
          5113 => x"59",
          5114 => x"05",
          5115 => x"87",
          5116 => x"88",
          5117 => x"88",
          5118 => x"56",
          5119 => x"13",
          5120 => x"13",
          5121 => x"d4",
          5122 => x"33",
          5123 => x"71",
          5124 => x"70",
          5125 => x"06",
          5126 => x"53",
          5127 => x"53",
          5128 => x"70",
          5129 => x"87",
          5130 => x"fa",
          5131 => x"a2",
          5132 => x"bb",
          5133 => x"83",
          5134 => x"70",
          5135 => x"33",
          5136 => x"07",
          5137 => x"15",
          5138 => x"12",
          5139 => x"2b",
          5140 => x"07",
          5141 => x"55",
          5142 => x"57",
          5143 => x"80",
          5144 => x"38",
          5145 => x"ab",
          5146 => x"d4",
          5147 => x"70",
          5148 => x"33",
          5149 => x"71",
          5150 => x"74",
          5151 => x"81",
          5152 => x"88",
          5153 => x"83",
          5154 => x"f8",
          5155 => x"54",
          5156 => x"58",
          5157 => x"74",
          5158 => x"52",
          5159 => x"34",
          5160 => x"34",
          5161 => x"08",
          5162 => x"33",
          5163 => x"71",
          5164 => x"83",
          5165 => x"59",
          5166 => x"05",
          5167 => x"12",
          5168 => x"2b",
          5169 => x"ff",
          5170 => x"88",
          5171 => x"52",
          5172 => x"74",
          5173 => x"15",
          5174 => x"0d",
          5175 => x"0d",
          5176 => x"08",
          5177 => x"9e",
          5178 => x"83",
          5179 => x"82",
          5180 => x"12",
          5181 => x"2b",
          5182 => x"07",
          5183 => x"52",
          5184 => x"05",
          5185 => x"13",
          5186 => x"2b",
          5187 => x"05",
          5188 => x"71",
          5189 => x"2a",
          5190 => x"53",
          5191 => x"34",
          5192 => x"34",
          5193 => x"08",
          5194 => x"33",
          5195 => x"71",
          5196 => x"83",
          5197 => x"59",
          5198 => x"05",
          5199 => x"83",
          5200 => x"88",
          5201 => x"88",
          5202 => x"56",
          5203 => x"13",
          5204 => x"13",
          5205 => x"d4",
          5206 => x"11",
          5207 => x"33",
          5208 => x"07",
          5209 => x"0c",
          5210 => x"3d",
          5211 => x"3d",
          5212 => x"bb",
          5213 => x"83",
          5214 => x"ff",
          5215 => x"53",
          5216 => x"a7",
          5217 => x"d4",
          5218 => x"2b",
          5219 => x"11",
          5220 => x"33",
          5221 => x"71",
          5222 => x"75",
          5223 => x"81",
          5224 => x"98",
          5225 => x"2b",
          5226 => x"40",
          5227 => x"58",
          5228 => x"72",
          5229 => x"38",
          5230 => x"52",
          5231 => x"9d",
          5232 => x"39",
          5233 => x"85",
          5234 => x"8b",
          5235 => x"2b",
          5236 => x"79",
          5237 => x"51",
          5238 => x"76",
          5239 => x"75",
          5240 => x"56",
          5241 => x"34",
          5242 => x"08",
          5243 => x"12",
          5244 => x"33",
          5245 => x"07",
          5246 => x"54",
          5247 => x"53",
          5248 => x"34",
          5249 => x"34",
          5250 => x"08",
          5251 => x"0b",
          5252 => x"80",
          5253 => x"34",
          5254 => x"08",
          5255 => x"14",
          5256 => x"14",
          5257 => x"d4",
          5258 => x"33",
          5259 => x"71",
          5260 => x"70",
          5261 => x"07",
          5262 => x"53",
          5263 => x"54",
          5264 => x"72",
          5265 => x"8b",
          5266 => x"ff",
          5267 => x"52",
          5268 => x"08",
          5269 => x"f2",
          5270 => x"2e",
          5271 => x"51",
          5272 => x"83",
          5273 => x"f5",
          5274 => x"7e",
          5275 => x"e2",
          5276 => x"dc",
          5277 => x"ff",
          5278 => x"d4",
          5279 => x"33",
          5280 => x"71",
          5281 => x"70",
          5282 => x"58",
          5283 => x"ff",
          5284 => x"2e",
          5285 => x"75",
          5286 => x"70",
          5287 => x"33",
          5288 => x"07",
          5289 => x"ff",
          5290 => x"70",
          5291 => x"06",
          5292 => x"52",
          5293 => x"59",
          5294 => x"27",
          5295 => x"80",
          5296 => x"75",
          5297 => x"84",
          5298 => x"16",
          5299 => x"2b",
          5300 => x"75",
          5301 => x"81",
          5302 => x"85",
          5303 => x"59",
          5304 => x"83",
          5305 => x"d4",
          5306 => x"33",
          5307 => x"71",
          5308 => x"70",
          5309 => x"06",
          5310 => x"56",
          5311 => x"75",
          5312 => x"81",
          5313 => x"79",
          5314 => x"cc",
          5315 => x"74",
          5316 => x"c4",
          5317 => x"2e",
          5318 => x"89",
          5319 => x"f8",
          5320 => x"ac",
          5321 => x"80",
          5322 => x"75",
          5323 => x"3f",
          5324 => x"08",
          5325 => x"11",
          5326 => x"33",
          5327 => x"71",
          5328 => x"53",
          5329 => x"74",
          5330 => x"70",
          5331 => x"06",
          5332 => x"5c",
          5333 => x"78",
          5334 => x"76",
          5335 => x"57",
          5336 => x"34",
          5337 => x"08",
          5338 => x"71",
          5339 => x"86",
          5340 => x"12",
          5341 => x"2b",
          5342 => x"2a",
          5343 => x"53",
          5344 => x"73",
          5345 => x"75",
          5346 => x"82",
          5347 => x"70",
          5348 => x"33",
          5349 => x"71",
          5350 => x"83",
          5351 => x"5d",
          5352 => x"05",
          5353 => x"15",
          5354 => x"15",
          5355 => x"d4",
          5356 => x"71",
          5357 => x"33",
          5358 => x"71",
          5359 => x"70",
          5360 => x"5a",
          5361 => x"54",
          5362 => x"34",
          5363 => x"34",
          5364 => x"08",
          5365 => x"54",
          5366 => x"dc",
          5367 => x"0d",
          5368 => x"0d",
          5369 => x"bb",
          5370 => x"38",
          5371 => x"71",
          5372 => x"2e",
          5373 => x"51",
          5374 => x"82",
          5375 => x"53",
          5376 => x"dc",
          5377 => x"0d",
          5378 => x"0d",
          5379 => x"5c",
          5380 => x"40",
          5381 => x"08",
          5382 => x"81",
          5383 => x"f4",
          5384 => x"8e",
          5385 => x"ff",
          5386 => x"bb",
          5387 => x"83",
          5388 => x"8b",
          5389 => x"fc",
          5390 => x"54",
          5391 => x"7e",
          5392 => x"3f",
          5393 => x"08",
          5394 => x"06",
          5395 => x"08",
          5396 => x"83",
          5397 => x"ff",
          5398 => x"83",
          5399 => x"70",
          5400 => x"33",
          5401 => x"07",
          5402 => x"70",
          5403 => x"06",
          5404 => x"fc",
          5405 => x"29",
          5406 => x"81",
          5407 => x"88",
          5408 => x"90",
          5409 => x"4e",
          5410 => x"52",
          5411 => x"41",
          5412 => x"5b",
          5413 => x"8f",
          5414 => x"ff",
          5415 => x"31",
          5416 => x"ff",
          5417 => x"82",
          5418 => x"17",
          5419 => x"2b",
          5420 => x"29",
          5421 => x"81",
          5422 => x"98",
          5423 => x"2b",
          5424 => x"45",
          5425 => x"73",
          5426 => x"38",
          5427 => x"70",
          5428 => x"06",
          5429 => x"7b",
          5430 => x"38",
          5431 => x"73",
          5432 => x"81",
          5433 => x"78",
          5434 => x"3f",
          5435 => x"ff",
          5436 => x"e5",
          5437 => x"38",
          5438 => x"89",
          5439 => x"f6",
          5440 => x"a5",
          5441 => x"55",
          5442 => x"80",
          5443 => x"1d",
          5444 => x"83",
          5445 => x"88",
          5446 => x"57",
          5447 => x"3f",
          5448 => x"51",
          5449 => x"82",
          5450 => x"83",
          5451 => x"7e",
          5452 => x"70",
          5453 => x"bb",
          5454 => x"84",
          5455 => x"59",
          5456 => x"3f",
          5457 => x"08",
          5458 => x"75",
          5459 => x"06",
          5460 => x"85",
          5461 => x"54",
          5462 => x"80",
          5463 => x"51",
          5464 => x"82",
          5465 => x"1d",
          5466 => x"83",
          5467 => x"88",
          5468 => x"43",
          5469 => x"3f",
          5470 => x"51",
          5471 => x"82",
          5472 => x"83",
          5473 => x"7e",
          5474 => x"70",
          5475 => x"bb",
          5476 => x"84",
          5477 => x"59",
          5478 => x"3f",
          5479 => x"08",
          5480 => x"60",
          5481 => x"55",
          5482 => x"ff",
          5483 => x"a9",
          5484 => x"52",
          5485 => x"3f",
          5486 => x"08",
          5487 => x"dc",
          5488 => x"93",
          5489 => x"73",
          5490 => x"dc",
          5491 => x"92",
          5492 => x"51",
          5493 => x"7a",
          5494 => x"27",
          5495 => x"53",
          5496 => x"51",
          5497 => x"7a",
          5498 => x"82",
          5499 => x"05",
          5500 => x"f6",
          5501 => x"54",
          5502 => x"dc",
          5503 => x"0d",
          5504 => x"0d",
          5505 => x"70",
          5506 => x"d5",
          5507 => x"dc",
          5508 => x"bb",
          5509 => x"2e",
          5510 => x"53",
          5511 => x"bb",
          5512 => x"ff",
          5513 => x"74",
          5514 => x"0c",
          5515 => x"04",
          5516 => x"02",
          5517 => x"51",
          5518 => x"72",
          5519 => x"82",
          5520 => x"33",
          5521 => x"bb",
          5522 => x"3d",
          5523 => x"3d",
          5524 => x"05",
          5525 => x"05",
          5526 => x"56",
          5527 => x"72",
          5528 => x"e0",
          5529 => x"2b",
          5530 => x"8c",
          5531 => x"88",
          5532 => x"2e",
          5533 => x"88",
          5534 => x"0c",
          5535 => x"8c",
          5536 => x"71",
          5537 => x"87",
          5538 => x"0c",
          5539 => x"08",
          5540 => x"51",
          5541 => x"2e",
          5542 => x"c0",
          5543 => x"51",
          5544 => x"71",
          5545 => x"80",
          5546 => x"92",
          5547 => x"98",
          5548 => x"70",
          5549 => x"38",
          5550 => x"d8",
          5551 => x"bb",
          5552 => x"51",
          5553 => x"dc",
          5554 => x"0d",
          5555 => x"0d",
          5556 => x"02",
          5557 => x"05",
          5558 => x"58",
          5559 => x"52",
          5560 => x"3f",
          5561 => x"08",
          5562 => x"54",
          5563 => x"be",
          5564 => x"75",
          5565 => x"c0",
          5566 => x"87",
          5567 => x"12",
          5568 => x"84",
          5569 => x"40",
          5570 => x"85",
          5571 => x"98",
          5572 => x"7d",
          5573 => x"0c",
          5574 => x"85",
          5575 => x"06",
          5576 => x"71",
          5577 => x"38",
          5578 => x"71",
          5579 => x"05",
          5580 => x"19",
          5581 => x"a2",
          5582 => x"71",
          5583 => x"38",
          5584 => x"83",
          5585 => x"38",
          5586 => x"8a",
          5587 => x"98",
          5588 => x"71",
          5589 => x"c0",
          5590 => x"52",
          5591 => x"87",
          5592 => x"80",
          5593 => x"81",
          5594 => x"c0",
          5595 => x"53",
          5596 => x"82",
          5597 => x"71",
          5598 => x"1a",
          5599 => x"84",
          5600 => x"19",
          5601 => x"06",
          5602 => x"79",
          5603 => x"38",
          5604 => x"80",
          5605 => x"87",
          5606 => x"26",
          5607 => x"73",
          5608 => x"06",
          5609 => x"2e",
          5610 => x"52",
          5611 => x"82",
          5612 => x"8f",
          5613 => x"f3",
          5614 => x"62",
          5615 => x"05",
          5616 => x"57",
          5617 => x"83",
          5618 => x"52",
          5619 => x"3f",
          5620 => x"08",
          5621 => x"54",
          5622 => x"2e",
          5623 => x"81",
          5624 => x"74",
          5625 => x"c0",
          5626 => x"87",
          5627 => x"12",
          5628 => x"84",
          5629 => x"5f",
          5630 => x"0b",
          5631 => x"8c",
          5632 => x"0c",
          5633 => x"80",
          5634 => x"70",
          5635 => x"81",
          5636 => x"54",
          5637 => x"8c",
          5638 => x"81",
          5639 => x"7c",
          5640 => x"58",
          5641 => x"70",
          5642 => x"52",
          5643 => x"8a",
          5644 => x"98",
          5645 => x"71",
          5646 => x"c0",
          5647 => x"52",
          5648 => x"87",
          5649 => x"80",
          5650 => x"81",
          5651 => x"c0",
          5652 => x"53",
          5653 => x"82",
          5654 => x"71",
          5655 => x"19",
          5656 => x"81",
          5657 => x"ff",
          5658 => x"19",
          5659 => x"78",
          5660 => x"38",
          5661 => x"80",
          5662 => x"87",
          5663 => x"26",
          5664 => x"73",
          5665 => x"06",
          5666 => x"2e",
          5667 => x"52",
          5668 => x"82",
          5669 => x"8f",
          5670 => x"fa",
          5671 => x"02",
          5672 => x"05",
          5673 => x"05",
          5674 => x"71",
          5675 => x"57",
          5676 => x"82",
          5677 => x"81",
          5678 => x"54",
          5679 => x"38",
          5680 => x"c0",
          5681 => x"81",
          5682 => x"2e",
          5683 => x"71",
          5684 => x"38",
          5685 => x"87",
          5686 => x"11",
          5687 => x"80",
          5688 => x"80",
          5689 => x"83",
          5690 => x"38",
          5691 => x"72",
          5692 => x"2a",
          5693 => x"51",
          5694 => x"80",
          5695 => x"87",
          5696 => x"08",
          5697 => x"38",
          5698 => x"8c",
          5699 => x"96",
          5700 => x"0c",
          5701 => x"8c",
          5702 => x"08",
          5703 => x"51",
          5704 => x"38",
          5705 => x"56",
          5706 => x"80",
          5707 => x"85",
          5708 => x"77",
          5709 => x"83",
          5710 => x"75",
          5711 => x"bb",
          5712 => x"3d",
          5713 => x"3d",
          5714 => x"11",
          5715 => x"71",
          5716 => x"82",
          5717 => x"53",
          5718 => x"0d",
          5719 => x"0d",
          5720 => x"33",
          5721 => x"71",
          5722 => x"88",
          5723 => x"14",
          5724 => x"07",
          5725 => x"33",
          5726 => x"bb",
          5727 => x"53",
          5728 => x"52",
          5729 => x"04",
          5730 => x"73",
          5731 => x"92",
          5732 => x"52",
          5733 => x"81",
          5734 => x"70",
          5735 => x"70",
          5736 => x"3d",
          5737 => x"3d",
          5738 => x"52",
          5739 => x"70",
          5740 => x"34",
          5741 => x"51",
          5742 => x"81",
          5743 => x"70",
          5744 => x"70",
          5745 => x"05",
          5746 => x"88",
          5747 => x"72",
          5748 => x"0d",
          5749 => x"0d",
          5750 => x"54",
          5751 => x"80",
          5752 => x"71",
          5753 => x"53",
          5754 => x"81",
          5755 => x"ff",
          5756 => x"39",
          5757 => x"04",
          5758 => x"75",
          5759 => x"52",
          5760 => x"70",
          5761 => x"34",
          5762 => x"70",
          5763 => x"3d",
          5764 => x"3d",
          5765 => x"79",
          5766 => x"74",
          5767 => x"56",
          5768 => x"81",
          5769 => x"71",
          5770 => x"16",
          5771 => x"52",
          5772 => x"86",
          5773 => x"2e",
          5774 => x"82",
          5775 => x"86",
          5776 => x"fe",
          5777 => x"76",
          5778 => x"39",
          5779 => x"8a",
          5780 => x"51",
          5781 => x"71",
          5782 => x"33",
          5783 => x"0c",
          5784 => x"04",
          5785 => x"bb",
          5786 => x"80",
          5787 => x"dc",
          5788 => x"3d",
          5789 => x"80",
          5790 => x"33",
          5791 => x"7a",
          5792 => x"38",
          5793 => x"16",
          5794 => x"16",
          5795 => x"17",
          5796 => x"fa",
          5797 => x"bb",
          5798 => x"2e",
          5799 => x"b7",
          5800 => x"dc",
          5801 => x"34",
          5802 => x"70",
          5803 => x"31",
          5804 => x"59",
          5805 => x"77",
          5806 => x"82",
          5807 => x"74",
          5808 => x"81",
          5809 => x"81",
          5810 => x"53",
          5811 => x"16",
          5812 => x"e3",
          5813 => x"81",
          5814 => x"bb",
          5815 => x"3d",
          5816 => x"3d",
          5817 => x"56",
          5818 => x"74",
          5819 => x"2e",
          5820 => x"51",
          5821 => x"82",
          5822 => x"57",
          5823 => x"08",
          5824 => x"54",
          5825 => x"16",
          5826 => x"33",
          5827 => x"3f",
          5828 => x"08",
          5829 => x"38",
          5830 => x"57",
          5831 => x"0c",
          5832 => x"dc",
          5833 => x"0d",
          5834 => x"0d",
          5835 => x"57",
          5836 => x"82",
          5837 => x"58",
          5838 => x"08",
          5839 => x"76",
          5840 => x"83",
          5841 => x"06",
          5842 => x"84",
          5843 => x"78",
          5844 => x"81",
          5845 => x"38",
          5846 => x"82",
          5847 => x"52",
          5848 => x"52",
          5849 => x"3f",
          5850 => x"52",
          5851 => x"51",
          5852 => x"84",
          5853 => x"d2",
          5854 => x"fc",
          5855 => x"8a",
          5856 => x"52",
          5857 => x"51",
          5858 => x"90",
          5859 => x"84",
          5860 => x"fc",
          5861 => x"17",
          5862 => x"a0",
          5863 => x"86",
          5864 => x"08",
          5865 => x"b0",
          5866 => x"55",
          5867 => x"81",
          5868 => x"f8",
          5869 => x"84",
          5870 => x"53",
          5871 => x"17",
          5872 => x"d7",
          5873 => x"dc",
          5874 => x"83",
          5875 => x"77",
          5876 => x"0c",
          5877 => x"04",
          5878 => x"77",
          5879 => x"12",
          5880 => x"55",
          5881 => x"56",
          5882 => x"8d",
          5883 => x"22",
          5884 => x"ac",
          5885 => x"57",
          5886 => x"bb",
          5887 => x"3d",
          5888 => x"3d",
          5889 => x"70",
          5890 => x"57",
          5891 => x"81",
          5892 => x"98",
          5893 => x"81",
          5894 => x"74",
          5895 => x"72",
          5896 => x"f5",
          5897 => x"24",
          5898 => x"81",
          5899 => x"81",
          5900 => x"83",
          5901 => x"38",
          5902 => x"76",
          5903 => x"70",
          5904 => x"16",
          5905 => x"74",
          5906 => x"96",
          5907 => x"dc",
          5908 => x"38",
          5909 => x"06",
          5910 => x"33",
          5911 => x"89",
          5912 => x"08",
          5913 => x"54",
          5914 => x"fc",
          5915 => x"bb",
          5916 => x"fe",
          5917 => x"ff",
          5918 => x"11",
          5919 => x"2b",
          5920 => x"81",
          5921 => x"2a",
          5922 => x"51",
          5923 => x"e2",
          5924 => x"ff",
          5925 => x"da",
          5926 => x"2a",
          5927 => x"05",
          5928 => x"fc",
          5929 => x"bb",
          5930 => x"c6",
          5931 => x"83",
          5932 => x"05",
          5933 => x"f9",
          5934 => x"bb",
          5935 => x"ff",
          5936 => x"ae",
          5937 => x"2a",
          5938 => x"05",
          5939 => x"fc",
          5940 => x"bb",
          5941 => x"38",
          5942 => x"83",
          5943 => x"05",
          5944 => x"f8",
          5945 => x"bb",
          5946 => x"0a",
          5947 => x"39",
          5948 => x"82",
          5949 => x"89",
          5950 => x"f8",
          5951 => x"7c",
          5952 => x"56",
          5953 => x"77",
          5954 => x"38",
          5955 => x"08",
          5956 => x"38",
          5957 => x"72",
          5958 => x"9d",
          5959 => x"24",
          5960 => x"81",
          5961 => x"82",
          5962 => x"83",
          5963 => x"38",
          5964 => x"76",
          5965 => x"70",
          5966 => x"18",
          5967 => x"76",
          5968 => x"9e",
          5969 => x"dc",
          5970 => x"bb",
          5971 => x"d9",
          5972 => x"ff",
          5973 => x"05",
          5974 => x"81",
          5975 => x"54",
          5976 => x"80",
          5977 => x"77",
          5978 => x"f0",
          5979 => x"8f",
          5980 => x"51",
          5981 => x"34",
          5982 => x"17",
          5983 => x"2a",
          5984 => x"05",
          5985 => x"fa",
          5986 => x"bb",
          5987 => x"82",
          5988 => x"81",
          5989 => x"83",
          5990 => x"b4",
          5991 => x"2a",
          5992 => x"8f",
          5993 => x"2a",
          5994 => x"f0",
          5995 => x"06",
          5996 => x"72",
          5997 => x"ec",
          5998 => x"2a",
          5999 => x"05",
          6000 => x"fa",
          6001 => x"bb",
          6002 => x"82",
          6003 => x"80",
          6004 => x"83",
          6005 => x"52",
          6006 => x"fe",
          6007 => x"b4",
          6008 => x"a4",
          6009 => x"76",
          6010 => x"17",
          6011 => x"75",
          6012 => x"3f",
          6013 => x"08",
          6014 => x"dc",
          6015 => x"77",
          6016 => x"77",
          6017 => x"fc",
          6018 => x"b4",
          6019 => x"51",
          6020 => x"c9",
          6021 => x"dc",
          6022 => x"06",
          6023 => x"72",
          6024 => x"3f",
          6025 => x"17",
          6026 => x"bb",
          6027 => x"3d",
          6028 => x"3d",
          6029 => x"7e",
          6030 => x"56",
          6031 => x"75",
          6032 => x"74",
          6033 => x"27",
          6034 => x"80",
          6035 => x"ff",
          6036 => x"75",
          6037 => x"3f",
          6038 => x"08",
          6039 => x"dc",
          6040 => x"38",
          6041 => x"54",
          6042 => x"81",
          6043 => x"39",
          6044 => x"08",
          6045 => x"39",
          6046 => x"51",
          6047 => x"82",
          6048 => x"58",
          6049 => x"08",
          6050 => x"c7",
          6051 => x"dc",
          6052 => x"d2",
          6053 => x"dc",
          6054 => x"cf",
          6055 => x"74",
          6056 => x"fc",
          6057 => x"bb",
          6058 => x"38",
          6059 => x"fe",
          6060 => x"08",
          6061 => x"74",
          6062 => x"38",
          6063 => x"17",
          6064 => x"33",
          6065 => x"73",
          6066 => x"77",
          6067 => x"26",
          6068 => x"80",
          6069 => x"bb",
          6070 => x"3d",
          6071 => x"3d",
          6072 => x"71",
          6073 => x"5b",
          6074 => x"8c",
          6075 => x"77",
          6076 => x"38",
          6077 => x"78",
          6078 => x"81",
          6079 => x"79",
          6080 => x"f9",
          6081 => x"55",
          6082 => x"dc",
          6083 => x"e0",
          6084 => x"dc",
          6085 => x"bb",
          6086 => x"2e",
          6087 => x"98",
          6088 => x"bb",
          6089 => x"82",
          6090 => x"58",
          6091 => x"70",
          6092 => x"80",
          6093 => x"38",
          6094 => x"09",
          6095 => x"e2",
          6096 => x"56",
          6097 => x"76",
          6098 => x"82",
          6099 => x"7a",
          6100 => x"3f",
          6101 => x"bb",
          6102 => x"2e",
          6103 => x"86",
          6104 => x"dc",
          6105 => x"bb",
          6106 => x"70",
          6107 => x"07",
          6108 => x"7c",
          6109 => x"dc",
          6110 => x"51",
          6111 => x"81",
          6112 => x"bb",
          6113 => x"2e",
          6114 => x"17",
          6115 => x"74",
          6116 => x"73",
          6117 => x"27",
          6118 => x"58",
          6119 => x"80",
          6120 => x"56",
          6121 => x"98",
          6122 => x"26",
          6123 => x"56",
          6124 => x"81",
          6125 => x"52",
          6126 => x"c6",
          6127 => x"dc",
          6128 => x"b8",
          6129 => x"82",
          6130 => x"81",
          6131 => x"06",
          6132 => x"bb",
          6133 => x"82",
          6134 => x"09",
          6135 => x"72",
          6136 => x"70",
          6137 => x"51",
          6138 => x"80",
          6139 => x"78",
          6140 => x"06",
          6141 => x"73",
          6142 => x"39",
          6143 => x"52",
          6144 => x"f7",
          6145 => x"dc",
          6146 => x"dc",
          6147 => x"82",
          6148 => x"07",
          6149 => x"55",
          6150 => x"2e",
          6151 => x"80",
          6152 => x"75",
          6153 => x"76",
          6154 => x"3f",
          6155 => x"08",
          6156 => x"38",
          6157 => x"0c",
          6158 => x"fe",
          6159 => x"08",
          6160 => x"74",
          6161 => x"ff",
          6162 => x"0c",
          6163 => x"81",
          6164 => x"84",
          6165 => x"39",
          6166 => x"81",
          6167 => x"8c",
          6168 => x"8c",
          6169 => x"dc",
          6170 => x"39",
          6171 => x"55",
          6172 => x"dc",
          6173 => x"0d",
          6174 => x"0d",
          6175 => x"55",
          6176 => x"82",
          6177 => x"58",
          6178 => x"bb",
          6179 => x"d8",
          6180 => x"74",
          6181 => x"3f",
          6182 => x"08",
          6183 => x"08",
          6184 => x"59",
          6185 => x"77",
          6186 => x"70",
          6187 => x"c8",
          6188 => x"84",
          6189 => x"56",
          6190 => x"58",
          6191 => x"97",
          6192 => x"75",
          6193 => x"52",
          6194 => x"51",
          6195 => x"82",
          6196 => x"80",
          6197 => x"8a",
          6198 => x"32",
          6199 => x"72",
          6200 => x"2a",
          6201 => x"56",
          6202 => x"dc",
          6203 => x"0d",
          6204 => x"0d",
          6205 => x"08",
          6206 => x"74",
          6207 => x"26",
          6208 => x"74",
          6209 => x"72",
          6210 => x"74",
          6211 => x"88",
          6212 => x"73",
          6213 => x"33",
          6214 => x"27",
          6215 => x"16",
          6216 => x"9b",
          6217 => x"2a",
          6218 => x"88",
          6219 => x"58",
          6220 => x"80",
          6221 => x"16",
          6222 => x"0c",
          6223 => x"8a",
          6224 => x"89",
          6225 => x"72",
          6226 => x"38",
          6227 => x"51",
          6228 => x"82",
          6229 => x"54",
          6230 => x"08",
          6231 => x"38",
          6232 => x"bb",
          6233 => x"8b",
          6234 => x"08",
          6235 => x"08",
          6236 => x"82",
          6237 => x"74",
          6238 => x"cb",
          6239 => x"75",
          6240 => x"3f",
          6241 => x"08",
          6242 => x"73",
          6243 => x"98",
          6244 => x"82",
          6245 => x"2e",
          6246 => x"39",
          6247 => x"39",
          6248 => x"13",
          6249 => x"74",
          6250 => x"16",
          6251 => x"18",
          6252 => x"77",
          6253 => x"0c",
          6254 => x"04",
          6255 => x"7a",
          6256 => x"12",
          6257 => x"59",
          6258 => x"80",
          6259 => x"86",
          6260 => x"98",
          6261 => x"14",
          6262 => x"55",
          6263 => x"81",
          6264 => x"83",
          6265 => x"77",
          6266 => x"81",
          6267 => x"0c",
          6268 => x"55",
          6269 => x"76",
          6270 => x"17",
          6271 => x"74",
          6272 => x"9b",
          6273 => x"39",
          6274 => x"ff",
          6275 => x"2a",
          6276 => x"81",
          6277 => x"52",
          6278 => x"e6",
          6279 => x"dc",
          6280 => x"55",
          6281 => x"bb",
          6282 => x"80",
          6283 => x"55",
          6284 => x"08",
          6285 => x"f4",
          6286 => x"08",
          6287 => x"08",
          6288 => x"38",
          6289 => x"77",
          6290 => x"84",
          6291 => x"39",
          6292 => x"52",
          6293 => x"86",
          6294 => x"dc",
          6295 => x"55",
          6296 => x"08",
          6297 => x"c4",
          6298 => x"82",
          6299 => x"81",
          6300 => x"81",
          6301 => x"dc",
          6302 => x"b0",
          6303 => x"dc",
          6304 => x"51",
          6305 => x"82",
          6306 => x"a0",
          6307 => x"15",
          6308 => x"75",
          6309 => x"3f",
          6310 => x"08",
          6311 => x"76",
          6312 => x"77",
          6313 => x"9c",
          6314 => x"55",
          6315 => x"dc",
          6316 => x"0d",
          6317 => x"0d",
          6318 => x"08",
          6319 => x"80",
          6320 => x"fc",
          6321 => x"bb",
          6322 => x"82",
          6323 => x"80",
          6324 => x"bb",
          6325 => x"98",
          6326 => x"78",
          6327 => x"3f",
          6328 => x"08",
          6329 => x"dc",
          6330 => x"38",
          6331 => x"08",
          6332 => x"70",
          6333 => x"58",
          6334 => x"2e",
          6335 => x"83",
          6336 => x"82",
          6337 => x"55",
          6338 => x"81",
          6339 => x"07",
          6340 => x"2e",
          6341 => x"16",
          6342 => x"2e",
          6343 => x"88",
          6344 => x"82",
          6345 => x"56",
          6346 => x"51",
          6347 => x"82",
          6348 => x"54",
          6349 => x"08",
          6350 => x"9b",
          6351 => x"2e",
          6352 => x"83",
          6353 => x"73",
          6354 => x"0c",
          6355 => x"04",
          6356 => x"76",
          6357 => x"54",
          6358 => x"82",
          6359 => x"83",
          6360 => x"76",
          6361 => x"53",
          6362 => x"2e",
          6363 => x"90",
          6364 => x"51",
          6365 => x"82",
          6366 => x"90",
          6367 => x"53",
          6368 => x"dc",
          6369 => x"0d",
          6370 => x"0d",
          6371 => x"83",
          6372 => x"54",
          6373 => x"55",
          6374 => x"3f",
          6375 => x"51",
          6376 => x"2e",
          6377 => x"8b",
          6378 => x"2a",
          6379 => x"51",
          6380 => x"86",
          6381 => x"f7",
          6382 => x"7d",
          6383 => x"75",
          6384 => x"98",
          6385 => x"2e",
          6386 => x"98",
          6387 => x"78",
          6388 => x"3f",
          6389 => x"08",
          6390 => x"dc",
          6391 => x"38",
          6392 => x"70",
          6393 => x"73",
          6394 => x"58",
          6395 => x"8b",
          6396 => x"bf",
          6397 => x"ff",
          6398 => x"53",
          6399 => x"34",
          6400 => x"08",
          6401 => x"e5",
          6402 => x"81",
          6403 => x"2e",
          6404 => x"70",
          6405 => x"57",
          6406 => x"9e",
          6407 => x"2e",
          6408 => x"bb",
          6409 => x"df",
          6410 => x"72",
          6411 => x"81",
          6412 => x"76",
          6413 => x"2e",
          6414 => x"52",
          6415 => x"fc",
          6416 => x"dc",
          6417 => x"bb",
          6418 => x"38",
          6419 => x"fe",
          6420 => x"39",
          6421 => x"16",
          6422 => x"bb",
          6423 => x"3d",
          6424 => x"3d",
          6425 => x"08",
          6426 => x"52",
          6427 => x"c5",
          6428 => x"dc",
          6429 => x"bb",
          6430 => x"38",
          6431 => x"52",
          6432 => x"de",
          6433 => x"dc",
          6434 => x"bb",
          6435 => x"38",
          6436 => x"bb",
          6437 => x"9c",
          6438 => x"ea",
          6439 => x"53",
          6440 => x"9c",
          6441 => x"ea",
          6442 => x"0b",
          6443 => x"74",
          6444 => x"0c",
          6445 => x"04",
          6446 => x"75",
          6447 => x"12",
          6448 => x"53",
          6449 => x"9a",
          6450 => x"dc",
          6451 => x"9c",
          6452 => x"e5",
          6453 => x"0b",
          6454 => x"85",
          6455 => x"fa",
          6456 => x"7a",
          6457 => x"0b",
          6458 => x"98",
          6459 => x"2e",
          6460 => x"80",
          6461 => x"55",
          6462 => x"17",
          6463 => x"33",
          6464 => x"51",
          6465 => x"2e",
          6466 => x"85",
          6467 => x"06",
          6468 => x"e5",
          6469 => x"2e",
          6470 => x"8b",
          6471 => x"70",
          6472 => x"34",
          6473 => x"71",
          6474 => x"05",
          6475 => x"15",
          6476 => x"27",
          6477 => x"15",
          6478 => x"80",
          6479 => x"34",
          6480 => x"52",
          6481 => x"88",
          6482 => x"17",
          6483 => x"52",
          6484 => x"3f",
          6485 => x"08",
          6486 => x"12",
          6487 => x"3f",
          6488 => x"08",
          6489 => x"98",
          6490 => x"da",
          6491 => x"dc",
          6492 => x"23",
          6493 => x"04",
          6494 => x"7f",
          6495 => x"5b",
          6496 => x"33",
          6497 => x"73",
          6498 => x"38",
          6499 => x"80",
          6500 => x"38",
          6501 => x"8c",
          6502 => x"08",
          6503 => x"aa",
          6504 => x"41",
          6505 => x"33",
          6506 => x"73",
          6507 => x"81",
          6508 => x"81",
          6509 => x"dc",
          6510 => x"70",
          6511 => x"07",
          6512 => x"73",
          6513 => x"88",
          6514 => x"70",
          6515 => x"73",
          6516 => x"38",
          6517 => x"ab",
          6518 => x"52",
          6519 => x"91",
          6520 => x"dc",
          6521 => x"98",
          6522 => x"61",
          6523 => x"5a",
          6524 => x"a0",
          6525 => x"e7",
          6526 => x"70",
          6527 => x"79",
          6528 => x"73",
          6529 => x"81",
          6530 => x"38",
          6531 => x"33",
          6532 => x"ae",
          6533 => x"70",
          6534 => x"82",
          6535 => x"51",
          6536 => x"54",
          6537 => x"79",
          6538 => x"74",
          6539 => x"57",
          6540 => x"af",
          6541 => x"70",
          6542 => x"51",
          6543 => x"dc",
          6544 => x"73",
          6545 => x"38",
          6546 => x"82",
          6547 => x"19",
          6548 => x"54",
          6549 => x"82",
          6550 => x"54",
          6551 => x"78",
          6552 => x"81",
          6553 => x"54",
          6554 => x"81",
          6555 => x"af",
          6556 => x"77",
          6557 => x"70",
          6558 => x"25",
          6559 => x"07",
          6560 => x"51",
          6561 => x"2e",
          6562 => x"39",
          6563 => x"80",
          6564 => x"33",
          6565 => x"73",
          6566 => x"81",
          6567 => x"81",
          6568 => x"dc",
          6569 => x"70",
          6570 => x"07",
          6571 => x"73",
          6572 => x"b5",
          6573 => x"2e",
          6574 => x"83",
          6575 => x"76",
          6576 => x"07",
          6577 => x"2e",
          6578 => x"8b",
          6579 => x"77",
          6580 => x"30",
          6581 => x"71",
          6582 => x"53",
          6583 => x"55",
          6584 => x"38",
          6585 => x"5c",
          6586 => x"75",
          6587 => x"73",
          6588 => x"38",
          6589 => x"06",
          6590 => x"11",
          6591 => x"75",
          6592 => x"3f",
          6593 => x"08",
          6594 => x"38",
          6595 => x"33",
          6596 => x"54",
          6597 => x"e6",
          6598 => x"bb",
          6599 => x"2e",
          6600 => x"ff",
          6601 => x"74",
          6602 => x"38",
          6603 => x"75",
          6604 => x"17",
          6605 => x"57",
          6606 => x"a7",
          6607 => x"82",
          6608 => x"e5",
          6609 => x"bb",
          6610 => x"38",
          6611 => x"54",
          6612 => x"89",
          6613 => x"70",
          6614 => x"57",
          6615 => x"54",
          6616 => x"81",
          6617 => x"f7",
          6618 => x"7e",
          6619 => x"2e",
          6620 => x"33",
          6621 => x"e5",
          6622 => x"06",
          6623 => x"7a",
          6624 => x"a0",
          6625 => x"38",
          6626 => x"55",
          6627 => x"84",
          6628 => x"39",
          6629 => x"8b",
          6630 => x"7b",
          6631 => x"7a",
          6632 => x"3f",
          6633 => x"08",
          6634 => x"dc",
          6635 => x"38",
          6636 => x"52",
          6637 => x"aa",
          6638 => x"dc",
          6639 => x"bb",
          6640 => x"c2",
          6641 => x"08",
          6642 => x"55",
          6643 => x"ff",
          6644 => x"15",
          6645 => x"54",
          6646 => x"34",
          6647 => x"70",
          6648 => x"81",
          6649 => x"58",
          6650 => x"8b",
          6651 => x"74",
          6652 => x"3f",
          6653 => x"08",
          6654 => x"38",
          6655 => x"51",
          6656 => x"ff",
          6657 => x"ab",
          6658 => x"55",
          6659 => x"bb",
          6660 => x"2e",
          6661 => x"80",
          6662 => x"85",
          6663 => x"06",
          6664 => x"58",
          6665 => x"80",
          6666 => x"75",
          6667 => x"73",
          6668 => x"b5",
          6669 => x"0b",
          6670 => x"80",
          6671 => x"39",
          6672 => x"54",
          6673 => x"85",
          6674 => x"75",
          6675 => x"81",
          6676 => x"73",
          6677 => x"1b",
          6678 => x"2a",
          6679 => x"51",
          6680 => x"80",
          6681 => x"90",
          6682 => x"ff",
          6683 => x"05",
          6684 => x"f5",
          6685 => x"bb",
          6686 => x"1c",
          6687 => x"39",
          6688 => x"dc",
          6689 => x"0d",
          6690 => x"0d",
          6691 => x"7b",
          6692 => x"73",
          6693 => x"55",
          6694 => x"2e",
          6695 => x"75",
          6696 => x"57",
          6697 => x"26",
          6698 => x"ba",
          6699 => x"70",
          6700 => x"ba",
          6701 => x"06",
          6702 => x"73",
          6703 => x"70",
          6704 => x"51",
          6705 => x"89",
          6706 => x"82",
          6707 => x"ff",
          6708 => x"56",
          6709 => x"2e",
          6710 => x"80",
          6711 => x"94",
          6712 => x"08",
          6713 => x"76",
          6714 => x"58",
          6715 => x"81",
          6716 => x"ff",
          6717 => x"53",
          6718 => x"26",
          6719 => x"13",
          6720 => x"06",
          6721 => x"9f",
          6722 => x"99",
          6723 => x"e0",
          6724 => x"ff",
          6725 => x"72",
          6726 => x"2a",
          6727 => x"72",
          6728 => x"06",
          6729 => x"ff",
          6730 => x"30",
          6731 => x"70",
          6732 => x"07",
          6733 => x"9f",
          6734 => x"54",
          6735 => x"80",
          6736 => x"81",
          6737 => x"59",
          6738 => x"25",
          6739 => x"8b",
          6740 => x"24",
          6741 => x"76",
          6742 => x"78",
          6743 => x"82",
          6744 => x"51",
          6745 => x"dc",
          6746 => x"0d",
          6747 => x"0d",
          6748 => x"0b",
          6749 => x"ff",
          6750 => x"0c",
          6751 => x"51",
          6752 => x"84",
          6753 => x"dc",
          6754 => x"38",
          6755 => x"51",
          6756 => x"82",
          6757 => x"83",
          6758 => x"54",
          6759 => x"82",
          6760 => x"09",
          6761 => x"e3",
          6762 => x"b4",
          6763 => x"57",
          6764 => x"2e",
          6765 => x"83",
          6766 => x"74",
          6767 => x"70",
          6768 => x"25",
          6769 => x"51",
          6770 => x"38",
          6771 => x"2e",
          6772 => x"b5",
          6773 => x"82",
          6774 => x"80",
          6775 => x"e0",
          6776 => x"bb",
          6777 => x"82",
          6778 => x"80",
          6779 => x"85",
          6780 => x"d8",
          6781 => x"16",
          6782 => x"3f",
          6783 => x"08",
          6784 => x"dc",
          6785 => x"83",
          6786 => x"74",
          6787 => x"0c",
          6788 => x"04",
          6789 => x"61",
          6790 => x"80",
          6791 => x"58",
          6792 => x"0c",
          6793 => x"e1",
          6794 => x"dc",
          6795 => x"56",
          6796 => x"bb",
          6797 => x"86",
          6798 => x"bb",
          6799 => x"29",
          6800 => x"05",
          6801 => x"53",
          6802 => x"80",
          6803 => x"38",
          6804 => x"76",
          6805 => x"74",
          6806 => x"72",
          6807 => x"38",
          6808 => x"51",
          6809 => x"82",
          6810 => x"81",
          6811 => x"81",
          6812 => x"72",
          6813 => x"80",
          6814 => x"38",
          6815 => x"70",
          6816 => x"53",
          6817 => x"86",
          6818 => x"a7",
          6819 => x"34",
          6820 => x"34",
          6821 => x"14",
          6822 => x"b2",
          6823 => x"dc",
          6824 => x"06",
          6825 => x"54",
          6826 => x"72",
          6827 => x"76",
          6828 => x"38",
          6829 => x"70",
          6830 => x"53",
          6831 => x"85",
          6832 => x"70",
          6833 => x"5b",
          6834 => x"82",
          6835 => x"81",
          6836 => x"76",
          6837 => x"81",
          6838 => x"38",
          6839 => x"56",
          6840 => x"83",
          6841 => x"70",
          6842 => x"80",
          6843 => x"83",
          6844 => x"dc",
          6845 => x"bb",
          6846 => x"76",
          6847 => x"05",
          6848 => x"16",
          6849 => x"56",
          6850 => x"d7",
          6851 => x"8d",
          6852 => x"72",
          6853 => x"54",
          6854 => x"57",
          6855 => x"95",
          6856 => x"73",
          6857 => x"3f",
          6858 => x"08",
          6859 => x"57",
          6860 => x"89",
          6861 => x"56",
          6862 => x"d7",
          6863 => x"76",
          6864 => x"f1",
          6865 => x"76",
          6866 => x"e9",
          6867 => x"51",
          6868 => x"82",
          6869 => x"83",
          6870 => x"53",
          6871 => x"2e",
          6872 => x"84",
          6873 => x"ca",
          6874 => x"da",
          6875 => x"dc",
          6876 => x"ff",
          6877 => x"8d",
          6878 => x"14",
          6879 => x"3f",
          6880 => x"08",
          6881 => x"15",
          6882 => x"14",
          6883 => x"34",
          6884 => x"33",
          6885 => x"81",
          6886 => x"54",
          6887 => x"72",
          6888 => x"91",
          6889 => x"ff",
          6890 => x"29",
          6891 => x"33",
          6892 => x"72",
          6893 => x"72",
          6894 => x"38",
          6895 => x"06",
          6896 => x"2e",
          6897 => x"56",
          6898 => x"80",
          6899 => x"da",
          6900 => x"bb",
          6901 => x"82",
          6902 => x"88",
          6903 => x"8f",
          6904 => x"56",
          6905 => x"38",
          6906 => x"51",
          6907 => x"82",
          6908 => x"83",
          6909 => x"55",
          6910 => x"80",
          6911 => x"da",
          6912 => x"bb",
          6913 => x"80",
          6914 => x"da",
          6915 => x"bb",
          6916 => x"ff",
          6917 => x"8d",
          6918 => x"2e",
          6919 => x"88",
          6920 => x"14",
          6921 => x"05",
          6922 => x"75",
          6923 => x"38",
          6924 => x"52",
          6925 => x"51",
          6926 => x"3f",
          6927 => x"08",
          6928 => x"dc",
          6929 => x"82",
          6930 => x"bb",
          6931 => x"ff",
          6932 => x"26",
          6933 => x"57",
          6934 => x"f5",
          6935 => x"82",
          6936 => x"f5",
          6937 => x"81",
          6938 => x"8d",
          6939 => x"2e",
          6940 => x"82",
          6941 => x"16",
          6942 => x"16",
          6943 => x"70",
          6944 => x"7a",
          6945 => x"0c",
          6946 => x"83",
          6947 => x"06",
          6948 => x"de",
          6949 => x"ae",
          6950 => x"dc",
          6951 => x"ff",
          6952 => x"56",
          6953 => x"38",
          6954 => x"38",
          6955 => x"51",
          6956 => x"82",
          6957 => x"a8",
          6958 => x"82",
          6959 => x"39",
          6960 => x"80",
          6961 => x"38",
          6962 => x"15",
          6963 => x"53",
          6964 => x"8d",
          6965 => x"15",
          6966 => x"76",
          6967 => x"51",
          6968 => x"13",
          6969 => x"8d",
          6970 => x"15",
          6971 => x"c5",
          6972 => x"90",
          6973 => x"0b",
          6974 => x"ff",
          6975 => x"15",
          6976 => x"2e",
          6977 => x"81",
          6978 => x"e4",
          6979 => x"b6",
          6980 => x"dc",
          6981 => x"ff",
          6982 => x"81",
          6983 => x"06",
          6984 => x"81",
          6985 => x"51",
          6986 => x"82",
          6987 => x"80",
          6988 => x"bb",
          6989 => x"15",
          6990 => x"14",
          6991 => x"3f",
          6992 => x"08",
          6993 => x"06",
          6994 => x"d4",
          6995 => x"81",
          6996 => x"38",
          6997 => x"d8",
          6998 => x"bb",
          6999 => x"8b",
          7000 => x"2e",
          7001 => x"b3",
          7002 => x"14",
          7003 => x"3f",
          7004 => x"08",
          7005 => x"e4",
          7006 => x"81",
          7007 => x"84",
          7008 => x"d7",
          7009 => x"bb",
          7010 => x"15",
          7011 => x"14",
          7012 => x"3f",
          7013 => x"08",
          7014 => x"76",
          7015 => x"d3",
          7016 => x"05",
          7017 => x"d3",
          7018 => x"86",
          7019 => x"0b",
          7020 => x"80",
          7021 => x"bb",
          7022 => x"3d",
          7023 => x"3d",
          7024 => x"89",
          7025 => x"2e",
          7026 => x"08",
          7027 => x"2e",
          7028 => x"33",
          7029 => x"2e",
          7030 => x"13",
          7031 => x"22",
          7032 => x"76",
          7033 => x"06",
          7034 => x"13",
          7035 => x"c0",
          7036 => x"dc",
          7037 => x"52",
          7038 => x"71",
          7039 => x"55",
          7040 => x"53",
          7041 => x"0c",
          7042 => x"bb",
          7043 => x"3d",
          7044 => x"3d",
          7045 => x"05",
          7046 => x"89",
          7047 => x"52",
          7048 => x"3f",
          7049 => x"0b",
          7050 => x"08",
          7051 => x"82",
          7052 => x"84",
          7053 => x"94",
          7054 => x"55",
          7055 => x"2e",
          7056 => x"74",
          7057 => x"73",
          7058 => x"38",
          7059 => x"78",
          7060 => x"54",
          7061 => x"92",
          7062 => x"89",
          7063 => x"84",
          7064 => x"b0",
          7065 => x"dc",
          7066 => x"82",
          7067 => x"88",
          7068 => x"eb",
          7069 => x"02",
          7070 => x"e7",
          7071 => x"59",
          7072 => x"80",
          7073 => x"38",
          7074 => x"70",
          7075 => x"d0",
          7076 => x"3d",
          7077 => x"58",
          7078 => x"82",
          7079 => x"55",
          7080 => x"08",
          7081 => x"7a",
          7082 => x"8c",
          7083 => x"56",
          7084 => x"82",
          7085 => x"55",
          7086 => x"08",
          7087 => x"80",
          7088 => x"70",
          7089 => x"57",
          7090 => x"83",
          7091 => x"77",
          7092 => x"73",
          7093 => x"ab",
          7094 => x"2e",
          7095 => x"84",
          7096 => x"06",
          7097 => x"51",
          7098 => x"82",
          7099 => x"55",
          7100 => x"b2",
          7101 => x"06",
          7102 => x"b8",
          7103 => x"2a",
          7104 => x"51",
          7105 => x"2e",
          7106 => x"55",
          7107 => x"77",
          7108 => x"74",
          7109 => x"77",
          7110 => x"81",
          7111 => x"73",
          7112 => x"af",
          7113 => x"7a",
          7114 => x"3f",
          7115 => x"08",
          7116 => x"b2",
          7117 => x"8e",
          7118 => x"ea",
          7119 => x"a0",
          7120 => x"34",
          7121 => x"52",
          7122 => x"bd",
          7123 => x"62",
          7124 => x"d4",
          7125 => x"54",
          7126 => x"15",
          7127 => x"2e",
          7128 => x"7a",
          7129 => x"51",
          7130 => x"75",
          7131 => x"d4",
          7132 => x"be",
          7133 => x"dc",
          7134 => x"bb",
          7135 => x"ca",
          7136 => x"74",
          7137 => x"02",
          7138 => x"70",
          7139 => x"81",
          7140 => x"56",
          7141 => x"86",
          7142 => x"82",
          7143 => x"81",
          7144 => x"06",
          7145 => x"80",
          7146 => x"75",
          7147 => x"73",
          7148 => x"38",
          7149 => x"92",
          7150 => x"7a",
          7151 => x"3f",
          7152 => x"08",
          7153 => x"8c",
          7154 => x"55",
          7155 => x"08",
          7156 => x"77",
          7157 => x"81",
          7158 => x"73",
          7159 => x"38",
          7160 => x"07",
          7161 => x"11",
          7162 => x"0c",
          7163 => x"0c",
          7164 => x"52",
          7165 => x"3f",
          7166 => x"08",
          7167 => x"08",
          7168 => x"63",
          7169 => x"5a",
          7170 => x"82",
          7171 => x"82",
          7172 => x"8c",
          7173 => x"7a",
          7174 => x"17",
          7175 => x"23",
          7176 => x"34",
          7177 => x"1a",
          7178 => x"9c",
          7179 => x"0b",
          7180 => x"77",
          7181 => x"81",
          7182 => x"73",
          7183 => x"8d",
          7184 => x"dc",
          7185 => x"81",
          7186 => x"bb",
          7187 => x"1a",
          7188 => x"22",
          7189 => x"7b",
          7190 => x"a8",
          7191 => x"78",
          7192 => x"3f",
          7193 => x"08",
          7194 => x"dc",
          7195 => x"83",
          7196 => x"82",
          7197 => x"ff",
          7198 => x"06",
          7199 => x"55",
          7200 => x"56",
          7201 => x"76",
          7202 => x"51",
          7203 => x"27",
          7204 => x"70",
          7205 => x"5a",
          7206 => x"76",
          7207 => x"74",
          7208 => x"83",
          7209 => x"73",
          7210 => x"38",
          7211 => x"51",
          7212 => x"82",
          7213 => x"85",
          7214 => x"8e",
          7215 => x"2a",
          7216 => x"08",
          7217 => x"0c",
          7218 => x"79",
          7219 => x"73",
          7220 => x"0c",
          7221 => x"04",
          7222 => x"60",
          7223 => x"40",
          7224 => x"80",
          7225 => x"3d",
          7226 => x"78",
          7227 => x"3f",
          7228 => x"08",
          7229 => x"dc",
          7230 => x"91",
          7231 => x"74",
          7232 => x"38",
          7233 => x"c4",
          7234 => x"33",
          7235 => x"87",
          7236 => x"2e",
          7237 => x"95",
          7238 => x"91",
          7239 => x"56",
          7240 => x"81",
          7241 => x"34",
          7242 => x"a0",
          7243 => x"08",
          7244 => x"31",
          7245 => x"27",
          7246 => x"5c",
          7247 => x"82",
          7248 => x"19",
          7249 => x"ff",
          7250 => x"74",
          7251 => x"7e",
          7252 => x"ff",
          7253 => x"2a",
          7254 => x"79",
          7255 => x"87",
          7256 => x"08",
          7257 => x"98",
          7258 => x"78",
          7259 => x"3f",
          7260 => x"08",
          7261 => x"27",
          7262 => x"74",
          7263 => x"a3",
          7264 => x"1a",
          7265 => x"08",
          7266 => x"d4",
          7267 => x"bb",
          7268 => x"2e",
          7269 => x"82",
          7270 => x"1a",
          7271 => x"59",
          7272 => x"2e",
          7273 => x"77",
          7274 => x"11",
          7275 => x"55",
          7276 => x"85",
          7277 => x"31",
          7278 => x"76",
          7279 => x"81",
          7280 => x"ca",
          7281 => x"bb",
          7282 => x"d7",
          7283 => x"11",
          7284 => x"74",
          7285 => x"38",
          7286 => x"77",
          7287 => x"78",
          7288 => x"84",
          7289 => x"16",
          7290 => x"08",
          7291 => x"2b",
          7292 => x"cf",
          7293 => x"89",
          7294 => x"39",
          7295 => x"0c",
          7296 => x"83",
          7297 => x"80",
          7298 => x"55",
          7299 => x"83",
          7300 => x"9c",
          7301 => x"7e",
          7302 => x"3f",
          7303 => x"08",
          7304 => x"75",
          7305 => x"08",
          7306 => x"1f",
          7307 => x"7c",
          7308 => x"3f",
          7309 => x"7e",
          7310 => x"0c",
          7311 => x"1b",
          7312 => x"1c",
          7313 => x"fd",
          7314 => x"56",
          7315 => x"dc",
          7316 => x"0d",
          7317 => x"0d",
          7318 => x"64",
          7319 => x"58",
          7320 => x"90",
          7321 => x"52",
          7322 => x"d2",
          7323 => x"dc",
          7324 => x"bb",
          7325 => x"38",
          7326 => x"55",
          7327 => x"86",
          7328 => x"83",
          7329 => x"18",
          7330 => x"2a",
          7331 => x"51",
          7332 => x"56",
          7333 => x"83",
          7334 => x"39",
          7335 => x"19",
          7336 => x"83",
          7337 => x"0b",
          7338 => x"81",
          7339 => x"39",
          7340 => x"7c",
          7341 => x"74",
          7342 => x"38",
          7343 => x"7b",
          7344 => x"ec",
          7345 => x"08",
          7346 => x"06",
          7347 => x"81",
          7348 => x"8a",
          7349 => x"05",
          7350 => x"06",
          7351 => x"bf",
          7352 => x"38",
          7353 => x"55",
          7354 => x"7a",
          7355 => x"98",
          7356 => x"77",
          7357 => x"3f",
          7358 => x"08",
          7359 => x"dc",
          7360 => x"82",
          7361 => x"81",
          7362 => x"38",
          7363 => x"ff",
          7364 => x"98",
          7365 => x"18",
          7366 => x"74",
          7367 => x"7e",
          7368 => x"08",
          7369 => x"2e",
          7370 => x"8d",
          7371 => x"ce",
          7372 => x"bb",
          7373 => x"ee",
          7374 => x"08",
          7375 => x"d1",
          7376 => x"bb",
          7377 => x"2e",
          7378 => x"82",
          7379 => x"1b",
          7380 => x"5a",
          7381 => x"2e",
          7382 => x"78",
          7383 => x"11",
          7384 => x"55",
          7385 => x"85",
          7386 => x"31",
          7387 => x"76",
          7388 => x"81",
          7389 => x"c8",
          7390 => x"bb",
          7391 => x"a6",
          7392 => x"11",
          7393 => x"56",
          7394 => x"27",
          7395 => x"80",
          7396 => x"08",
          7397 => x"2b",
          7398 => x"b4",
          7399 => x"b5",
          7400 => x"80",
          7401 => x"34",
          7402 => x"56",
          7403 => x"8c",
          7404 => x"19",
          7405 => x"38",
          7406 => x"b6",
          7407 => x"dc",
          7408 => x"38",
          7409 => x"12",
          7410 => x"9c",
          7411 => x"18",
          7412 => x"06",
          7413 => x"31",
          7414 => x"76",
          7415 => x"7b",
          7416 => x"08",
          7417 => x"cd",
          7418 => x"bb",
          7419 => x"b6",
          7420 => x"7c",
          7421 => x"08",
          7422 => x"1f",
          7423 => x"cb",
          7424 => x"55",
          7425 => x"16",
          7426 => x"31",
          7427 => x"7f",
          7428 => x"94",
          7429 => x"70",
          7430 => x"8c",
          7431 => x"58",
          7432 => x"76",
          7433 => x"75",
          7434 => x"19",
          7435 => x"39",
          7436 => x"80",
          7437 => x"74",
          7438 => x"80",
          7439 => x"bb",
          7440 => x"3d",
          7441 => x"3d",
          7442 => x"3d",
          7443 => x"70",
          7444 => x"ea",
          7445 => x"dc",
          7446 => x"bb",
          7447 => x"fb",
          7448 => x"33",
          7449 => x"70",
          7450 => x"55",
          7451 => x"2e",
          7452 => x"a0",
          7453 => x"78",
          7454 => x"3f",
          7455 => x"08",
          7456 => x"dc",
          7457 => x"38",
          7458 => x"8b",
          7459 => x"07",
          7460 => x"8b",
          7461 => x"16",
          7462 => x"52",
          7463 => x"dd",
          7464 => x"16",
          7465 => x"15",
          7466 => x"3f",
          7467 => x"0a",
          7468 => x"51",
          7469 => x"76",
          7470 => x"51",
          7471 => x"78",
          7472 => x"83",
          7473 => x"51",
          7474 => x"82",
          7475 => x"90",
          7476 => x"bf",
          7477 => x"73",
          7478 => x"76",
          7479 => x"0c",
          7480 => x"04",
          7481 => x"76",
          7482 => x"fe",
          7483 => x"bb",
          7484 => x"82",
          7485 => x"9c",
          7486 => x"fc",
          7487 => x"51",
          7488 => x"82",
          7489 => x"53",
          7490 => x"08",
          7491 => x"bb",
          7492 => x"0c",
          7493 => x"dc",
          7494 => x"0d",
          7495 => x"0d",
          7496 => x"e6",
          7497 => x"52",
          7498 => x"bb",
          7499 => x"8b",
          7500 => x"dc",
          7501 => x"a8",
          7502 => x"71",
          7503 => x"0c",
          7504 => x"04",
          7505 => x"80",
          7506 => x"d0",
          7507 => x"3d",
          7508 => x"3f",
          7509 => x"08",
          7510 => x"dc",
          7511 => x"38",
          7512 => x"52",
          7513 => x"05",
          7514 => x"3f",
          7515 => x"08",
          7516 => x"dc",
          7517 => x"02",
          7518 => x"33",
          7519 => x"55",
          7520 => x"25",
          7521 => x"7a",
          7522 => x"54",
          7523 => x"a2",
          7524 => x"84",
          7525 => x"06",
          7526 => x"73",
          7527 => x"38",
          7528 => x"70",
          7529 => x"a8",
          7530 => x"dc",
          7531 => x"0c",
          7532 => x"bb",
          7533 => x"2e",
          7534 => x"83",
          7535 => x"74",
          7536 => x"0c",
          7537 => x"04",
          7538 => x"6f",
          7539 => x"80",
          7540 => x"53",
          7541 => x"b8",
          7542 => x"3d",
          7543 => x"3f",
          7544 => x"08",
          7545 => x"dc",
          7546 => x"38",
          7547 => x"7c",
          7548 => x"47",
          7549 => x"54",
          7550 => x"81",
          7551 => x"52",
          7552 => x"52",
          7553 => x"3f",
          7554 => x"08",
          7555 => x"dc",
          7556 => x"38",
          7557 => x"51",
          7558 => x"82",
          7559 => x"57",
          7560 => x"08",
          7561 => x"69",
          7562 => x"da",
          7563 => x"bb",
          7564 => x"76",
          7565 => x"d5",
          7566 => x"bb",
          7567 => x"82",
          7568 => x"82",
          7569 => x"52",
          7570 => x"eb",
          7571 => x"dc",
          7572 => x"bb",
          7573 => x"38",
          7574 => x"51",
          7575 => x"73",
          7576 => x"08",
          7577 => x"76",
          7578 => x"d6",
          7579 => x"bb",
          7580 => x"82",
          7581 => x"80",
          7582 => x"76",
          7583 => x"81",
          7584 => x"82",
          7585 => x"39",
          7586 => x"38",
          7587 => x"bc",
          7588 => x"51",
          7589 => x"76",
          7590 => x"11",
          7591 => x"51",
          7592 => x"73",
          7593 => x"38",
          7594 => x"55",
          7595 => x"16",
          7596 => x"56",
          7597 => x"38",
          7598 => x"73",
          7599 => x"90",
          7600 => x"2e",
          7601 => x"16",
          7602 => x"ff",
          7603 => x"ff",
          7604 => x"58",
          7605 => x"74",
          7606 => x"75",
          7607 => x"18",
          7608 => x"58",
          7609 => x"fe",
          7610 => x"7b",
          7611 => x"06",
          7612 => x"18",
          7613 => x"58",
          7614 => x"80",
          7615 => x"a8",
          7616 => x"29",
          7617 => x"05",
          7618 => x"33",
          7619 => x"56",
          7620 => x"2e",
          7621 => x"16",
          7622 => x"33",
          7623 => x"73",
          7624 => x"16",
          7625 => x"26",
          7626 => x"55",
          7627 => x"91",
          7628 => x"54",
          7629 => x"70",
          7630 => x"34",
          7631 => x"ec",
          7632 => x"70",
          7633 => x"34",
          7634 => x"09",
          7635 => x"38",
          7636 => x"39",
          7637 => x"19",
          7638 => x"33",
          7639 => x"05",
          7640 => x"78",
          7641 => x"80",
          7642 => x"82",
          7643 => x"9e",
          7644 => x"f7",
          7645 => x"7d",
          7646 => x"05",
          7647 => x"57",
          7648 => x"3f",
          7649 => x"08",
          7650 => x"dc",
          7651 => x"38",
          7652 => x"53",
          7653 => x"38",
          7654 => x"54",
          7655 => x"92",
          7656 => x"33",
          7657 => x"70",
          7658 => x"54",
          7659 => x"38",
          7660 => x"15",
          7661 => x"70",
          7662 => x"58",
          7663 => x"82",
          7664 => x"8a",
          7665 => x"89",
          7666 => x"53",
          7667 => x"b7",
          7668 => x"ff",
          7669 => x"d7",
          7670 => x"bb",
          7671 => x"15",
          7672 => x"53",
          7673 => x"d7",
          7674 => x"bb",
          7675 => x"26",
          7676 => x"30",
          7677 => x"70",
          7678 => x"77",
          7679 => x"18",
          7680 => x"51",
          7681 => x"88",
          7682 => x"73",
          7683 => x"52",
          7684 => x"ca",
          7685 => x"dc",
          7686 => x"bb",
          7687 => x"2e",
          7688 => x"82",
          7689 => x"ff",
          7690 => x"38",
          7691 => x"08",
          7692 => x"73",
          7693 => x"73",
          7694 => x"9c",
          7695 => x"27",
          7696 => x"75",
          7697 => x"16",
          7698 => x"17",
          7699 => x"33",
          7700 => x"70",
          7701 => x"55",
          7702 => x"80",
          7703 => x"73",
          7704 => x"cc",
          7705 => x"bb",
          7706 => x"82",
          7707 => x"94",
          7708 => x"dc",
          7709 => x"39",
          7710 => x"51",
          7711 => x"82",
          7712 => x"54",
          7713 => x"be",
          7714 => x"27",
          7715 => x"53",
          7716 => x"08",
          7717 => x"73",
          7718 => x"ff",
          7719 => x"15",
          7720 => x"16",
          7721 => x"ff",
          7722 => x"80",
          7723 => x"73",
          7724 => x"c6",
          7725 => x"bb",
          7726 => x"38",
          7727 => x"16",
          7728 => x"80",
          7729 => x"0b",
          7730 => x"81",
          7731 => x"75",
          7732 => x"bb",
          7733 => x"58",
          7734 => x"54",
          7735 => x"74",
          7736 => x"73",
          7737 => x"90",
          7738 => x"c0",
          7739 => x"90",
          7740 => x"83",
          7741 => x"72",
          7742 => x"38",
          7743 => x"08",
          7744 => x"77",
          7745 => x"80",
          7746 => x"bb",
          7747 => x"3d",
          7748 => x"3d",
          7749 => x"89",
          7750 => x"2e",
          7751 => x"80",
          7752 => x"fc",
          7753 => x"3d",
          7754 => x"e1",
          7755 => x"bb",
          7756 => x"82",
          7757 => x"80",
          7758 => x"76",
          7759 => x"75",
          7760 => x"3f",
          7761 => x"08",
          7762 => x"dc",
          7763 => x"38",
          7764 => x"70",
          7765 => x"57",
          7766 => x"a2",
          7767 => x"33",
          7768 => x"70",
          7769 => x"55",
          7770 => x"2e",
          7771 => x"16",
          7772 => x"51",
          7773 => x"82",
          7774 => x"88",
          7775 => x"54",
          7776 => x"84",
          7777 => x"52",
          7778 => x"e5",
          7779 => x"dc",
          7780 => x"84",
          7781 => x"06",
          7782 => x"55",
          7783 => x"80",
          7784 => x"80",
          7785 => x"54",
          7786 => x"dc",
          7787 => x"0d",
          7788 => x"0d",
          7789 => x"fc",
          7790 => x"52",
          7791 => x"3f",
          7792 => x"08",
          7793 => x"bb",
          7794 => x"0c",
          7795 => x"04",
          7796 => x"77",
          7797 => x"fc",
          7798 => x"53",
          7799 => x"de",
          7800 => x"dc",
          7801 => x"bb",
          7802 => x"df",
          7803 => x"38",
          7804 => x"08",
          7805 => x"cd",
          7806 => x"bb",
          7807 => x"80",
          7808 => x"bb",
          7809 => x"73",
          7810 => x"3f",
          7811 => x"08",
          7812 => x"dc",
          7813 => x"09",
          7814 => x"38",
          7815 => x"39",
          7816 => x"08",
          7817 => x"52",
          7818 => x"b3",
          7819 => x"73",
          7820 => x"3f",
          7821 => x"08",
          7822 => x"30",
          7823 => x"9f",
          7824 => x"bb",
          7825 => x"51",
          7826 => x"72",
          7827 => x"0c",
          7828 => x"04",
          7829 => x"65",
          7830 => x"89",
          7831 => x"96",
          7832 => x"df",
          7833 => x"bb",
          7834 => x"82",
          7835 => x"b2",
          7836 => x"75",
          7837 => x"3f",
          7838 => x"08",
          7839 => x"dc",
          7840 => x"02",
          7841 => x"33",
          7842 => x"55",
          7843 => x"25",
          7844 => x"55",
          7845 => x"80",
          7846 => x"76",
          7847 => x"d4",
          7848 => x"82",
          7849 => x"94",
          7850 => x"f0",
          7851 => x"65",
          7852 => x"53",
          7853 => x"05",
          7854 => x"51",
          7855 => x"82",
          7856 => x"5b",
          7857 => x"08",
          7858 => x"7c",
          7859 => x"08",
          7860 => x"fe",
          7861 => x"08",
          7862 => x"55",
          7863 => x"91",
          7864 => x"0c",
          7865 => x"81",
          7866 => x"39",
          7867 => x"c7",
          7868 => x"dc",
          7869 => x"55",
          7870 => x"2e",
          7871 => x"bf",
          7872 => x"5f",
          7873 => x"92",
          7874 => x"51",
          7875 => x"82",
          7876 => x"ff",
          7877 => x"82",
          7878 => x"81",
          7879 => x"82",
          7880 => x"30",
          7881 => x"dc",
          7882 => x"25",
          7883 => x"19",
          7884 => x"5a",
          7885 => x"08",
          7886 => x"38",
          7887 => x"a4",
          7888 => x"bb",
          7889 => x"58",
          7890 => x"77",
          7891 => x"7d",
          7892 => x"bf",
          7893 => x"bb",
          7894 => x"82",
          7895 => x"80",
          7896 => x"70",
          7897 => x"ff",
          7898 => x"56",
          7899 => x"2e",
          7900 => x"9e",
          7901 => x"51",
          7902 => x"3f",
          7903 => x"08",
          7904 => x"06",
          7905 => x"80",
          7906 => x"19",
          7907 => x"54",
          7908 => x"14",
          7909 => x"c5",
          7910 => x"dc",
          7911 => x"06",
          7912 => x"80",
          7913 => x"19",
          7914 => x"54",
          7915 => x"06",
          7916 => x"79",
          7917 => x"78",
          7918 => x"79",
          7919 => x"84",
          7920 => x"07",
          7921 => x"84",
          7922 => x"82",
          7923 => x"92",
          7924 => x"f9",
          7925 => x"8a",
          7926 => x"53",
          7927 => x"e3",
          7928 => x"bb",
          7929 => x"82",
          7930 => x"81",
          7931 => x"17",
          7932 => x"81",
          7933 => x"17",
          7934 => x"2a",
          7935 => x"51",
          7936 => x"55",
          7937 => x"81",
          7938 => x"17",
          7939 => x"8c",
          7940 => x"81",
          7941 => x"9b",
          7942 => x"dc",
          7943 => x"17",
          7944 => x"51",
          7945 => x"82",
          7946 => x"74",
          7947 => x"56",
          7948 => x"98",
          7949 => x"76",
          7950 => x"c6",
          7951 => x"dc",
          7952 => x"09",
          7953 => x"38",
          7954 => x"bb",
          7955 => x"2e",
          7956 => x"85",
          7957 => x"a3",
          7958 => x"38",
          7959 => x"bb",
          7960 => x"15",
          7961 => x"38",
          7962 => x"53",
          7963 => x"08",
          7964 => x"c3",
          7965 => x"bb",
          7966 => x"94",
          7967 => x"18",
          7968 => x"33",
          7969 => x"54",
          7970 => x"34",
          7971 => x"85",
          7972 => x"18",
          7973 => x"74",
          7974 => x"0c",
          7975 => x"04",
          7976 => x"82",
          7977 => x"ff",
          7978 => x"a1",
          7979 => x"e4",
          7980 => x"dc",
          7981 => x"bb",
          7982 => x"f5",
          7983 => x"a1",
          7984 => x"95",
          7985 => x"58",
          7986 => x"82",
          7987 => x"55",
          7988 => x"08",
          7989 => x"02",
          7990 => x"33",
          7991 => x"70",
          7992 => x"55",
          7993 => x"73",
          7994 => x"75",
          7995 => x"80",
          7996 => x"bd",
          7997 => x"d6",
          7998 => x"81",
          7999 => x"87",
          8000 => x"ad",
          8001 => x"78",
          8002 => x"3f",
          8003 => x"08",
          8004 => x"70",
          8005 => x"55",
          8006 => x"2e",
          8007 => x"78",
          8008 => x"dc",
          8009 => x"08",
          8010 => x"38",
          8011 => x"bb",
          8012 => x"76",
          8013 => x"70",
          8014 => x"b5",
          8015 => x"dc",
          8016 => x"bb",
          8017 => x"e9",
          8018 => x"dc",
          8019 => x"51",
          8020 => x"82",
          8021 => x"55",
          8022 => x"08",
          8023 => x"55",
          8024 => x"82",
          8025 => x"84",
          8026 => x"82",
          8027 => x"80",
          8028 => x"51",
          8029 => x"82",
          8030 => x"82",
          8031 => x"30",
          8032 => x"dc",
          8033 => x"25",
          8034 => x"75",
          8035 => x"38",
          8036 => x"8f",
          8037 => x"75",
          8038 => x"c1",
          8039 => x"bb",
          8040 => x"74",
          8041 => x"51",
          8042 => x"3f",
          8043 => x"08",
          8044 => x"bb",
          8045 => x"3d",
          8046 => x"3d",
          8047 => x"99",
          8048 => x"52",
          8049 => x"d8",
          8050 => x"bb",
          8051 => x"82",
          8052 => x"82",
          8053 => x"5e",
          8054 => x"3d",
          8055 => x"cf",
          8056 => x"bb",
          8057 => x"82",
          8058 => x"86",
          8059 => x"82",
          8060 => x"bb",
          8061 => x"2e",
          8062 => x"82",
          8063 => x"80",
          8064 => x"70",
          8065 => x"06",
          8066 => x"54",
          8067 => x"38",
          8068 => x"52",
          8069 => x"52",
          8070 => x"3f",
          8071 => x"08",
          8072 => x"82",
          8073 => x"83",
          8074 => x"82",
          8075 => x"81",
          8076 => x"06",
          8077 => x"54",
          8078 => x"08",
          8079 => x"81",
          8080 => x"81",
          8081 => x"39",
          8082 => x"38",
          8083 => x"08",
          8084 => x"c4",
          8085 => x"bb",
          8086 => x"82",
          8087 => x"81",
          8088 => x"53",
          8089 => x"19",
          8090 => x"8c",
          8091 => x"ae",
          8092 => x"34",
          8093 => x"0b",
          8094 => x"82",
          8095 => x"52",
          8096 => x"51",
          8097 => x"3f",
          8098 => x"b4",
          8099 => x"c9",
          8100 => x"53",
          8101 => x"53",
          8102 => x"51",
          8103 => x"3f",
          8104 => x"0b",
          8105 => x"34",
          8106 => x"80",
          8107 => x"51",
          8108 => x"78",
          8109 => x"83",
          8110 => x"51",
          8111 => x"82",
          8112 => x"54",
          8113 => x"08",
          8114 => x"88",
          8115 => x"64",
          8116 => x"ff",
          8117 => x"75",
          8118 => x"78",
          8119 => x"3f",
          8120 => x"0b",
          8121 => x"78",
          8122 => x"83",
          8123 => x"51",
          8124 => x"3f",
          8125 => x"08",
          8126 => x"80",
          8127 => x"76",
          8128 => x"ae",
          8129 => x"bb",
          8130 => x"3d",
          8131 => x"3d",
          8132 => x"84",
          8133 => x"f1",
          8134 => x"a8",
          8135 => x"05",
          8136 => x"51",
          8137 => x"82",
          8138 => x"55",
          8139 => x"08",
          8140 => x"78",
          8141 => x"08",
          8142 => x"70",
          8143 => x"b8",
          8144 => x"dc",
          8145 => x"bb",
          8146 => x"b9",
          8147 => x"9b",
          8148 => x"a0",
          8149 => x"55",
          8150 => x"38",
          8151 => x"3d",
          8152 => x"3d",
          8153 => x"51",
          8154 => x"3f",
          8155 => x"52",
          8156 => x"52",
          8157 => x"dd",
          8158 => x"08",
          8159 => x"cb",
          8160 => x"bb",
          8161 => x"82",
          8162 => x"95",
          8163 => x"2e",
          8164 => x"88",
          8165 => x"3d",
          8166 => x"38",
          8167 => x"e5",
          8168 => x"dc",
          8169 => x"09",
          8170 => x"b8",
          8171 => x"c9",
          8172 => x"bb",
          8173 => x"82",
          8174 => x"81",
          8175 => x"56",
          8176 => x"3d",
          8177 => x"52",
          8178 => x"ff",
          8179 => x"02",
          8180 => x"8b",
          8181 => x"16",
          8182 => x"2a",
          8183 => x"51",
          8184 => x"89",
          8185 => x"07",
          8186 => x"17",
          8187 => x"81",
          8188 => x"34",
          8189 => x"70",
          8190 => x"81",
          8191 => x"55",
          8192 => x"80",
          8193 => x"64",
          8194 => x"38",
          8195 => x"51",
          8196 => x"82",
          8197 => x"52",
          8198 => x"b7",
          8199 => x"55",
          8200 => x"08",
          8201 => x"dd",
          8202 => x"dc",
          8203 => x"51",
          8204 => x"3f",
          8205 => x"08",
          8206 => x"11",
          8207 => x"82",
          8208 => x"80",
          8209 => x"16",
          8210 => x"ae",
          8211 => x"06",
          8212 => x"53",
          8213 => x"51",
          8214 => x"78",
          8215 => x"83",
          8216 => x"39",
          8217 => x"08",
          8218 => x"51",
          8219 => x"82",
          8220 => x"55",
          8221 => x"08",
          8222 => x"51",
          8223 => x"3f",
          8224 => x"08",
          8225 => x"bb",
          8226 => x"3d",
          8227 => x"3d",
          8228 => x"db",
          8229 => x"84",
          8230 => x"05",
          8231 => x"82",
          8232 => x"d0",
          8233 => x"3d",
          8234 => x"3f",
          8235 => x"08",
          8236 => x"dc",
          8237 => x"38",
          8238 => x"52",
          8239 => x"05",
          8240 => x"3f",
          8241 => x"08",
          8242 => x"dc",
          8243 => x"02",
          8244 => x"33",
          8245 => x"54",
          8246 => x"aa",
          8247 => x"06",
          8248 => x"8b",
          8249 => x"06",
          8250 => x"07",
          8251 => x"56",
          8252 => x"34",
          8253 => x"0b",
          8254 => x"78",
          8255 => x"a9",
          8256 => x"dc",
          8257 => x"82",
          8258 => x"95",
          8259 => x"ef",
          8260 => x"56",
          8261 => x"3d",
          8262 => x"94",
          8263 => x"f4",
          8264 => x"dc",
          8265 => x"bb",
          8266 => x"cb",
          8267 => x"63",
          8268 => x"d4",
          8269 => x"c0",
          8270 => x"dc",
          8271 => x"bb",
          8272 => x"38",
          8273 => x"05",
          8274 => x"06",
          8275 => x"73",
          8276 => x"16",
          8277 => x"22",
          8278 => x"07",
          8279 => x"1f",
          8280 => x"c2",
          8281 => x"81",
          8282 => x"34",
          8283 => x"b3",
          8284 => x"bb",
          8285 => x"74",
          8286 => x"0c",
          8287 => x"04",
          8288 => x"69",
          8289 => x"80",
          8290 => x"d0",
          8291 => x"3d",
          8292 => x"3f",
          8293 => x"08",
          8294 => x"08",
          8295 => x"bb",
          8296 => x"80",
          8297 => x"57",
          8298 => x"81",
          8299 => x"70",
          8300 => x"55",
          8301 => x"80",
          8302 => x"5d",
          8303 => x"52",
          8304 => x"52",
          8305 => x"a9",
          8306 => x"dc",
          8307 => x"bb",
          8308 => x"d1",
          8309 => x"73",
          8310 => x"3f",
          8311 => x"08",
          8312 => x"dc",
          8313 => x"82",
          8314 => x"82",
          8315 => x"65",
          8316 => x"78",
          8317 => x"7b",
          8318 => x"55",
          8319 => x"34",
          8320 => x"8a",
          8321 => x"38",
          8322 => x"1a",
          8323 => x"34",
          8324 => x"9e",
          8325 => x"70",
          8326 => x"51",
          8327 => x"a0",
          8328 => x"8e",
          8329 => x"2e",
          8330 => x"86",
          8331 => x"34",
          8332 => x"30",
          8333 => x"80",
          8334 => x"7a",
          8335 => x"c1",
          8336 => x"2e",
          8337 => x"a0",
          8338 => x"51",
          8339 => x"3f",
          8340 => x"08",
          8341 => x"dc",
          8342 => x"7b",
          8343 => x"55",
          8344 => x"73",
          8345 => x"38",
          8346 => x"73",
          8347 => x"38",
          8348 => x"15",
          8349 => x"ff",
          8350 => x"82",
          8351 => x"7b",
          8352 => x"bb",
          8353 => x"3d",
          8354 => x"3d",
          8355 => x"9c",
          8356 => x"05",
          8357 => x"51",
          8358 => x"82",
          8359 => x"82",
          8360 => x"56",
          8361 => x"dc",
          8362 => x"38",
          8363 => x"52",
          8364 => x"52",
          8365 => x"c0",
          8366 => x"70",
          8367 => x"ff",
          8368 => x"55",
          8369 => x"27",
          8370 => x"78",
          8371 => x"ff",
          8372 => x"05",
          8373 => x"55",
          8374 => x"3f",
          8375 => x"08",
          8376 => x"38",
          8377 => x"70",
          8378 => x"ff",
          8379 => x"82",
          8380 => x"80",
          8381 => x"74",
          8382 => x"07",
          8383 => x"4e",
          8384 => x"82",
          8385 => x"55",
          8386 => x"70",
          8387 => x"06",
          8388 => x"99",
          8389 => x"e0",
          8390 => x"ff",
          8391 => x"54",
          8392 => x"27",
          8393 => x"b4",
          8394 => x"55",
          8395 => x"a3",
          8396 => x"82",
          8397 => x"ff",
          8398 => x"82",
          8399 => x"93",
          8400 => x"75",
          8401 => x"76",
          8402 => x"38",
          8403 => x"77",
          8404 => x"86",
          8405 => x"39",
          8406 => x"27",
          8407 => x"88",
          8408 => x"78",
          8409 => x"5a",
          8410 => x"57",
          8411 => x"81",
          8412 => x"81",
          8413 => x"33",
          8414 => x"06",
          8415 => x"57",
          8416 => x"fe",
          8417 => x"3d",
          8418 => x"55",
          8419 => x"2e",
          8420 => x"76",
          8421 => x"38",
          8422 => x"55",
          8423 => x"33",
          8424 => x"a0",
          8425 => x"06",
          8426 => x"17",
          8427 => x"38",
          8428 => x"43",
          8429 => x"3d",
          8430 => x"ff",
          8431 => x"82",
          8432 => x"54",
          8433 => x"08",
          8434 => x"81",
          8435 => x"ff",
          8436 => x"82",
          8437 => x"54",
          8438 => x"08",
          8439 => x"80",
          8440 => x"54",
          8441 => x"80",
          8442 => x"bb",
          8443 => x"2e",
          8444 => x"80",
          8445 => x"54",
          8446 => x"80",
          8447 => x"52",
          8448 => x"bd",
          8449 => x"bb",
          8450 => x"82",
          8451 => x"b1",
          8452 => x"82",
          8453 => x"52",
          8454 => x"ab",
          8455 => x"54",
          8456 => x"15",
          8457 => x"78",
          8458 => x"ff",
          8459 => x"79",
          8460 => x"83",
          8461 => x"51",
          8462 => x"3f",
          8463 => x"08",
          8464 => x"74",
          8465 => x"0c",
          8466 => x"04",
          8467 => x"60",
          8468 => x"05",
          8469 => x"33",
          8470 => x"05",
          8471 => x"40",
          8472 => x"da",
          8473 => x"dc",
          8474 => x"bb",
          8475 => x"bd",
          8476 => x"33",
          8477 => x"b5",
          8478 => x"2e",
          8479 => x"1a",
          8480 => x"90",
          8481 => x"33",
          8482 => x"70",
          8483 => x"55",
          8484 => x"38",
          8485 => x"97",
          8486 => x"82",
          8487 => x"58",
          8488 => x"7e",
          8489 => x"70",
          8490 => x"55",
          8491 => x"56",
          8492 => x"d2",
          8493 => x"7d",
          8494 => x"70",
          8495 => x"2a",
          8496 => x"08",
          8497 => x"08",
          8498 => x"5d",
          8499 => x"77",
          8500 => x"98",
          8501 => x"26",
          8502 => x"57",
          8503 => x"59",
          8504 => x"52",
          8505 => x"ae",
          8506 => x"15",
          8507 => x"98",
          8508 => x"26",
          8509 => x"55",
          8510 => x"08",
          8511 => x"99",
          8512 => x"dc",
          8513 => x"ff",
          8514 => x"bb",
          8515 => x"38",
          8516 => x"75",
          8517 => x"81",
          8518 => x"93",
          8519 => x"80",
          8520 => x"2e",
          8521 => x"ff",
          8522 => x"58",
          8523 => x"7d",
          8524 => x"38",
          8525 => x"55",
          8526 => x"b4",
          8527 => x"56",
          8528 => x"09",
          8529 => x"38",
          8530 => x"53",
          8531 => x"51",
          8532 => x"3f",
          8533 => x"08",
          8534 => x"dc",
          8535 => x"38",
          8536 => x"ff",
          8537 => x"5c",
          8538 => x"84",
          8539 => x"5c",
          8540 => x"12",
          8541 => x"80",
          8542 => x"78",
          8543 => x"7c",
          8544 => x"90",
          8545 => x"c0",
          8546 => x"90",
          8547 => x"15",
          8548 => x"90",
          8549 => x"54",
          8550 => x"91",
          8551 => x"31",
          8552 => x"84",
          8553 => x"07",
          8554 => x"16",
          8555 => x"73",
          8556 => x"0c",
          8557 => x"04",
          8558 => x"6b",
          8559 => x"05",
          8560 => x"33",
          8561 => x"5a",
          8562 => x"bd",
          8563 => x"80",
          8564 => x"dc",
          8565 => x"f8",
          8566 => x"dc",
          8567 => x"82",
          8568 => x"70",
          8569 => x"74",
          8570 => x"38",
          8571 => x"82",
          8572 => x"81",
          8573 => x"81",
          8574 => x"ff",
          8575 => x"82",
          8576 => x"81",
          8577 => x"81",
          8578 => x"83",
          8579 => x"c0",
          8580 => x"2a",
          8581 => x"51",
          8582 => x"74",
          8583 => x"99",
          8584 => x"53",
          8585 => x"51",
          8586 => x"3f",
          8587 => x"08",
          8588 => x"55",
          8589 => x"92",
          8590 => x"80",
          8591 => x"38",
          8592 => x"06",
          8593 => x"2e",
          8594 => x"48",
          8595 => x"87",
          8596 => x"79",
          8597 => x"78",
          8598 => x"26",
          8599 => x"19",
          8600 => x"74",
          8601 => x"38",
          8602 => x"e4",
          8603 => x"2a",
          8604 => x"70",
          8605 => x"59",
          8606 => x"7a",
          8607 => x"56",
          8608 => x"80",
          8609 => x"51",
          8610 => x"74",
          8611 => x"99",
          8612 => x"53",
          8613 => x"51",
          8614 => x"3f",
          8615 => x"bb",
          8616 => x"ac",
          8617 => x"2a",
          8618 => x"82",
          8619 => x"43",
          8620 => x"83",
          8621 => x"66",
          8622 => x"60",
          8623 => x"90",
          8624 => x"31",
          8625 => x"80",
          8626 => x"8a",
          8627 => x"56",
          8628 => x"26",
          8629 => x"77",
          8630 => x"81",
          8631 => x"74",
          8632 => x"38",
          8633 => x"55",
          8634 => x"83",
          8635 => x"81",
          8636 => x"80",
          8637 => x"38",
          8638 => x"55",
          8639 => x"5e",
          8640 => x"89",
          8641 => x"5a",
          8642 => x"09",
          8643 => x"e1",
          8644 => x"38",
          8645 => x"57",
          8646 => x"b6",
          8647 => x"5a",
          8648 => x"9d",
          8649 => x"26",
          8650 => x"b6",
          8651 => x"10",
          8652 => x"22",
          8653 => x"74",
          8654 => x"38",
          8655 => x"ee",
          8656 => x"66",
          8657 => x"be",
          8658 => x"dc",
          8659 => x"84",
          8660 => x"89",
          8661 => x"a0",
          8662 => x"82",
          8663 => x"fc",
          8664 => x"56",
          8665 => x"f0",
          8666 => x"80",
          8667 => x"d3",
          8668 => x"38",
          8669 => x"57",
          8670 => x"b6",
          8671 => x"5a",
          8672 => x"9d",
          8673 => x"26",
          8674 => x"b6",
          8675 => x"10",
          8676 => x"22",
          8677 => x"74",
          8678 => x"38",
          8679 => x"ee",
          8680 => x"66",
          8681 => x"de",
          8682 => x"dc",
          8683 => x"05",
          8684 => x"dc",
          8685 => x"26",
          8686 => x"0b",
          8687 => x"08",
          8688 => x"dc",
          8689 => x"11",
          8690 => x"05",
          8691 => x"83",
          8692 => x"2a",
          8693 => x"a0",
          8694 => x"7d",
          8695 => x"69",
          8696 => x"05",
          8697 => x"72",
          8698 => x"5c",
          8699 => x"59",
          8700 => x"2e",
          8701 => x"89",
          8702 => x"60",
          8703 => x"84",
          8704 => x"5d",
          8705 => x"18",
          8706 => x"68",
          8707 => x"74",
          8708 => x"af",
          8709 => x"31",
          8710 => x"53",
          8711 => x"52",
          8712 => x"e2",
          8713 => x"dc",
          8714 => x"83",
          8715 => x"06",
          8716 => x"bb",
          8717 => x"ff",
          8718 => x"dd",
          8719 => x"83",
          8720 => x"2a",
          8721 => x"be",
          8722 => x"39",
          8723 => x"09",
          8724 => x"c5",
          8725 => x"f5",
          8726 => x"dc",
          8727 => x"38",
          8728 => x"79",
          8729 => x"80",
          8730 => x"38",
          8731 => x"96",
          8732 => x"06",
          8733 => x"2e",
          8734 => x"5e",
          8735 => x"82",
          8736 => x"9f",
          8737 => x"38",
          8738 => x"38",
          8739 => x"81",
          8740 => x"fc",
          8741 => x"ab",
          8742 => x"7d",
          8743 => x"81",
          8744 => x"7d",
          8745 => x"78",
          8746 => x"74",
          8747 => x"8e",
          8748 => x"9c",
          8749 => x"53",
          8750 => x"51",
          8751 => x"3f",
          8752 => x"b4",
          8753 => x"51",
          8754 => x"3f",
          8755 => x"8b",
          8756 => x"a1",
          8757 => x"8d",
          8758 => x"83",
          8759 => x"52",
          8760 => x"ff",
          8761 => x"81",
          8762 => x"34",
          8763 => x"70",
          8764 => x"2a",
          8765 => x"54",
          8766 => x"1b",
          8767 => x"88",
          8768 => x"74",
          8769 => x"26",
          8770 => x"83",
          8771 => x"52",
          8772 => x"ff",
          8773 => x"8a",
          8774 => x"a0",
          8775 => x"a1",
          8776 => x"0b",
          8777 => x"bf",
          8778 => x"51",
          8779 => x"3f",
          8780 => x"9a",
          8781 => x"a0",
          8782 => x"52",
          8783 => x"ff",
          8784 => x"7d",
          8785 => x"81",
          8786 => x"38",
          8787 => x"0a",
          8788 => x"1b",
          8789 => x"ce",
          8790 => x"a4",
          8791 => x"a0",
          8792 => x"52",
          8793 => x"ff",
          8794 => x"81",
          8795 => x"51",
          8796 => x"3f",
          8797 => x"1b",
          8798 => x"8c",
          8799 => x"0b",
          8800 => x"34",
          8801 => x"c2",
          8802 => x"53",
          8803 => x"52",
          8804 => x"51",
          8805 => x"88",
          8806 => x"a7",
          8807 => x"a0",
          8808 => x"83",
          8809 => x"52",
          8810 => x"ff",
          8811 => x"ff",
          8812 => x"1c",
          8813 => x"a6",
          8814 => x"53",
          8815 => x"52",
          8816 => x"ff",
          8817 => x"82",
          8818 => x"83",
          8819 => x"52",
          8820 => x"b4",
          8821 => x"60",
          8822 => x"7e",
          8823 => x"d7",
          8824 => x"82",
          8825 => x"83",
          8826 => x"83",
          8827 => x"06",
          8828 => x"75",
          8829 => x"05",
          8830 => x"7e",
          8831 => x"b7",
          8832 => x"53",
          8833 => x"51",
          8834 => x"3f",
          8835 => x"a4",
          8836 => x"51",
          8837 => x"3f",
          8838 => x"e4",
          8839 => x"e4",
          8840 => x"9f",
          8841 => x"18",
          8842 => x"1b",
          8843 => x"f6",
          8844 => x"83",
          8845 => x"ff",
          8846 => x"82",
          8847 => x"78",
          8848 => x"c4",
          8849 => x"60",
          8850 => x"7a",
          8851 => x"ff",
          8852 => x"75",
          8853 => x"53",
          8854 => x"51",
          8855 => x"3f",
          8856 => x"52",
          8857 => x"9f",
          8858 => x"56",
          8859 => x"83",
          8860 => x"06",
          8861 => x"52",
          8862 => x"9e",
          8863 => x"52",
          8864 => x"ff",
          8865 => x"f0",
          8866 => x"1b",
          8867 => x"87",
          8868 => x"55",
          8869 => x"83",
          8870 => x"74",
          8871 => x"ff",
          8872 => x"7c",
          8873 => x"74",
          8874 => x"38",
          8875 => x"54",
          8876 => x"52",
          8877 => x"99",
          8878 => x"bb",
          8879 => x"87",
          8880 => x"53",
          8881 => x"08",
          8882 => x"ff",
          8883 => x"76",
          8884 => x"31",
          8885 => x"cd",
          8886 => x"58",
          8887 => x"ff",
          8888 => x"55",
          8889 => x"83",
          8890 => x"61",
          8891 => x"26",
          8892 => x"57",
          8893 => x"53",
          8894 => x"51",
          8895 => x"3f",
          8896 => x"08",
          8897 => x"76",
          8898 => x"31",
          8899 => x"db",
          8900 => x"7d",
          8901 => x"38",
          8902 => x"83",
          8903 => x"8a",
          8904 => x"7d",
          8905 => x"38",
          8906 => x"81",
          8907 => x"80",
          8908 => x"80",
          8909 => x"7a",
          8910 => x"bc",
          8911 => x"d5",
          8912 => x"ff",
          8913 => x"83",
          8914 => x"77",
          8915 => x"0b",
          8916 => x"81",
          8917 => x"34",
          8918 => x"34",
          8919 => x"34",
          8920 => x"56",
          8921 => x"52",
          8922 => x"b0",
          8923 => x"0b",
          8924 => x"82",
          8925 => x"82",
          8926 => x"56",
          8927 => x"34",
          8928 => x"08",
          8929 => x"60",
          8930 => x"1b",
          8931 => x"96",
          8932 => x"83",
          8933 => x"ff",
          8934 => x"81",
          8935 => x"7a",
          8936 => x"ff",
          8937 => x"81",
          8938 => x"dc",
          8939 => x"80",
          8940 => x"7e",
          8941 => x"e3",
          8942 => x"82",
          8943 => x"90",
          8944 => x"8e",
          8945 => x"81",
          8946 => x"82",
          8947 => x"56",
          8948 => x"dc",
          8949 => x"0d",
          8950 => x"0d",
          8951 => x"59",
          8952 => x"ff",
          8953 => x"57",
          8954 => x"b4",
          8955 => x"f8",
          8956 => x"81",
          8957 => x"52",
          8958 => x"dc",
          8959 => x"2e",
          8960 => x"9c",
          8961 => x"33",
          8962 => x"2e",
          8963 => x"76",
          8964 => x"58",
          8965 => x"57",
          8966 => x"09",
          8967 => x"38",
          8968 => x"78",
          8969 => x"38",
          8970 => x"82",
          8971 => x"8d",
          8972 => x"f7",
          8973 => x"02",
          8974 => x"05",
          8975 => x"77",
          8976 => x"81",
          8977 => x"8d",
          8978 => x"e7",
          8979 => x"08",
          8980 => x"24",
          8981 => x"17",
          8982 => x"8c",
          8983 => x"77",
          8984 => x"16",
          8985 => x"25",
          8986 => x"3d",
          8987 => x"75",
          8988 => x"52",
          8989 => x"cb",
          8990 => x"76",
          8991 => x"70",
          8992 => x"2a",
          8993 => x"51",
          8994 => x"84",
          8995 => x"19",
          8996 => x"8b",
          8997 => x"f9",
          8998 => x"84",
          8999 => x"56",
          9000 => x"a7",
          9001 => x"fc",
          9002 => x"53",
          9003 => x"75",
          9004 => x"a1",
          9005 => x"dc",
          9006 => x"84",
          9007 => x"2e",
          9008 => x"87",
          9009 => x"08",
          9010 => x"ff",
          9011 => x"bb",
          9012 => x"3d",
          9013 => x"3d",
          9014 => x"80",
          9015 => x"52",
          9016 => x"9a",
          9017 => x"74",
          9018 => x"0d",
          9019 => x"0d",
          9020 => x"05",
          9021 => x"86",
          9022 => x"54",
          9023 => x"73",
          9024 => x"fe",
          9025 => x"51",
          9026 => x"98",
          9027 => x"00",
          9028 => x"ff",
          9029 => x"ff",
          9030 => x"ff",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"00",
          9136 => x"00",
          9137 => x"00",
          9138 => x"00",
          9139 => x"00",
          9140 => x"00",
          9141 => x"00",
          9142 => x"00",
          9143 => x"00",
          9144 => x"00",
          9145 => x"00",
          9146 => x"00",
          9147 => x"00",
          9148 => x"00",
          9149 => x"00",
          9150 => x"00",
          9151 => x"00",
          9152 => x"00",
          9153 => x"00",
          9154 => x"00",
          9155 => x"00",
          9156 => x"00",
          9157 => x"00",
          9158 => x"00",
          9159 => x"00",
          9160 => x"00",
          9161 => x"00",
          9162 => x"00",
          9163 => x"00",
          9164 => x"00",
          9165 => x"00",
          9166 => x"00",
          9167 => x"64",
          9168 => x"74",
          9169 => x"64",
          9170 => x"74",
          9171 => x"66",
          9172 => x"74",
          9173 => x"66",
          9174 => x"64",
          9175 => x"66",
          9176 => x"63",
          9177 => x"6d",
          9178 => x"61",
          9179 => x"6d",
          9180 => x"79",
          9181 => x"6d",
          9182 => x"66",
          9183 => x"6d",
          9184 => x"70",
          9185 => x"6d",
          9186 => x"6d",
          9187 => x"6d",
          9188 => x"68",
          9189 => x"68",
          9190 => x"68",
          9191 => x"68",
          9192 => x"63",
          9193 => x"00",
          9194 => x"6a",
          9195 => x"72",
          9196 => x"61",
          9197 => x"72",
          9198 => x"74",
          9199 => x"69",
          9200 => x"00",
          9201 => x"74",
          9202 => x"00",
          9203 => x"74",
          9204 => x"69",
          9205 => x"6d",
          9206 => x"69",
          9207 => x"6b",
          9208 => x"00",
          9209 => x"65",
          9210 => x"44",
          9211 => x"20",
          9212 => x"6f",
          9213 => x"49",
          9214 => x"72",
          9215 => x"20",
          9216 => x"6f",
          9217 => x"44",
          9218 => x"20",
          9219 => x"20",
          9220 => x"64",
          9221 => x"4e",
          9222 => x"69",
          9223 => x"66",
          9224 => x"64",
          9225 => x"4e",
          9226 => x"61",
          9227 => x"66",
          9228 => x"64",
          9229 => x"49",
          9230 => x"6c",
          9231 => x"66",
          9232 => x"6e",
          9233 => x"2e",
          9234 => x"41",
          9235 => x"73",
          9236 => x"65",
          9237 => x"64",
          9238 => x"46",
          9239 => x"20",
          9240 => x"65",
          9241 => x"20",
          9242 => x"73",
          9243 => x"00",
          9244 => x"46",
          9245 => x"20",
          9246 => x"64",
          9247 => x"69",
          9248 => x"6c",
          9249 => x"00",
          9250 => x"53",
          9251 => x"73",
          9252 => x"69",
          9253 => x"70",
          9254 => x"65",
          9255 => x"64",
          9256 => x"44",
          9257 => x"65",
          9258 => x"6d",
          9259 => x"20",
          9260 => x"69",
          9261 => x"6c",
          9262 => x"00",
          9263 => x"44",
          9264 => x"20",
          9265 => x"20",
          9266 => x"62",
          9267 => x"2e",
          9268 => x"4e",
          9269 => x"6f",
          9270 => x"74",
          9271 => x"65",
          9272 => x"6c",
          9273 => x"73",
          9274 => x"20",
          9275 => x"6e",
          9276 => x"6e",
          9277 => x"73",
          9278 => x"46",
          9279 => x"61",
          9280 => x"62",
          9281 => x"65",
          9282 => x"54",
          9283 => x"6f",
          9284 => x"20",
          9285 => x"72",
          9286 => x"6f",
          9287 => x"61",
          9288 => x"6c",
          9289 => x"2e",
          9290 => x"46",
          9291 => x"20",
          9292 => x"6c",
          9293 => x"65",
          9294 => x"49",
          9295 => x"66",
          9296 => x"69",
          9297 => x"20",
          9298 => x"6f",
          9299 => x"00",
          9300 => x"54",
          9301 => x"6d",
          9302 => x"20",
          9303 => x"6e",
          9304 => x"6c",
          9305 => x"00",
          9306 => x"50",
          9307 => x"6d",
          9308 => x"72",
          9309 => x"6e",
          9310 => x"72",
          9311 => x"2e",
          9312 => x"53",
          9313 => x"65",
          9314 => x"00",
          9315 => x"55",
          9316 => x"6f",
          9317 => x"65",
          9318 => x"72",
          9319 => x"0a",
          9320 => x"20",
          9321 => x"65",
          9322 => x"73",
          9323 => x"20",
          9324 => x"20",
          9325 => x"65",
          9326 => x"65",
          9327 => x"00",
          9328 => x"72",
          9329 => x"00",
          9330 => x"25",
          9331 => x"58",
          9332 => x"3a",
          9333 => x"25",
          9334 => x"00",
          9335 => x"20",
          9336 => x"20",
          9337 => x"00",
          9338 => x"25",
          9339 => x"00",
          9340 => x"20",
          9341 => x"20",
          9342 => x"7c",
          9343 => x"5a",
          9344 => x"41",
          9345 => x"0a",
          9346 => x"25",
          9347 => x"00",
          9348 => x"30",
          9349 => x"35",
          9350 => x"32",
          9351 => x"76",
          9352 => x"32",
          9353 => x"20",
          9354 => x"2c",
          9355 => x"76",
          9356 => x"32",
          9357 => x"25",
          9358 => x"73",
          9359 => x"0a",
          9360 => x"5a",
          9361 => x"41",
          9362 => x"74",
          9363 => x"75",
          9364 => x"48",
          9365 => x"6c",
          9366 => x"54",
          9367 => x"72",
          9368 => x"74",
          9369 => x"75",
          9370 => x"50",
          9371 => x"69",
          9372 => x"72",
          9373 => x"74",
          9374 => x"49",
          9375 => x"4c",
          9376 => x"20",
          9377 => x"65",
          9378 => x"70",
          9379 => x"49",
          9380 => x"4c",
          9381 => x"20",
          9382 => x"65",
          9383 => x"70",
          9384 => x"55",
          9385 => x"30",
          9386 => x"20",
          9387 => x"65",
          9388 => x"70",
          9389 => x"55",
          9390 => x"30",
          9391 => x"20",
          9392 => x"65",
          9393 => x"70",
          9394 => x"55",
          9395 => x"31",
          9396 => x"20",
          9397 => x"65",
          9398 => x"70",
          9399 => x"55",
          9400 => x"31",
          9401 => x"20",
          9402 => x"65",
          9403 => x"70",
          9404 => x"53",
          9405 => x"69",
          9406 => x"75",
          9407 => x"69",
          9408 => x"2e",
          9409 => x"45",
          9410 => x"6c",
          9411 => x"20",
          9412 => x"65",
          9413 => x"2e",
          9414 => x"61",
          9415 => x"65",
          9416 => x"2e",
          9417 => x"00",
          9418 => x"7a",
          9419 => x"61",
          9420 => x"74",
          9421 => x"30",
          9422 => x"46",
          9423 => x"65",
          9424 => x"6f",
          9425 => x"69",
          9426 => x"6c",
          9427 => x"20",
          9428 => x"63",
          9429 => x"20",
          9430 => x"70",
          9431 => x"73",
          9432 => x"6e",
          9433 => x"6d",
          9434 => x"61",
          9435 => x"2e",
          9436 => x"2a",
          9437 => x"42",
          9438 => x"64",
          9439 => x"20",
          9440 => x"00",
          9441 => x"49",
          9442 => x"69",
          9443 => x"73",
          9444 => x"00",
          9445 => x"46",
          9446 => x"65",
          9447 => x"6f",
          9448 => x"69",
          9449 => x"6c",
          9450 => x"2e",
          9451 => x"72",
          9452 => x"64",
          9453 => x"25",
          9454 => x"43",
          9455 => x"72",
          9456 => x"2e",
          9457 => x"00",
          9458 => x"43",
          9459 => x"69",
          9460 => x"2e",
          9461 => x"43",
          9462 => x"61",
          9463 => x"67",
          9464 => x"00",
          9465 => x"25",
          9466 => x"78",
          9467 => x"38",
          9468 => x"3e",
          9469 => x"6c",
          9470 => x"30",
          9471 => x"0a",
          9472 => x"44",
          9473 => x"20",
          9474 => x"6f",
          9475 => x"0a",
          9476 => x"70",
          9477 => x"65",
          9478 => x"25",
          9479 => x"58",
          9480 => x"32",
          9481 => x"3f",
          9482 => x"25",
          9483 => x"58",
          9484 => x"34",
          9485 => x"25",
          9486 => x"58",
          9487 => x"38",
          9488 => x"00",
          9489 => x"44",
          9490 => x"62",
          9491 => x"67",
          9492 => x"74",
          9493 => x"75",
          9494 => x"00",
          9495 => x"45",
          9496 => x"6c",
          9497 => x"20",
          9498 => x"65",
          9499 => x"70",
          9500 => x"44",
          9501 => x"62",
          9502 => x"20",
          9503 => x"74",
          9504 => x"66",
          9505 => x"45",
          9506 => x"6c",
          9507 => x"20",
          9508 => x"74",
          9509 => x"66",
          9510 => x"45",
          9511 => x"75",
          9512 => x"67",
          9513 => x"64",
          9514 => x"20",
          9515 => x"6c",
          9516 => x"2e",
          9517 => x"43",
          9518 => x"69",
          9519 => x"63",
          9520 => x"20",
          9521 => x"30",
          9522 => x"20",
          9523 => x"0a",
          9524 => x"43",
          9525 => x"20",
          9526 => x"75",
          9527 => x"64",
          9528 => x"64",
          9529 => x"25",
          9530 => x"0a",
          9531 => x"52",
          9532 => x"61",
          9533 => x"6e",
          9534 => x"70",
          9535 => x"63",
          9536 => x"6f",
          9537 => x"2e",
          9538 => x"43",
          9539 => x"20",
          9540 => x"6f",
          9541 => x"6e",
          9542 => x"2e",
          9543 => x"5a",
          9544 => x"62",
          9545 => x"25",
          9546 => x"25",
          9547 => x"73",
          9548 => x"00",
          9549 => x"25",
          9550 => x"25",
          9551 => x"73",
          9552 => x"25",
          9553 => x"25",
          9554 => x"42",
          9555 => x"63",
          9556 => x"61",
          9557 => x"00",
          9558 => x"52",
          9559 => x"69",
          9560 => x"2e",
          9561 => x"45",
          9562 => x"6c",
          9563 => x"20",
          9564 => x"65",
          9565 => x"70",
          9566 => x"2e",
          9567 => x"25",
          9568 => x"64",
          9569 => x"20",
          9570 => x"25",
          9571 => x"64",
          9572 => x"25",
          9573 => x"53",
          9574 => x"43",
          9575 => x"69",
          9576 => x"61",
          9577 => x"6e",
          9578 => x"20",
          9579 => x"6f",
          9580 => x"6f",
          9581 => x"6f",
          9582 => x"67",
          9583 => x"3a",
          9584 => x"76",
          9585 => x"73",
          9586 => x"70",
          9587 => x"65",
          9588 => x"64",
          9589 => x"20",
          9590 => x"57",
          9591 => x"44",
          9592 => x"20",
          9593 => x"30",
          9594 => x"25",
          9595 => x"29",
          9596 => x"20",
          9597 => x"53",
          9598 => x"4d",
          9599 => x"20",
          9600 => x"30",
          9601 => x"25",
          9602 => x"29",
          9603 => x"20",
          9604 => x"49",
          9605 => x"20",
          9606 => x"4d",
          9607 => x"30",
          9608 => x"25",
          9609 => x"29",
          9610 => x"20",
          9611 => x"42",
          9612 => x"20",
          9613 => x"20",
          9614 => x"30",
          9615 => x"25",
          9616 => x"29",
          9617 => x"20",
          9618 => x"52",
          9619 => x"20",
          9620 => x"20",
          9621 => x"30",
          9622 => x"25",
          9623 => x"29",
          9624 => x"20",
          9625 => x"53",
          9626 => x"41",
          9627 => x"20",
          9628 => x"65",
          9629 => x"65",
          9630 => x"25",
          9631 => x"29",
          9632 => x"20",
          9633 => x"54",
          9634 => x"52",
          9635 => x"20",
          9636 => x"69",
          9637 => x"73",
          9638 => x"25",
          9639 => x"29",
          9640 => x"20",
          9641 => x"49",
          9642 => x"20",
          9643 => x"4c",
          9644 => x"68",
          9645 => x"65",
          9646 => x"25",
          9647 => x"29",
          9648 => x"20",
          9649 => x"57",
          9650 => x"42",
          9651 => x"20",
          9652 => x"0a",
          9653 => x"20",
          9654 => x"57",
          9655 => x"32",
          9656 => x"20",
          9657 => x"49",
          9658 => x"4c",
          9659 => x"20",
          9660 => x"50",
          9661 => x"00",
          9662 => x"20",
          9663 => x"53",
          9664 => x"00",
          9665 => x"41",
          9666 => x"65",
          9667 => x"73",
          9668 => x"20",
          9669 => x"43",
          9670 => x"52",
          9671 => x"74",
          9672 => x"63",
          9673 => x"20",
          9674 => x"72",
          9675 => x"20",
          9676 => x"30",
          9677 => x"00",
          9678 => x"20",
          9679 => x"43",
          9680 => x"4d",
          9681 => x"72",
          9682 => x"74",
          9683 => x"20",
          9684 => x"72",
          9685 => x"20",
          9686 => x"30",
          9687 => x"00",
          9688 => x"20",
          9689 => x"53",
          9690 => x"6b",
          9691 => x"61",
          9692 => x"41",
          9693 => x"65",
          9694 => x"20",
          9695 => x"20",
          9696 => x"30",
          9697 => x"00",
          9698 => x"4d",
          9699 => x"3a",
          9700 => x"20",
          9701 => x"5a",
          9702 => x"49",
          9703 => x"20",
          9704 => x"20",
          9705 => x"20",
          9706 => x"20",
          9707 => x"20",
          9708 => x"30",
          9709 => x"00",
          9710 => x"20",
          9711 => x"53",
          9712 => x"65",
          9713 => x"6c",
          9714 => x"20",
          9715 => x"71",
          9716 => x"20",
          9717 => x"20",
          9718 => x"64",
          9719 => x"34",
          9720 => x"7a",
          9721 => x"20",
          9722 => x"53",
          9723 => x"4d",
          9724 => x"6f",
          9725 => x"46",
          9726 => x"20",
          9727 => x"20",
          9728 => x"20",
          9729 => x"64",
          9730 => x"34",
          9731 => x"7a",
          9732 => x"20",
          9733 => x"57",
          9734 => x"62",
          9735 => x"20",
          9736 => x"41",
          9737 => x"6c",
          9738 => x"20",
          9739 => x"71",
          9740 => x"64",
          9741 => x"34",
          9742 => x"7a",
          9743 => x"53",
          9744 => x"6c",
          9745 => x"4d",
          9746 => x"75",
          9747 => x"46",
          9748 => x"00",
          9749 => x"45",
          9750 => x"45",
          9751 => x"69",
          9752 => x"55",
          9753 => x"6f",
          9754 => x"00",
          9755 => x"01",
          9756 => x"00",
          9757 => x"00",
          9758 => x"01",
          9759 => x"00",
          9760 => x"00",
          9761 => x"01",
          9762 => x"00",
          9763 => x"00",
          9764 => x"01",
          9765 => x"00",
          9766 => x"00",
          9767 => x"01",
          9768 => x"00",
          9769 => x"00",
          9770 => x"01",
          9771 => x"00",
          9772 => x"00",
          9773 => x"01",
          9774 => x"00",
          9775 => x"00",
          9776 => x"01",
          9777 => x"00",
          9778 => x"00",
          9779 => x"01",
          9780 => x"00",
          9781 => x"00",
          9782 => x"01",
          9783 => x"00",
          9784 => x"00",
          9785 => x"01",
          9786 => x"00",
          9787 => x"00",
          9788 => x"04",
          9789 => x"00",
          9790 => x"00",
          9791 => x"04",
          9792 => x"00",
          9793 => x"00",
          9794 => x"04",
          9795 => x"00",
          9796 => x"00",
          9797 => x"03",
          9798 => x"00",
          9799 => x"00",
          9800 => x"04",
          9801 => x"00",
          9802 => x"00",
          9803 => x"04",
          9804 => x"00",
          9805 => x"00",
          9806 => x"04",
          9807 => x"00",
          9808 => x"00",
          9809 => x"03",
          9810 => x"00",
          9811 => x"00",
          9812 => x"03",
          9813 => x"00",
          9814 => x"00",
          9815 => x"03",
          9816 => x"00",
          9817 => x"00",
          9818 => x"03",
          9819 => x"00",
          9820 => x"1b",
          9821 => x"1b",
          9822 => x"1b",
          9823 => x"1b",
          9824 => x"1b",
          9825 => x"1b",
          9826 => x"1b",
          9827 => x"1b",
          9828 => x"1b",
          9829 => x"1b",
          9830 => x"1b",
          9831 => x"10",
          9832 => x"0e",
          9833 => x"0d",
          9834 => x"0b",
          9835 => x"08",
          9836 => x"06",
          9837 => x"05",
          9838 => x"04",
          9839 => x"03",
          9840 => x"02",
          9841 => x"01",
          9842 => x"68",
          9843 => x"6f",
          9844 => x"68",
          9845 => x"00",
          9846 => x"21",
          9847 => x"25",
          9848 => x"75",
          9849 => x"73",
          9850 => x"46",
          9851 => x"65",
          9852 => x"6f",
          9853 => x"73",
          9854 => x"74",
          9855 => x"68",
          9856 => x"6f",
          9857 => x"66",
          9858 => x"20",
          9859 => x"45",
          9860 => x"00",
          9861 => x"43",
          9862 => x"6f",
          9863 => x"70",
          9864 => x"63",
          9865 => x"74",
          9866 => x"69",
          9867 => x"72",
          9868 => x"69",
          9869 => x"20",
          9870 => x"61",
          9871 => x"6e",
          9872 => x"53",
          9873 => x"22",
          9874 => x"3a",
          9875 => x"3e",
          9876 => x"7c",
          9877 => x"46",
          9878 => x"46",
          9879 => x"32",
          9880 => x"eb",
          9881 => x"53",
          9882 => x"35",
          9883 => x"4e",
          9884 => x"41",
          9885 => x"20",
          9886 => x"41",
          9887 => x"20",
          9888 => x"4e",
          9889 => x"41",
          9890 => x"20",
          9891 => x"41",
          9892 => x"20",
          9893 => x"00",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"80",
          9898 => x"8e",
          9899 => x"45",
          9900 => x"49",
          9901 => x"90",
          9902 => x"99",
          9903 => x"59",
          9904 => x"9c",
          9905 => x"41",
          9906 => x"a5",
          9907 => x"a8",
          9908 => x"ac",
          9909 => x"b0",
          9910 => x"b4",
          9911 => x"b8",
          9912 => x"bc",
          9913 => x"c0",
          9914 => x"c4",
          9915 => x"c8",
          9916 => x"cc",
          9917 => x"d0",
          9918 => x"d4",
          9919 => x"d8",
          9920 => x"dc",
          9921 => x"e0",
          9922 => x"e4",
          9923 => x"e8",
          9924 => x"ec",
          9925 => x"f0",
          9926 => x"f4",
          9927 => x"f8",
          9928 => x"fc",
          9929 => x"2b",
          9930 => x"3d",
          9931 => x"5c",
          9932 => x"3c",
          9933 => x"7f",
          9934 => x"00",
          9935 => x"00",
          9936 => x"01",
          9937 => x"00",
          9938 => x"00",
          9939 => x"00",
          9940 => x"00",
          9941 => x"00",
          9942 => x"00",
          9943 => x"00",
          9944 => x"01",
          9945 => x"00",
          9946 => x"00",
          9947 => x"00",
          9948 => x"01",
          9949 => x"00",
          9950 => x"00",
          9951 => x"00",
          9952 => x"01",
          9953 => x"00",
          9954 => x"00",
          9955 => x"00",
          9956 => x"01",
          9957 => x"00",
          9958 => x"00",
          9959 => x"00",
          9960 => x"01",
          9961 => x"00",
          9962 => x"00",
          9963 => x"00",
          9964 => x"01",
          9965 => x"00",
          9966 => x"00",
          9967 => x"00",
          9968 => x"01",
          9969 => x"00",
          9970 => x"00",
          9971 => x"00",
          9972 => x"01",
          9973 => x"00",
          9974 => x"00",
          9975 => x"00",
          9976 => x"01",
          9977 => x"00",
          9978 => x"00",
          9979 => x"00",
          9980 => x"01",
          9981 => x"00",
          9982 => x"00",
          9983 => x"00",
          9984 => x"01",
          9985 => x"00",
          9986 => x"00",
          9987 => x"00",
          9988 => x"01",
          9989 => x"00",
          9990 => x"00",
          9991 => x"00",
          9992 => x"01",
          9993 => x"00",
          9994 => x"00",
          9995 => x"00",
          9996 => x"01",
          9997 => x"00",
          9998 => x"00",
          9999 => x"00",
         10000 => x"01",
         10001 => x"00",
         10002 => x"00",
         10003 => x"00",
         10004 => x"01",
         10005 => x"00",
         10006 => x"00",
         10007 => x"00",
         10008 => x"01",
         10009 => x"00",
         10010 => x"00",
         10011 => x"00",
         10012 => x"01",
         10013 => x"00",
         10014 => x"00",
         10015 => x"00",
         10016 => x"01",
         10017 => x"00",
         10018 => x"00",
         10019 => x"00",
         10020 => x"01",
         10021 => x"00",
         10022 => x"00",
         10023 => x"00",
         10024 => x"01",
         10025 => x"00",
         10026 => x"00",
         10027 => x"00",
         10028 => x"01",
         10029 => x"00",
         10030 => x"00",
         10031 => x"00",
         10032 => x"01",
         10033 => x"00",
         10034 => x"00",
         10035 => x"00",
         10036 => x"01",
         10037 => x"00",
         10038 => x"00",
         10039 => x"00",
         10040 => x"01",
         10041 => x"00",
         10042 => x"00",
         10043 => x"00",
         10044 => x"01",
         10045 => x"00",
         10046 => x"00",
         10047 => x"00",
         10048 => x"00",
         10049 => x"00",
         10050 => x"00",
         10051 => x"00",
         10052 => x"00",
         10053 => x"00",
         10054 => x"00",
         10055 => x"00",
         10056 => x"01",
         10057 => x"01",
         10058 => x"00",
         10059 => x"00",
         10060 => x"00",
         10061 => x"00",
         10062 => x"05",
         10063 => x"05",
         10064 => x"05",
         10065 => x"00",
         10066 => x"01",
         10067 => x"01",
         10068 => x"01",
         10069 => x"01",
         10070 => x"00",
         10071 => x"00",
         10072 => x"00",
         10073 => x"00",
         10074 => x"00",
         10075 => x"00",
         10076 => x"00",
         10077 => x"00",
         10078 => x"00",
         10079 => x"00",
         10080 => x"00",
         10081 => x"00",
         10082 => x"00",
         10083 => x"00",
         10084 => x"00",
         10085 => x"00",
         10086 => x"00",
         10087 => x"00",
         10088 => x"00",
         10089 => x"00",
         10090 => x"00",
         10091 => x"00",
         10092 => x"00",
         10093 => x"00",
         10094 => x"00",
         10095 => x"01",
         10096 => x"00",
         10097 => x"01",
         10098 => x"00",
         10099 => x"02",
         10100 => x"00",
         10101 => x"00",
         10102 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
