-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"ff",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"fe",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"99",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"cf",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"d1",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"a4",
           386 => x"f5",
           387 => x"a4",
           388 => x"90",
           389 => x"a4",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"82",
           395 => x"82",
           396 => x"82",
           397 => x"b4",
           398 => x"bb",
           399 => x"e0",
           400 => x"bb",
           401 => x"ab",
           402 => x"a4",
           403 => x"90",
           404 => x"a4",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"82",
           410 => x"82",
           411 => x"82",
           412 => x"af",
           413 => x"bb",
           414 => x"e0",
           415 => x"bb",
           416 => x"d6",
           417 => x"a4",
           418 => x"90",
           419 => x"a4",
           420 => x"2d",
           421 => x"08",
           422 => x"04",
           423 => x"0c",
           424 => x"82",
           425 => x"82",
           426 => x"82",
           427 => x"80",
           428 => x"82",
           429 => x"82",
           430 => x"82",
           431 => x"80",
           432 => x"82",
           433 => x"82",
           434 => x"82",
           435 => x"80",
           436 => x"82",
           437 => x"82",
           438 => x"82",
           439 => x"80",
           440 => x"82",
           441 => x"82",
           442 => x"82",
           443 => x"80",
           444 => x"82",
           445 => x"82",
           446 => x"82",
           447 => x"81",
           448 => x"82",
           449 => x"82",
           450 => x"82",
           451 => x"81",
           452 => x"82",
           453 => x"82",
           454 => x"82",
           455 => x"81",
           456 => x"82",
           457 => x"82",
           458 => x"82",
           459 => x"81",
           460 => x"82",
           461 => x"82",
           462 => x"82",
           463 => x"81",
           464 => x"82",
           465 => x"82",
           466 => x"82",
           467 => x"81",
           468 => x"82",
           469 => x"82",
           470 => x"82",
           471 => x"81",
           472 => x"82",
           473 => x"82",
           474 => x"82",
           475 => x"81",
           476 => x"82",
           477 => x"82",
           478 => x"82",
           479 => x"81",
           480 => x"82",
           481 => x"82",
           482 => x"82",
           483 => x"81",
           484 => x"82",
           485 => x"82",
           486 => x"82",
           487 => x"81",
           488 => x"82",
           489 => x"82",
           490 => x"82",
           491 => x"81",
           492 => x"82",
           493 => x"82",
           494 => x"82",
           495 => x"81",
           496 => x"82",
           497 => x"82",
           498 => x"82",
           499 => x"81",
           500 => x"82",
           501 => x"82",
           502 => x"82",
           503 => x"82",
           504 => x"82",
           505 => x"82",
           506 => x"82",
           507 => x"82",
           508 => x"82",
           509 => x"82",
           510 => x"82",
           511 => x"81",
           512 => x"82",
           513 => x"82",
           514 => x"82",
           515 => x"81",
           516 => x"82",
           517 => x"82",
           518 => x"82",
           519 => x"81",
           520 => x"82",
           521 => x"82",
           522 => x"82",
           523 => x"81",
           524 => x"82",
           525 => x"82",
           526 => x"82",
           527 => x"82",
           528 => x"82",
           529 => x"82",
           530 => x"82",
           531 => x"82",
           532 => x"82",
           533 => x"82",
           534 => x"82",
           535 => x"82",
           536 => x"82",
           537 => x"82",
           538 => x"82",
           539 => x"81",
           540 => x"82",
           541 => x"82",
           542 => x"82",
           543 => x"82",
           544 => x"82",
           545 => x"82",
           546 => x"82",
           547 => x"82",
           548 => x"82",
           549 => x"82",
           550 => x"82",
           551 => x"82",
           552 => x"82",
           553 => x"82",
           554 => x"82",
           555 => x"81",
           556 => x"82",
           557 => x"82",
           558 => x"82",
           559 => x"81",
           560 => x"82",
           561 => x"82",
           562 => x"82",
           563 => x"81",
           564 => x"82",
           565 => x"82",
           566 => x"82",
           567 => x"80",
           568 => x"82",
           569 => x"82",
           570 => x"82",
           571 => x"80",
           572 => x"82",
           573 => x"82",
           574 => x"82",
           575 => x"80",
           576 => x"82",
           577 => x"82",
           578 => x"82",
           579 => x"80",
           580 => x"82",
           581 => x"82",
           582 => x"82",
           583 => x"81",
           584 => x"82",
           585 => x"82",
           586 => x"82",
           587 => x"81",
           588 => x"82",
           589 => x"82",
           590 => x"82",
           591 => x"81",
           592 => x"82",
           593 => x"82",
           594 => x"82",
           595 => x"81",
           596 => x"82",
           597 => x"82",
           598 => x"3c",
           599 => x"10",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"51",
           608 => x"73",
           609 => x"73",
           610 => x"81",
           611 => x"10",
           612 => x"07",
           613 => x"0c",
           614 => x"72",
           615 => x"81",
           616 => x"09",
           617 => x"71",
           618 => x"0a",
           619 => x"72",
           620 => x"51",
           621 => x"82",
           622 => x"82",
           623 => x"8e",
           624 => x"70",
           625 => x"0c",
           626 => x"93",
           627 => x"81",
           628 => x"fe",
           629 => x"bb",
           630 => x"82",
           631 => x"fb",
           632 => x"bb",
           633 => x"05",
           634 => x"a4",
           635 => x"0c",
           636 => x"08",
           637 => x"54",
           638 => x"08",
           639 => x"53",
           640 => x"08",
           641 => x"9a",
           642 => x"98",
           643 => x"bb",
           644 => x"05",
           645 => x"a4",
           646 => x"08",
           647 => x"98",
           648 => x"87",
           649 => x"bb",
           650 => x"82",
           651 => x"02",
           652 => x"0c",
           653 => x"82",
           654 => x"90",
           655 => x"11",
           656 => x"32",
           657 => x"51",
           658 => x"71",
           659 => x"0b",
           660 => x"08",
           661 => x"25",
           662 => x"39",
           663 => x"bb",
           664 => x"05",
           665 => x"39",
           666 => x"08",
           667 => x"ff",
           668 => x"a4",
           669 => x"0c",
           670 => x"bb",
           671 => x"05",
           672 => x"a4",
           673 => x"08",
           674 => x"08",
           675 => x"82",
           676 => x"f8",
           677 => x"2e",
           678 => x"80",
           679 => x"a4",
           680 => x"08",
           681 => x"38",
           682 => x"08",
           683 => x"51",
           684 => x"82",
           685 => x"70",
           686 => x"08",
           687 => x"52",
           688 => x"08",
           689 => x"ff",
           690 => x"06",
           691 => x"0b",
           692 => x"08",
           693 => x"80",
           694 => x"bb",
           695 => x"05",
           696 => x"a4",
           697 => x"08",
           698 => x"73",
           699 => x"a4",
           700 => x"08",
           701 => x"bb",
           702 => x"05",
           703 => x"a4",
           704 => x"08",
           705 => x"bb",
           706 => x"05",
           707 => x"39",
           708 => x"08",
           709 => x"52",
           710 => x"82",
           711 => x"88",
           712 => x"82",
           713 => x"f4",
           714 => x"82",
           715 => x"f4",
           716 => x"bb",
           717 => x"3d",
           718 => x"a4",
           719 => x"bb",
           720 => x"82",
           721 => x"f4",
           722 => x"0b",
           723 => x"08",
           724 => x"82",
           725 => x"88",
           726 => x"bb",
           727 => x"05",
           728 => x"0b",
           729 => x"08",
           730 => x"82",
           731 => x"90",
           732 => x"bb",
           733 => x"05",
           734 => x"a4",
           735 => x"08",
           736 => x"a4",
           737 => x"08",
           738 => x"a4",
           739 => x"70",
           740 => x"81",
           741 => x"bb",
           742 => x"82",
           743 => x"dc",
           744 => x"bb",
           745 => x"05",
           746 => x"a4",
           747 => x"08",
           748 => x"80",
           749 => x"bb",
           750 => x"05",
           751 => x"bb",
           752 => x"8e",
           753 => x"bb",
           754 => x"82",
           755 => x"02",
           756 => x"0c",
           757 => x"82",
           758 => x"90",
           759 => x"bb",
           760 => x"05",
           761 => x"a4",
           762 => x"08",
           763 => x"a4",
           764 => x"08",
           765 => x"a4",
           766 => x"08",
           767 => x"3f",
           768 => x"08",
           769 => x"a4",
           770 => x"0c",
           771 => x"08",
           772 => x"70",
           773 => x"0c",
           774 => x"3d",
           775 => x"a4",
           776 => x"bb",
           777 => x"82",
           778 => x"ed",
           779 => x"0b",
           780 => x"08",
           781 => x"82",
           782 => x"88",
           783 => x"80",
           784 => x"0c",
           785 => x"08",
           786 => x"85",
           787 => x"81",
           788 => x"32",
           789 => x"51",
           790 => x"53",
           791 => x"8d",
           792 => x"82",
           793 => x"e0",
           794 => x"ac",
           795 => x"a4",
           796 => x"08",
           797 => x"53",
           798 => x"a4",
           799 => x"34",
           800 => x"06",
           801 => x"2e",
           802 => x"82",
           803 => x"8c",
           804 => x"05",
           805 => x"08",
           806 => x"82",
           807 => x"e4",
           808 => x"81",
           809 => x"72",
           810 => x"8b",
           811 => x"a4",
           812 => x"33",
           813 => x"27",
           814 => x"82",
           815 => x"f8",
           816 => x"72",
           817 => x"ee",
           818 => x"a4",
           819 => x"33",
           820 => x"2e",
           821 => x"80",
           822 => x"bb",
           823 => x"05",
           824 => x"2b",
           825 => x"51",
           826 => x"b2",
           827 => x"a4",
           828 => x"22",
           829 => x"70",
           830 => x"81",
           831 => x"51",
           832 => x"2e",
           833 => x"bb",
           834 => x"05",
           835 => x"80",
           836 => x"72",
           837 => x"08",
           838 => x"fe",
           839 => x"bb",
           840 => x"05",
           841 => x"2b",
           842 => x"70",
           843 => x"72",
           844 => x"51",
           845 => x"51",
           846 => x"82",
           847 => x"e8",
           848 => x"bb",
           849 => x"05",
           850 => x"bb",
           851 => x"05",
           852 => x"d0",
           853 => x"53",
           854 => x"a4",
           855 => x"34",
           856 => x"08",
           857 => x"70",
           858 => x"98",
           859 => x"53",
           860 => x"8b",
           861 => x"0b",
           862 => x"08",
           863 => x"82",
           864 => x"e4",
           865 => x"83",
           866 => x"06",
           867 => x"72",
           868 => x"82",
           869 => x"e8",
           870 => x"88",
           871 => x"2b",
           872 => x"70",
           873 => x"51",
           874 => x"72",
           875 => x"08",
           876 => x"fd",
           877 => x"bb",
           878 => x"05",
           879 => x"2a",
           880 => x"51",
           881 => x"80",
           882 => x"82",
           883 => x"e8",
           884 => x"98",
           885 => x"2c",
           886 => x"72",
           887 => x"0b",
           888 => x"08",
           889 => x"82",
           890 => x"f8",
           891 => x"11",
           892 => x"08",
           893 => x"53",
           894 => x"08",
           895 => x"80",
           896 => x"94",
           897 => x"a4",
           898 => x"08",
           899 => x"82",
           900 => x"70",
           901 => x"51",
           902 => x"82",
           903 => x"e4",
           904 => x"90",
           905 => x"72",
           906 => x"08",
           907 => x"82",
           908 => x"e4",
           909 => x"a0",
           910 => x"72",
           911 => x"08",
           912 => x"fc",
           913 => x"bb",
           914 => x"05",
           915 => x"80",
           916 => x"72",
           917 => x"08",
           918 => x"fc",
           919 => x"bb",
           920 => x"05",
           921 => x"c0",
           922 => x"72",
           923 => x"08",
           924 => x"fb",
           925 => x"bb",
           926 => x"05",
           927 => x"07",
           928 => x"82",
           929 => x"e4",
           930 => x"0b",
           931 => x"08",
           932 => x"fb",
           933 => x"bb",
           934 => x"05",
           935 => x"07",
           936 => x"82",
           937 => x"e4",
           938 => x"c1",
           939 => x"82",
           940 => x"fc",
           941 => x"bb",
           942 => x"05",
           943 => x"51",
           944 => x"bb",
           945 => x"05",
           946 => x"0b",
           947 => x"08",
           948 => x"8d",
           949 => x"bb",
           950 => x"05",
           951 => x"a4",
           952 => x"08",
           953 => x"bb",
           954 => x"05",
           955 => x"51",
           956 => x"bb",
           957 => x"05",
           958 => x"a4",
           959 => x"22",
           960 => x"53",
           961 => x"a4",
           962 => x"23",
           963 => x"82",
           964 => x"90",
           965 => x"bb",
           966 => x"05",
           967 => x"82",
           968 => x"90",
           969 => x"08",
           970 => x"08",
           971 => x"82",
           972 => x"e4",
           973 => x"83",
           974 => x"06",
           975 => x"53",
           976 => x"ab",
           977 => x"a4",
           978 => x"33",
           979 => x"53",
           980 => x"53",
           981 => x"08",
           982 => x"52",
           983 => x"3f",
           984 => x"08",
           985 => x"bb",
           986 => x"05",
           987 => x"82",
           988 => x"fc",
           989 => x"a8",
           990 => x"bb",
           991 => x"72",
           992 => x"08",
           993 => x"82",
           994 => x"ec",
           995 => x"82",
           996 => x"f4",
           997 => x"71",
           998 => x"72",
           999 => x"08",
          1000 => x"8b",
          1001 => x"bb",
          1002 => x"05",
          1003 => x"a4",
          1004 => x"08",
          1005 => x"bb",
          1006 => x"05",
          1007 => x"82",
          1008 => x"fc",
          1009 => x"bb",
          1010 => x"05",
          1011 => x"2a",
          1012 => x"51",
          1013 => x"72",
          1014 => x"38",
          1015 => x"08",
          1016 => x"70",
          1017 => x"72",
          1018 => x"82",
          1019 => x"fc",
          1020 => x"53",
          1021 => x"82",
          1022 => x"53",
          1023 => x"a4",
          1024 => x"23",
          1025 => x"bb",
          1026 => x"05",
          1027 => x"95",
          1028 => x"98",
          1029 => x"82",
          1030 => x"f4",
          1031 => x"bb",
          1032 => x"05",
          1033 => x"bb",
          1034 => x"05",
          1035 => x"31",
          1036 => x"82",
          1037 => x"ec",
          1038 => x"c1",
          1039 => x"a4",
          1040 => x"22",
          1041 => x"70",
          1042 => x"51",
          1043 => x"2e",
          1044 => x"bb",
          1045 => x"05",
          1046 => x"a4",
          1047 => x"08",
          1048 => x"bb",
          1049 => x"05",
          1050 => x"82",
          1051 => x"dc",
          1052 => x"a2",
          1053 => x"a4",
          1054 => x"08",
          1055 => x"08",
          1056 => x"84",
          1057 => x"a4",
          1058 => x"0c",
          1059 => x"bb",
          1060 => x"05",
          1061 => x"bb",
          1062 => x"05",
          1063 => x"a4",
          1064 => x"0c",
          1065 => x"08",
          1066 => x"80",
          1067 => x"82",
          1068 => x"e4",
          1069 => x"82",
          1070 => x"72",
          1071 => x"08",
          1072 => x"82",
          1073 => x"fc",
          1074 => x"82",
          1075 => x"fc",
          1076 => x"bb",
          1077 => x"05",
          1078 => x"bf",
          1079 => x"72",
          1080 => x"08",
          1081 => x"81",
          1082 => x"0b",
          1083 => x"08",
          1084 => x"a9",
          1085 => x"a4",
          1086 => x"22",
          1087 => x"07",
          1088 => x"82",
          1089 => x"e4",
          1090 => x"f8",
          1091 => x"a4",
          1092 => x"34",
          1093 => x"bb",
          1094 => x"05",
          1095 => x"a4",
          1096 => x"22",
          1097 => x"70",
          1098 => x"51",
          1099 => x"2e",
          1100 => x"bb",
          1101 => x"05",
          1102 => x"a4",
          1103 => x"08",
          1104 => x"bb",
          1105 => x"05",
          1106 => x"82",
          1107 => x"d8",
          1108 => x"a2",
          1109 => x"a4",
          1110 => x"08",
          1111 => x"08",
          1112 => x"84",
          1113 => x"a4",
          1114 => x"0c",
          1115 => x"bb",
          1116 => x"05",
          1117 => x"bb",
          1118 => x"05",
          1119 => x"a4",
          1120 => x"0c",
          1121 => x"08",
          1122 => x"70",
          1123 => x"53",
          1124 => x"a4",
          1125 => x"23",
          1126 => x"0b",
          1127 => x"08",
          1128 => x"82",
          1129 => x"f0",
          1130 => x"bb",
          1131 => x"05",
          1132 => x"a4",
          1133 => x"08",
          1134 => x"54",
          1135 => x"af",
          1136 => x"bb",
          1137 => x"72",
          1138 => x"bb",
          1139 => x"05",
          1140 => x"a4",
          1141 => x"0c",
          1142 => x"08",
          1143 => x"70",
          1144 => x"89",
          1145 => x"38",
          1146 => x"08",
          1147 => x"53",
          1148 => x"82",
          1149 => x"f8",
          1150 => x"15",
          1151 => x"51",
          1152 => x"bb",
          1153 => x"05",
          1154 => x"82",
          1155 => x"f0",
          1156 => x"72",
          1157 => x"51",
          1158 => x"bb",
          1159 => x"05",
          1160 => x"a4",
          1161 => x"08",
          1162 => x"a4",
          1163 => x"33",
          1164 => x"bb",
          1165 => x"05",
          1166 => x"82",
          1167 => x"f0",
          1168 => x"bb",
          1169 => x"05",
          1170 => x"82",
          1171 => x"fc",
          1172 => x"53",
          1173 => x"82",
          1174 => x"70",
          1175 => x"08",
          1176 => x"53",
          1177 => x"08",
          1178 => x"80",
          1179 => x"fe",
          1180 => x"bb",
          1181 => x"05",
          1182 => x"a8",
          1183 => x"54",
          1184 => x"31",
          1185 => x"82",
          1186 => x"fc",
          1187 => x"bb",
          1188 => x"05",
          1189 => x"06",
          1190 => x"80",
          1191 => x"82",
          1192 => x"ec",
          1193 => x"11",
          1194 => x"82",
          1195 => x"ec",
          1196 => x"bb",
          1197 => x"05",
          1198 => x"2a",
          1199 => x"51",
          1200 => x"80",
          1201 => x"38",
          1202 => x"08",
          1203 => x"70",
          1204 => x"bb",
          1205 => x"05",
          1206 => x"a4",
          1207 => x"08",
          1208 => x"bb",
          1209 => x"05",
          1210 => x"a4",
          1211 => x"22",
          1212 => x"90",
          1213 => x"06",
          1214 => x"bb",
          1215 => x"05",
          1216 => x"53",
          1217 => x"a4",
          1218 => x"23",
          1219 => x"bb",
          1220 => x"05",
          1221 => x"53",
          1222 => x"a4",
          1223 => x"23",
          1224 => x"08",
          1225 => x"82",
          1226 => x"ec",
          1227 => x"bb",
          1228 => x"05",
          1229 => x"2a",
          1230 => x"51",
          1231 => x"80",
          1232 => x"38",
          1233 => x"08",
          1234 => x"70",
          1235 => x"98",
          1236 => x"a4",
          1237 => x"33",
          1238 => x"53",
          1239 => x"97",
          1240 => x"a4",
          1241 => x"22",
          1242 => x"51",
          1243 => x"bb",
          1244 => x"05",
          1245 => x"82",
          1246 => x"e8",
          1247 => x"82",
          1248 => x"fc",
          1249 => x"71",
          1250 => x"72",
          1251 => x"08",
          1252 => x"82",
          1253 => x"e4",
          1254 => x"83",
          1255 => x"06",
          1256 => x"72",
          1257 => x"38",
          1258 => x"08",
          1259 => x"70",
          1260 => x"90",
          1261 => x"2c",
          1262 => x"51",
          1263 => x"53",
          1264 => x"bb",
          1265 => x"05",
          1266 => x"31",
          1267 => x"82",
          1268 => x"ec",
          1269 => x"39",
          1270 => x"08",
          1271 => x"70",
          1272 => x"90",
          1273 => x"2c",
          1274 => x"51",
          1275 => x"53",
          1276 => x"bb",
          1277 => x"05",
          1278 => x"31",
          1279 => x"82",
          1280 => x"ec",
          1281 => x"bb",
          1282 => x"05",
          1283 => x"80",
          1284 => x"72",
          1285 => x"bb",
          1286 => x"05",
          1287 => x"54",
          1288 => x"bb",
          1289 => x"05",
          1290 => x"2b",
          1291 => x"51",
          1292 => x"25",
          1293 => x"bb",
          1294 => x"05",
          1295 => x"51",
          1296 => x"d2",
          1297 => x"a4",
          1298 => x"22",
          1299 => x"70",
          1300 => x"51",
          1301 => x"2e",
          1302 => x"bb",
          1303 => x"05",
          1304 => x"51",
          1305 => x"80",
          1306 => x"bb",
          1307 => x"05",
          1308 => x"2a",
          1309 => x"51",
          1310 => x"80",
          1311 => x"82",
          1312 => x"88",
          1313 => x"ab",
          1314 => x"3f",
          1315 => x"bb",
          1316 => x"05",
          1317 => x"2a",
          1318 => x"51",
          1319 => x"80",
          1320 => x"82",
          1321 => x"88",
          1322 => x"a0",
          1323 => x"3f",
          1324 => x"08",
          1325 => x"70",
          1326 => x"81",
          1327 => x"53",
          1328 => x"b1",
          1329 => x"a4",
          1330 => x"08",
          1331 => x"95",
          1332 => x"bb",
          1333 => x"05",
          1334 => x"90",
          1335 => x"06",
          1336 => x"bb",
          1337 => x"05",
          1338 => x"bb",
          1339 => x"05",
          1340 => x"de",
          1341 => x"a4",
          1342 => x"22",
          1343 => x"70",
          1344 => x"51",
          1345 => x"2e",
          1346 => x"bb",
          1347 => x"05",
          1348 => x"54",
          1349 => x"bb",
          1350 => x"05",
          1351 => x"2b",
          1352 => x"51",
          1353 => x"25",
          1354 => x"bb",
          1355 => x"05",
          1356 => x"51",
          1357 => x"d2",
          1358 => x"a4",
          1359 => x"22",
          1360 => x"70",
          1361 => x"51",
          1362 => x"2e",
          1363 => x"bb",
          1364 => x"05",
          1365 => x"54",
          1366 => x"bb",
          1367 => x"05",
          1368 => x"2b",
          1369 => x"51",
          1370 => x"25",
          1371 => x"bb",
          1372 => x"05",
          1373 => x"51",
          1374 => x"d2",
          1375 => x"a4",
          1376 => x"22",
          1377 => x"70",
          1378 => x"51",
          1379 => x"38",
          1380 => x"08",
          1381 => x"ff",
          1382 => x"72",
          1383 => x"08",
          1384 => x"73",
          1385 => x"90",
          1386 => x"80",
          1387 => x"38",
          1388 => x"08",
          1389 => x"52",
          1390 => x"96",
          1391 => x"82",
          1392 => x"f8",
          1393 => x"72",
          1394 => x"09",
          1395 => x"38",
          1396 => x"08",
          1397 => x"52",
          1398 => x"08",
          1399 => x"51",
          1400 => x"81",
          1401 => x"bb",
          1402 => x"05",
          1403 => x"80",
          1404 => x"81",
          1405 => x"38",
          1406 => x"08",
          1407 => x"ff",
          1408 => x"72",
          1409 => x"08",
          1410 => x"72",
          1411 => x"06",
          1412 => x"ff",
          1413 => x"bb",
          1414 => x"a4",
          1415 => x"08",
          1416 => x"a4",
          1417 => x"08",
          1418 => x"82",
          1419 => x"fc",
          1420 => x"05",
          1421 => x"08",
          1422 => x"53",
          1423 => x"ff",
          1424 => x"bb",
          1425 => x"05",
          1426 => x"80",
          1427 => x"81",
          1428 => x"38",
          1429 => x"08",
          1430 => x"ff",
          1431 => x"72",
          1432 => x"08",
          1433 => x"72",
          1434 => x"06",
          1435 => x"ff",
          1436 => x"df",
          1437 => x"a4",
          1438 => x"08",
          1439 => x"a4",
          1440 => x"08",
          1441 => x"53",
          1442 => x"82",
          1443 => x"fc",
          1444 => x"05",
          1445 => x"08",
          1446 => x"ff",
          1447 => x"bb",
          1448 => x"05",
          1449 => x"a8",
          1450 => x"82",
          1451 => x"88",
          1452 => x"82",
          1453 => x"f0",
          1454 => x"05",
          1455 => x"08",
          1456 => x"82",
          1457 => x"f0",
          1458 => x"33",
          1459 => x"82",
          1460 => x"82",
          1461 => x"e4",
          1462 => x"87",
          1463 => x"06",
          1464 => x"72",
          1465 => x"c3",
          1466 => x"a4",
          1467 => x"22",
          1468 => x"54",
          1469 => x"a4",
          1470 => x"23",
          1471 => x"70",
          1472 => x"53",
          1473 => x"a3",
          1474 => x"a4",
          1475 => x"08",
          1476 => x"90",
          1477 => x"39",
          1478 => x"08",
          1479 => x"52",
          1480 => x"08",
          1481 => x"51",
          1482 => x"80",
          1483 => x"a4",
          1484 => x"23",
          1485 => x"82",
          1486 => x"f8",
          1487 => x"72",
          1488 => x"81",
          1489 => x"81",
          1490 => x"a4",
          1491 => x"23",
          1492 => x"bb",
          1493 => x"05",
          1494 => x"82",
          1495 => x"e8",
          1496 => x"0b",
          1497 => x"08",
          1498 => x"ea",
          1499 => x"bb",
          1500 => x"05",
          1501 => x"bb",
          1502 => x"05",
          1503 => x"d2",
          1504 => x"39",
          1505 => x"08",
          1506 => x"8c",
          1507 => x"82",
          1508 => x"e0",
          1509 => x"53",
          1510 => x"08",
          1511 => x"82",
          1512 => x"95",
          1513 => x"bb",
          1514 => x"82",
          1515 => x"02",
          1516 => x"0c",
          1517 => x"80",
          1518 => x"a4",
          1519 => x"34",
          1520 => x"08",
          1521 => x"53",
          1522 => x"82",
          1523 => x"88",
          1524 => x"08",
          1525 => x"33",
          1526 => x"bb",
          1527 => x"05",
          1528 => x"ff",
          1529 => x"a0",
          1530 => x"06",
          1531 => x"bb",
          1532 => x"05",
          1533 => x"81",
          1534 => x"53",
          1535 => x"bb",
          1536 => x"05",
          1537 => x"ad",
          1538 => x"06",
          1539 => x"0b",
          1540 => x"08",
          1541 => x"82",
          1542 => x"88",
          1543 => x"08",
          1544 => x"0c",
          1545 => x"53",
          1546 => x"bb",
          1547 => x"05",
          1548 => x"a4",
          1549 => x"33",
          1550 => x"2e",
          1551 => x"81",
          1552 => x"bb",
          1553 => x"05",
          1554 => x"81",
          1555 => x"70",
          1556 => x"72",
          1557 => x"a4",
          1558 => x"34",
          1559 => x"08",
          1560 => x"82",
          1561 => x"e8",
          1562 => x"bb",
          1563 => x"05",
          1564 => x"2e",
          1565 => x"bb",
          1566 => x"05",
          1567 => x"2e",
          1568 => x"cd",
          1569 => x"82",
          1570 => x"f4",
          1571 => x"bb",
          1572 => x"05",
          1573 => x"81",
          1574 => x"70",
          1575 => x"72",
          1576 => x"a4",
          1577 => x"34",
          1578 => x"82",
          1579 => x"a4",
          1580 => x"34",
          1581 => x"08",
          1582 => x"70",
          1583 => x"71",
          1584 => x"51",
          1585 => x"82",
          1586 => x"f8",
          1587 => x"fe",
          1588 => x"a4",
          1589 => x"33",
          1590 => x"26",
          1591 => x"0b",
          1592 => x"08",
          1593 => x"83",
          1594 => x"bb",
          1595 => x"05",
          1596 => x"73",
          1597 => x"82",
          1598 => x"f8",
          1599 => x"72",
          1600 => x"38",
          1601 => x"0b",
          1602 => x"08",
          1603 => x"82",
          1604 => x"0b",
          1605 => x"08",
          1606 => x"b2",
          1607 => x"a4",
          1608 => x"33",
          1609 => x"27",
          1610 => x"bb",
          1611 => x"05",
          1612 => x"b9",
          1613 => x"8d",
          1614 => x"82",
          1615 => x"ec",
          1616 => x"a5",
          1617 => x"82",
          1618 => x"f4",
          1619 => x"0b",
          1620 => x"08",
          1621 => x"82",
          1622 => x"f8",
          1623 => x"a0",
          1624 => x"cf",
          1625 => x"a4",
          1626 => x"33",
          1627 => x"73",
          1628 => x"82",
          1629 => x"f8",
          1630 => x"11",
          1631 => x"82",
          1632 => x"f8",
          1633 => x"bb",
          1634 => x"05",
          1635 => x"51",
          1636 => x"bb",
          1637 => x"05",
          1638 => x"a4",
          1639 => x"33",
          1640 => x"27",
          1641 => x"bb",
          1642 => x"05",
          1643 => x"51",
          1644 => x"bb",
          1645 => x"05",
          1646 => x"a4",
          1647 => x"33",
          1648 => x"26",
          1649 => x"0b",
          1650 => x"08",
          1651 => x"81",
          1652 => x"bb",
          1653 => x"05",
          1654 => x"a4",
          1655 => x"33",
          1656 => x"74",
          1657 => x"80",
          1658 => x"a4",
          1659 => x"0c",
          1660 => x"82",
          1661 => x"f4",
          1662 => x"82",
          1663 => x"fc",
          1664 => x"82",
          1665 => x"f8",
          1666 => x"12",
          1667 => x"08",
          1668 => x"82",
          1669 => x"88",
          1670 => x"08",
          1671 => x"0c",
          1672 => x"51",
          1673 => x"72",
          1674 => x"a4",
          1675 => x"34",
          1676 => x"82",
          1677 => x"f0",
          1678 => x"72",
          1679 => x"38",
          1680 => x"08",
          1681 => x"30",
          1682 => x"08",
          1683 => x"82",
          1684 => x"8c",
          1685 => x"bb",
          1686 => x"05",
          1687 => x"53",
          1688 => x"bb",
          1689 => x"05",
          1690 => x"a4",
          1691 => x"08",
          1692 => x"0c",
          1693 => x"82",
          1694 => x"04",
          1695 => x"08",
          1696 => x"a4",
          1697 => x"0d",
          1698 => x"08",
          1699 => x"a4",
          1700 => x"08",
          1701 => x"a4",
          1702 => x"08",
          1703 => x"3f",
          1704 => x"08",
          1705 => x"98",
          1706 => x"3d",
          1707 => x"a4",
          1708 => x"bb",
          1709 => x"82",
          1710 => x"f7",
          1711 => x"0b",
          1712 => x"08",
          1713 => x"82",
          1714 => x"8c",
          1715 => x"80",
          1716 => x"bb",
          1717 => x"05",
          1718 => x"51",
          1719 => x"53",
          1720 => x"a4",
          1721 => x"34",
          1722 => x"06",
          1723 => x"2e",
          1724 => x"91",
          1725 => x"a4",
          1726 => x"08",
          1727 => x"05",
          1728 => x"ce",
          1729 => x"a4",
          1730 => x"33",
          1731 => x"2e",
          1732 => x"a4",
          1733 => x"82",
          1734 => x"f0",
          1735 => x"bb",
          1736 => x"05",
          1737 => x"81",
          1738 => x"70",
          1739 => x"72",
          1740 => x"a4",
          1741 => x"34",
          1742 => x"08",
          1743 => x"53",
          1744 => x"09",
          1745 => x"dc",
          1746 => x"a4",
          1747 => x"08",
          1748 => x"05",
          1749 => x"08",
          1750 => x"33",
          1751 => x"08",
          1752 => x"82",
          1753 => x"f8",
          1754 => x"bb",
          1755 => x"05",
          1756 => x"a4",
          1757 => x"08",
          1758 => x"b6",
          1759 => x"a4",
          1760 => x"08",
          1761 => x"84",
          1762 => x"39",
          1763 => x"bb",
          1764 => x"05",
          1765 => x"a4",
          1766 => x"08",
          1767 => x"05",
          1768 => x"08",
          1769 => x"33",
          1770 => x"08",
          1771 => x"81",
          1772 => x"0b",
          1773 => x"08",
          1774 => x"82",
          1775 => x"88",
          1776 => x"08",
          1777 => x"0c",
          1778 => x"53",
          1779 => x"bb",
          1780 => x"05",
          1781 => x"39",
          1782 => x"08",
          1783 => x"53",
          1784 => x"8d",
          1785 => x"82",
          1786 => x"ec",
          1787 => x"80",
          1788 => x"a4",
          1789 => x"33",
          1790 => x"27",
          1791 => x"bb",
          1792 => x"05",
          1793 => x"b9",
          1794 => x"8d",
          1795 => x"82",
          1796 => x"ec",
          1797 => x"d8",
          1798 => x"82",
          1799 => x"f4",
          1800 => x"39",
          1801 => x"08",
          1802 => x"53",
          1803 => x"90",
          1804 => x"a4",
          1805 => x"33",
          1806 => x"26",
          1807 => x"39",
          1808 => x"bb",
          1809 => x"05",
          1810 => x"39",
          1811 => x"bb",
          1812 => x"05",
          1813 => x"82",
          1814 => x"fc",
          1815 => x"bb",
          1816 => x"05",
          1817 => x"73",
          1818 => x"38",
          1819 => x"08",
          1820 => x"53",
          1821 => x"27",
          1822 => x"bb",
          1823 => x"05",
          1824 => x"51",
          1825 => x"bb",
          1826 => x"05",
          1827 => x"a4",
          1828 => x"33",
          1829 => x"53",
          1830 => x"a4",
          1831 => x"34",
          1832 => x"08",
          1833 => x"53",
          1834 => x"ad",
          1835 => x"a4",
          1836 => x"33",
          1837 => x"53",
          1838 => x"a4",
          1839 => x"34",
          1840 => x"08",
          1841 => x"53",
          1842 => x"8d",
          1843 => x"82",
          1844 => x"ec",
          1845 => x"98",
          1846 => x"a4",
          1847 => x"33",
          1848 => x"08",
          1849 => x"54",
          1850 => x"26",
          1851 => x"0b",
          1852 => x"08",
          1853 => x"80",
          1854 => x"bb",
          1855 => x"05",
          1856 => x"bb",
          1857 => x"05",
          1858 => x"bb",
          1859 => x"05",
          1860 => x"82",
          1861 => x"fc",
          1862 => x"bb",
          1863 => x"05",
          1864 => x"81",
          1865 => x"70",
          1866 => x"52",
          1867 => x"33",
          1868 => x"08",
          1869 => x"fe",
          1870 => x"bb",
          1871 => x"05",
          1872 => x"80",
          1873 => x"82",
          1874 => x"fc",
          1875 => x"82",
          1876 => x"fc",
          1877 => x"bb",
          1878 => x"05",
          1879 => x"a4",
          1880 => x"08",
          1881 => x"81",
          1882 => x"a4",
          1883 => x"0c",
          1884 => x"08",
          1885 => x"82",
          1886 => x"8b",
          1887 => x"bb",
          1888 => x"82",
          1889 => x"02",
          1890 => x"0c",
          1891 => x"80",
          1892 => x"a4",
          1893 => x"0c",
          1894 => x"08",
          1895 => x"70",
          1896 => x"81",
          1897 => x"06",
          1898 => x"51",
          1899 => x"2e",
          1900 => x"0b",
          1901 => x"08",
          1902 => x"81",
          1903 => x"bb",
          1904 => x"05",
          1905 => x"33",
          1906 => x"08",
          1907 => x"81",
          1908 => x"a4",
          1909 => x"0c",
          1910 => x"bb",
          1911 => x"05",
          1912 => x"ff",
          1913 => x"80",
          1914 => x"82",
          1915 => x"82",
          1916 => x"53",
          1917 => x"08",
          1918 => x"52",
          1919 => x"51",
          1920 => x"82",
          1921 => x"53",
          1922 => x"ff",
          1923 => x"0b",
          1924 => x"08",
          1925 => x"ff",
          1926 => x"d2",
          1927 => x"d2",
          1928 => x"53",
          1929 => x"13",
          1930 => x"2d",
          1931 => x"08",
          1932 => x"2e",
          1933 => x"0b",
          1934 => x"08",
          1935 => x"82",
          1936 => x"f8",
          1937 => x"82",
          1938 => x"f4",
          1939 => x"82",
          1940 => x"f4",
          1941 => x"bb",
          1942 => x"3d",
          1943 => x"a4",
          1944 => x"bb",
          1945 => x"82",
          1946 => x"fb",
          1947 => x"0b",
          1948 => x"08",
          1949 => x"82",
          1950 => x"8c",
          1951 => x"11",
          1952 => x"2a",
          1953 => x"70",
          1954 => x"51",
          1955 => x"72",
          1956 => x"38",
          1957 => x"bb",
          1958 => x"05",
          1959 => x"39",
          1960 => x"08",
          1961 => x"53",
          1962 => x"bb",
          1963 => x"05",
          1964 => x"82",
          1965 => x"88",
          1966 => x"72",
          1967 => x"08",
          1968 => x"72",
          1969 => x"53",
          1970 => x"b6",
          1971 => x"a4",
          1972 => x"08",
          1973 => x"08",
          1974 => x"53",
          1975 => x"08",
          1976 => x"52",
          1977 => x"51",
          1978 => x"82",
          1979 => x"53",
          1980 => x"ff",
          1981 => x"0b",
          1982 => x"08",
          1983 => x"ff",
          1984 => x"bb",
          1985 => x"05",
          1986 => x"bb",
          1987 => x"05",
          1988 => x"bb",
          1989 => x"05",
          1990 => x"98",
          1991 => x"0d",
          1992 => x"0c",
          1993 => x"a4",
          1994 => x"bb",
          1995 => x"3d",
          1996 => x"ec",
          1997 => x"bb",
          1998 => x"05",
          1999 => x"3f",
          2000 => x"08",
          2001 => x"98",
          2002 => x"3d",
          2003 => x"a4",
          2004 => x"bb",
          2005 => x"82",
          2006 => x"fb",
          2007 => x"bb",
          2008 => x"05",
          2009 => x"33",
          2010 => x"70",
          2011 => x"81",
          2012 => x"51",
          2013 => x"80",
          2014 => x"ff",
          2015 => x"a4",
          2016 => x"0c",
          2017 => x"82",
          2018 => x"8c",
          2019 => x"11",
          2020 => x"2a",
          2021 => x"51",
          2022 => x"72",
          2023 => x"db",
          2024 => x"a4",
          2025 => x"08",
          2026 => x"08",
          2027 => x"54",
          2028 => x"08",
          2029 => x"25",
          2030 => x"bb",
          2031 => x"05",
          2032 => x"70",
          2033 => x"08",
          2034 => x"52",
          2035 => x"72",
          2036 => x"08",
          2037 => x"0c",
          2038 => x"08",
          2039 => x"8c",
          2040 => x"05",
          2041 => x"82",
          2042 => x"88",
          2043 => x"82",
          2044 => x"fc",
          2045 => x"53",
          2046 => x"82",
          2047 => x"8c",
          2048 => x"bb",
          2049 => x"05",
          2050 => x"bb",
          2051 => x"05",
          2052 => x"ff",
          2053 => x"12",
          2054 => x"54",
          2055 => x"bb",
          2056 => x"72",
          2057 => x"bb",
          2058 => x"05",
          2059 => x"08",
          2060 => x"12",
          2061 => x"a4",
          2062 => x"08",
          2063 => x"a4",
          2064 => x"0c",
          2065 => x"39",
          2066 => x"bb",
          2067 => x"05",
          2068 => x"a4",
          2069 => x"08",
          2070 => x"0c",
          2071 => x"82",
          2072 => x"04",
          2073 => x"08",
          2074 => x"a4",
          2075 => x"0d",
          2076 => x"08",
          2077 => x"85",
          2078 => x"81",
          2079 => x"06",
          2080 => x"52",
          2081 => x"8d",
          2082 => x"82",
          2083 => x"f8",
          2084 => x"94",
          2085 => x"a4",
          2086 => x"08",
          2087 => x"70",
          2088 => x"81",
          2089 => x"51",
          2090 => x"2e",
          2091 => x"82",
          2092 => x"88",
          2093 => x"bb",
          2094 => x"05",
          2095 => x"85",
          2096 => x"ff",
          2097 => x"52",
          2098 => x"34",
          2099 => x"08",
          2100 => x"8c",
          2101 => x"05",
          2102 => x"82",
          2103 => x"88",
          2104 => x"11",
          2105 => x"bb",
          2106 => x"05",
          2107 => x"52",
          2108 => x"82",
          2109 => x"88",
          2110 => x"11",
          2111 => x"2a",
          2112 => x"51",
          2113 => x"71",
          2114 => x"d7",
          2115 => x"a4",
          2116 => x"08",
          2117 => x"33",
          2118 => x"08",
          2119 => x"51",
          2120 => x"a4",
          2121 => x"08",
          2122 => x"bb",
          2123 => x"05",
          2124 => x"a4",
          2125 => x"08",
          2126 => x"12",
          2127 => x"07",
          2128 => x"85",
          2129 => x"0b",
          2130 => x"08",
          2131 => x"81",
          2132 => x"bb",
          2133 => x"05",
          2134 => x"81",
          2135 => x"52",
          2136 => x"82",
          2137 => x"88",
          2138 => x"bb",
          2139 => x"05",
          2140 => x"11",
          2141 => x"71",
          2142 => x"98",
          2143 => x"bb",
          2144 => x"05",
          2145 => x"bb",
          2146 => x"05",
          2147 => x"80",
          2148 => x"bb",
          2149 => x"05",
          2150 => x"a4",
          2151 => x"0c",
          2152 => x"08",
          2153 => x"85",
          2154 => x"bb",
          2155 => x"05",
          2156 => x"bb",
          2157 => x"05",
          2158 => x"09",
          2159 => x"38",
          2160 => x"08",
          2161 => x"90",
          2162 => x"82",
          2163 => x"ec",
          2164 => x"39",
          2165 => x"08",
          2166 => x"a0",
          2167 => x"82",
          2168 => x"ec",
          2169 => x"bb",
          2170 => x"05",
          2171 => x"bb",
          2172 => x"05",
          2173 => x"34",
          2174 => x"bb",
          2175 => x"05",
          2176 => x"82",
          2177 => x"88",
          2178 => x"11",
          2179 => x"8c",
          2180 => x"bb",
          2181 => x"05",
          2182 => x"ff",
          2183 => x"bb",
          2184 => x"05",
          2185 => x"52",
          2186 => x"08",
          2187 => x"82",
          2188 => x"89",
          2189 => x"bb",
          2190 => x"82",
          2191 => x"02",
          2192 => x"0c",
          2193 => x"82",
          2194 => x"88",
          2195 => x"bb",
          2196 => x"05",
          2197 => x"a4",
          2198 => x"08",
          2199 => x"08",
          2200 => x"82",
          2201 => x"90",
          2202 => x"2e",
          2203 => x"82",
          2204 => x"f8",
          2205 => x"bb",
          2206 => x"05",
          2207 => x"ac",
          2208 => x"a4",
          2209 => x"08",
          2210 => x"08",
          2211 => x"05",
          2212 => x"a4",
          2213 => x"08",
          2214 => x"90",
          2215 => x"a4",
          2216 => x"08",
          2217 => x"08",
          2218 => x"05",
          2219 => x"08",
          2220 => x"82",
          2221 => x"f8",
          2222 => x"bb",
          2223 => x"05",
          2224 => x"bb",
          2225 => x"05",
          2226 => x"a4",
          2227 => x"08",
          2228 => x"bb",
          2229 => x"05",
          2230 => x"a4",
          2231 => x"08",
          2232 => x"bb",
          2233 => x"05",
          2234 => x"a4",
          2235 => x"08",
          2236 => x"9c",
          2237 => x"a4",
          2238 => x"08",
          2239 => x"bb",
          2240 => x"05",
          2241 => x"a4",
          2242 => x"08",
          2243 => x"bb",
          2244 => x"05",
          2245 => x"a4",
          2246 => x"08",
          2247 => x"08",
          2248 => x"53",
          2249 => x"71",
          2250 => x"39",
          2251 => x"08",
          2252 => x"81",
          2253 => x"a4",
          2254 => x"0c",
          2255 => x"08",
          2256 => x"ff",
          2257 => x"a4",
          2258 => x"0c",
          2259 => x"08",
          2260 => x"80",
          2261 => x"82",
          2262 => x"f8",
          2263 => x"70",
          2264 => x"a4",
          2265 => x"08",
          2266 => x"bb",
          2267 => x"05",
          2268 => x"a4",
          2269 => x"08",
          2270 => x"71",
          2271 => x"a4",
          2272 => x"08",
          2273 => x"bb",
          2274 => x"05",
          2275 => x"39",
          2276 => x"08",
          2277 => x"70",
          2278 => x"0c",
          2279 => x"0d",
          2280 => x"0c",
          2281 => x"a4",
          2282 => x"bb",
          2283 => x"3d",
          2284 => x"a4",
          2285 => x"08",
          2286 => x"08",
          2287 => x"82",
          2288 => x"fc",
          2289 => x"71",
          2290 => x"a4",
          2291 => x"08",
          2292 => x"bb",
          2293 => x"05",
          2294 => x"ff",
          2295 => x"70",
          2296 => x"38",
          2297 => x"bb",
          2298 => x"05",
          2299 => x"82",
          2300 => x"fc",
          2301 => x"bb",
          2302 => x"05",
          2303 => x"a4",
          2304 => x"08",
          2305 => x"bb",
          2306 => x"84",
          2307 => x"bb",
          2308 => x"82",
          2309 => x"02",
          2310 => x"0c",
          2311 => x"82",
          2312 => x"88",
          2313 => x"bb",
          2314 => x"05",
          2315 => x"a4",
          2316 => x"08",
          2317 => x"82",
          2318 => x"8c",
          2319 => x"05",
          2320 => x"08",
          2321 => x"82",
          2322 => x"fc",
          2323 => x"51",
          2324 => x"82",
          2325 => x"fc",
          2326 => x"05",
          2327 => x"08",
          2328 => x"70",
          2329 => x"51",
          2330 => x"84",
          2331 => x"39",
          2332 => x"08",
          2333 => x"70",
          2334 => x"0c",
          2335 => x"0d",
          2336 => x"0c",
          2337 => x"a4",
          2338 => x"bb",
          2339 => x"3d",
          2340 => x"a4",
          2341 => x"08",
          2342 => x"08",
          2343 => x"82",
          2344 => x"8c",
          2345 => x"bb",
          2346 => x"05",
          2347 => x"a4",
          2348 => x"08",
          2349 => x"e5",
          2350 => x"a4",
          2351 => x"08",
          2352 => x"bb",
          2353 => x"05",
          2354 => x"a4",
          2355 => x"08",
          2356 => x"bb",
          2357 => x"05",
          2358 => x"a4",
          2359 => x"08",
          2360 => x"38",
          2361 => x"08",
          2362 => x"51",
          2363 => x"bb",
          2364 => x"05",
          2365 => x"82",
          2366 => x"f8",
          2367 => x"bb",
          2368 => x"05",
          2369 => x"71",
          2370 => x"bb",
          2371 => x"05",
          2372 => x"82",
          2373 => x"fc",
          2374 => x"ad",
          2375 => x"a4",
          2376 => x"08",
          2377 => x"98",
          2378 => x"3d",
          2379 => x"a4",
          2380 => x"bb",
          2381 => x"82",
          2382 => x"fd",
          2383 => x"bb",
          2384 => x"05",
          2385 => x"81",
          2386 => x"bb",
          2387 => x"05",
          2388 => x"33",
          2389 => x"08",
          2390 => x"81",
          2391 => x"a4",
          2392 => x"0c",
          2393 => x"08",
          2394 => x"70",
          2395 => x"ff",
          2396 => x"54",
          2397 => x"2e",
          2398 => x"ce",
          2399 => x"a4",
          2400 => x"08",
          2401 => x"82",
          2402 => x"88",
          2403 => x"05",
          2404 => x"08",
          2405 => x"70",
          2406 => x"51",
          2407 => x"38",
          2408 => x"bb",
          2409 => x"05",
          2410 => x"39",
          2411 => x"08",
          2412 => x"ff",
          2413 => x"a4",
          2414 => x"0c",
          2415 => x"08",
          2416 => x"80",
          2417 => x"ff",
          2418 => x"bb",
          2419 => x"05",
          2420 => x"80",
          2421 => x"bb",
          2422 => x"05",
          2423 => x"52",
          2424 => x"38",
          2425 => x"bb",
          2426 => x"05",
          2427 => x"39",
          2428 => x"08",
          2429 => x"ff",
          2430 => x"a4",
          2431 => x"0c",
          2432 => x"08",
          2433 => x"70",
          2434 => x"70",
          2435 => x"0b",
          2436 => x"08",
          2437 => x"ae",
          2438 => x"a4",
          2439 => x"08",
          2440 => x"bb",
          2441 => x"05",
          2442 => x"72",
          2443 => x"82",
          2444 => x"fc",
          2445 => x"55",
          2446 => x"8a",
          2447 => x"82",
          2448 => x"fc",
          2449 => x"bb",
          2450 => x"05",
          2451 => x"98",
          2452 => x"0d",
          2453 => x"0c",
          2454 => x"a4",
          2455 => x"bb",
          2456 => x"3d",
          2457 => x"a4",
          2458 => x"08",
          2459 => x"08",
          2460 => x"82",
          2461 => x"8c",
          2462 => x"38",
          2463 => x"bb",
          2464 => x"05",
          2465 => x"39",
          2466 => x"08",
          2467 => x"52",
          2468 => x"bb",
          2469 => x"05",
          2470 => x"82",
          2471 => x"f8",
          2472 => x"81",
          2473 => x"51",
          2474 => x"9f",
          2475 => x"a4",
          2476 => x"08",
          2477 => x"bb",
          2478 => x"05",
          2479 => x"a4",
          2480 => x"08",
          2481 => x"38",
          2482 => x"82",
          2483 => x"f8",
          2484 => x"05",
          2485 => x"08",
          2486 => x"82",
          2487 => x"f8",
          2488 => x"bb",
          2489 => x"05",
          2490 => x"82",
          2491 => x"fc",
          2492 => x"82",
          2493 => x"fc",
          2494 => x"bb",
          2495 => x"3d",
          2496 => x"a4",
          2497 => x"bb",
          2498 => x"82",
          2499 => x"fe",
          2500 => x"bb",
          2501 => x"05",
          2502 => x"a4",
          2503 => x"0c",
          2504 => x"08",
          2505 => x"80",
          2506 => x"38",
          2507 => x"08",
          2508 => x"81",
          2509 => x"a4",
          2510 => x"0c",
          2511 => x"08",
          2512 => x"ff",
          2513 => x"a4",
          2514 => x"0c",
          2515 => x"08",
          2516 => x"80",
          2517 => x"82",
          2518 => x"8c",
          2519 => x"70",
          2520 => x"08",
          2521 => x"52",
          2522 => x"34",
          2523 => x"08",
          2524 => x"81",
          2525 => x"a4",
          2526 => x"0c",
          2527 => x"82",
          2528 => x"88",
          2529 => x"82",
          2530 => x"51",
          2531 => x"82",
          2532 => x"04",
          2533 => x"08",
          2534 => x"a4",
          2535 => x"0d",
          2536 => x"bb",
          2537 => x"05",
          2538 => x"a4",
          2539 => x"08",
          2540 => x"38",
          2541 => x"08",
          2542 => x"30",
          2543 => x"08",
          2544 => x"80",
          2545 => x"a4",
          2546 => x"0c",
          2547 => x"08",
          2548 => x"8a",
          2549 => x"82",
          2550 => x"f4",
          2551 => x"bb",
          2552 => x"05",
          2553 => x"a4",
          2554 => x"0c",
          2555 => x"08",
          2556 => x"80",
          2557 => x"82",
          2558 => x"8c",
          2559 => x"82",
          2560 => x"8c",
          2561 => x"0b",
          2562 => x"08",
          2563 => x"82",
          2564 => x"fc",
          2565 => x"38",
          2566 => x"bb",
          2567 => x"05",
          2568 => x"a4",
          2569 => x"08",
          2570 => x"08",
          2571 => x"80",
          2572 => x"a4",
          2573 => x"08",
          2574 => x"a4",
          2575 => x"08",
          2576 => x"3f",
          2577 => x"08",
          2578 => x"a4",
          2579 => x"0c",
          2580 => x"a4",
          2581 => x"08",
          2582 => x"38",
          2583 => x"08",
          2584 => x"30",
          2585 => x"08",
          2586 => x"82",
          2587 => x"f8",
          2588 => x"82",
          2589 => x"54",
          2590 => x"82",
          2591 => x"04",
          2592 => x"08",
          2593 => x"a4",
          2594 => x"0d",
          2595 => x"bb",
          2596 => x"05",
          2597 => x"a4",
          2598 => x"08",
          2599 => x"38",
          2600 => x"08",
          2601 => x"30",
          2602 => x"08",
          2603 => x"81",
          2604 => x"a4",
          2605 => x"0c",
          2606 => x"08",
          2607 => x"80",
          2608 => x"82",
          2609 => x"8c",
          2610 => x"82",
          2611 => x"8c",
          2612 => x"53",
          2613 => x"08",
          2614 => x"52",
          2615 => x"08",
          2616 => x"51",
          2617 => x"82",
          2618 => x"70",
          2619 => x"08",
          2620 => x"54",
          2621 => x"08",
          2622 => x"80",
          2623 => x"82",
          2624 => x"f8",
          2625 => x"82",
          2626 => x"f8",
          2627 => x"bb",
          2628 => x"05",
          2629 => x"bb",
          2630 => x"87",
          2631 => x"bb",
          2632 => x"82",
          2633 => x"02",
          2634 => x"0c",
          2635 => x"80",
          2636 => x"a4",
          2637 => x"08",
          2638 => x"a4",
          2639 => x"08",
          2640 => x"3f",
          2641 => x"08",
          2642 => x"98",
          2643 => x"3d",
          2644 => x"a4",
          2645 => x"bb",
          2646 => x"82",
          2647 => x"fd",
          2648 => x"53",
          2649 => x"08",
          2650 => x"52",
          2651 => x"08",
          2652 => x"51",
          2653 => x"bb",
          2654 => x"82",
          2655 => x"54",
          2656 => x"82",
          2657 => x"04",
          2658 => x"08",
          2659 => x"a4",
          2660 => x"0d",
          2661 => x"bb",
          2662 => x"05",
          2663 => x"82",
          2664 => x"f8",
          2665 => x"bb",
          2666 => x"05",
          2667 => x"a4",
          2668 => x"08",
          2669 => x"82",
          2670 => x"fc",
          2671 => x"2e",
          2672 => x"0b",
          2673 => x"08",
          2674 => x"24",
          2675 => x"bb",
          2676 => x"05",
          2677 => x"bb",
          2678 => x"05",
          2679 => x"a4",
          2680 => x"08",
          2681 => x"a4",
          2682 => x"0c",
          2683 => x"82",
          2684 => x"fc",
          2685 => x"2e",
          2686 => x"82",
          2687 => x"8c",
          2688 => x"bb",
          2689 => x"05",
          2690 => x"38",
          2691 => x"08",
          2692 => x"82",
          2693 => x"8c",
          2694 => x"82",
          2695 => x"88",
          2696 => x"bb",
          2697 => x"05",
          2698 => x"a4",
          2699 => x"08",
          2700 => x"a4",
          2701 => x"0c",
          2702 => x"08",
          2703 => x"81",
          2704 => x"a4",
          2705 => x"0c",
          2706 => x"08",
          2707 => x"81",
          2708 => x"a4",
          2709 => x"0c",
          2710 => x"82",
          2711 => x"90",
          2712 => x"2e",
          2713 => x"bb",
          2714 => x"05",
          2715 => x"bb",
          2716 => x"05",
          2717 => x"39",
          2718 => x"08",
          2719 => x"70",
          2720 => x"08",
          2721 => x"51",
          2722 => x"08",
          2723 => x"82",
          2724 => x"85",
          2725 => x"bb",
          2726 => x"f9",
          2727 => x"70",
          2728 => x"56",
          2729 => x"2e",
          2730 => x"95",
          2731 => x"51",
          2732 => x"82",
          2733 => x"15",
          2734 => x"16",
          2735 => x"cd",
          2736 => x"54",
          2737 => x"09",
          2738 => x"38",
          2739 => x"f1",
          2740 => x"76",
          2741 => x"b6",
          2742 => x"08",
          2743 => x"c5",
          2744 => x"98",
          2745 => x"52",
          2746 => x"f4",
          2747 => x"bb",
          2748 => x"38",
          2749 => x"54",
          2750 => x"ff",
          2751 => x"17",
          2752 => x"06",
          2753 => x"77",
          2754 => x"ff",
          2755 => x"bb",
          2756 => x"3d",
          2757 => x"3d",
          2758 => x"71",
          2759 => x"8e",
          2760 => x"29",
          2761 => x"05",
          2762 => x"04",
          2763 => x"51",
          2764 => x"82",
          2765 => x"80",
          2766 => x"9f",
          2767 => x"f2",
          2768 => x"b0",
          2769 => x"39",
          2770 => x"51",
          2771 => x"82",
          2772 => x"80",
          2773 => x"9f",
          2774 => x"d6",
          2775 => x"f4",
          2776 => x"39",
          2777 => x"51",
          2778 => x"82",
          2779 => x"80",
          2780 => x"a0",
          2781 => x"39",
          2782 => x"51",
          2783 => x"a0",
          2784 => x"39",
          2785 => x"51",
          2786 => x"a1",
          2787 => x"39",
          2788 => x"51",
          2789 => x"a1",
          2790 => x"39",
          2791 => x"51",
          2792 => x"a2",
          2793 => x"39",
          2794 => x"51",
          2795 => x"a2",
          2796 => x"cf",
          2797 => x"0d",
          2798 => x"0d",
          2799 => x"56",
          2800 => x"26",
          2801 => x"52",
          2802 => x"29",
          2803 => x"87",
          2804 => x"51",
          2805 => x"82",
          2806 => x"52",
          2807 => x"c3",
          2808 => x"98",
          2809 => x"53",
          2810 => x"a2",
          2811 => x"bb",
          2812 => x"3d",
          2813 => x"3d",
          2814 => x"84",
          2815 => x"05",
          2816 => x"80",
          2817 => x"70",
          2818 => x"25",
          2819 => x"59",
          2820 => x"87",
          2821 => x"38",
          2822 => x"76",
          2823 => x"ff",
          2824 => x"93",
          2825 => x"82",
          2826 => x"76",
          2827 => x"70",
          2828 => x"83",
          2829 => x"bb",
          2830 => x"82",
          2831 => x"b9",
          2832 => x"98",
          2833 => x"98",
          2834 => x"bb",
          2835 => x"96",
          2836 => x"54",
          2837 => x"77",
          2838 => x"81",
          2839 => x"82",
          2840 => x"57",
          2841 => x"08",
          2842 => x"55",
          2843 => x"89",
          2844 => x"75",
          2845 => x"d7",
          2846 => x"d8",
          2847 => x"8f",
          2848 => x"30",
          2849 => x"80",
          2850 => x"70",
          2851 => x"06",
          2852 => x"56",
          2853 => x"90",
          2854 => x"e8",
          2855 => x"98",
          2856 => x"78",
          2857 => x"3f",
          2858 => x"82",
          2859 => x"96",
          2860 => x"f8",
          2861 => x"02",
          2862 => x"05",
          2863 => x"ff",
          2864 => x"7b",
          2865 => x"fe",
          2866 => x"bb",
          2867 => x"38",
          2868 => x"88",
          2869 => x"2e",
          2870 => x"39",
          2871 => x"55",
          2872 => x"bb",
          2873 => x"52",
          2874 => x"2d",
          2875 => x"08",
          2876 => x"78",
          2877 => x"bb",
          2878 => x"3d",
          2879 => x"3d",
          2880 => x"63",
          2881 => x"80",
          2882 => x"73",
          2883 => x"41",
          2884 => x"5e",
          2885 => x"52",
          2886 => x"51",
          2887 => x"3f",
          2888 => x"51",
          2889 => x"80",
          2890 => x"27",
          2891 => x"7b",
          2892 => x"38",
          2893 => x"a6",
          2894 => x"39",
          2895 => x"72",
          2896 => x"38",
          2897 => x"82",
          2898 => x"ff",
          2899 => x"88",
          2900 => x"88",
          2901 => x"3f",
          2902 => x"80",
          2903 => x"18",
          2904 => x"27",
          2905 => x"08",
          2906 => x"f0",
          2907 => x"e6",
          2908 => x"82",
          2909 => x"e0",
          2910 => x"15",
          2911 => x"74",
          2912 => x"7a",
          2913 => x"72",
          2914 => x"a3",
          2915 => x"b8",
          2916 => x"39",
          2917 => x"51",
          2918 => x"81",
          2919 => x"d2",
          2920 => x"a0",
          2921 => x"3f",
          2922 => x"82",
          2923 => x"df",
          2924 => x"55",
          2925 => x"80",
          2926 => x"18",
          2927 => x"53",
          2928 => x"7a",
          2929 => x"81",
          2930 => x"9f",
          2931 => x"38",
          2932 => x"73",
          2933 => x"ff",
          2934 => x"72",
          2935 => x"38",
          2936 => x"26",
          2937 => x"d2",
          2938 => x"73",
          2939 => x"82",
          2940 => x"52",
          2941 => x"da",
          2942 => x"55",
          2943 => x"82",
          2944 => x"de",
          2945 => x"18",
          2946 => x"58",
          2947 => x"82",
          2948 => x"98",
          2949 => x"2c",
          2950 => x"a0",
          2951 => x"06",
          2952 => x"d9",
          2953 => x"98",
          2954 => x"70",
          2955 => x"a0",
          2956 => x"72",
          2957 => x"30",
          2958 => x"73",
          2959 => x"51",
          2960 => x"57",
          2961 => x"73",
          2962 => x"76",
          2963 => x"81",
          2964 => x"80",
          2965 => x"7c",
          2966 => x"78",
          2967 => x"38",
          2968 => x"82",
          2969 => x"8f",
          2970 => x"fc",
          2971 => x"9b",
          2972 => x"a3",
          2973 => x"a3",
          2974 => x"ff",
          2975 => x"82",
          2976 => x"51",
          2977 => x"82",
          2978 => x"82",
          2979 => x"82",
          2980 => x"52",
          2981 => x"51",
          2982 => x"3f",
          2983 => x"84",
          2984 => x"3f",
          2985 => x"04",
          2986 => x"87",
          2987 => x"08",
          2988 => x"3f",
          2989 => x"b2",
          2990 => x"e8",
          2991 => x"3f",
          2992 => x"a6",
          2993 => x"2a",
          2994 => x"51",
          2995 => x"2e",
          2996 => x"51",
          2997 => x"82",
          2998 => x"9d",
          2999 => x"51",
          3000 => x"72",
          3001 => x"81",
          3002 => x"71",
          3003 => x"38",
          3004 => x"f6",
          3005 => x"98",
          3006 => x"3f",
          3007 => x"ea",
          3008 => x"2a",
          3009 => x"51",
          3010 => x"2e",
          3011 => x"51",
          3012 => x"82",
          3013 => x"9c",
          3014 => x"51",
          3015 => x"72",
          3016 => x"81",
          3017 => x"71",
          3018 => x"38",
          3019 => x"ba",
          3020 => x"bc",
          3021 => x"3f",
          3022 => x"ae",
          3023 => x"2a",
          3024 => x"51",
          3025 => x"2e",
          3026 => x"51",
          3027 => x"82",
          3028 => x"9c",
          3029 => x"51",
          3030 => x"72",
          3031 => x"81",
          3032 => x"71",
          3033 => x"38",
          3034 => x"fe",
          3035 => x"e4",
          3036 => x"3f",
          3037 => x"f2",
          3038 => x"2a",
          3039 => x"51",
          3040 => x"2e",
          3041 => x"51",
          3042 => x"82",
          3043 => x"9b",
          3044 => x"51",
          3045 => x"72",
          3046 => x"81",
          3047 => x"71",
          3048 => x"38",
          3049 => x"c2",
          3050 => x"8c",
          3051 => x"3f",
          3052 => x"b6",
          3053 => x"3f",
          3054 => x"04",
          3055 => x"77",
          3056 => x"a3",
          3057 => x"55",
          3058 => x"52",
          3059 => x"b6",
          3060 => x"82",
          3061 => x"54",
          3062 => x"81",
          3063 => x"cc",
          3064 => x"98",
          3065 => x"9c",
          3066 => x"98",
          3067 => x"82",
          3068 => x"07",
          3069 => x"71",
          3070 => x"54",
          3071 => x"82",
          3072 => x"0b",
          3073 => x"94",
          3074 => x"81",
          3075 => x"06",
          3076 => x"d2",
          3077 => x"52",
          3078 => x"b6",
          3079 => x"bb",
          3080 => x"2e",
          3081 => x"bb",
          3082 => x"da",
          3083 => x"39",
          3084 => x"51",
          3085 => x"3f",
          3086 => x"0b",
          3087 => x"34",
          3088 => x"b6",
          3089 => x"73",
          3090 => x"81",
          3091 => x"82",
          3092 => x"74",
          3093 => x"ae",
          3094 => x"0b",
          3095 => x"0c",
          3096 => x"04",
          3097 => x"80",
          3098 => x"d2",
          3099 => x"5e",
          3100 => x"51",
          3101 => x"3f",
          3102 => x"08",
          3103 => x"5a",
          3104 => x"09",
          3105 => x"38",
          3106 => x"83",
          3107 => x"e8",
          3108 => x"e7",
          3109 => x"53",
          3110 => x"bc",
          3111 => x"fa",
          3112 => x"bb",
          3113 => x"2e",
          3114 => x"a5",
          3115 => x"c8",
          3116 => x"40",
          3117 => x"a4",
          3118 => x"3f",
          3119 => x"47",
          3120 => x"52",
          3121 => x"f4",
          3122 => x"ff",
          3123 => x"f3",
          3124 => x"bb",
          3125 => x"2b",
          3126 => x"51",
          3127 => x"c1",
          3128 => x"38",
          3129 => x"24",
          3130 => x"79",
          3131 => x"b9",
          3132 => x"24",
          3133 => x"82",
          3134 => x"38",
          3135 => x"8a",
          3136 => x"2e",
          3137 => x"8e",
          3138 => x"84",
          3139 => x"38",
          3140 => x"82",
          3141 => x"de",
          3142 => x"2e",
          3143 => x"79",
          3144 => x"38",
          3145 => x"83",
          3146 => x"bc",
          3147 => x"38",
          3148 => x"79",
          3149 => x"c6",
          3150 => x"c0",
          3151 => x"38",
          3152 => x"79",
          3153 => x"8d",
          3154 => x"80",
          3155 => x"38",
          3156 => x"2e",
          3157 => x"79",
          3158 => x"92",
          3159 => x"c2",
          3160 => x"38",
          3161 => x"2e",
          3162 => x"8e",
          3163 => x"80",
          3164 => x"ba",
          3165 => x"d4",
          3166 => x"38",
          3167 => x"79",
          3168 => x"8d",
          3169 => x"81",
          3170 => x"38",
          3171 => x"2e",
          3172 => x"79",
          3173 => x"8d",
          3174 => x"da",
          3175 => x"83",
          3176 => x"38",
          3177 => x"2e",
          3178 => x"8d",
          3179 => x"3d",
          3180 => x"53",
          3181 => x"51",
          3182 => x"82",
          3183 => x"88",
          3184 => x"a8",
          3185 => x"39",
          3186 => x"fc",
          3187 => x"84",
          3188 => x"de",
          3189 => x"98",
          3190 => x"88",
          3191 => x"25",
          3192 => x"44",
          3193 => x"05",
          3194 => x"80",
          3195 => x"51",
          3196 => x"3f",
          3197 => x"08",
          3198 => x"5a",
          3199 => x"82",
          3200 => x"d6",
          3201 => x"5f",
          3202 => x"82",
          3203 => x"8e",
          3204 => x"3d",
          3205 => x"53",
          3206 => x"51",
          3207 => x"82",
          3208 => x"80",
          3209 => x"38",
          3210 => x"52",
          3211 => x"05",
          3212 => x"cb",
          3213 => x"bb",
          3214 => x"82",
          3215 => x"8c",
          3216 => x"3d",
          3217 => x"53",
          3218 => x"51",
          3219 => x"82",
          3220 => x"80",
          3221 => x"64",
          3222 => x"d9",
          3223 => x"fe",
          3224 => x"ff",
          3225 => x"d0",
          3226 => x"bb",
          3227 => x"38",
          3228 => x"08",
          3229 => x"82",
          3230 => x"7a",
          3231 => x"be",
          3232 => x"cf",
          3233 => x"7a",
          3234 => x"b4",
          3235 => x"c4",
          3236 => x"f6",
          3237 => x"bb",
          3238 => x"90",
          3239 => x"b8",
          3240 => x"3f",
          3241 => x"8d",
          3242 => x"ff",
          3243 => x"8f",
          3244 => x"bb",
          3245 => x"3d",
          3246 => x"52",
          3247 => x"3f",
          3248 => x"bb",
          3249 => x"7b",
          3250 => x"3f",
          3251 => x"b5",
          3252 => x"05",
          3253 => x"3f",
          3254 => x"08",
          3255 => x"84",
          3256 => x"90",
          3257 => x"bb",
          3258 => x"3d",
          3259 => x"52",
          3260 => x"3f",
          3261 => x"08",
          3262 => x"84",
          3263 => x"90",
          3264 => x"d2",
          3265 => x"b9",
          3266 => x"bb",
          3267 => x"56",
          3268 => x"bb",
          3269 => x"ff",
          3270 => x"53",
          3271 => x"51",
          3272 => x"82",
          3273 => x"80",
          3274 => x"38",
          3275 => x"08",
          3276 => x"3f",
          3277 => x"b5",
          3278 => x"11",
          3279 => x"05",
          3280 => x"3f",
          3281 => x"08",
          3282 => x"e9",
          3283 => x"fe",
          3284 => x"ff",
          3285 => x"ce",
          3286 => x"bb",
          3287 => x"2e",
          3288 => x"b5",
          3289 => x"11",
          3290 => x"05",
          3291 => x"3f",
          3292 => x"08",
          3293 => x"bb",
          3294 => x"82",
          3295 => x"d4",
          3296 => x"64",
          3297 => x"7c",
          3298 => x"38",
          3299 => x"7b",
          3300 => x"5d",
          3301 => x"26",
          3302 => x"d9",
          3303 => x"ff",
          3304 => x"ff",
          3305 => x"ce",
          3306 => x"bb",
          3307 => x"2e",
          3308 => x"b5",
          3309 => x"11",
          3310 => x"05",
          3311 => x"3f",
          3312 => x"08",
          3313 => x"ed",
          3314 => x"fe",
          3315 => x"ff",
          3316 => x"cd",
          3317 => x"bb",
          3318 => x"2e",
          3319 => x"82",
          3320 => x"d3",
          3321 => x"5b",
          3322 => x"81",
          3323 => x"5a",
          3324 => x"05",
          3325 => x"34",
          3326 => x"43",
          3327 => x"3d",
          3328 => x"53",
          3329 => x"51",
          3330 => x"82",
          3331 => x"80",
          3332 => x"38",
          3333 => x"fc",
          3334 => x"84",
          3335 => x"92",
          3336 => x"98",
          3337 => x"f9",
          3338 => x"3d",
          3339 => x"53",
          3340 => x"51",
          3341 => x"82",
          3342 => x"80",
          3343 => x"38",
          3344 => x"51",
          3345 => x"64",
          3346 => x"27",
          3347 => x"70",
          3348 => x"5f",
          3349 => x"7d",
          3350 => x"79",
          3351 => x"7a",
          3352 => x"52",
          3353 => x"51",
          3354 => x"3f",
          3355 => x"81",
          3356 => x"d5",
          3357 => x"b0",
          3358 => x"39",
          3359 => x"80",
          3360 => x"84",
          3361 => x"aa",
          3362 => x"98",
          3363 => x"38",
          3364 => x"33",
          3365 => x"2e",
          3366 => x"b9",
          3367 => x"80",
          3368 => x"ba",
          3369 => x"79",
          3370 => x"38",
          3371 => x"08",
          3372 => x"82",
          3373 => x"5a",
          3374 => x"88",
          3375 => x"cc",
          3376 => x"39",
          3377 => x"33",
          3378 => x"2e",
          3379 => x"b9",
          3380 => x"9a",
          3381 => x"82",
          3382 => x"80",
          3383 => x"82",
          3384 => x"45",
          3385 => x"b9",
          3386 => x"80",
          3387 => x"3d",
          3388 => x"53",
          3389 => x"51",
          3390 => x"82",
          3391 => x"80",
          3392 => x"ba",
          3393 => x"79",
          3394 => x"38",
          3395 => x"08",
          3396 => x"39",
          3397 => x"33",
          3398 => x"2e",
          3399 => x"b9",
          3400 => x"bb",
          3401 => x"86",
          3402 => x"80",
          3403 => x"82",
          3404 => x"44",
          3405 => x"ba",
          3406 => x"79",
          3407 => x"38",
          3408 => x"08",
          3409 => x"82",
          3410 => x"5a",
          3411 => x"88",
          3412 => x"e0",
          3413 => x"39",
          3414 => x"08",
          3415 => x"b5",
          3416 => x"11",
          3417 => x"05",
          3418 => x"3f",
          3419 => x"08",
          3420 => x"38",
          3421 => x"5d",
          3422 => x"83",
          3423 => x"7b",
          3424 => x"30",
          3425 => x"9f",
          3426 => x"06",
          3427 => x"5b",
          3428 => x"88",
          3429 => x"2e",
          3430 => x"43",
          3431 => x"51",
          3432 => x"a0",
          3433 => x"62",
          3434 => x"64",
          3435 => x"3f",
          3436 => x"51",
          3437 => x"b5",
          3438 => x"11",
          3439 => x"05",
          3440 => x"3f",
          3441 => x"08",
          3442 => x"e9",
          3443 => x"fe",
          3444 => x"ff",
          3445 => x"c9",
          3446 => x"bb",
          3447 => x"2e",
          3448 => x"5a",
          3449 => x"05",
          3450 => x"64",
          3451 => x"b5",
          3452 => x"11",
          3453 => x"05",
          3454 => x"3f",
          3455 => x"08",
          3456 => x"b1",
          3457 => x"33",
          3458 => x"a7",
          3459 => x"a7",
          3460 => x"f8",
          3461 => x"c8",
          3462 => x"46",
          3463 => x"79",
          3464 => x"91",
          3465 => x"27",
          3466 => x"3d",
          3467 => x"53",
          3468 => x"51",
          3469 => x"82",
          3470 => x"80",
          3471 => x"64",
          3472 => x"cf",
          3473 => x"34",
          3474 => x"45",
          3475 => x"82",
          3476 => x"ce",
          3477 => x"ad",
          3478 => x"fe",
          3479 => x"ff",
          3480 => x"c2",
          3481 => x"bb",
          3482 => x"2e",
          3483 => x"b5",
          3484 => x"11",
          3485 => x"05",
          3486 => x"3f",
          3487 => x"08",
          3488 => x"38",
          3489 => x"80",
          3490 => x"7a",
          3491 => x"5c",
          3492 => x"b5",
          3493 => x"11",
          3494 => x"05",
          3495 => x"3f",
          3496 => x"08",
          3497 => x"8d",
          3498 => x"22",
          3499 => x"a7",
          3500 => x"a6",
          3501 => x"f8",
          3502 => x"c7",
          3503 => x"46",
          3504 => x"79",
          3505 => x"ed",
          3506 => x"26",
          3507 => x"82",
          3508 => x"39",
          3509 => x"f0",
          3510 => x"84",
          3511 => x"cb",
          3512 => x"98",
          3513 => x"93",
          3514 => x"02",
          3515 => x"22",
          3516 => x"05",
          3517 => x"42",
          3518 => x"82",
          3519 => x"cd",
          3520 => x"a5",
          3521 => x"fe",
          3522 => x"ff",
          3523 => x"c1",
          3524 => x"bb",
          3525 => x"2e",
          3526 => x"b5",
          3527 => x"11",
          3528 => x"05",
          3529 => x"3f",
          3530 => x"08",
          3531 => x"38",
          3532 => x"0c",
          3533 => x"05",
          3534 => x"fe",
          3535 => x"ff",
          3536 => x"c0",
          3537 => x"bb",
          3538 => x"38",
          3539 => x"61",
          3540 => x"52",
          3541 => x"51",
          3542 => x"3f",
          3543 => x"7a",
          3544 => x"3f",
          3545 => x"33",
          3546 => x"2e",
          3547 => x"9f",
          3548 => x"38",
          3549 => x"f0",
          3550 => x"84",
          3551 => x"ab",
          3552 => x"98",
          3553 => x"8d",
          3554 => x"71",
          3555 => x"84",
          3556 => x"bb",
          3557 => x"dc",
          3558 => x"3f",
          3559 => x"82",
          3560 => x"cb",
          3561 => x"51",
          3562 => x"f2",
          3563 => x"a8",
          3564 => x"cf",
          3565 => x"97",
          3566 => x"f9",
          3567 => x"ac",
          3568 => x"3f",
          3569 => x"0b",
          3570 => x"84",
          3571 => x"81",
          3572 => x"94",
          3573 => x"dd",
          3574 => x"c0",
          3575 => x"3f",
          3576 => x"0b",
          3577 => x"84",
          3578 => x"83",
          3579 => x"94",
          3580 => x"c1",
          3581 => x"ff",
          3582 => x"ff",
          3583 => x"c5",
          3584 => x"bb",
          3585 => x"2e",
          3586 => x"64",
          3587 => x"d4",
          3588 => x"c2",
          3589 => x"79",
          3590 => x"ff",
          3591 => x"ff",
          3592 => x"c5",
          3593 => x"bb",
          3594 => x"2e",
          3595 => x"64",
          3596 => x"f0",
          3597 => x"9e",
          3598 => x"79",
          3599 => x"98",
          3600 => x"f0",
          3601 => x"bb",
          3602 => x"82",
          3603 => x"ff",
          3604 => x"f0",
          3605 => x"a9",
          3606 => x"a7",
          3607 => x"d7",
          3608 => x"39",
          3609 => x"51",
          3610 => x"80",
          3611 => x"39",
          3612 => x"f0",
          3613 => x"46",
          3614 => x"79",
          3615 => x"b5",
          3616 => x"06",
          3617 => x"2e",
          3618 => x"b5",
          3619 => x"05",
          3620 => x"3f",
          3621 => x"08",
          3622 => x"7c",
          3623 => x"38",
          3624 => x"89",
          3625 => x"2e",
          3626 => x"cd",
          3627 => x"2e",
          3628 => x"c5",
          3629 => x"d8",
          3630 => x"82",
          3631 => x"80",
          3632 => x"e0",
          3633 => x"ff",
          3634 => x"ff",
          3635 => x"bb",
          3636 => x"80",
          3637 => x"ff",
          3638 => x"ff",
          3639 => x"ab",
          3640 => x"82",
          3641 => x"80",
          3642 => x"f0",
          3643 => x"ff",
          3644 => x"ff",
          3645 => x"93",
          3646 => x"80",
          3647 => x"fc",
          3648 => x"ff",
          3649 => x"ff",
          3650 => x"82",
          3651 => x"82",
          3652 => x"82",
          3653 => x"80",
          3654 => x"80",
          3655 => x"80",
          3656 => x"80",
          3657 => x"ff",
          3658 => x"e7",
          3659 => x"bb",
          3660 => x"bb",
          3661 => x"70",
          3662 => x"07",
          3663 => x"5c",
          3664 => x"5b",
          3665 => x"83",
          3666 => x"79",
          3667 => x"79",
          3668 => x"38",
          3669 => x"81",
          3670 => x"5a",
          3671 => x"38",
          3672 => x"7e",
          3673 => x"5a",
          3674 => x"7f",
          3675 => x"81",
          3676 => x"38",
          3677 => x"51",
          3678 => x"ee",
          3679 => x"3d",
          3680 => x"82",
          3681 => x"87",
          3682 => x"70",
          3683 => x"87",
          3684 => x"72",
          3685 => x"3f",
          3686 => x"08",
          3687 => x"08",
          3688 => x"84",
          3689 => x"51",
          3690 => x"72",
          3691 => x"08",
          3692 => x"87",
          3693 => x"70",
          3694 => x"87",
          3695 => x"72",
          3696 => x"3f",
          3697 => x"08",
          3698 => x"08",
          3699 => x"84",
          3700 => x"51",
          3701 => x"72",
          3702 => x"08",
          3703 => x"8c",
          3704 => x"87",
          3705 => x"0c",
          3706 => x"0b",
          3707 => x"94",
          3708 => x"82",
          3709 => x"ee",
          3710 => x"84",
          3711 => x"34",
          3712 => x"d2",
          3713 => x"3d",
          3714 => x"0c",
          3715 => x"82",
          3716 => x"54",
          3717 => x"93",
          3718 => x"aa",
          3719 => x"e3",
          3720 => x"a0",
          3721 => x"3f",
          3722 => x"51",
          3723 => x"81",
          3724 => x"3f",
          3725 => x"80",
          3726 => x"0d",
          3727 => x"53",
          3728 => x"52",
          3729 => x"82",
          3730 => x"81",
          3731 => x"07",
          3732 => x"52",
          3733 => x"e8",
          3734 => x"bb",
          3735 => x"3d",
          3736 => x"3d",
          3737 => x"08",
          3738 => x"73",
          3739 => x"74",
          3740 => x"38",
          3741 => x"70",
          3742 => x"81",
          3743 => x"81",
          3744 => x"39",
          3745 => x"70",
          3746 => x"81",
          3747 => x"81",
          3748 => x"54",
          3749 => x"81",
          3750 => x"06",
          3751 => x"39",
          3752 => x"80",
          3753 => x"54",
          3754 => x"83",
          3755 => x"70",
          3756 => x"38",
          3757 => x"98",
          3758 => x"52",
          3759 => x"52",
          3760 => x"2e",
          3761 => x"54",
          3762 => x"84",
          3763 => x"38",
          3764 => x"52",
          3765 => x"2e",
          3766 => x"83",
          3767 => x"70",
          3768 => x"30",
          3769 => x"76",
          3770 => x"51",
          3771 => x"88",
          3772 => x"70",
          3773 => x"34",
          3774 => x"72",
          3775 => x"bb",
          3776 => x"3d",
          3777 => x"3d",
          3778 => x"72",
          3779 => x"92",
          3780 => x"fc",
          3781 => x"51",
          3782 => x"3f",
          3783 => x"08",
          3784 => x"53",
          3785 => x"53",
          3786 => x"98",
          3787 => x"0d",
          3788 => x"0d",
          3789 => x"33",
          3790 => x"53",
          3791 => x"8b",
          3792 => x"38",
          3793 => x"ff",
          3794 => x"52",
          3795 => x"81",
          3796 => x"13",
          3797 => x"52",
          3798 => x"80",
          3799 => x"13",
          3800 => x"52",
          3801 => x"80",
          3802 => x"13",
          3803 => x"52",
          3804 => x"80",
          3805 => x"13",
          3806 => x"52",
          3807 => x"26",
          3808 => x"8a",
          3809 => x"87",
          3810 => x"e7",
          3811 => x"38",
          3812 => x"c0",
          3813 => x"72",
          3814 => x"98",
          3815 => x"13",
          3816 => x"98",
          3817 => x"13",
          3818 => x"98",
          3819 => x"13",
          3820 => x"98",
          3821 => x"13",
          3822 => x"98",
          3823 => x"13",
          3824 => x"98",
          3825 => x"87",
          3826 => x"0c",
          3827 => x"98",
          3828 => x"0b",
          3829 => x"9c",
          3830 => x"71",
          3831 => x"0c",
          3832 => x"04",
          3833 => x"7f",
          3834 => x"98",
          3835 => x"7d",
          3836 => x"98",
          3837 => x"7d",
          3838 => x"c0",
          3839 => x"5a",
          3840 => x"34",
          3841 => x"b4",
          3842 => x"83",
          3843 => x"c0",
          3844 => x"5a",
          3845 => x"34",
          3846 => x"ac",
          3847 => x"85",
          3848 => x"c0",
          3849 => x"5a",
          3850 => x"34",
          3851 => x"a4",
          3852 => x"88",
          3853 => x"c0",
          3854 => x"5a",
          3855 => x"23",
          3856 => x"79",
          3857 => x"06",
          3858 => x"ff",
          3859 => x"86",
          3860 => x"85",
          3861 => x"84",
          3862 => x"83",
          3863 => x"82",
          3864 => x"7d",
          3865 => x"06",
          3866 => x"b8",
          3867 => x"e6",
          3868 => x"0d",
          3869 => x"0d",
          3870 => x"33",
          3871 => x"33",
          3872 => x"06",
          3873 => x"87",
          3874 => x"51",
          3875 => x"86",
          3876 => x"94",
          3877 => x"08",
          3878 => x"70",
          3879 => x"54",
          3880 => x"2e",
          3881 => x"91",
          3882 => x"06",
          3883 => x"d7",
          3884 => x"32",
          3885 => x"51",
          3886 => x"2e",
          3887 => x"93",
          3888 => x"06",
          3889 => x"ff",
          3890 => x"81",
          3891 => x"87",
          3892 => x"52",
          3893 => x"86",
          3894 => x"94",
          3895 => x"72",
          3896 => x"bb",
          3897 => x"3d",
          3898 => x"3d",
          3899 => x"05",
          3900 => x"70",
          3901 => x"52",
          3902 => x"b9",
          3903 => x"3d",
          3904 => x"3d",
          3905 => x"05",
          3906 => x"8a",
          3907 => x"06",
          3908 => x"52",
          3909 => x"3f",
          3910 => x"33",
          3911 => x"06",
          3912 => x"c0",
          3913 => x"76",
          3914 => x"38",
          3915 => x"94",
          3916 => x"70",
          3917 => x"81",
          3918 => x"54",
          3919 => x"8c",
          3920 => x"2a",
          3921 => x"51",
          3922 => x"38",
          3923 => x"70",
          3924 => x"53",
          3925 => x"8d",
          3926 => x"2a",
          3927 => x"51",
          3928 => x"be",
          3929 => x"ff",
          3930 => x"c0",
          3931 => x"72",
          3932 => x"38",
          3933 => x"90",
          3934 => x"0c",
          3935 => x"bb",
          3936 => x"3d",
          3937 => x"3d",
          3938 => x"80",
          3939 => x"81",
          3940 => x"53",
          3941 => x"2e",
          3942 => x"71",
          3943 => x"81",
          3944 => x"b8",
          3945 => x"ff",
          3946 => x"55",
          3947 => x"94",
          3948 => x"80",
          3949 => x"87",
          3950 => x"51",
          3951 => x"96",
          3952 => x"06",
          3953 => x"70",
          3954 => x"38",
          3955 => x"70",
          3956 => x"51",
          3957 => x"72",
          3958 => x"81",
          3959 => x"70",
          3960 => x"38",
          3961 => x"70",
          3962 => x"51",
          3963 => x"38",
          3964 => x"06",
          3965 => x"94",
          3966 => x"80",
          3967 => x"87",
          3968 => x"52",
          3969 => x"81",
          3970 => x"70",
          3971 => x"53",
          3972 => x"ff",
          3973 => x"82",
          3974 => x"89",
          3975 => x"fe",
          3976 => x"b9",
          3977 => x"81",
          3978 => x"52",
          3979 => x"84",
          3980 => x"2e",
          3981 => x"c0",
          3982 => x"70",
          3983 => x"2a",
          3984 => x"51",
          3985 => x"80",
          3986 => x"71",
          3987 => x"51",
          3988 => x"80",
          3989 => x"2e",
          3990 => x"c0",
          3991 => x"71",
          3992 => x"ff",
          3993 => x"98",
          3994 => x"3d",
          3995 => x"af",
          3996 => x"98",
          3997 => x"06",
          3998 => x"0c",
          3999 => x"0d",
          4000 => x"33",
          4001 => x"06",
          4002 => x"c0",
          4003 => x"70",
          4004 => x"38",
          4005 => x"94",
          4006 => x"70",
          4007 => x"81",
          4008 => x"51",
          4009 => x"80",
          4010 => x"72",
          4011 => x"51",
          4012 => x"80",
          4013 => x"2e",
          4014 => x"c0",
          4015 => x"71",
          4016 => x"2b",
          4017 => x"51",
          4018 => x"82",
          4019 => x"84",
          4020 => x"ff",
          4021 => x"c0",
          4022 => x"70",
          4023 => x"06",
          4024 => x"80",
          4025 => x"38",
          4026 => x"a4",
          4027 => x"bc",
          4028 => x"9e",
          4029 => x"b9",
          4030 => x"c0",
          4031 => x"82",
          4032 => x"87",
          4033 => x"08",
          4034 => x"0c",
          4035 => x"9c",
          4036 => x"cc",
          4037 => x"9e",
          4038 => x"b9",
          4039 => x"c0",
          4040 => x"82",
          4041 => x"87",
          4042 => x"08",
          4043 => x"0c",
          4044 => x"b4",
          4045 => x"dc",
          4046 => x"9e",
          4047 => x"b9",
          4048 => x"c0",
          4049 => x"82",
          4050 => x"87",
          4051 => x"08",
          4052 => x"0c",
          4053 => x"c4",
          4054 => x"ec",
          4055 => x"9e",
          4056 => x"70",
          4057 => x"23",
          4058 => x"84",
          4059 => x"f4",
          4060 => x"9e",
          4061 => x"b9",
          4062 => x"c0",
          4063 => x"82",
          4064 => x"81",
          4065 => x"80",
          4066 => x"87",
          4067 => x"08",
          4068 => x"0a",
          4069 => x"52",
          4070 => x"83",
          4071 => x"71",
          4072 => x"34",
          4073 => x"c0",
          4074 => x"70",
          4075 => x"06",
          4076 => x"70",
          4077 => x"38",
          4078 => x"82",
          4079 => x"80",
          4080 => x"9e",
          4081 => x"90",
          4082 => x"51",
          4083 => x"80",
          4084 => x"81",
          4085 => x"ba",
          4086 => x"0b",
          4087 => x"90",
          4088 => x"80",
          4089 => x"52",
          4090 => x"2e",
          4091 => x"52",
          4092 => x"84",
          4093 => x"87",
          4094 => x"08",
          4095 => x"80",
          4096 => x"52",
          4097 => x"83",
          4098 => x"71",
          4099 => x"34",
          4100 => x"c0",
          4101 => x"70",
          4102 => x"06",
          4103 => x"70",
          4104 => x"38",
          4105 => x"82",
          4106 => x"80",
          4107 => x"9e",
          4108 => x"84",
          4109 => x"51",
          4110 => x"80",
          4111 => x"81",
          4112 => x"ba",
          4113 => x"0b",
          4114 => x"90",
          4115 => x"80",
          4116 => x"52",
          4117 => x"2e",
          4118 => x"52",
          4119 => x"88",
          4120 => x"87",
          4121 => x"08",
          4122 => x"80",
          4123 => x"52",
          4124 => x"83",
          4125 => x"71",
          4126 => x"34",
          4127 => x"c0",
          4128 => x"70",
          4129 => x"06",
          4130 => x"70",
          4131 => x"38",
          4132 => x"82",
          4133 => x"80",
          4134 => x"9e",
          4135 => x"a0",
          4136 => x"52",
          4137 => x"2e",
          4138 => x"52",
          4139 => x"8b",
          4140 => x"9e",
          4141 => x"98",
          4142 => x"8a",
          4143 => x"51",
          4144 => x"8c",
          4145 => x"87",
          4146 => x"08",
          4147 => x"06",
          4148 => x"70",
          4149 => x"38",
          4150 => x"82",
          4151 => x"87",
          4152 => x"08",
          4153 => x"06",
          4154 => x"51",
          4155 => x"82",
          4156 => x"80",
          4157 => x"9e",
          4158 => x"88",
          4159 => x"52",
          4160 => x"83",
          4161 => x"71",
          4162 => x"34",
          4163 => x"90",
          4164 => x"06",
          4165 => x"82",
          4166 => x"83",
          4167 => x"fb",
          4168 => x"aa",
          4169 => x"b8",
          4170 => x"ba",
          4171 => x"73",
          4172 => x"38",
          4173 => x"51",
          4174 => x"3f",
          4175 => x"51",
          4176 => x"3f",
          4177 => x"33",
          4178 => x"2e",
          4179 => x"b9",
          4180 => x"b9",
          4181 => x"54",
          4182 => x"90",
          4183 => x"f6",
          4184 => x"87",
          4185 => x"80",
          4186 => x"82",
          4187 => x"82",
          4188 => x"11",
          4189 => x"ab",
          4190 => x"90",
          4191 => x"ba",
          4192 => x"73",
          4193 => x"38",
          4194 => x"08",
          4195 => x"08",
          4196 => x"82",
          4197 => x"ff",
          4198 => x"82",
          4199 => x"54",
          4200 => x"94",
          4201 => x"c4",
          4202 => x"c8",
          4203 => x"52",
          4204 => x"51",
          4205 => x"3f",
          4206 => x"33",
          4207 => x"2e",
          4208 => x"b9",
          4209 => x"b9",
          4210 => x"54",
          4211 => x"80",
          4212 => x"82",
          4213 => x"8b",
          4214 => x"80",
          4215 => x"82",
          4216 => x"52",
          4217 => x"51",
          4218 => x"3f",
          4219 => x"33",
          4220 => x"2e",
          4221 => x"ba",
          4222 => x"82",
          4223 => x"ff",
          4224 => x"82",
          4225 => x"54",
          4226 => x"8e",
          4227 => x"8e",
          4228 => x"ac",
          4229 => x"8f",
          4230 => x"ba",
          4231 => x"73",
          4232 => x"38",
          4233 => x"51",
          4234 => x"3f",
          4235 => x"33",
          4236 => x"2e",
          4237 => x"ad",
          4238 => x"b6",
          4239 => x"ba",
          4240 => x"73",
          4241 => x"38",
          4242 => x"51",
          4243 => x"3f",
          4244 => x"33",
          4245 => x"2e",
          4246 => x"ad",
          4247 => x"b6",
          4248 => x"ba",
          4249 => x"73",
          4250 => x"38",
          4251 => x"51",
          4252 => x"3f",
          4253 => x"51",
          4254 => x"3f",
          4255 => x"08",
          4256 => x"cc",
          4257 => x"ce",
          4258 => x"e8",
          4259 => x"ad",
          4260 => x"8e",
          4261 => x"b9",
          4262 => x"82",
          4263 => x"ff",
          4264 => x"82",
          4265 => x"ff",
          4266 => x"82",
          4267 => x"52",
          4268 => x"51",
          4269 => x"3f",
          4270 => x"08",
          4271 => x"c0",
          4272 => x"cc",
          4273 => x"bb",
          4274 => x"84",
          4275 => x"71",
          4276 => x"82",
          4277 => x"52",
          4278 => x"51",
          4279 => x"3f",
          4280 => x"33",
          4281 => x"2e",
          4282 => x"b9",
          4283 => x"bd",
          4284 => x"75",
          4285 => x"3f",
          4286 => x"08",
          4287 => x"29",
          4288 => x"54",
          4289 => x"98",
          4290 => x"af",
          4291 => x"8d",
          4292 => x"ba",
          4293 => x"73",
          4294 => x"38",
          4295 => x"08",
          4296 => x"c0",
          4297 => x"cb",
          4298 => x"bb",
          4299 => x"84",
          4300 => x"71",
          4301 => x"82",
          4302 => x"52",
          4303 => x"51",
          4304 => x"3f",
          4305 => x"51",
          4306 => x"3f",
          4307 => x"04",
          4308 => x"02",
          4309 => x"ff",
          4310 => x"84",
          4311 => x"71",
          4312 => x"9a",
          4313 => x"71",
          4314 => x"af",
          4315 => x"39",
          4316 => x"51",
          4317 => x"b0",
          4318 => x"39",
          4319 => x"51",
          4320 => x"b0",
          4321 => x"39",
          4322 => x"51",
          4323 => x"3f",
          4324 => x"04",
          4325 => x"0c",
          4326 => x"0d",
          4327 => x"84",
          4328 => x"52",
          4329 => x"70",
          4330 => x"82",
          4331 => x"72",
          4332 => x"0d",
          4333 => x"0d",
          4334 => x"84",
          4335 => x"ba",
          4336 => x"80",
          4337 => x"09",
          4338 => x"94",
          4339 => x"82",
          4340 => x"73",
          4341 => x"3d",
          4342 => x"0b",
          4343 => x"84",
          4344 => x"ba",
          4345 => x"c0",
          4346 => x"04",
          4347 => x"76",
          4348 => x"98",
          4349 => x"2b",
          4350 => x"72",
          4351 => x"82",
          4352 => x"51",
          4353 => x"80",
          4354 => x"a8",
          4355 => x"53",
          4356 => x"9c",
          4357 => x"a4",
          4358 => x"02",
          4359 => x"05",
          4360 => x"52",
          4361 => x"72",
          4362 => x"06",
          4363 => x"53",
          4364 => x"98",
          4365 => x"0d",
          4366 => x"0d",
          4367 => x"05",
          4368 => x"71",
          4369 => x"53",
          4370 => x"a2",
          4371 => x"ff",
          4372 => x"a0",
          4373 => x"cd",
          4374 => x"ff",
          4375 => x"72",
          4376 => x"52",
          4377 => x"71",
          4378 => x"52",
          4379 => x"51",
          4380 => x"3f",
          4381 => x"86",
          4382 => x"f6",
          4383 => x"02",
          4384 => x"05",
          4385 => x"05",
          4386 => x"82",
          4387 => x"70",
          4388 => x"ba",
          4389 => x"08",
          4390 => x"5a",
          4391 => x"80",
          4392 => x"74",
          4393 => x"3f",
          4394 => x"33",
          4395 => x"82",
          4396 => x"81",
          4397 => x"58",
          4398 => x"b6",
          4399 => x"98",
          4400 => x"82",
          4401 => x"70",
          4402 => x"ba",
          4403 => x"08",
          4404 => x"74",
          4405 => x"38",
          4406 => x"52",
          4407 => x"bf",
          4408 => x"ba",
          4409 => x"05",
          4410 => x"ba",
          4411 => x"81",
          4412 => x"93",
          4413 => x"38",
          4414 => x"ba",
          4415 => x"80",
          4416 => x"82",
          4417 => x"56",
          4418 => x"ac",
          4419 => x"e8",
          4420 => x"a4",
          4421 => x"fc",
          4422 => x"53",
          4423 => x"51",
          4424 => x"3f",
          4425 => x"08",
          4426 => x"81",
          4427 => x"82",
          4428 => x"51",
          4429 => x"3f",
          4430 => x"04",
          4431 => x"82",
          4432 => x"93",
          4433 => x"52",
          4434 => x"89",
          4435 => x"99",
          4436 => x"73",
          4437 => x"84",
          4438 => x"73",
          4439 => x"38",
          4440 => x"ba",
          4441 => x"ba",
          4442 => x"71",
          4443 => x"38",
          4444 => x"de",
          4445 => x"ba",
          4446 => x"98",
          4447 => x"0b",
          4448 => x"0c",
          4449 => x"04",
          4450 => x"81",
          4451 => x"82",
          4452 => x"51",
          4453 => x"3f",
          4454 => x"08",
          4455 => x"82",
          4456 => x"53",
          4457 => x"88",
          4458 => x"56",
          4459 => x"3f",
          4460 => x"08",
          4461 => x"38",
          4462 => x"bb",
          4463 => x"bb",
          4464 => x"80",
          4465 => x"98",
          4466 => x"38",
          4467 => x"08",
          4468 => x"17",
          4469 => x"74",
          4470 => x"76",
          4471 => x"82",
          4472 => x"57",
          4473 => x"3f",
          4474 => x"09",
          4475 => x"af",
          4476 => x"0d",
          4477 => x"0d",
          4478 => x"ad",
          4479 => x"5a",
          4480 => x"58",
          4481 => x"ba",
          4482 => x"80",
          4483 => x"82",
          4484 => x"81",
          4485 => x"0b",
          4486 => x"08",
          4487 => x"f8",
          4488 => x"70",
          4489 => x"8a",
          4490 => x"bb",
          4491 => x"2e",
          4492 => x"51",
          4493 => x"3f",
          4494 => x"08",
          4495 => x"55",
          4496 => x"bb",
          4497 => x"8e",
          4498 => x"98",
          4499 => x"70",
          4500 => x"80",
          4501 => x"09",
          4502 => x"72",
          4503 => x"51",
          4504 => x"77",
          4505 => x"73",
          4506 => x"82",
          4507 => x"8c",
          4508 => x"51",
          4509 => x"3f",
          4510 => x"08",
          4511 => x"38",
          4512 => x"51",
          4513 => x"3f",
          4514 => x"09",
          4515 => x"38",
          4516 => x"51",
          4517 => x"3f",
          4518 => x"ba",
          4519 => x"3d",
          4520 => x"bb",
          4521 => x"34",
          4522 => x"82",
          4523 => x"a9",
          4524 => x"f6",
          4525 => x"7e",
          4526 => x"72",
          4527 => x"5a",
          4528 => x"2e",
          4529 => x"a2",
          4530 => x"78",
          4531 => x"76",
          4532 => x"81",
          4533 => x"70",
          4534 => x"58",
          4535 => x"2e",
          4536 => x"86",
          4537 => x"26",
          4538 => x"54",
          4539 => x"82",
          4540 => x"70",
          4541 => x"ff",
          4542 => x"82",
          4543 => x"53",
          4544 => x"08",
          4545 => x"aa",
          4546 => x"98",
          4547 => x"38",
          4548 => x"55",
          4549 => x"88",
          4550 => x"2e",
          4551 => x"39",
          4552 => x"ad",
          4553 => x"5a",
          4554 => x"11",
          4555 => x"51",
          4556 => x"3f",
          4557 => x"08",
          4558 => x"38",
          4559 => x"78",
          4560 => x"fd",
          4561 => x"bb",
          4562 => x"ff",
          4563 => x"85",
          4564 => x"91",
          4565 => x"70",
          4566 => x"51",
          4567 => x"27",
          4568 => x"80",
          4569 => x"bb",
          4570 => x"3d",
          4571 => x"3d",
          4572 => x"08",
          4573 => x"b4",
          4574 => x"5f",
          4575 => x"af",
          4576 => x"ba",
          4577 => x"ba",
          4578 => x"5b",
          4579 => x"38",
          4580 => x"e8",
          4581 => x"73",
          4582 => x"55",
          4583 => x"81",
          4584 => x"70",
          4585 => x"56",
          4586 => x"81",
          4587 => x"51",
          4588 => x"82",
          4589 => x"82",
          4590 => x"82",
          4591 => x"80",
          4592 => x"38",
          4593 => x"52",
          4594 => x"08",
          4595 => x"b4",
          4596 => x"98",
          4597 => x"8c",
          4598 => x"d0",
          4599 => x"a3",
          4600 => x"39",
          4601 => x"08",
          4602 => x"ec",
          4603 => x"f8",
          4604 => x"70",
          4605 => x"86",
          4606 => x"bb",
          4607 => x"82",
          4608 => x"74",
          4609 => x"06",
          4610 => x"82",
          4611 => x"51",
          4612 => x"3f",
          4613 => x"08",
          4614 => x"82",
          4615 => x"25",
          4616 => x"bb",
          4617 => x"05",
          4618 => x"55",
          4619 => x"80",
          4620 => x"ff",
          4621 => x"51",
          4622 => x"81",
          4623 => x"ff",
          4624 => x"93",
          4625 => x"38",
          4626 => x"ff",
          4627 => x"06",
          4628 => x"86",
          4629 => x"ba",
          4630 => x"8c",
          4631 => x"ec",
          4632 => x"84",
          4633 => x"3f",
          4634 => x"ec",
          4635 => x"bb",
          4636 => x"2b",
          4637 => x"51",
          4638 => x"2e",
          4639 => x"81",
          4640 => x"d2",
          4641 => x"98",
          4642 => x"2c",
          4643 => x"33",
          4644 => x"70",
          4645 => x"98",
          4646 => x"84",
          4647 => x"a4",
          4648 => x"15",
          4649 => x"51",
          4650 => x"59",
          4651 => x"58",
          4652 => x"78",
          4653 => x"38",
          4654 => x"b4",
          4655 => x"80",
          4656 => x"ff",
          4657 => x"98",
          4658 => x"80",
          4659 => x"ce",
          4660 => x"74",
          4661 => x"f6",
          4662 => x"bb",
          4663 => x"ff",
          4664 => x"80",
          4665 => x"74",
          4666 => x"34",
          4667 => x"39",
          4668 => x"0a",
          4669 => x"0a",
          4670 => x"2c",
          4671 => x"06",
          4672 => x"73",
          4673 => x"38",
          4674 => x"52",
          4675 => x"dc",
          4676 => x"98",
          4677 => x"06",
          4678 => x"38",
          4679 => x"56",
          4680 => x"80",
          4681 => x"1c",
          4682 => x"d2",
          4683 => x"98",
          4684 => x"2c",
          4685 => x"33",
          4686 => x"70",
          4687 => x"10",
          4688 => x"2b",
          4689 => x"11",
          4690 => x"51",
          4691 => x"51",
          4692 => x"2e",
          4693 => x"fe",
          4694 => x"b0",
          4695 => x"7d",
          4696 => x"82",
          4697 => x"80",
          4698 => x"c0",
          4699 => x"75",
          4700 => x"34",
          4701 => x"c0",
          4702 => x"3d",
          4703 => x"0c",
          4704 => x"95",
          4705 => x"38",
          4706 => x"82",
          4707 => x"54",
          4708 => x"82",
          4709 => x"54",
          4710 => x"fd",
          4711 => x"d2",
          4712 => x"73",
          4713 => x"38",
          4714 => x"70",
          4715 => x"55",
          4716 => x"9e",
          4717 => x"54",
          4718 => x"15",
          4719 => x"80",
          4720 => x"ff",
          4721 => x"98",
          4722 => x"cc",
          4723 => x"55",
          4724 => x"d2",
          4725 => x"11",
          4726 => x"82",
          4727 => x"73",
          4728 => x"3d",
          4729 => x"82",
          4730 => x"54",
          4731 => x"89",
          4732 => x"54",
          4733 => x"c8",
          4734 => x"cc",
          4735 => x"80",
          4736 => x"ff",
          4737 => x"98",
          4738 => x"c8",
          4739 => x"56",
          4740 => x"25",
          4741 => x"1a",
          4742 => x"54",
          4743 => x"3f",
          4744 => x"0a",
          4745 => x"0a",
          4746 => x"2c",
          4747 => x"33",
          4748 => x"73",
          4749 => x"38",
          4750 => x"33",
          4751 => x"70",
          4752 => x"d2",
          4753 => x"51",
          4754 => x"77",
          4755 => x"38",
          4756 => x"a9",
          4757 => x"81",
          4758 => x"81",
          4759 => x"70",
          4760 => x"d2",
          4761 => x"51",
          4762 => x"24",
          4763 => x"f8",
          4764 => x"34",
          4765 => x"1b",
          4766 => x"cc",
          4767 => x"82",
          4768 => x"f3",
          4769 => x"e4",
          4770 => x"cc",
          4771 => x"ff",
          4772 => x"73",
          4773 => x"d0",
          4774 => x"c8",
          4775 => x"54",
          4776 => x"c8",
          4777 => x"54",
          4778 => x"cc",
          4779 => x"ff",
          4780 => x"82",
          4781 => x"70",
          4782 => x"98",
          4783 => x"c8",
          4784 => x"56",
          4785 => x"25",
          4786 => x"1a",
          4787 => x"33",
          4788 => x"33",
          4789 => x"cd",
          4790 => x"80",
          4791 => x"80",
          4792 => x"98",
          4793 => x"c8",
          4794 => x"55",
          4795 => x"da",
          4796 => x"ff",
          4797 => x"82",
          4798 => x"70",
          4799 => x"98",
          4800 => x"c8",
          4801 => x"56",
          4802 => x"24",
          4803 => x"88",
          4804 => x"91",
          4805 => x"80",
          4806 => x"80",
          4807 => x"98",
          4808 => x"c8",
          4809 => x"55",
          4810 => x"e3",
          4811 => x"39",
          4812 => x"33",
          4813 => x"80",
          4814 => x"51",
          4815 => x"3f",
          4816 => x"52",
          4817 => x"eb",
          4818 => x"98",
          4819 => x"06",
          4820 => x"38",
          4821 => x"33",
          4822 => x"2e",
          4823 => x"53",
          4824 => x"51",
          4825 => x"84",
          4826 => x"34",
          4827 => x"d2",
          4828 => x"0b",
          4829 => x"34",
          4830 => x"98",
          4831 => x"0d",
          4832 => x"cc",
          4833 => x"80",
          4834 => x"38",
          4835 => x"a7",
          4836 => x"d2",
          4837 => x"05",
          4838 => x"d2",
          4839 => x"81",
          4840 => x"e2",
          4841 => x"cc",
          4842 => x"c8",
          4843 => x"73",
          4844 => x"b4",
          4845 => x"54",
          4846 => x"c8",
          4847 => x"2b",
          4848 => x"75",
          4849 => x"56",
          4850 => x"74",
          4851 => x"74",
          4852 => x"14",
          4853 => x"73",
          4854 => x"a6",
          4855 => x"81",
          4856 => x"81",
          4857 => x"70",
          4858 => x"d2",
          4859 => x"51",
          4860 => x"24",
          4861 => x"51",
          4862 => x"3f",
          4863 => x"33",
          4864 => x"70",
          4865 => x"d2",
          4866 => x"51",
          4867 => x"74",
          4868 => x"38",
          4869 => x"a6",
          4870 => x"81",
          4871 => x"81",
          4872 => x"70",
          4873 => x"d2",
          4874 => x"51",
          4875 => x"25",
          4876 => x"b4",
          4877 => x"cc",
          4878 => x"ff",
          4879 => x"c8",
          4880 => x"54",
          4881 => x"f8",
          4882 => x"14",
          4883 => x"d2",
          4884 => x"1a",
          4885 => x"54",
          4886 => x"3f",
          4887 => x"33",
          4888 => x"06",
          4889 => x"33",
          4890 => x"75",
          4891 => x"38",
          4892 => x"82",
          4893 => x"80",
          4894 => x"88",
          4895 => x"3f",
          4896 => x"d2",
          4897 => x"0b",
          4898 => x"34",
          4899 => x"7a",
          4900 => x"ba",
          4901 => x"74",
          4902 => x"38",
          4903 => x"ae",
          4904 => x"bb",
          4905 => x"d2",
          4906 => x"bb",
          4907 => x"ff",
          4908 => x"53",
          4909 => x"51",
          4910 => x"3f",
          4911 => x"c0",
          4912 => x"29",
          4913 => x"05",
          4914 => x"56",
          4915 => x"2e",
          4916 => x"51",
          4917 => x"3f",
          4918 => x"08",
          4919 => x"34",
          4920 => x"08",
          4921 => x"81",
          4922 => x"52",
          4923 => x"af",
          4924 => x"1b",
          4925 => x"39",
          4926 => x"74",
          4927 => x"e8",
          4928 => x"ff",
          4929 => x"99",
          4930 => x"2e",
          4931 => x"ae",
          4932 => x"98",
          4933 => x"80",
          4934 => x"74",
          4935 => x"85",
          4936 => x"98",
          4937 => x"c8",
          4938 => x"98",
          4939 => x"06",
          4940 => x"74",
          4941 => x"ff",
          4942 => x"80",
          4943 => x"84",
          4944 => x"9c",
          4945 => x"56",
          4946 => x"2e",
          4947 => x"51",
          4948 => x"3f",
          4949 => x"08",
          4950 => x"34",
          4951 => x"08",
          4952 => x"81",
          4953 => x"52",
          4954 => x"ae",
          4955 => x"1b",
          4956 => x"ff",
          4957 => x"39",
          4958 => x"c8",
          4959 => x"34",
          4960 => x"53",
          4961 => x"33",
          4962 => x"ed",
          4963 => x"d8",
          4964 => x"cc",
          4965 => x"ff",
          4966 => x"c8",
          4967 => x"54",
          4968 => x"f5",
          4969 => x"14",
          4970 => x"d2",
          4971 => x"1a",
          4972 => x"54",
          4973 => x"3f",
          4974 => x"82",
          4975 => x"54",
          4976 => x"f5",
          4977 => x"51",
          4978 => x"3f",
          4979 => x"33",
          4980 => x"73",
          4981 => x"34",
          4982 => x"f9",
          4983 => x"c0",
          4984 => x"bb",
          4985 => x"80",
          4986 => x"8c",
          4987 => x"53",
          4988 => x"c0",
          4989 => x"b2",
          4990 => x"bb",
          4991 => x"80",
          4992 => x"34",
          4993 => x"81",
          4994 => x"bb",
          4995 => x"77",
          4996 => x"76",
          4997 => x"82",
          4998 => x"54",
          4999 => x"34",
          5000 => x"34",
          5001 => x"08",
          5002 => x"22",
          5003 => x"80",
          5004 => x"83",
          5005 => x"70",
          5006 => x"51",
          5007 => x"88",
          5008 => x"89",
          5009 => x"bb",
          5010 => x"88",
          5011 => x"90",
          5012 => x"11",
          5013 => x"77",
          5014 => x"76",
          5015 => x"89",
          5016 => x"ff",
          5017 => x"52",
          5018 => x"72",
          5019 => x"fb",
          5020 => x"82",
          5021 => x"ff",
          5022 => x"51",
          5023 => x"bb",
          5024 => x"3d",
          5025 => x"3d",
          5026 => x"05",
          5027 => x"05",
          5028 => x"71",
          5029 => x"90",
          5030 => x"2b",
          5031 => x"83",
          5032 => x"70",
          5033 => x"33",
          5034 => x"07",
          5035 => x"ae",
          5036 => x"81",
          5037 => x"07",
          5038 => x"53",
          5039 => x"54",
          5040 => x"53",
          5041 => x"77",
          5042 => x"18",
          5043 => x"90",
          5044 => x"88",
          5045 => x"70",
          5046 => x"74",
          5047 => x"82",
          5048 => x"70",
          5049 => x"81",
          5050 => x"88",
          5051 => x"83",
          5052 => x"f8",
          5053 => x"56",
          5054 => x"73",
          5055 => x"06",
          5056 => x"54",
          5057 => x"82",
          5058 => x"81",
          5059 => x"72",
          5060 => x"82",
          5061 => x"16",
          5062 => x"34",
          5063 => x"34",
          5064 => x"04",
          5065 => x"82",
          5066 => x"02",
          5067 => x"05",
          5068 => x"2b",
          5069 => x"11",
          5070 => x"33",
          5071 => x"71",
          5072 => x"58",
          5073 => x"55",
          5074 => x"84",
          5075 => x"13",
          5076 => x"2b",
          5077 => x"2a",
          5078 => x"52",
          5079 => x"34",
          5080 => x"34",
          5081 => x"08",
          5082 => x"11",
          5083 => x"33",
          5084 => x"71",
          5085 => x"56",
          5086 => x"72",
          5087 => x"33",
          5088 => x"71",
          5089 => x"70",
          5090 => x"56",
          5091 => x"86",
          5092 => x"87",
          5093 => x"bb",
          5094 => x"70",
          5095 => x"33",
          5096 => x"07",
          5097 => x"ff",
          5098 => x"2a",
          5099 => x"53",
          5100 => x"34",
          5101 => x"34",
          5102 => x"04",
          5103 => x"02",
          5104 => x"82",
          5105 => x"71",
          5106 => x"11",
          5107 => x"12",
          5108 => x"2b",
          5109 => x"29",
          5110 => x"81",
          5111 => x"98",
          5112 => x"2b",
          5113 => x"53",
          5114 => x"56",
          5115 => x"71",
          5116 => x"f6",
          5117 => x"fe",
          5118 => x"bb",
          5119 => x"16",
          5120 => x"12",
          5121 => x"2b",
          5122 => x"07",
          5123 => x"33",
          5124 => x"71",
          5125 => x"70",
          5126 => x"ff",
          5127 => x"52",
          5128 => x"5a",
          5129 => x"05",
          5130 => x"54",
          5131 => x"13",
          5132 => x"13",
          5133 => x"90",
          5134 => x"70",
          5135 => x"33",
          5136 => x"71",
          5137 => x"56",
          5138 => x"72",
          5139 => x"81",
          5140 => x"88",
          5141 => x"81",
          5142 => x"70",
          5143 => x"51",
          5144 => x"72",
          5145 => x"81",
          5146 => x"3d",
          5147 => x"3d",
          5148 => x"90",
          5149 => x"05",
          5150 => x"70",
          5151 => x"11",
          5152 => x"83",
          5153 => x"8b",
          5154 => x"2b",
          5155 => x"59",
          5156 => x"73",
          5157 => x"81",
          5158 => x"88",
          5159 => x"8c",
          5160 => x"22",
          5161 => x"88",
          5162 => x"53",
          5163 => x"73",
          5164 => x"14",
          5165 => x"90",
          5166 => x"70",
          5167 => x"33",
          5168 => x"71",
          5169 => x"56",
          5170 => x"72",
          5171 => x"33",
          5172 => x"71",
          5173 => x"70",
          5174 => x"55",
          5175 => x"82",
          5176 => x"83",
          5177 => x"bb",
          5178 => x"82",
          5179 => x"12",
          5180 => x"2b",
          5181 => x"98",
          5182 => x"87",
          5183 => x"f7",
          5184 => x"82",
          5185 => x"31",
          5186 => x"83",
          5187 => x"70",
          5188 => x"fd",
          5189 => x"bb",
          5190 => x"83",
          5191 => x"82",
          5192 => x"12",
          5193 => x"2b",
          5194 => x"07",
          5195 => x"33",
          5196 => x"71",
          5197 => x"90",
          5198 => x"42",
          5199 => x"5b",
          5200 => x"54",
          5201 => x"8d",
          5202 => x"80",
          5203 => x"fe",
          5204 => x"84",
          5205 => x"33",
          5206 => x"71",
          5207 => x"83",
          5208 => x"11",
          5209 => x"53",
          5210 => x"55",
          5211 => x"34",
          5212 => x"06",
          5213 => x"14",
          5214 => x"90",
          5215 => x"84",
          5216 => x"13",
          5217 => x"2b",
          5218 => x"2a",
          5219 => x"56",
          5220 => x"16",
          5221 => x"16",
          5222 => x"90",
          5223 => x"80",
          5224 => x"34",
          5225 => x"14",
          5226 => x"90",
          5227 => x"84",
          5228 => x"85",
          5229 => x"bb",
          5230 => x"70",
          5231 => x"33",
          5232 => x"07",
          5233 => x"80",
          5234 => x"2a",
          5235 => x"56",
          5236 => x"34",
          5237 => x"34",
          5238 => x"04",
          5239 => x"73",
          5240 => x"90",
          5241 => x"f7",
          5242 => x"80",
          5243 => x"71",
          5244 => x"3f",
          5245 => x"04",
          5246 => x"80",
          5247 => x"f8",
          5248 => x"bb",
          5249 => x"ff",
          5250 => x"bb",
          5251 => x"11",
          5252 => x"33",
          5253 => x"07",
          5254 => x"56",
          5255 => x"ff",
          5256 => x"78",
          5257 => x"38",
          5258 => x"17",
          5259 => x"12",
          5260 => x"2b",
          5261 => x"ff",
          5262 => x"31",
          5263 => x"ff",
          5264 => x"27",
          5265 => x"56",
          5266 => x"79",
          5267 => x"73",
          5268 => x"38",
          5269 => x"5b",
          5270 => x"85",
          5271 => x"88",
          5272 => x"54",
          5273 => x"78",
          5274 => x"2e",
          5275 => x"79",
          5276 => x"76",
          5277 => x"bb",
          5278 => x"70",
          5279 => x"33",
          5280 => x"07",
          5281 => x"ff",
          5282 => x"5a",
          5283 => x"73",
          5284 => x"38",
          5285 => x"54",
          5286 => x"81",
          5287 => x"54",
          5288 => x"81",
          5289 => x"7a",
          5290 => x"06",
          5291 => x"51",
          5292 => x"81",
          5293 => x"80",
          5294 => x"52",
          5295 => x"c6",
          5296 => x"90",
          5297 => x"86",
          5298 => x"12",
          5299 => x"2b",
          5300 => x"07",
          5301 => x"55",
          5302 => x"17",
          5303 => x"ff",
          5304 => x"2a",
          5305 => x"54",
          5306 => x"34",
          5307 => x"06",
          5308 => x"15",
          5309 => x"90",
          5310 => x"2b",
          5311 => x"1e",
          5312 => x"87",
          5313 => x"88",
          5314 => x"88",
          5315 => x"5e",
          5316 => x"54",
          5317 => x"34",
          5318 => x"34",
          5319 => x"08",
          5320 => x"11",
          5321 => x"33",
          5322 => x"71",
          5323 => x"53",
          5324 => x"74",
          5325 => x"86",
          5326 => x"87",
          5327 => x"bb",
          5328 => x"16",
          5329 => x"11",
          5330 => x"33",
          5331 => x"07",
          5332 => x"53",
          5333 => x"56",
          5334 => x"16",
          5335 => x"16",
          5336 => x"90",
          5337 => x"05",
          5338 => x"bb",
          5339 => x"3d",
          5340 => x"3d",
          5341 => x"82",
          5342 => x"84",
          5343 => x"3f",
          5344 => x"80",
          5345 => x"71",
          5346 => x"3f",
          5347 => x"08",
          5348 => x"bb",
          5349 => x"3d",
          5350 => x"3d",
          5351 => x"40",
          5352 => x"42",
          5353 => x"90",
          5354 => x"09",
          5355 => x"38",
          5356 => x"7b",
          5357 => x"51",
          5358 => x"82",
          5359 => x"54",
          5360 => x"7e",
          5361 => x"51",
          5362 => x"7e",
          5363 => x"39",
          5364 => x"8f",
          5365 => x"98",
          5366 => x"ff",
          5367 => x"90",
          5368 => x"31",
          5369 => x"83",
          5370 => x"70",
          5371 => x"11",
          5372 => x"12",
          5373 => x"2b",
          5374 => x"31",
          5375 => x"ff",
          5376 => x"29",
          5377 => x"88",
          5378 => x"33",
          5379 => x"71",
          5380 => x"70",
          5381 => x"44",
          5382 => x"41",
          5383 => x"5b",
          5384 => x"5b",
          5385 => x"25",
          5386 => x"81",
          5387 => x"75",
          5388 => x"ff",
          5389 => x"54",
          5390 => x"83",
          5391 => x"88",
          5392 => x"88",
          5393 => x"33",
          5394 => x"71",
          5395 => x"90",
          5396 => x"47",
          5397 => x"54",
          5398 => x"8b",
          5399 => x"31",
          5400 => x"ff",
          5401 => x"77",
          5402 => x"fe",
          5403 => x"54",
          5404 => x"09",
          5405 => x"38",
          5406 => x"c0",
          5407 => x"ff",
          5408 => x"81",
          5409 => x"8e",
          5410 => x"24",
          5411 => x"51",
          5412 => x"81",
          5413 => x"18",
          5414 => x"24",
          5415 => x"79",
          5416 => x"33",
          5417 => x"71",
          5418 => x"53",
          5419 => x"f4",
          5420 => x"78",
          5421 => x"3f",
          5422 => x"08",
          5423 => x"06",
          5424 => x"53",
          5425 => x"82",
          5426 => x"11",
          5427 => x"55",
          5428 => x"e7",
          5429 => x"90",
          5430 => x"05",
          5431 => x"ff",
          5432 => x"81",
          5433 => x"15",
          5434 => x"24",
          5435 => x"78",
          5436 => x"3f",
          5437 => x"08",
          5438 => x"33",
          5439 => x"71",
          5440 => x"53",
          5441 => x"9c",
          5442 => x"78",
          5443 => x"3f",
          5444 => x"08",
          5445 => x"06",
          5446 => x"53",
          5447 => x"82",
          5448 => x"11",
          5449 => x"55",
          5450 => x"8f",
          5451 => x"90",
          5452 => x"05",
          5453 => x"19",
          5454 => x"83",
          5455 => x"58",
          5456 => x"7f",
          5457 => x"b0",
          5458 => x"98",
          5459 => x"bb",
          5460 => x"2e",
          5461 => x"53",
          5462 => x"bb",
          5463 => x"ff",
          5464 => x"73",
          5465 => x"3f",
          5466 => x"78",
          5467 => x"80",
          5468 => x"78",
          5469 => x"3f",
          5470 => x"2b",
          5471 => x"08",
          5472 => x"51",
          5473 => x"7b",
          5474 => x"bb",
          5475 => x"3d",
          5476 => x"3d",
          5477 => x"29",
          5478 => x"fb",
          5479 => x"bb",
          5480 => x"82",
          5481 => x"80",
          5482 => x"73",
          5483 => x"82",
          5484 => x"51",
          5485 => x"3f",
          5486 => x"98",
          5487 => x"0d",
          5488 => x"0d",
          5489 => x"33",
          5490 => x"70",
          5491 => x"38",
          5492 => x"11",
          5493 => x"82",
          5494 => x"83",
          5495 => x"fc",
          5496 => x"9b",
          5497 => x"84",
          5498 => x"33",
          5499 => x"51",
          5500 => x"80",
          5501 => x"84",
          5502 => x"92",
          5503 => x"51",
          5504 => x"80",
          5505 => x"81",
          5506 => x"72",
          5507 => x"92",
          5508 => x"81",
          5509 => x"0b",
          5510 => x"8c",
          5511 => x"71",
          5512 => x"06",
          5513 => x"80",
          5514 => x"87",
          5515 => x"08",
          5516 => x"38",
          5517 => x"80",
          5518 => x"71",
          5519 => x"c0",
          5520 => x"51",
          5521 => x"87",
          5522 => x"bb",
          5523 => x"82",
          5524 => x"33",
          5525 => x"bb",
          5526 => x"3d",
          5527 => x"3d",
          5528 => x"64",
          5529 => x"bf",
          5530 => x"40",
          5531 => x"74",
          5532 => x"cd",
          5533 => x"98",
          5534 => x"7a",
          5535 => x"81",
          5536 => x"72",
          5537 => x"87",
          5538 => x"11",
          5539 => x"8c",
          5540 => x"92",
          5541 => x"5a",
          5542 => x"58",
          5543 => x"c0",
          5544 => x"76",
          5545 => x"76",
          5546 => x"70",
          5547 => x"81",
          5548 => x"54",
          5549 => x"8e",
          5550 => x"52",
          5551 => x"81",
          5552 => x"81",
          5553 => x"74",
          5554 => x"53",
          5555 => x"83",
          5556 => x"78",
          5557 => x"8f",
          5558 => x"2e",
          5559 => x"c0",
          5560 => x"52",
          5561 => x"87",
          5562 => x"08",
          5563 => x"2e",
          5564 => x"84",
          5565 => x"38",
          5566 => x"87",
          5567 => x"15",
          5568 => x"70",
          5569 => x"52",
          5570 => x"ff",
          5571 => x"39",
          5572 => x"81",
          5573 => x"ff",
          5574 => x"57",
          5575 => x"90",
          5576 => x"80",
          5577 => x"71",
          5578 => x"78",
          5579 => x"38",
          5580 => x"80",
          5581 => x"80",
          5582 => x"81",
          5583 => x"72",
          5584 => x"0c",
          5585 => x"04",
          5586 => x"60",
          5587 => x"8c",
          5588 => x"33",
          5589 => x"5b",
          5590 => x"74",
          5591 => x"e1",
          5592 => x"98",
          5593 => x"79",
          5594 => x"78",
          5595 => x"06",
          5596 => x"77",
          5597 => x"87",
          5598 => x"11",
          5599 => x"8c",
          5600 => x"92",
          5601 => x"59",
          5602 => x"85",
          5603 => x"98",
          5604 => x"7d",
          5605 => x"0c",
          5606 => x"08",
          5607 => x"70",
          5608 => x"53",
          5609 => x"2e",
          5610 => x"70",
          5611 => x"33",
          5612 => x"18",
          5613 => x"2a",
          5614 => x"51",
          5615 => x"2e",
          5616 => x"c0",
          5617 => x"52",
          5618 => x"87",
          5619 => x"08",
          5620 => x"2e",
          5621 => x"84",
          5622 => x"38",
          5623 => x"87",
          5624 => x"15",
          5625 => x"70",
          5626 => x"52",
          5627 => x"ff",
          5628 => x"39",
          5629 => x"81",
          5630 => x"80",
          5631 => x"52",
          5632 => x"90",
          5633 => x"80",
          5634 => x"71",
          5635 => x"7a",
          5636 => x"38",
          5637 => x"80",
          5638 => x"80",
          5639 => x"81",
          5640 => x"72",
          5641 => x"0c",
          5642 => x"04",
          5643 => x"7a",
          5644 => x"a3",
          5645 => x"88",
          5646 => x"33",
          5647 => x"56",
          5648 => x"3f",
          5649 => x"08",
          5650 => x"83",
          5651 => x"fe",
          5652 => x"87",
          5653 => x"0c",
          5654 => x"76",
          5655 => x"38",
          5656 => x"93",
          5657 => x"2b",
          5658 => x"8c",
          5659 => x"71",
          5660 => x"38",
          5661 => x"71",
          5662 => x"c6",
          5663 => x"39",
          5664 => x"81",
          5665 => x"06",
          5666 => x"71",
          5667 => x"38",
          5668 => x"8c",
          5669 => x"e8",
          5670 => x"98",
          5671 => x"71",
          5672 => x"73",
          5673 => x"92",
          5674 => x"72",
          5675 => x"06",
          5676 => x"f7",
          5677 => x"80",
          5678 => x"88",
          5679 => x"0c",
          5680 => x"80",
          5681 => x"56",
          5682 => x"56",
          5683 => x"82",
          5684 => x"88",
          5685 => x"fe",
          5686 => x"81",
          5687 => x"33",
          5688 => x"07",
          5689 => x"0c",
          5690 => x"3d",
          5691 => x"3d",
          5692 => x"11",
          5693 => x"33",
          5694 => x"71",
          5695 => x"81",
          5696 => x"72",
          5697 => x"75",
          5698 => x"82",
          5699 => x"52",
          5700 => x"54",
          5701 => x"0d",
          5702 => x"0d",
          5703 => x"05",
          5704 => x"52",
          5705 => x"70",
          5706 => x"34",
          5707 => x"51",
          5708 => x"83",
          5709 => x"ff",
          5710 => x"75",
          5711 => x"72",
          5712 => x"54",
          5713 => x"2a",
          5714 => x"70",
          5715 => x"34",
          5716 => x"51",
          5717 => x"81",
          5718 => x"70",
          5719 => x"70",
          5720 => x"3d",
          5721 => x"3d",
          5722 => x"77",
          5723 => x"70",
          5724 => x"38",
          5725 => x"05",
          5726 => x"70",
          5727 => x"34",
          5728 => x"eb",
          5729 => x"0d",
          5730 => x"0d",
          5731 => x"54",
          5732 => x"72",
          5733 => x"54",
          5734 => x"51",
          5735 => x"84",
          5736 => x"fc",
          5737 => x"77",
          5738 => x"53",
          5739 => x"05",
          5740 => x"70",
          5741 => x"33",
          5742 => x"ff",
          5743 => x"52",
          5744 => x"2e",
          5745 => x"80",
          5746 => x"71",
          5747 => x"0c",
          5748 => x"04",
          5749 => x"74",
          5750 => x"89",
          5751 => x"2e",
          5752 => x"11",
          5753 => x"52",
          5754 => x"70",
          5755 => x"98",
          5756 => x"0d",
          5757 => x"82",
          5758 => x"04",
          5759 => x"bb",
          5760 => x"f7",
          5761 => x"56",
          5762 => x"17",
          5763 => x"74",
          5764 => x"d6",
          5765 => x"b0",
          5766 => x"b4",
          5767 => x"81",
          5768 => x"59",
          5769 => x"82",
          5770 => x"7a",
          5771 => x"06",
          5772 => x"bb",
          5773 => x"17",
          5774 => x"08",
          5775 => x"08",
          5776 => x"08",
          5777 => x"74",
          5778 => x"38",
          5779 => x"55",
          5780 => x"09",
          5781 => x"38",
          5782 => x"18",
          5783 => x"81",
          5784 => x"f9",
          5785 => x"39",
          5786 => x"82",
          5787 => x"8b",
          5788 => x"fa",
          5789 => x"7a",
          5790 => x"57",
          5791 => x"08",
          5792 => x"75",
          5793 => x"3f",
          5794 => x"08",
          5795 => x"98",
          5796 => x"81",
          5797 => x"b4",
          5798 => x"16",
          5799 => x"be",
          5800 => x"98",
          5801 => x"85",
          5802 => x"81",
          5803 => x"17",
          5804 => x"bb",
          5805 => x"3d",
          5806 => x"3d",
          5807 => x"52",
          5808 => x"3f",
          5809 => x"08",
          5810 => x"98",
          5811 => x"38",
          5812 => x"74",
          5813 => x"81",
          5814 => x"38",
          5815 => x"59",
          5816 => x"09",
          5817 => x"e3",
          5818 => x"53",
          5819 => x"08",
          5820 => x"70",
          5821 => x"91",
          5822 => x"d5",
          5823 => x"17",
          5824 => x"3f",
          5825 => x"a4",
          5826 => x"51",
          5827 => x"86",
          5828 => x"f2",
          5829 => x"17",
          5830 => x"3f",
          5831 => x"52",
          5832 => x"51",
          5833 => x"8c",
          5834 => x"84",
          5835 => x"fc",
          5836 => x"17",
          5837 => x"70",
          5838 => x"79",
          5839 => x"52",
          5840 => x"51",
          5841 => x"77",
          5842 => x"80",
          5843 => x"81",
          5844 => x"f9",
          5845 => x"bb",
          5846 => x"2e",
          5847 => x"58",
          5848 => x"98",
          5849 => x"0d",
          5850 => x"0d",
          5851 => x"98",
          5852 => x"05",
          5853 => x"80",
          5854 => x"27",
          5855 => x"14",
          5856 => x"29",
          5857 => x"05",
          5858 => x"82",
          5859 => x"87",
          5860 => x"f9",
          5861 => x"7a",
          5862 => x"54",
          5863 => x"27",
          5864 => x"76",
          5865 => x"27",
          5866 => x"ff",
          5867 => x"58",
          5868 => x"80",
          5869 => x"82",
          5870 => x"72",
          5871 => x"38",
          5872 => x"72",
          5873 => x"8e",
          5874 => x"39",
          5875 => x"17",
          5876 => x"a4",
          5877 => x"53",
          5878 => x"fd",
          5879 => x"bb",
          5880 => x"9f",
          5881 => x"ff",
          5882 => x"11",
          5883 => x"70",
          5884 => x"18",
          5885 => x"76",
          5886 => x"53",
          5887 => x"82",
          5888 => x"80",
          5889 => x"83",
          5890 => x"b4",
          5891 => x"88",
          5892 => x"79",
          5893 => x"84",
          5894 => x"58",
          5895 => x"80",
          5896 => x"9f",
          5897 => x"80",
          5898 => x"88",
          5899 => x"08",
          5900 => x"51",
          5901 => x"82",
          5902 => x"80",
          5903 => x"10",
          5904 => x"74",
          5905 => x"51",
          5906 => x"82",
          5907 => x"83",
          5908 => x"58",
          5909 => x"87",
          5910 => x"08",
          5911 => x"51",
          5912 => x"82",
          5913 => x"9b",
          5914 => x"2b",
          5915 => x"74",
          5916 => x"51",
          5917 => x"82",
          5918 => x"f0",
          5919 => x"83",
          5920 => x"77",
          5921 => x"0c",
          5922 => x"04",
          5923 => x"7a",
          5924 => x"58",
          5925 => x"81",
          5926 => x"9e",
          5927 => x"17",
          5928 => x"96",
          5929 => x"53",
          5930 => x"81",
          5931 => x"79",
          5932 => x"72",
          5933 => x"38",
          5934 => x"72",
          5935 => x"b8",
          5936 => x"39",
          5937 => x"17",
          5938 => x"a4",
          5939 => x"53",
          5940 => x"fb",
          5941 => x"bb",
          5942 => x"82",
          5943 => x"81",
          5944 => x"83",
          5945 => x"b4",
          5946 => x"78",
          5947 => x"56",
          5948 => x"76",
          5949 => x"38",
          5950 => x"9f",
          5951 => x"33",
          5952 => x"07",
          5953 => x"74",
          5954 => x"83",
          5955 => x"89",
          5956 => x"08",
          5957 => x"51",
          5958 => x"82",
          5959 => x"59",
          5960 => x"08",
          5961 => x"74",
          5962 => x"16",
          5963 => x"84",
          5964 => x"76",
          5965 => x"88",
          5966 => x"81",
          5967 => x"8f",
          5968 => x"53",
          5969 => x"80",
          5970 => x"88",
          5971 => x"08",
          5972 => x"51",
          5973 => x"82",
          5974 => x"59",
          5975 => x"08",
          5976 => x"77",
          5977 => x"06",
          5978 => x"83",
          5979 => x"05",
          5980 => x"f7",
          5981 => x"39",
          5982 => x"a4",
          5983 => x"52",
          5984 => x"ef",
          5985 => x"98",
          5986 => x"bb",
          5987 => x"38",
          5988 => x"06",
          5989 => x"83",
          5990 => x"18",
          5991 => x"54",
          5992 => x"f6",
          5993 => x"bb",
          5994 => x"0a",
          5995 => x"52",
          5996 => x"83",
          5997 => x"83",
          5998 => x"82",
          5999 => x"8a",
          6000 => x"f8",
          6001 => x"7c",
          6002 => x"59",
          6003 => x"81",
          6004 => x"38",
          6005 => x"08",
          6006 => x"73",
          6007 => x"38",
          6008 => x"52",
          6009 => x"a4",
          6010 => x"98",
          6011 => x"bb",
          6012 => x"f2",
          6013 => x"82",
          6014 => x"39",
          6015 => x"e6",
          6016 => x"98",
          6017 => x"de",
          6018 => x"78",
          6019 => x"3f",
          6020 => x"08",
          6021 => x"98",
          6022 => x"80",
          6023 => x"bb",
          6024 => x"2e",
          6025 => x"bb",
          6026 => x"2e",
          6027 => x"53",
          6028 => x"51",
          6029 => x"82",
          6030 => x"c5",
          6031 => x"08",
          6032 => x"18",
          6033 => x"57",
          6034 => x"90",
          6035 => x"90",
          6036 => x"16",
          6037 => x"54",
          6038 => x"34",
          6039 => x"78",
          6040 => x"38",
          6041 => x"82",
          6042 => x"8a",
          6043 => x"f6",
          6044 => x"7e",
          6045 => x"5b",
          6046 => x"38",
          6047 => x"58",
          6048 => x"88",
          6049 => x"08",
          6050 => x"38",
          6051 => x"39",
          6052 => x"51",
          6053 => x"81",
          6054 => x"bb",
          6055 => x"82",
          6056 => x"bb",
          6057 => x"82",
          6058 => x"ff",
          6059 => x"38",
          6060 => x"82",
          6061 => x"26",
          6062 => x"79",
          6063 => x"08",
          6064 => x"73",
          6065 => x"b9",
          6066 => x"2e",
          6067 => x"80",
          6068 => x"1a",
          6069 => x"08",
          6070 => x"38",
          6071 => x"52",
          6072 => x"af",
          6073 => x"82",
          6074 => x"81",
          6075 => x"06",
          6076 => x"bb",
          6077 => x"82",
          6078 => x"09",
          6079 => x"72",
          6080 => x"70",
          6081 => x"bb",
          6082 => x"51",
          6083 => x"73",
          6084 => x"82",
          6085 => x"80",
          6086 => x"8c",
          6087 => x"81",
          6088 => x"38",
          6089 => x"08",
          6090 => x"73",
          6091 => x"75",
          6092 => x"77",
          6093 => x"56",
          6094 => x"76",
          6095 => x"82",
          6096 => x"26",
          6097 => x"75",
          6098 => x"f8",
          6099 => x"bb",
          6100 => x"2e",
          6101 => x"59",
          6102 => x"08",
          6103 => x"81",
          6104 => x"82",
          6105 => x"59",
          6106 => x"08",
          6107 => x"70",
          6108 => x"25",
          6109 => x"51",
          6110 => x"73",
          6111 => x"75",
          6112 => x"81",
          6113 => x"38",
          6114 => x"f5",
          6115 => x"75",
          6116 => x"f9",
          6117 => x"bb",
          6118 => x"bb",
          6119 => x"70",
          6120 => x"08",
          6121 => x"51",
          6122 => x"80",
          6123 => x"73",
          6124 => x"38",
          6125 => x"52",
          6126 => x"d0",
          6127 => x"98",
          6128 => x"a5",
          6129 => x"18",
          6130 => x"08",
          6131 => x"18",
          6132 => x"74",
          6133 => x"38",
          6134 => x"18",
          6135 => x"33",
          6136 => x"73",
          6137 => x"97",
          6138 => x"74",
          6139 => x"38",
          6140 => x"55",
          6141 => x"bb",
          6142 => x"85",
          6143 => x"75",
          6144 => x"bb",
          6145 => x"3d",
          6146 => x"3d",
          6147 => x"52",
          6148 => x"3f",
          6149 => x"08",
          6150 => x"82",
          6151 => x"80",
          6152 => x"52",
          6153 => x"c1",
          6154 => x"98",
          6155 => x"98",
          6156 => x"0c",
          6157 => x"53",
          6158 => x"15",
          6159 => x"f2",
          6160 => x"56",
          6161 => x"16",
          6162 => x"22",
          6163 => x"27",
          6164 => x"54",
          6165 => x"76",
          6166 => x"33",
          6167 => x"3f",
          6168 => x"08",
          6169 => x"38",
          6170 => x"76",
          6171 => x"70",
          6172 => x"9f",
          6173 => x"56",
          6174 => x"bb",
          6175 => x"3d",
          6176 => x"3d",
          6177 => x"71",
          6178 => x"57",
          6179 => x"0a",
          6180 => x"38",
          6181 => x"53",
          6182 => x"38",
          6183 => x"0c",
          6184 => x"54",
          6185 => x"75",
          6186 => x"73",
          6187 => x"a8",
          6188 => x"73",
          6189 => x"85",
          6190 => x"0b",
          6191 => x"5a",
          6192 => x"27",
          6193 => x"a8",
          6194 => x"18",
          6195 => x"39",
          6196 => x"70",
          6197 => x"58",
          6198 => x"b2",
          6199 => x"76",
          6200 => x"3f",
          6201 => x"08",
          6202 => x"98",
          6203 => x"bd",
          6204 => x"82",
          6205 => x"27",
          6206 => x"16",
          6207 => x"98",
          6208 => x"38",
          6209 => x"39",
          6210 => x"55",
          6211 => x"52",
          6212 => x"d5",
          6213 => x"98",
          6214 => x"0c",
          6215 => x"0c",
          6216 => x"53",
          6217 => x"80",
          6218 => x"85",
          6219 => x"94",
          6220 => x"2a",
          6221 => x"0c",
          6222 => x"06",
          6223 => x"9c",
          6224 => x"58",
          6225 => x"98",
          6226 => x"0d",
          6227 => x"0d",
          6228 => x"90",
          6229 => x"05",
          6230 => x"f0",
          6231 => x"27",
          6232 => x"0b",
          6233 => x"98",
          6234 => x"84",
          6235 => x"2e",
          6236 => x"76",
          6237 => x"58",
          6238 => x"38",
          6239 => x"15",
          6240 => x"08",
          6241 => x"38",
          6242 => x"88",
          6243 => x"53",
          6244 => x"81",
          6245 => x"c0",
          6246 => x"22",
          6247 => x"89",
          6248 => x"72",
          6249 => x"74",
          6250 => x"f3",
          6251 => x"bb",
          6252 => x"82",
          6253 => x"82",
          6254 => x"27",
          6255 => x"81",
          6256 => x"98",
          6257 => x"80",
          6258 => x"16",
          6259 => x"98",
          6260 => x"ca",
          6261 => x"38",
          6262 => x"0c",
          6263 => x"dd",
          6264 => x"08",
          6265 => x"f9",
          6266 => x"bb",
          6267 => x"87",
          6268 => x"98",
          6269 => x"80",
          6270 => x"55",
          6271 => x"08",
          6272 => x"38",
          6273 => x"bb",
          6274 => x"2e",
          6275 => x"bb",
          6276 => x"75",
          6277 => x"3f",
          6278 => x"08",
          6279 => x"94",
          6280 => x"52",
          6281 => x"c1",
          6282 => x"98",
          6283 => x"0c",
          6284 => x"0c",
          6285 => x"05",
          6286 => x"80",
          6287 => x"bb",
          6288 => x"3d",
          6289 => x"3d",
          6290 => x"71",
          6291 => x"57",
          6292 => x"51",
          6293 => x"82",
          6294 => x"54",
          6295 => x"08",
          6296 => x"82",
          6297 => x"56",
          6298 => x"52",
          6299 => x"83",
          6300 => x"98",
          6301 => x"bb",
          6302 => x"d2",
          6303 => x"98",
          6304 => x"08",
          6305 => x"54",
          6306 => x"e5",
          6307 => x"06",
          6308 => x"58",
          6309 => x"08",
          6310 => x"38",
          6311 => x"75",
          6312 => x"80",
          6313 => x"81",
          6314 => x"7a",
          6315 => x"06",
          6316 => x"39",
          6317 => x"08",
          6318 => x"76",
          6319 => x"3f",
          6320 => x"08",
          6321 => x"98",
          6322 => x"ff",
          6323 => x"84",
          6324 => x"06",
          6325 => x"54",
          6326 => x"98",
          6327 => x"0d",
          6328 => x"0d",
          6329 => x"52",
          6330 => x"3f",
          6331 => x"08",
          6332 => x"06",
          6333 => x"51",
          6334 => x"83",
          6335 => x"06",
          6336 => x"14",
          6337 => x"3f",
          6338 => x"08",
          6339 => x"07",
          6340 => x"bb",
          6341 => x"3d",
          6342 => x"3d",
          6343 => x"70",
          6344 => x"06",
          6345 => x"53",
          6346 => x"ed",
          6347 => x"33",
          6348 => x"83",
          6349 => x"06",
          6350 => x"90",
          6351 => x"15",
          6352 => x"3f",
          6353 => x"04",
          6354 => x"7b",
          6355 => x"84",
          6356 => x"58",
          6357 => x"80",
          6358 => x"38",
          6359 => x"52",
          6360 => x"8f",
          6361 => x"98",
          6362 => x"bb",
          6363 => x"f5",
          6364 => x"08",
          6365 => x"53",
          6366 => x"84",
          6367 => x"39",
          6368 => x"70",
          6369 => x"81",
          6370 => x"51",
          6371 => x"16",
          6372 => x"98",
          6373 => x"81",
          6374 => x"38",
          6375 => x"ae",
          6376 => x"81",
          6377 => x"54",
          6378 => x"2e",
          6379 => x"8f",
          6380 => x"82",
          6381 => x"76",
          6382 => x"54",
          6383 => x"09",
          6384 => x"38",
          6385 => x"7a",
          6386 => x"80",
          6387 => x"fa",
          6388 => x"bb",
          6389 => x"82",
          6390 => x"89",
          6391 => x"08",
          6392 => x"86",
          6393 => x"98",
          6394 => x"82",
          6395 => x"8b",
          6396 => x"fb",
          6397 => x"70",
          6398 => x"81",
          6399 => x"fc",
          6400 => x"bb",
          6401 => x"82",
          6402 => x"b4",
          6403 => x"08",
          6404 => x"ec",
          6405 => x"bb",
          6406 => x"82",
          6407 => x"a0",
          6408 => x"82",
          6409 => x"52",
          6410 => x"51",
          6411 => x"8b",
          6412 => x"52",
          6413 => x"51",
          6414 => x"81",
          6415 => x"34",
          6416 => x"98",
          6417 => x"0d",
          6418 => x"0d",
          6419 => x"98",
          6420 => x"70",
          6421 => x"ec",
          6422 => x"bb",
          6423 => x"38",
          6424 => x"53",
          6425 => x"81",
          6426 => x"34",
          6427 => x"04",
          6428 => x"78",
          6429 => x"80",
          6430 => x"34",
          6431 => x"80",
          6432 => x"38",
          6433 => x"18",
          6434 => x"9c",
          6435 => x"70",
          6436 => x"56",
          6437 => x"a0",
          6438 => x"71",
          6439 => x"81",
          6440 => x"81",
          6441 => x"89",
          6442 => x"06",
          6443 => x"73",
          6444 => x"55",
          6445 => x"55",
          6446 => x"81",
          6447 => x"81",
          6448 => x"74",
          6449 => x"75",
          6450 => x"52",
          6451 => x"13",
          6452 => x"08",
          6453 => x"33",
          6454 => x"9c",
          6455 => x"11",
          6456 => x"8a",
          6457 => x"98",
          6458 => x"96",
          6459 => x"e7",
          6460 => x"98",
          6461 => x"23",
          6462 => x"e7",
          6463 => x"bb",
          6464 => x"17",
          6465 => x"0d",
          6466 => x"0d",
          6467 => x"5e",
          6468 => x"70",
          6469 => x"55",
          6470 => x"83",
          6471 => x"73",
          6472 => x"91",
          6473 => x"2e",
          6474 => x"1d",
          6475 => x"0c",
          6476 => x"15",
          6477 => x"70",
          6478 => x"56",
          6479 => x"09",
          6480 => x"38",
          6481 => x"80",
          6482 => x"30",
          6483 => x"78",
          6484 => x"54",
          6485 => x"73",
          6486 => x"60",
          6487 => x"54",
          6488 => x"96",
          6489 => x"0b",
          6490 => x"80",
          6491 => x"f6",
          6492 => x"bb",
          6493 => x"85",
          6494 => x"3d",
          6495 => x"5c",
          6496 => x"53",
          6497 => x"51",
          6498 => x"80",
          6499 => x"88",
          6500 => x"5c",
          6501 => x"09",
          6502 => x"d4",
          6503 => x"70",
          6504 => x"71",
          6505 => x"30",
          6506 => x"73",
          6507 => x"51",
          6508 => x"57",
          6509 => x"38",
          6510 => x"75",
          6511 => x"17",
          6512 => x"75",
          6513 => x"30",
          6514 => x"51",
          6515 => x"80",
          6516 => x"38",
          6517 => x"87",
          6518 => x"26",
          6519 => x"77",
          6520 => x"a4",
          6521 => x"27",
          6522 => x"a0",
          6523 => x"39",
          6524 => x"33",
          6525 => x"57",
          6526 => x"27",
          6527 => x"75",
          6528 => x"30",
          6529 => x"32",
          6530 => x"80",
          6531 => x"25",
          6532 => x"56",
          6533 => x"80",
          6534 => x"84",
          6535 => x"58",
          6536 => x"70",
          6537 => x"55",
          6538 => x"09",
          6539 => x"38",
          6540 => x"80",
          6541 => x"30",
          6542 => x"77",
          6543 => x"54",
          6544 => x"81",
          6545 => x"ae",
          6546 => x"06",
          6547 => x"54",
          6548 => x"74",
          6549 => x"80",
          6550 => x"7b",
          6551 => x"30",
          6552 => x"70",
          6553 => x"25",
          6554 => x"07",
          6555 => x"51",
          6556 => x"a7",
          6557 => x"8b",
          6558 => x"39",
          6559 => x"54",
          6560 => x"8c",
          6561 => x"ff",
          6562 => x"e0",
          6563 => x"54",
          6564 => x"e1",
          6565 => x"98",
          6566 => x"b2",
          6567 => x"70",
          6568 => x"71",
          6569 => x"54",
          6570 => x"82",
          6571 => x"80",
          6572 => x"38",
          6573 => x"76",
          6574 => x"df",
          6575 => x"54",
          6576 => x"81",
          6577 => x"55",
          6578 => x"34",
          6579 => x"52",
          6580 => x"51",
          6581 => x"82",
          6582 => x"bf",
          6583 => x"16",
          6584 => x"26",
          6585 => x"16",
          6586 => x"06",
          6587 => x"17",
          6588 => x"34",
          6589 => x"fd",
          6590 => x"19",
          6591 => x"80",
          6592 => x"79",
          6593 => x"81",
          6594 => x"81",
          6595 => x"85",
          6596 => x"54",
          6597 => x"8f",
          6598 => x"86",
          6599 => x"39",
          6600 => x"f3",
          6601 => x"73",
          6602 => x"80",
          6603 => x"52",
          6604 => x"ce",
          6605 => x"98",
          6606 => x"bb",
          6607 => x"d7",
          6608 => x"08",
          6609 => x"e6",
          6610 => x"bb",
          6611 => x"82",
          6612 => x"80",
          6613 => x"1b",
          6614 => x"55",
          6615 => x"2e",
          6616 => x"8b",
          6617 => x"06",
          6618 => x"1c",
          6619 => x"33",
          6620 => x"70",
          6621 => x"55",
          6622 => x"38",
          6623 => x"52",
          6624 => x"9f",
          6625 => x"98",
          6626 => x"8b",
          6627 => x"7a",
          6628 => x"3f",
          6629 => x"75",
          6630 => x"57",
          6631 => x"2e",
          6632 => x"84",
          6633 => x"06",
          6634 => x"75",
          6635 => x"81",
          6636 => x"2a",
          6637 => x"73",
          6638 => x"38",
          6639 => x"54",
          6640 => x"fb",
          6641 => x"80",
          6642 => x"34",
          6643 => x"c1",
          6644 => x"06",
          6645 => x"38",
          6646 => x"39",
          6647 => x"70",
          6648 => x"54",
          6649 => x"86",
          6650 => x"84",
          6651 => x"06",
          6652 => x"73",
          6653 => x"38",
          6654 => x"83",
          6655 => x"b4",
          6656 => x"51",
          6657 => x"82",
          6658 => x"88",
          6659 => x"ea",
          6660 => x"bb",
          6661 => x"3d",
          6662 => x"3d",
          6663 => x"ff",
          6664 => x"71",
          6665 => x"5c",
          6666 => x"80",
          6667 => x"38",
          6668 => x"05",
          6669 => x"a0",
          6670 => x"71",
          6671 => x"38",
          6672 => x"71",
          6673 => x"81",
          6674 => x"38",
          6675 => x"11",
          6676 => x"06",
          6677 => x"70",
          6678 => x"38",
          6679 => x"81",
          6680 => x"05",
          6681 => x"76",
          6682 => x"38",
          6683 => x"b4",
          6684 => x"77",
          6685 => x"57",
          6686 => x"05",
          6687 => x"70",
          6688 => x"33",
          6689 => x"53",
          6690 => x"99",
          6691 => x"e0",
          6692 => x"ff",
          6693 => x"ff",
          6694 => x"70",
          6695 => x"38",
          6696 => x"81",
          6697 => x"51",
          6698 => x"9f",
          6699 => x"72",
          6700 => x"81",
          6701 => x"70",
          6702 => x"72",
          6703 => x"32",
          6704 => x"72",
          6705 => x"73",
          6706 => x"53",
          6707 => x"70",
          6708 => x"38",
          6709 => x"19",
          6710 => x"75",
          6711 => x"38",
          6712 => x"83",
          6713 => x"74",
          6714 => x"59",
          6715 => x"39",
          6716 => x"33",
          6717 => x"bb",
          6718 => x"3d",
          6719 => x"3d",
          6720 => x"80",
          6721 => x"34",
          6722 => x"17",
          6723 => x"75",
          6724 => x"3f",
          6725 => x"bb",
          6726 => x"80",
          6727 => x"16",
          6728 => x"3f",
          6729 => x"08",
          6730 => x"06",
          6731 => x"73",
          6732 => x"2e",
          6733 => x"80",
          6734 => x"0b",
          6735 => x"56",
          6736 => x"e9",
          6737 => x"06",
          6738 => x"57",
          6739 => x"32",
          6740 => x"80",
          6741 => x"51",
          6742 => x"8a",
          6743 => x"e8",
          6744 => x"06",
          6745 => x"53",
          6746 => x"52",
          6747 => x"51",
          6748 => x"82",
          6749 => x"55",
          6750 => x"08",
          6751 => x"38",
          6752 => x"b4",
          6753 => x"86",
          6754 => x"97",
          6755 => x"98",
          6756 => x"bb",
          6757 => x"2e",
          6758 => x"55",
          6759 => x"98",
          6760 => x"0d",
          6761 => x"0d",
          6762 => x"05",
          6763 => x"33",
          6764 => x"75",
          6765 => x"fc",
          6766 => x"bb",
          6767 => x"8b",
          6768 => x"82",
          6769 => x"24",
          6770 => x"82",
          6771 => x"84",
          6772 => x"d0",
          6773 => x"55",
          6774 => x"73",
          6775 => x"e6",
          6776 => x"0c",
          6777 => x"06",
          6778 => x"57",
          6779 => x"ae",
          6780 => x"33",
          6781 => x"3f",
          6782 => x"08",
          6783 => x"70",
          6784 => x"55",
          6785 => x"76",
          6786 => x"b8",
          6787 => x"2a",
          6788 => x"51",
          6789 => x"72",
          6790 => x"86",
          6791 => x"74",
          6792 => x"15",
          6793 => x"81",
          6794 => x"d7",
          6795 => x"bb",
          6796 => x"ff",
          6797 => x"06",
          6798 => x"56",
          6799 => x"38",
          6800 => x"8f",
          6801 => x"2a",
          6802 => x"51",
          6803 => x"72",
          6804 => x"80",
          6805 => x"52",
          6806 => x"3f",
          6807 => x"08",
          6808 => x"57",
          6809 => x"09",
          6810 => x"e2",
          6811 => x"74",
          6812 => x"56",
          6813 => x"33",
          6814 => x"72",
          6815 => x"38",
          6816 => x"51",
          6817 => x"82",
          6818 => x"57",
          6819 => x"84",
          6820 => x"ff",
          6821 => x"56",
          6822 => x"25",
          6823 => x"0b",
          6824 => x"56",
          6825 => x"05",
          6826 => x"83",
          6827 => x"2e",
          6828 => x"52",
          6829 => x"c6",
          6830 => x"98",
          6831 => x"06",
          6832 => x"27",
          6833 => x"16",
          6834 => x"27",
          6835 => x"56",
          6836 => x"84",
          6837 => x"56",
          6838 => x"84",
          6839 => x"14",
          6840 => x"3f",
          6841 => x"08",
          6842 => x"06",
          6843 => x"80",
          6844 => x"06",
          6845 => x"80",
          6846 => x"db",
          6847 => x"bb",
          6848 => x"ff",
          6849 => x"77",
          6850 => x"d8",
          6851 => x"de",
          6852 => x"98",
          6853 => x"9c",
          6854 => x"c4",
          6855 => x"15",
          6856 => x"14",
          6857 => x"70",
          6858 => x"51",
          6859 => x"56",
          6860 => x"84",
          6861 => x"81",
          6862 => x"71",
          6863 => x"16",
          6864 => x"53",
          6865 => x"23",
          6866 => x"8b",
          6867 => x"73",
          6868 => x"80",
          6869 => x"8d",
          6870 => x"39",
          6871 => x"51",
          6872 => x"82",
          6873 => x"53",
          6874 => x"08",
          6875 => x"72",
          6876 => x"8d",
          6877 => x"ce",
          6878 => x"14",
          6879 => x"3f",
          6880 => x"08",
          6881 => x"06",
          6882 => x"38",
          6883 => x"51",
          6884 => x"82",
          6885 => x"55",
          6886 => x"51",
          6887 => x"82",
          6888 => x"83",
          6889 => x"53",
          6890 => x"80",
          6891 => x"38",
          6892 => x"78",
          6893 => x"2a",
          6894 => x"78",
          6895 => x"86",
          6896 => x"22",
          6897 => x"31",
          6898 => x"d7",
          6899 => x"98",
          6900 => x"bb",
          6901 => x"2e",
          6902 => x"82",
          6903 => x"80",
          6904 => x"f5",
          6905 => x"83",
          6906 => x"ff",
          6907 => x"38",
          6908 => x"9f",
          6909 => x"38",
          6910 => x"39",
          6911 => x"80",
          6912 => x"38",
          6913 => x"98",
          6914 => x"a0",
          6915 => x"1c",
          6916 => x"0c",
          6917 => x"17",
          6918 => x"76",
          6919 => x"81",
          6920 => x"80",
          6921 => x"d9",
          6922 => x"bb",
          6923 => x"ff",
          6924 => x"8d",
          6925 => x"8e",
          6926 => x"8a",
          6927 => x"14",
          6928 => x"3f",
          6929 => x"08",
          6930 => x"74",
          6931 => x"a2",
          6932 => x"79",
          6933 => x"ee",
          6934 => x"a8",
          6935 => x"15",
          6936 => x"2e",
          6937 => x"10",
          6938 => x"2a",
          6939 => x"05",
          6940 => x"ff",
          6941 => x"53",
          6942 => x"9c",
          6943 => x"81",
          6944 => x"0b",
          6945 => x"ff",
          6946 => x"0c",
          6947 => x"84",
          6948 => x"83",
          6949 => x"06",
          6950 => x"80",
          6951 => x"d8",
          6952 => x"bb",
          6953 => x"ff",
          6954 => x"72",
          6955 => x"81",
          6956 => x"38",
          6957 => x"73",
          6958 => x"3f",
          6959 => x"08",
          6960 => x"82",
          6961 => x"84",
          6962 => x"b2",
          6963 => x"87",
          6964 => x"98",
          6965 => x"ff",
          6966 => x"82",
          6967 => x"09",
          6968 => x"c8",
          6969 => x"51",
          6970 => x"82",
          6971 => x"84",
          6972 => x"d2",
          6973 => x"06",
          6974 => x"98",
          6975 => x"ee",
          6976 => x"98",
          6977 => x"85",
          6978 => x"09",
          6979 => x"38",
          6980 => x"51",
          6981 => x"82",
          6982 => x"90",
          6983 => x"a0",
          6984 => x"ca",
          6985 => x"98",
          6986 => x"0c",
          6987 => x"82",
          6988 => x"81",
          6989 => x"82",
          6990 => x"72",
          6991 => x"80",
          6992 => x"0c",
          6993 => x"82",
          6994 => x"90",
          6995 => x"fb",
          6996 => x"54",
          6997 => x"80",
          6998 => x"73",
          6999 => x"80",
          7000 => x"72",
          7001 => x"80",
          7002 => x"86",
          7003 => x"15",
          7004 => x"71",
          7005 => x"81",
          7006 => x"81",
          7007 => x"d0",
          7008 => x"bb",
          7009 => x"06",
          7010 => x"38",
          7011 => x"54",
          7012 => x"80",
          7013 => x"71",
          7014 => x"82",
          7015 => x"87",
          7016 => x"fa",
          7017 => x"ab",
          7018 => x"58",
          7019 => x"05",
          7020 => x"e6",
          7021 => x"80",
          7022 => x"98",
          7023 => x"38",
          7024 => x"08",
          7025 => x"d2",
          7026 => x"08",
          7027 => x"80",
          7028 => x"80",
          7029 => x"54",
          7030 => x"84",
          7031 => x"34",
          7032 => x"75",
          7033 => x"2e",
          7034 => x"53",
          7035 => x"53",
          7036 => x"f7",
          7037 => x"bb",
          7038 => x"73",
          7039 => x"0c",
          7040 => x"04",
          7041 => x"67",
          7042 => x"80",
          7043 => x"59",
          7044 => x"78",
          7045 => x"c8",
          7046 => x"06",
          7047 => x"3d",
          7048 => x"99",
          7049 => x"52",
          7050 => x"3f",
          7051 => x"08",
          7052 => x"98",
          7053 => x"38",
          7054 => x"52",
          7055 => x"52",
          7056 => x"3f",
          7057 => x"08",
          7058 => x"98",
          7059 => x"02",
          7060 => x"33",
          7061 => x"55",
          7062 => x"25",
          7063 => x"55",
          7064 => x"54",
          7065 => x"81",
          7066 => x"80",
          7067 => x"74",
          7068 => x"81",
          7069 => x"75",
          7070 => x"3f",
          7071 => x"08",
          7072 => x"02",
          7073 => x"91",
          7074 => x"81",
          7075 => x"82",
          7076 => x"06",
          7077 => x"80",
          7078 => x"88",
          7079 => x"39",
          7080 => x"58",
          7081 => x"38",
          7082 => x"70",
          7083 => x"54",
          7084 => x"81",
          7085 => x"52",
          7086 => x"a5",
          7087 => x"98",
          7088 => x"88",
          7089 => x"62",
          7090 => x"d4",
          7091 => x"54",
          7092 => x"15",
          7093 => x"62",
          7094 => x"e8",
          7095 => x"52",
          7096 => x"51",
          7097 => x"7a",
          7098 => x"83",
          7099 => x"80",
          7100 => x"38",
          7101 => x"08",
          7102 => x"53",
          7103 => x"3d",
          7104 => x"dd",
          7105 => x"bb",
          7106 => x"82",
          7107 => x"82",
          7108 => x"39",
          7109 => x"38",
          7110 => x"33",
          7111 => x"70",
          7112 => x"55",
          7113 => x"2e",
          7114 => x"55",
          7115 => x"77",
          7116 => x"81",
          7117 => x"73",
          7118 => x"38",
          7119 => x"54",
          7120 => x"a0",
          7121 => x"82",
          7122 => x"52",
          7123 => x"a3",
          7124 => x"98",
          7125 => x"18",
          7126 => x"55",
          7127 => x"98",
          7128 => x"38",
          7129 => x"70",
          7130 => x"54",
          7131 => x"86",
          7132 => x"c0",
          7133 => x"b0",
          7134 => x"1b",
          7135 => x"1b",
          7136 => x"70",
          7137 => x"d9",
          7138 => x"98",
          7139 => x"98",
          7140 => x"0c",
          7141 => x"52",
          7142 => x"3f",
          7143 => x"08",
          7144 => x"08",
          7145 => x"77",
          7146 => x"86",
          7147 => x"1a",
          7148 => x"1a",
          7149 => x"91",
          7150 => x"0b",
          7151 => x"80",
          7152 => x"0c",
          7153 => x"70",
          7154 => x"54",
          7155 => x"81",
          7156 => x"bb",
          7157 => x"2e",
          7158 => x"82",
          7159 => x"94",
          7160 => x"17",
          7161 => x"2b",
          7162 => x"57",
          7163 => x"52",
          7164 => x"9f",
          7165 => x"98",
          7166 => x"bb",
          7167 => x"26",
          7168 => x"55",
          7169 => x"08",
          7170 => x"81",
          7171 => x"79",
          7172 => x"31",
          7173 => x"70",
          7174 => x"25",
          7175 => x"76",
          7176 => x"81",
          7177 => x"55",
          7178 => x"38",
          7179 => x"0c",
          7180 => x"75",
          7181 => x"54",
          7182 => x"a2",
          7183 => x"7a",
          7184 => x"3f",
          7185 => x"08",
          7186 => x"55",
          7187 => x"89",
          7188 => x"98",
          7189 => x"1a",
          7190 => x"80",
          7191 => x"54",
          7192 => x"98",
          7193 => x"0d",
          7194 => x"0d",
          7195 => x"64",
          7196 => x"59",
          7197 => x"90",
          7198 => x"52",
          7199 => x"cf",
          7200 => x"98",
          7201 => x"bb",
          7202 => x"38",
          7203 => x"55",
          7204 => x"86",
          7205 => x"82",
          7206 => x"19",
          7207 => x"55",
          7208 => x"80",
          7209 => x"38",
          7210 => x"0b",
          7211 => x"82",
          7212 => x"39",
          7213 => x"1a",
          7214 => x"82",
          7215 => x"19",
          7216 => x"08",
          7217 => x"7c",
          7218 => x"74",
          7219 => x"2e",
          7220 => x"94",
          7221 => x"83",
          7222 => x"56",
          7223 => x"38",
          7224 => x"22",
          7225 => x"89",
          7226 => x"55",
          7227 => x"75",
          7228 => x"19",
          7229 => x"39",
          7230 => x"52",
          7231 => x"93",
          7232 => x"98",
          7233 => x"75",
          7234 => x"38",
          7235 => x"ff",
          7236 => x"98",
          7237 => x"19",
          7238 => x"51",
          7239 => x"82",
          7240 => x"80",
          7241 => x"38",
          7242 => x"08",
          7243 => x"2a",
          7244 => x"80",
          7245 => x"38",
          7246 => x"8a",
          7247 => x"5c",
          7248 => x"27",
          7249 => x"7a",
          7250 => x"54",
          7251 => x"52",
          7252 => x"51",
          7253 => x"82",
          7254 => x"fe",
          7255 => x"83",
          7256 => x"56",
          7257 => x"9f",
          7258 => x"08",
          7259 => x"74",
          7260 => x"38",
          7261 => x"b4",
          7262 => x"16",
          7263 => x"89",
          7264 => x"51",
          7265 => x"77",
          7266 => x"b9",
          7267 => x"1a",
          7268 => x"08",
          7269 => x"84",
          7270 => x"57",
          7271 => x"27",
          7272 => x"56",
          7273 => x"52",
          7274 => x"c7",
          7275 => x"98",
          7276 => x"38",
          7277 => x"19",
          7278 => x"06",
          7279 => x"52",
          7280 => x"a2",
          7281 => x"31",
          7282 => x"7f",
          7283 => x"94",
          7284 => x"94",
          7285 => x"5c",
          7286 => x"80",
          7287 => x"bb",
          7288 => x"3d",
          7289 => x"3d",
          7290 => x"65",
          7291 => x"5d",
          7292 => x"0c",
          7293 => x"05",
          7294 => x"f6",
          7295 => x"bb",
          7296 => x"82",
          7297 => x"8a",
          7298 => x"33",
          7299 => x"2e",
          7300 => x"56",
          7301 => x"90",
          7302 => x"81",
          7303 => x"06",
          7304 => x"87",
          7305 => x"2e",
          7306 => x"95",
          7307 => x"91",
          7308 => x"56",
          7309 => x"81",
          7310 => x"34",
          7311 => x"8e",
          7312 => x"08",
          7313 => x"56",
          7314 => x"84",
          7315 => x"5c",
          7316 => x"82",
          7317 => x"18",
          7318 => x"ff",
          7319 => x"74",
          7320 => x"7e",
          7321 => x"ff",
          7322 => x"2a",
          7323 => x"7a",
          7324 => x"8c",
          7325 => x"08",
          7326 => x"38",
          7327 => x"39",
          7328 => x"52",
          7329 => x"e7",
          7330 => x"98",
          7331 => x"bb",
          7332 => x"2e",
          7333 => x"74",
          7334 => x"91",
          7335 => x"2e",
          7336 => x"74",
          7337 => x"88",
          7338 => x"38",
          7339 => x"0c",
          7340 => x"15",
          7341 => x"08",
          7342 => x"06",
          7343 => x"51",
          7344 => x"82",
          7345 => x"fe",
          7346 => x"18",
          7347 => x"51",
          7348 => x"82",
          7349 => x"80",
          7350 => x"38",
          7351 => x"08",
          7352 => x"2a",
          7353 => x"80",
          7354 => x"38",
          7355 => x"8a",
          7356 => x"5b",
          7357 => x"27",
          7358 => x"7b",
          7359 => x"54",
          7360 => x"52",
          7361 => x"51",
          7362 => x"82",
          7363 => x"fe",
          7364 => x"b0",
          7365 => x"31",
          7366 => x"79",
          7367 => x"84",
          7368 => x"16",
          7369 => x"89",
          7370 => x"52",
          7371 => x"cc",
          7372 => x"55",
          7373 => x"16",
          7374 => x"2b",
          7375 => x"39",
          7376 => x"94",
          7377 => x"93",
          7378 => x"cd",
          7379 => x"bb",
          7380 => x"e3",
          7381 => x"b0",
          7382 => x"76",
          7383 => x"94",
          7384 => x"ff",
          7385 => x"71",
          7386 => x"7b",
          7387 => x"38",
          7388 => x"18",
          7389 => x"51",
          7390 => x"82",
          7391 => x"fd",
          7392 => x"53",
          7393 => x"18",
          7394 => x"06",
          7395 => x"51",
          7396 => x"7e",
          7397 => x"83",
          7398 => x"76",
          7399 => x"17",
          7400 => x"1e",
          7401 => x"18",
          7402 => x"0c",
          7403 => x"58",
          7404 => x"74",
          7405 => x"38",
          7406 => x"8c",
          7407 => x"90",
          7408 => x"33",
          7409 => x"55",
          7410 => x"34",
          7411 => x"82",
          7412 => x"90",
          7413 => x"f8",
          7414 => x"8b",
          7415 => x"53",
          7416 => x"f2",
          7417 => x"bb",
          7418 => x"82",
          7419 => x"80",
          7420 => x"16",
          7421 => x"2a",
          7422 => x"51",
          7423 => x"80",
          7424 => x"38",
          7425 => x"52",
          7426 => x"e7",
          7427 => x"98",
          7428 => x"bb",
          7429 => x"d4",
          7430 => x"08",
          7431 => x"a0",
          7432 => x"73",
          7433 => x"88",
          7434 => x"74",
          7435 => x"51",
          7436 => x"8c",
          7437 => x"9c",
          7438 => x"fb",
          7439 => x"b2",
          7440 => x"15",
          7441 => x"3f",
          7442 => x"15",
          7443 => x"3f",
          7444 => x"0b",
          7445 => x"78",
          7446 => x"3f",
          7447 => x"08",
          7448 => x"81",
          7449 => x"57",
          7450 => x"34",
          7451 => x"98",
          7452 => x"0d",
          7453 => x"0d",
          7454 => x"54",
          7455 => x"82",
          7456 => x"53",
          7457 => x"08",
          7458 => x"3d",
          7459 => x"73",
          7460 => x"3f",
          7461 => x"08",
          7462 => x"98",
          7463 => x"82",
          7464 => x"74",
          7465 => x"bb",
          7466 => x"3d",
          7467 => x"3d",
          7468 => x"51",
          7469 => x"8b",
          7470 => x"82",
          7471 => x"24",
          7472 => x"bb",
          7473 => x"d2",
          7474 => x"52",
          7475 => x"98",
          7476 => x"0d",
          7477 => x"0d",
          7478 => x"3d",
          7479 => x"94",
          7480 => x"c1",
          7481 => x"98",
          7482 => x"bb",
          7483 => x"e0",
          7484 => x"63",
          7485 => x"d4",
          7486 => x"8d",
          7487 => x"98",
          7488 => x"bb",
          7489 => x"38",
          7490 => x"05",
          7491 => x"2b",
          7492 => x"80",
          7493 => x"76",
          7494 => x"0c",
          7495 => x"02",
          7496 => x"70",
          7497 => x"81",
          7498 => x"56",
          7499 => x"9e",
          7500 => x"53",
          7501 => x"db",
          7502 => x"bb",
          7503 => x"15",
          7504 => x"82",
          7505 => x"84",
          7506 => x"06",
          7507 => x"55",
          7508 => x"98",
          7509 => x"0d",
          7510 => x"0d",
          7511 => x"5b",
          7512 => x"80",
          7513 => x"ff",
          7514 => x"9f",
          7515 => x"b5",
          7516 => x"98",
          7517 => x"bb",
          7518 => x"fc",
          7519 => x"7a",
          7520 => x"08",
          7521 => x"64",
          7522 => x"2e",
          7523 => x"a0",
          7524 => x"70",
          7525 => x"ea",
          7526 => x"98",
          7527 => x"bb",
          7528 => x"d4",
          7529 => x"7b",
          7530 => x"3f",
          7531 => x"08",
          7532 => x"98",
          7533 => x"38",
          7534 => x"51",
          7535 => x"82",
          7536 => x"45",
          7537 => x"51",
          7538 => x"82",
          7539 => x"57",
          7540 => x"08",
          7541 => x"80",
          7542 => x"da",
          7543 => x"bb",
          7544 => x"82",
          7545 => x"a4",
          7546 => x"7b",
          7547 => x"3f",
          7548 => x"98",
          7549 => x"38",
          7550 => x"51",
          7551 => x"82",
          7552 => x"57",
          7553 => x"08",
          7554 => x"38",
          7555 => x"09",
          7556 => x"38",
          7557 => x"e0",
          7558 => x"dc",
          7559 => x"ff",
          7560 => x"74",
          7561 => x"3f",
          7562 => x"78",
          7563 => x"33",
          7564 => x"56",
          7565 => x"91",
          7566 => x"05",
          7567 => x"81",
          7568 => x"56",
          7569 => x"f5",
          7570 => x"54",
          7571 => x"81",
          7572 => x"80",
          7573 => x"78",
          7574 => x"55",
          7575 => x"11",
          7576 => x"18",
          7577 => x"58",
          7578 => x"34",
          7579 => x"ff",
          7580 => x"55",
          7581 => x"34",
          7582 => x"77",
          7583 => x"81",
          7584 => x"ff",
          7585 => x"55",
          7586 => x"34",
          7587 => x"d2",
          7588 => x"84",
          7589 => x"d0",
          7590 => x"70",
          7591 => x"56",
          7592 => x"76",
          7593 => x"81",
          7594 => x"70",
          7595 => x"56",
          7596 => x"82",
          7597 => x"78",
          7598 => x"80",
          7599 => x"27",
          7600 => x"19",
          7601 => x"7a",
          7602 => x"5c",
          7603 => x"55",
          7604 => x"7a",
          7605 => x"5c",
          7606 => x"2e",
          7607 => x"85",
          7608 => x"94",
          7609 => x"81",
          7610 => x"73",
          7611 => x"81",
          7612 => x"7a",
          7613 => x"38",
          7614 => x"76",
          7615 => x"0c",
          7616 => x"04",
          7617 => x"7b",
          7618 => x"fc",
          7619 => x"53",
          7620 => x"bb",
          7621 => x"98",
          7622 => x"bb",
          7623 => x"fa",
          7624 => x"33",
          7625 => x"f2",
          7626 => x"08",
          7627 => x"27",
          7628 => x"15",
          7629 => x"2a",
          7630 => x"51",
          7631 => x"83",
          7632 => x"94",
          7633 => x"80",
          7634 => x"0c",
          7635 => x"2e",
          7636 => x"79",
          7637 => x"70",
          7638 => x"51",
          7639 => x"2e",
          7640 => x"52",
          7641 => x"fe",
          7642 => x"82",
          7643 => x"ff",
          7644 => x"70",
          7645 => x"fe",
          7646 => x"82",
          7647 => x"73",
          7648 => x"76",
          7649 => x"06",
          7650 => x"0c",
          7651 => x"98",
          7652 => x"58",
          7653 => x"39",
          7654 => x"54",
          7655 => x"73",
          7656 => x"cd",
          7657 => x"bb",
          7658 => x"82",
          7659 => x"81",
          7660 => x"38",
          7661 => x"08",
          7662 => x"9b",
          7663 => x"98",
          7664 => x"0c",
          7665 => x"0c",
          7666 => x"81",
          7667 => x"76",
          7668 => x"38",
          7669 => x"94",
          7670 => x"94",
          7671 => x"16",
          7672 => x"2a",
          7673 => x"51",
          7674 => x"72",
          7675 => x"38",
          7676 => x"51",
          7677 => x"82",
          7678 => x"54",
          7679 => x"08",
          7680 => x"bb",
          7681 => x"a7",
          7682 => x"74",
          7683 => x"3f",
          7684 => x"08",
          7685 => x"2e",
          7686 => x"74",
          7687 => x"79",
          7688 => x"14",
          7689 => x"38",
          7690 => x"0c",
          7691 => x"94",
          7692 => x"94",
          7693 => x"83",
          7694 => x"72",
          7695 => x"38",
          7696 => x"51",
          7697 => x"82",
          7698 => x"94",
          7699 => x"91",
          7700 => x"53",
          7701 => x"81",
          7702 => x"34",
          7703 => x"39",
          7704 => x"82",
          7705 => x"05",
          7706 => x"08",
          7707 => x"08",
          7708 => x"38",
          7709 => x"0c",
          7710 => x"80",
          7711 => x"72",
          7712 => x"73",
          7713 => x"53",
          7714 => x"8c",
          7715 => x"16",
          7716 => x"38",
          7717 => x"0c",
          7718 => x"82",
          7719 => x"8b",
          7720 => x"f9",
          7721 => x"56",
          7722 => x"80",
          7723 => x"38",
          7724 => x"3d",
          7725 => x"8a",
          7726 => x"51",
          7727 => x"82",
          7728 => x"55",
          7729 => x"08",
          7730 => x"77",
          7731 => x"52",
          7732 => x"b5",
          7733 => x"98",
          7734 => x"bb",
          7735 => x"c3",
          7736 => x"33",
          7737 => x"55",
          7738 => x"24",
          7739 => x"16",
          7740 => x"2a",
          7741 => x"51",
          7742 => x"80",
          7743 => x"9c",
          7744 => x"77",
          7745 => x"3f",
          7746 => x"08",
          7747 => x"77",
          7748 => x"22",
          7749 => x"74",
          7750 => x"ce",
          7751 => x"bb",
          7752 => x"74",
          7753 => x"81",
          7754 => x"85",
          7755 => x"74",
          7756 => x"38",
          7757 => x"74",
          7758 => x"bb",
          7759 => x"3d",
          7760 => x"3d",
          7761 => x"3d",
          7762 => x"70",
          7763 => x"ff",
          7764 => x"98",
          7765 => x"82",
          7766 => x"73",
          7767 => x"0d",
          7768 => x"0d",
          7769 => x"3d",
          7770 => x"71",
          7771 => x"e7",
          7772 => x"bb",
          7773 => x"82",
          7774 => x"80",
          7775 => x"93",
          7776 => x"98",
          7777 => x"51",
          7778 => x"82",
          7779 => x"53",
          7780 => x"82",
          7781 => x"52",
          7782 => x"ac",
          7783 => x"98",
          7784 => x"bb",
          7785 => x"2e",
          7786 => x"85",
          7787 => x"87",
          7788 => x"98",
          7789 => x"74",
          7790 => x"d5",
          7791 => x"52",
          7792 => x"89",
          7793 => x"98",
          7794 => x"70",
          7795 => x"07",
          7796 => x"82",
          7797 => x"06",
          7798 => x"54",
          7799 => x"98",
          7800 => x"0d",
          7801 => x"0d",
          7802 => x"53",
          7803 => x"53",
          7804 => x"56",
          7805 => x"82",
          7806 => x"55",
          7807 => x"08",
          7808 => x"52",
          7809 => x"81",
          7810 => x"98",
          7811 => x"bb",
          7812 => x"38",
          7813 => x"05",
          7814 => x"2b",
          7815 => x"80",
          7816 => x"86",
          7817 => x"76",
          7818 => x"38",
          7819 => x"51",
          7820 => x"74",
          7821 => x"0c",
          7822 => x"04",
          7823 => x"63",
          7824 => x"80",
          7825 => x"ec",
          7826 => x"3d",
          7827 => x"3f",
          7828 => x"08",
          7829 => x"98",
          7830 => x"38",
          7831 => x"73",
          7832 => x"08",
          7833 => x"13",
          7834 => x"58",
          7835 => x"26",
          7836 => x"7c",
          7837 => x"39",
          7838 => x"cc",
          7839 => x"81",
          7840 => x"bb",
          7841 => x"33",
          7842 => x"81",
          7843 => x"06",
          7844 => x"75",
          7845 => x"52",
          7846 => x"05",
          7847 => x"3f",
          7848 => x"08",
          7849 => x"38",
          7850 => x"08",
          7851 => x"38",
          7852 => x"08",
          7853 => x"bb",
          7854 => x"80",
          7855 => x"81",
          7856 => x"59",
          7857 => x"14",
          7858 => x"ca",
          7859 => x"39",
          7860 => x"82",
          7861 => x"57",
          7862 => x"38",
          7863 => x"18",
          7864 => x"ff",
          7865 => x"82",
          7866 => x"5b",
          7867 => x"08",
          7868 => x"7c",
          7869 => x"12",
          7870 => x"52",
          7871 => x"82",
          7872 => x"06",
          7873 => x"14",
          7874 => x"cb",
          7875 => x"98",
          7876 => x"ff",
          7877 => x"70",
          7878 => x"82",
          7879 => x"51",
          7880 => x"b4",
          7881 => x"bb",
          7882 => x"bb",
          7883 => x"0a",
          7884 => x"70",
          7885 => x"84",
          7886 => x"51",
          7887 => x"ff",
          7888 => x"56",
          7889 => x"38",
          7890 => x"7c",
          7891 => x"0c",
          7892 => x"81",
          7893 => x"74",
          7894 => x"7a",
          7895 => x"0c",
          7896 => x"04",
          7897 => x"79",
          7898 => x"05",
          7899 => x"57",
          7900 => x"82",
          7901 => x"56",
          7902 => x"08",
          7903 => x"91",
          7904 => x"75",
          7905 => x"90",
          7906 => x"81",
          7907 => x"06",
          7908 => x"87",
          7909 => x"2e",
          7910 => x"94",
          7911 => x"73",
          7912 => x"27",
          7913 => x"73",
          7914 => x"bb",
          7915 => x"88",
          7916 => x"76",
          7917 => x"3f",
          7918 => x"08",
          7919 => x"0c",
          7920 => x"39",
          7921 => x"52",
          7922 => x"bf",
          7923 => x"bb",
          7924 => x"2e",
          7925 => x"83",
          7926 => x"82",
          7927 => x"81",
          7928 => x"06",
          7929 => x"56",
          7930 => x"a0",
          7931 => x"82",
          7932 => x"98",
          7933 => x"94",
          7934 => x"08",
          7935 => x"98",
          7936 => x"51",
          7937 => x"82",
          7938 => x"56",
          7939 => x"8c",
          7940 => x"17",
          7941 => x"07",
          7942 => x"18",
          7943 => x"2e",
          7944 => x"91",
          7945 => x"55",
          7946 => x"98",
          7947 => x"0d",
          7948 => x"0d",
          7949 => x"3d",
          7950 => x"52",
          7951 => x"da",
          7952 => x"bb",
          7953 => x"82",
          7954 => x"81",
          7955 => x"45",
          7956 => x"52",
          7957 => x"52",
          7958 => x"3f",
          7959 => x"08",
          7960 => x"98",
          7961 => x"38",
          7962 => x"05",
          7963 => x"2a",
          7964 => x"51",
          7965 => x"55",
          7966 => x"38",
          7967 => x"54",
          7968 => x"81",
          7969 => x"80",
          7970 => x"70",
          7971 => x"54",
          7972 => x"81",
          7973 => x"52",
          7974 => x"c5",
          7975 => x"98",
          7976 => x"2a",
          7977 => x"51",
          7978 => x"80",
          7979 => x"38",
          7980 => x"bb",
          7981 => x"15",
          7982 => x"86",
          7983 => x"82",
          7984 => x"5c",
          7985 => x"3d",
          7986 => x"c7",
          7987 => x"bb",
          7988 => x"82",
          7989 => x"80",
          7990 => x"bb",
          7991 => x"73",
          7992 => x"3f",
          7993 => x"08",
          7994 => x"98",
          7995 => x"87",
          7996 => x"39",
          7997 => x"08",
          7998 => x"38",
          7999 => x"08",
          8000 => x"77",
          8001 => x"3f",
          8002 => x"08",
          8003 => x"08",
          8004 => x"bb",
          8005 => x"80",
          8006 => x"55",
          8007 => x"94",
          8008 => x"2e",
          8009 => x"53",
          8010 => x"51",
          8011 => x"82",
          8012 => x"55",
          8013 => x"78",
          8014 => x"fe",
          8015 => x"98",
          8016 => x"82",
          8017 => x"a0",
          8018 => x"e9",
          8019 => x"53",
          8020 => x"05",
          8021 => x"51",
          8022 => x"82",
          8023 => x"54",
          8024 => x"08",
          8025 => x"78",
          8026 => x"8e",
          8027 => x"58",
          8028 => x"82",
          8029 => x"54",
          8030 => x"08",
          8031 => x"54",
          8032 => x"82",
          8033 => x"84",
          8034 => x"06",
          8035 => x"02",
          8036 => x"33",
          8037 => x"81",
          8038 => x"86",
          8039 => x"f6",
          8040 => x"74",
          8041 => x"70",
          8042 => x"c3",
          8043 => x"98",
          8044 => x"56",
          8045 => x"08",
          8046 => x"54",
          8047 => x"08",
          8048 => x"81",
          8049 => x"82",
          8050 => x"98",
          8051 => x"09",
          8052 => x"38",
          8053 => x"b4",
          8054 => x"b0",
          8055 => x"98",
          8056 => x"51",
          8057 => x"82",
          8058 => x"54",
          8059 => x"08",
          8060 => x"8b",
          8061 => x"b4",
          8062 => x"b7",
          8063 => x"54",
          8064 => x"15",
          8065 => x"90",
          8066 => x"34",
          8067 => x"0a",
          8068 => x"19",
          8069 => x"9f",
          8070 => x"78",
          8071 => x"51",
          8072 => x"a0",
          8073 => x"11",
          8074 => x"05",
          8075 => x"b6",
          8076 => x"ae",
          8077 => x"15",
          8078 => x"78",
          8079 => x"53",
          8080 => x"3f",
          8081 => x"0b",
          8082 => x"77",
          8083 => x"3f",
          8084 => x"08",
          8085 => x"98",
          8086 => x"82",
          8087 => x"52",
          8088 => x"51",
          8089 => x"3f",
          8090 => x"52",
          8091 => x"aa",
          8092 => x"90",
          8093 => x"34",
          8094 => x"0b",
          8095 => x"78",
          8096 => x"b6",
          8097 => x"98",
          8098 => x"39",
          8099 => x"52",
          8100 => x"be",
          8101 => x"82",
          8102 => x"99",
          8103 => x"da",
          8104 => x"3d",
          8105 => x"d2",
          8106 => x"53",
          8107 => x"84",
          8108 => x"3d",
          8109 => x"3f",
          8110 => x"08",
          8111 => x"98",
          8112 => x"38",
          8113 => x"3d",
          8114 => x"3d",
          8115 => x"cc",
          8116 => x"bb",
          8117 => x"82",
          8118 => x"82",
          8119 => x"81",
          8120 => x"81",
          8121 => x"86",
          8122 => x"aa",
          8123 => x"a4",
          8124 => x"a8",
          8125 => x"05",
          8126 => x"ea",
          8127 => x"77",
          8128 => x"70",
          8129 => x"b4",
          8130 => x"3d",
          8131 => x"51",
          8132 => x"82",
          8133 => x"55",
          8134 => x"08",
          8135 => x"6f",
          8136 => x"06",
          8137 => x"a2",
          8138 => x"92",
          8139 => x"81",
          8140 => x"bb",
          8141 => x"2e",
          8142 => x"81",
          8143 => x"51",
          8144 => x"82",
          8145 => x"55",
          8146 => x"08",
          8147 => x"68",
          8148 => x"a8",
          8149 => x"05",
          8150 => x"51",
          8151 => x"3f",
          8152 => x"33",
          8153 => x"8b",
          8154 => x"84",
          8155 => x"06",
          8156 => x"73",
          8157 => x"a0",
          8158 => x"8b",
          8159 => x"54",
          8160 => x"15",
          8161 => x"33",
          8162 => x"70",
          8163 => x"55",
          8164 => x"2e",
          8165 => x"6e",
          8166 => x"df",
          8167 => x"78",
          8168 => x"3f",
          8169 => x"08",
          8170 => x"ff",
          8171 => x"82",
          8172 => x"98",
          8173 => x"80",
          8174 => x"bb",
          8175 => x"78",
          8176 => x"af",
          8177 => x"98",
          8178 => x"d4",
          8179 => x"55",
          8180 => x"08",
          8181 => x"81",
          8182 => x"73",
          8183 => x"81",
          8184 => x"63",
          8185 => x"76",
          8186 => x"3f",
          8187 => x"0b",
          8188 => x"87",
          8189 => x"98",
          8190 => x"77",
          8191 => x"3f",
          8192 => x"08",
          8193 => x"98",
          8194 => x"78",
          8195 => x"aa",
          8196 => x"98",
          8197 => x"82",
          8198 => x"a8",
          8199 => x"ed",
          8200 => x"80",
          8201 => x"02",
          8202 => x"df",
          8203 => x"57",
          8204 => x"3d",
          8205 => x"96",
          8206 => x"e9",
          8207 => x"98",
          8208 => x"bb",
          8209 => x"cf",
          8210 => x"65",
          8211 => x"d4",
          8212 => x"b5",
          8213 => x"98",
          8214 => x"bb",
          8215 => x"38",
          8216 => x"05",
          8217 => x"06",
          8218 => x"73",
          8219 => x"a7",
          8220 => x"09",
          8221 => x"71",
          8222 => x"06",
          8223 => x"55",
          8224 => x"15",
          8225 => x"81",
          8226 => x"34",
          8227 => x"b4",
          8228 => x"bb",
          8229 => x"74",
          8230 => x"0c",
          8231 => x"04",
          8232 => x"64",
          8233 => x"93",
          8234 => x"52",
          8235 => x"d1",
          8236 => x"bb",
          8237 => x"82",
          8238 => x"80",
          8239 => x"58",
          8240 => x"3d",
          8241 => x"c8",
          8242 => x"bb",
          8243 => x"82",
          8244 => x"b4",
          8245 => x"c7",
          8246 => x"a0",
          8247 => x"55",
          8248 => x"84",
          8249 => x"17",
          8250 => x"2b",
          8251 => x"96",
          8252 => x"b0",
          8253 => x"54",
          8254 => x"15",
          8255 => x"ff",
          8256 => x"82",
          8257 => x"55",
          8258 => x"98",
          8259 => x"0d",
          8260 => x"0d",
          8261 => x"5a",
          8262 => x"3d",
          8263 => x"99",
          8264 => x"81",
          8265 => x"98",
          8266 => x"98",
          8267 => x"82",
          8268 => x"07",
          8269 => x"55",
          8270 => x"2e",
          8271 => x"81",
          8272 => x"55",
          8273 => x"2e",
          8274 => x"7b",
          8275 => x"80",
          8276 => x"70",
          8277 => x"be",
          8278 => x"bb",
          8279 => x"82",
          8280 => x"80",
          8281 => x"52",
          8282 => x"dc",
          8283 => x"98",
          8284 => x"bb",
          8285 => x"38",
          8286 => x"08",
          8287 => x"08",
          8288 => x"56",
          8289 => x"19",
          8290 => x"59",
          8291 => x"74",
          8292 => x"56",
          8293 => x"ec",
          8294 => x"75",
          8295 => x"74",
          8296 => x"2e",
          8297 => x"16",
          8298 => x"33",
          8299 => x"73",
          8300 => x"38",
          8301 => x"84",
          8302 => x"06",
          8303 => x"7a",
          8304 => x"76",
          8305 => x"07",
          8306 => x"54",
          8307 => x"80",
          8308 => x"80",
          8309 => x"7b",
          8310 => x"53",
          8311 => x"93",
          8312 => x"98",
          8313 => x"bb",
          8314 => x"38",
          8315 => x"55",
          8316 => x"56",
          8317 => x"8b",
          8318 => x"56",
          8319 => x"83",
          8320 => x"75",
          8321 => x"51",
          8322 => x"3f",
          8323 => x"08",
          8324 => x"82",
          8325 => x"98",
          8326 => x"e6",
          8327 => x"53",
          8328 => x"b8",
          8329 => x"3d",
          8330 => x"3f",
          8331 => x"08",
          8332 => x"08",
          8333 => x"bb",
          8334 => x"98",
          8335 => x"a0",
          8336 => x"70",
          8337 => x"ae",
          8338 => x"6d",
          8339 => x"81",
          8340 => x"57",
          8341 => x"74",
          8342 => x"38",
          8343 => x"81",
          8344 => x"81",
          8345 => x"52",
          8346 => x"89",
          8347 => x"98",
          8348 => x"a5",
          8349 => x"33",
          8350 => x"54",
          8351 => x"3f",
          8352 => x"08",
          8353 => x"38",
          8354 => x"76",
          8355 => x"05",
          8356 => x"39",
          8357 => x"08",
          8358 => x"15",
          8359 => x"ff",
          8360 => x"73",
          8361 => x"38",
          8362 => x"83",
          8363 => x"56",
          8364 => x"75",
          8365 => x"82",
          8366 => x"33",
          8367 => x"2e",
          8368 => x"52",
          8369 => x"51",
          8370 => x"3f",
          8371 => x"08",
          8372 => x"ff",
          8373 => x"38",
          8374 => x"88",
          8375 => x"8a",
          8376 => x"38",
          8377 => x"ec",
          8378 => x"75",
          8379 => x"74",
          8380 => x"73",
          8381 => x"05",
          8382 => x"17",
          8383 => x"70",
          8384 => x"34",
          8385 => x"70",
          8386 => x"ff",
          8387 => x"55",
          8388 => x"26",
          8389 => x"8b",
          8390 => x"86",
          8391 => x"e5",
          8392 => x"38",
          8393 => x"99",
          8394 => x"05",
          8395 => x"70",
          8396 => x"73",
          8397 => x"81",
          8398 => x"ff",
          8399 => x"ed",
          8400 => x"80",
          8401 => x"91",
          8402 => x"55",
          8403 => x"3f",
          8404 => x"08",
          8405 => x"98",
          8406 => x"38",
          8407 => x"51",
          8408 => x"3f",
          8409 => x"08",
          8410 => x"98",
          8411 => x"76",
          8412 => x"67",
          8413 => x"34",
          8414 => x"82",
          8415 => x"84",
          8416 => x"06",
          8417 => x"80",
          8418 => x"2e",
          8419 => x"81",
          8420 => x"ff",
          8421 => x"82",
          8422 => x"54",
          8423 => x"08",
          8424 => x"53",
          8425 => x"08",
          8426 => x"ff",
          8427 => x"67",
          8428 => x"8b",
          8429 => x"53",
          8430 => x"51",
          8431 => x"3f",
          8432 => x"0b",
          8433 => x"79",
          8434 => x"ee",
          8435 => x"98",
          8436 => x"55",
          8437 => x"98",
          8438 => x"0d",
          8439 => x"0d",
          8440 => x"88",
          8441 => x"05",
          8442 => x"fc",
          8443 => x"54",
          8444 => x"d2",
          8445 => x"bb",
          8446 => x"82",
          8447 => x"82",
          8448 => x"1a",
          8449 => x"82",
          8450 => x"80",
          8451 => x"8c",
          8452 => x"78",
          8453 => x"1a",
          8454 => x"2a",
          8455 => x"51",
          8456 => x"90",
          8457 => x"82",
          8458 => x"58",
          8459 => x"81",
          8460 => x"39",
          8461 => x"22",
          8462 => x"70",
          8463 => x"56",
          8464 => x"c9",
          8465 => x"14",
          8466 => x"30",
          8467 => x"9f",
          8468 => x"98",
          8469 => x"19",
          8470 => x"5a",
          8471 => x"81",
          8472 => x"38",
          8473 => x"77",
          8474 => x"82",
          8475 => x"56",
          8476 => x"74",
          8477 => x"ff",
          8478 => x"81",
          8479 => x"55",
          8480 => x"75",
          8481 => x"82",
          8482 => x"98",
          8483 => x"ff",
          8484 => x"bb",
          8485 => x"2e",
          8486 => x"82",
          8487 => x"8e",
          8488 => x"56",
          8489 => x"09",
          8490 => x"38",
          8491 => x"59",
          8492 => x"77",
          8493 => x"06",
          8494 => x"87",
          8495 => x"39",
          8496 => x"ba",
          8497 => x"55",
          8498 => x"2e",
          8499 => x"15",
          8500 => x"2e",
          8501 => x"83",
          8502 => x"75",
          8503 => x"7e",
          8504 => x"a8",
          8505 => x"98",
          8506 => x"bb",
          8507 => x"ce",
          8508 => x"16",
          8509 => x"56",
          8510 => x"38",
          8511 => x"19",
          8512 => x"8c",
          8513 => x"7d",
          8514 => x"38",
          8515 => x"0c",
          8516 => x"0c",
          8517 => x"80",
          8518 => x"73",
          8519 => x"98",
          8520 => x"05",
          8521 => x"57",
          8522 => x"26",
          8523 => x"7b",
          8524 => x"0c",
          8525 => x"81",
          8526 => x"84",
          8527 => x"54",
          8528 => x"98",
          8529 => x"0d",
          8530 => x"0d",
          8531 => x"88",
          8532 => x"05",
          8533 => x"54",
          8534 => x"c5",
          8535 => x"56",
          8536 => x"bb",
          8537 => x"8b",
          8538 => x"bb",
          8539 => x"29",
          8540 => x"05",
          8541 => x"55",
          8542 => x"84",
          8543 => x"34",
          8544 => x"08",
          8545 => x"5f",
          8546 => x"51",
          8547 => x"3f",
          8548 => x"08",
          8549 => x"70",
          8550 => x"57",
          8551 => x"8b",
          8552 => x"82",
          8553 => x"06",
          8554 => x"56",
          8555 => x"38",
          8556 => x"05",
          8557 => x"7e",
          8558 => x"f0",
          8559 => x"98",
          8560 => x"67",
          8561 => x"2e",
          8562 => x"82",
          8563 => x"8b",
          8564 => x"75",
          8565 => x"80",
          8566 => x"81",
          8567 => x"2e",
          8568 => x"80",
          8569 => x"38",
          8570 => x"0a",
          8571 => x"ff",
          8572 => x"55",
          8573 => x"86",
          8574 => x"8a",
          8575 => x"89",
          8576 => x"2a",
          8577 => x"77",
          8578 => x"59",
          8579 => x"81",
          8580 => x"70",
          8581 => x"07",
          8582 => x"56",
          8583 => x"38",
          8584 => x"05",
          8585 => x"7e",
          8586 => x"80",
          8587 => x"82",
          8588 => x"8a",
          8589 => x"83",
          8590 => x"06",
          8591 => x"08",
          8592 => x"74",
          8593 => x"41",
          8594 => x"56",
          8595 => x"8a",
          8596 => x"61",
          8597 => x"55",
          8598 => x"27",
          8599 => x"93",
          8600 => x"80",
          8601 => x"38",
          8602 => x"70",
          8603 => x"43",
          8604 => x"95",
          8605 => x"06",
          8606 => x"2e",
          8607 => x"77",
          8608 => x"74",
          8609 => x"83",
          8610 => x"06",
          8611 => x"82",
          8612 => x"2e",
          8613 => x"78",
          8614 => x"2e",
          8615 => x"80",
          8616 => x"ae",
          8617 => x"2a",
          8618 => x"82",
          8619 => x"56",
          8620 => x"2e",
          8621 => x"77",
          8622 => x"82",
          8623 => x"79",
          8624 => x"70",
          8625 => x"5a",
          8626 => x"86",
          8627 => x"27",
          8628 => x"52",
          8629 => x"c4",
          8630 => x"bb",
          8631 => x"29",
          8632 => x"70",
          8633 => x"55",
          8634 => x"0b",
          8635 => x"08",
          8636 => x"05",
          8637 => x"ff",
          8638 => x"27",
          8639 => x"88",
          8640 => x"ae",
          8641 => x"2a",
          8642 => x"82",
          8643 => x"56",
          8644 => x"2e",
          8645 => x"77",
          8646 => x"82",
          8647 => x"79",
          8648 => x"70",
          8649 => x"5a",
          8650 => x"86",
          8651 => x"27",
          8652 => x"52",
          8653 => x"c3",
          8654 => x"bb",
          8655 => x"84",
          8656 => x"bb",
          8657 => x"f5",
          8658 => x"81",
          8659 => x"98",
          8660 => x"bb",
          8661 => x"71",
          8662 => x"83",
          8663 => x"5e",
          8664 => x"89",
          8665 => x"5c",
          8666 => x"1c",
          8667 => x"05",
          8668 => x"ff",
          8669 => x"70",
          8670 => x"31",
          8671 => x"57",
          8672 => x"83",
          8673 => x"06",
          8674 => x"1c",
          8675 => x"5c",
          8676 => x"1d",
          8677 => x"29",
          8678 => x"31",
          8679 => x"55",
          8680 => x"87",
          8681 => x"7c",
          8682 => x"7a",
          8683 => x"31",
          8684 => x"c2",
          8685 => x"bb",
          8686 => x"7d",
          8687 => x"81",
          8688 => x"82",
          8689 => x"83",
          8690 => x"80",
          8691 => x"87",
          8692 => x"81",
          8693 => x"fd",
          8694 => x"f8",
          8695 => x"2e",
          8696 => x"80",
          8697 => x"ff",
          8698 => x"bb",
          8699 => x"a0",
          8700 => x"38",
          8701 => x"74",
          8702 => x"86",
          8703 => x"fd",
          8704 => x"81",
          8705 => x"80",
          8706 => x"83",
          8707 => x"39",
          8708 => x"08",
          8709 => x"92",
          8710 => x"b8",
          8711 => x"59",
          8712 => x"27",
          8713 => x"86",
          8714 => x"55",
          8715 => x"09",
          8716 => x"38",
          8717 => x"f5",
          8718 => x"38",
          8719 => x"55",
          8720 => x"86",
          8721 => x"80",
          8722 => x"7a",
          8723 => x"b9",
          8724 => x"82",
          8725 => x"7a",
          8726 => x"8a",
          8727 => x"52",
          8728 => x"ff",
          8729 => x"79",
          8730 => x"7b",
          8731 => x"06",
          8732 => x"51",
          8733 => x"3f",
          8734 => x"1c",
          8735 => x"32",
          8736 => x"96",
          8737 => x"06",
          8738 => x"91",
          8739 => x"a1",
          8740 => x"55",
          8741 => x"ff",
          8742 => x"74",
          8743 => x"06",
          8744 => x"51",
          8745 => x"3f",
          8746 => x"52",
          8747 => x"ff",
          8748 => x"f8",
          8749 => x"34",
          8750 => x"1b",
          8751 => x"d9",
          8752 => x"52",
          8753 => x"ff",
          8754 => x"60",
          8755 => x"51",
          8756 => x"3f",
          8757 => x"09",
          8758 => x"cb",
          8759 => x"b2",
          8760 => x"c3",
          8761 => x"a0",
          8762 => x"52",
          8763 => x"ff",
          8764 => x"82",
          8765 => x"51",
          8766 => x"3f",
          8767 => x"1b",
          8768 => x"95",
          8769 => x"b2",
          8770 => x"a0",
          8771 => x"80",
          8772 => x"1c",
          8773 => x"80",
          8774 => x"93",
          8775 => x"a8",
          8776 => x"1b",
          8777 => x"82",
          8778 => x"52",
          8779 => x"ff",
          8780 => x"7c",
          8781 => x"06",
          8782 => x"51",
          8783 => x"3f",
          8784 => x"a4",
          8785 => x"0b",
          8786 => x"93",
          8787 => x"bc",
          8788 => x"51",
          8789 => x"3f",
          8790 => x"52",
          8791 => x"70",
          8792 => x"9f",
          8793 => x"54",
          8794 => x"52",
          8795 => x"9b",
          8796 => x"56",
          8797 => x"08",
          8798 => x"7d",
          8799 => x"81",
          8800 => x"38",
          8801 => x"86",
          8802 => x"52",
          8803 => x"9b",
          8804 => x"80",
          8805 => x"7a",
          8806 => x"ed",
          8807 => x"85",
          8808 => x"7a",
          8809 => x"8f",
          8810 => x"85",
          8811 => x"83",
          8812 => x"ff",
          8813 => x"ff",
          8814 => x"e8",
          8815 => x"9e",
          8816 => x"52",
          8817 => x"51",
          8818 => x"3f",
          8819 => x"52",
          8820 => x"9e",
          8821 => x"54",
          8822 => x"53",
          8823 => x"51",
          8824 => x"3f",
          8825 => x"16",
          8826 => x"7e",
          8827 => x"d8",
          8828 => x"80",
          8829 => x"ff",
          8830 => x"7f",
          8831 => x"7d",
          8832 => x"81",
          8833 => x"f8",
          8834 => x"ff",
          8835 => x"ff",
          8836 => x"51",
          8837 => x"3f",
          8838 => x"88",
          8839 => x"39",
          8840 => x"f8",
          8841 => x"2e",
          8842 => x"55",
          8843 => x"51",
          8844 => x"3f",
          8845 => x"57",
          8846 => x"83",
          8847 => x"76",
          8848 => x"7a",
          8849 => x"ff",
          8850 => x"82",
          8851 => x"82",
          8852 => x"80",
          8853 => x"98",
          8854 => x"51",
          8855 => x"3f",
          8856 => x"78",
          8857 => x"74",
          8858 => x"18",
          8859 => x"2e",
          8860 => x"79",
          8861 => x"2e",
          8862 => x"55",
          8863 => x"62",
          8864 => x"74",
          8865 => x"75",
          8866 => x"7e",
          8867 => x"b8",
          8868 => x"98",
          8869 => x"38",
          8870 => x"78",
          8871 => x"74",
          8872 => x"56",
          8873 => x"93",
          8874 => x"66",
          8875 => x"26",
          8876 => x"56",
          8877 => x"83",
          8878 => x"64",
          8879 => x"77",
          8880 => x"84",
          8881 => x"52",
          8882 => x"9d",
          8883 => x"d4",
          8884 => x"51",
          8885 => x"3f",
          8886 => x"55",
          8887 => x"81",
          8888 => x"34",
          8889 => x"16",
          8890 => x"16",
          8891 => x"16",
          8892 => x"05",
          8893 => x"c1",
          8894 => x"fe",
          8895 => x"fe",
          8896 => x"34",
          8897 => x"08",
          8898 => x"07",
          8899 => x"16",
          8900 => x"98",
          8901 => x"34",
          8902 => x"c6",
          8903 => x"9c",
          8904 => x"52",
          8905 => x"51",
          8906 => x"3f",
          8907 => x"53",
          8908 => x"51",
          8909 => x"3f",
          8910 => x"bb",
          8911 => x"38",
          8912 => x"52",
          8913 => x"99",
          8914 => x"56",
          8915 => x"08",
          8916 => x"39",
          8917 => x"39",
          8918 => x"39",
          8919 => x"08",
          8920 => x"bb",
          8921 => x"3d",
          8922 => x"3d",
          8923 => x"5b",
          8924 => x"60",
          8925 => x"57",
          8926 => x"25",
          8927 => x"3d",
          8928 => x"55",
          8929 => x"15",
          8930 => x"c9",
          8931 => x"81",
          8932 => x"06",
          8933 => x"3d",
          8934 => x"8d",
          8935 => x"74",
          8936 => x"05",
          8937 => x"17",
          8938 => x"2e",
          8939 => x"c9",
          8940 => x"34",
          8941 => x"83",
          8942 => x"74",
          8943 => x"0c",
          8944 => x"04",
          8945 => x"7b",
          8946 => x"b3",
          8947 => x"57",
          8948 => x"09",
          8949 => x"38",
          8950 => x"51",
          8951 => x"17",
          8952 => x"76",
          8953 => x"88",
          8954 => x"17",
          8955 => x"59",
          8956 => x"81",
          8957 => x"76",
          8958 => x"8b",
          8959 => x"54",
          8960 => x"17",
          8961 => x"51",
          8962 => x"79",
          8963 => x"30",
          8964 => x"9f",
          8965 => x"53",
          8966 => x"75",
          8967 => x"81",
          8968 => x"0c",
          8969 => x"04",
          8970 => x"79",
          8971 => x"56",
          8972 => x"24",
          8973 => x"3d",
          8974 => x"74",
          8975 => x"52",
          8976 => x"cb",
          8977 => x"bb",
          8978 => x"38",
          8979 => x"78",
          8980 => x"06",
          8981 => x"16",
          8982 => x"39",
          8983 => x"82",
          8984 => x"89",
          8985 => x"fd",
          8986 => x"54",
          8987 => x"80",
          8988 => x"ff",
          8989 => x"76",
          8990 => x"3d",
          8991 => x"3d",
          8992 => x"e3",
          8993 => x"53",
          8994 => x"53",
          8995 => x"3f",
          8996 => x"51",
          8997 => x"72",
          8998 => x"3f",
          8999 => x"04",
          9000 => x"ff",
          9001 => x"ff",
          9002 => x"ff",
          9003 => x"00",
          9004 => x"a8",
          9005 => x"2c",
          9006 => x"33",
          9007 => x"3a",
          9008 => x"41",
          9009 => x"48",
          9010 => x"4f",
          9011 => x"56",
          9012 => x"5d",
          9013 => x"64",
          9014 => x"6b",
          9015 => x"72",
          9016 => x"78",
          9017 => x"7e",
          9018 => x"84",
          9019 => x"8a",
          9020 => x"90",
          9021 => x"96",
          9022 => x"9c",
          9023 => x"a2",
          9024 => x"6a",
          9025 => x"70",
          9026 => x"76",
          9027 => x"7c",
          9028 => x"82",
          9029 => x"93",
          9030 => x"89",
          9031 => x"81",
          9032 => x"bb",
          9033 => x"71",
          9034 => x"68",
          9035 => x"35",
          9036 => x"91",
          9037 => x"73",
          9038 => x"09",
          9039 => x"8f",
          9040 => x"30",
          9041 => x"68",
          9042 => x"81",
          9043 => x"a5",
          9044 => x"35",
          9045 => x"68",
          9046 => x"68",
          9047 => x"8f",
          9048 => x"09",
          9049 => x"91",
          9050 => x"bb",
          9051 => x"2f",
          9052 => x"18",
          9053 => x"18",
          9054 => x"5e",
          9055 => x"18",
          9056 => x"18",
          9057 => x"18",
          9058 => x"18",
          9059 => x"18",
          9060 => x"18",
          9061 => x"18",
          9062 => x"1b",
          9063 => x"18",
          9064 => x"46",
          9065 => x"76",
          9066 => x"18",
          9067 => x"18",
          9068 => x"18",
          9069 => x"18",
          9070 => x"18",
          9071 => x"18",
          9072 => x"18",
          9073 => x"18",
          9074 => x"18",
          9075 => x"18",
          9076 => x"18",
          9077 => x"18",
          9078 => x"18",
          9079 => x"18",
          9080 => x"18",
          9081 => x"18",
          9082 => x"18",
          9083 => x"18",
          9084 => x"18",
          9085 => x"18",
          9086 => x"18",
          9087 => x"18",
          9088 => x"18",
          9089 => x"18",
          9090 => x"18",
          9091 => x"18",
          9092 => x"18",
          9093 => x"18",
          9094 => x"18",
          9095 => x"18",
          9096 => x"18",
          9097 => x"18",
          9098 => x"18",
          9099 => x"18",
          9100 => x"18",
          9101 => x"18",
          9102 => x"a6",
          9103 => x"18",
          9104 => x"18",
          9105 => x"18",
          9106 => x"18",
          9107 => x"14",
          9108 => x"18",
          9109 => x"18",
          9110 => x"18",
          9111 => x"18",
          9112 => x"18",
          9113 => x"18",
          9114 => x"18",
          9115 => x"18",
          9116 => x"18",
          9117 => x"18",
          9118 => x"d6",
          9119 => x"3d",
          9120 => x"ad",
          9121 => x"ad",
          9122 => x"ad",
          9123 => x"18",
          9124 => x"3d",
          9125 => x"18",
          9126 => x"18",
          9127 => x"96",
          9128 => x"18",
          9129 => x"18",
          9130 => x"ea",
          9131 => x"f5",
          9132 => x"18",
          9133 => x"18",
          9134 => x"0f",
          9135 => x"18",
          9136 => x"1d",
          9137 => x"18",
          9138 => x"18",
          9139 => x"14",
          9140 => x"69",
          9141 => x"00",
          9142 => x"63",
          9143 => x"00",
          9144 => x"69",
          9145 => x"00",
          9146 => x"61",
          9147 => x"00",
          9148 => x"65",
          9149 => x"00",
          9150 => x"65",
          9151 => x"00",
          9152 => x"70",
          9153 => x"00",
          9154 => x"66",
          9155 => x"00",
          9156 => x"6d",
          9157 => x"00",
          9158 => x"00",
          9159 => x"00",
          9160 => x"00",
          9161 => x"00",
          9162 => x"00",
          9163 => x"00",
          9164 => x"00",
          9165 => x"6c",
          9166 => x"00",
          9167 => x"00",
          9168 => x"74",
          9169 => x"00",
          9170 => x"65",
          9171 => x"00",
          9172 => x"6f",
          9173 => x"00",
          9174 => x"74",
          9175 => x"00",
          9176 => x"73",
          9177 => x"00",
          9178 => x"73",
          9179 => x"00",
          9180 => x"6f",
          9181 => x"00",
          9182 => x"00",
          9183 => x"6b",
          9184 => x"72",
          9185 => x"00",
          9186 => x"65",
          9187 => x"6c",
          9188 => x"72",
          9189 => x"0a",
          9190 => x"00",
          9191 => x"6b",
          9192 => x"74",
          9193 => x"61",
          9194 => x"0a",
          9195 => x"00",
          9196 => x"66",
          9197 => x"20",
          9198 => x"6e",
          9199 => x"00",
          9200 => x"70",
          9201 => x"20",
          9202 => x"6e",
          9203 => x"00",
          9204 => x"61",
          9205 => x"20",
          9206 => x"65",
          9207 => x"65",
          9208 => x"00",
          9209 => x"65",
          9210 => x"64",
          9211 => x"65",
          9212 => x"00",
          9213 => x"65",
          9214 => x"72",
          9215 => x"79",
          9216 => x"69",
          9217 => x"2e",
          9218 => x"00",
          9219 => x"65",
          9220 => x"6e",
          9221 => x"20",
          9222 => x"61",
          9223 => x"2e",
          9224 => x"00",
          9225 => x"69",
          9226 => x"72",
          9227 => x"20",
          9228 => x"74",
          9229 => x"65",
          9230 => x"00",
          9231 => x"76",
          9232 => x"75",
          9233 => x"72",
          9234 => x"20",
          9235 => x"61",
          9236 => x"2e",
          9237 => x"00",
          9238 => x"6b",
          9239 => x"74",
          9240 => x"61",
          9241 => x"64",
          9242 => x"00",
          9243 => x"63",
          9244 => x"61",
          9245 => x"6c",
          9246 => x"69",
          9247 => x"79",
          9248 => x"6d",
          9249 => x"75",
          9250 => x"6f",
          9251 => x"69",
          9252 => x"0a",
          9253 => x"00",
          9254 => x"6d",
          9255 => x"61",
          9256 => x"74",
          9257 => x"0a",
          9258 => x"00",
          9259 => x"65",
          9260 => x"2c",
          9261 => x"65",
          9262 => x"69",
          9263 => x"63",
          9264 => x"65",
          9265 => x"64",
          9266 => x"00",
          9267 => x"65",
          9268 => x"20",
          9269 => x"6b",
          9270 => x"0a",
          9271 => x"00",
          9272 => x"75",
          9273 => x"63",
          9274 => x"74",
          9275 => x"6d",
          9276 => x"2e",
          9277 => x"00",
          9278 => x"20",
          9279 => x"79",
          9280 => x"65",
          9281 => x"69",
          9282 => x"2e",
          9283 => x"00",
          9284 => x"61",
          9285 => x"65",
          9286 => x"69",
          9287 => x"72",
          9288 => x"74",
          9289 => x"00",
          9290 => x"63",
          9291 => x"2e",
          9292 => x"00",
          9293 => x"6e",
          9294 => x"20",
          9295 => x"6f",
          9296 => x"00",
          9297 => x"75",
          9298 => x"74",
          9299 => x"25",
          9300 => x"74",
          9301 => x"75",
          9302 => x"74",
          9303 => x"73",
          9304 => x"0a",
          9305 => x"00",
          9306 => x"64",
          9307 => x"00",
          9308 => x"58",
          9309 => x"00",
          9310 => x"00",
          9311 => x"58",
          9312 => x"00",
          9313 => x"20",
          9314 => x"20",
          9315 => x"00",
          9316 => x"58",
          9317 => x"00",
          9318 => x"00",
          9319 => x"00",
          9320 => x"00",
          9321 => x"54",
          9322 => x"00",
          9323 => x"20",
          9324 => x"28",
          9325 => x"00",
          9326 => x"30",
          9327 => x"30",
          9328 => x"00",
          9329 => x"35",
          9330 => x"00",
          9331 => x"55",
          9332 => x"65",
          9333 => x"30",
          9334 => x"20",
          9335 => x"25",
          9336 => x"2a",
          9337 => x"00",
          9338 => x"54",
          9339 => x"6e",
          9340 => x"72",
          9341 => x"20",
          9342 => x"64",
          9343 => x"0a",
          9344 => x"00",
          9345 => x"65",
          9346 => x"6e",
          9347 => x"72",
          9348 => x"0a",
          9349 => x"00",
          9350 => x"20",
          9351 => x"65",
          9352 => x"70",
          9353 => x"00",
          9354 => x"54",
          9355 => x"44",
          9356 => x"74",
          9357 => x"75",
          9358 => x"00",
          9359 => x"54",
          9360 => x"52",
          9361 => x"74",
          9362 => x"75",
          9363 => x"00",
          9364 => x"54",
          9365 => x"58",
          9366 => x"74",
          9367 => x"75",
          9368 => x"00",
          9369 => x"54",
          9370 => x"58",
          9371 => x"74",
          9372 => x"75",
          9373 => x"00",
          9374 => x"54",
          9375 => x"58",
          9376 => x"74",
          9377 => x"75",
          9378 => x"00",
          9379 => x"54",
          9380 => x"58",
          9381 => x"74",
          9382 => x"75",
          9383 => x"00",
          9384 => x"74",
          9385 => x"20",
          9386 => x"74",
          9387 => x"72",
          9388 => x"0a",
          9389 => x"00",
          9390 => x"62",
          9391 => x"67",
          9392 => x"6d",
          9393 => x"2e",
          9394 => x"00",
          9395 => x"6f",
          9396 => x"63",
          9397 => x"74",
          9398 => x"00",
          9399 => x"74",
          9400 => x"73",
          9401 => x"00",
          9402 => x"00",
          9403 => x"6c",
          9404 => x"74",
          9405 => x"6e",
          9406 => x"61",
          9407 => x"65",
          9408 => x"20",
          9409 => x"64",
          9410 => x"20",
          9411 => x"61",
          9412 => x"69",
          9413 => x"20",
          9414 => x"75",
          9415 => x"79",
          9416 => x"00",
          9417 => x"00",
          9418 => x"20",
          9419 => x"6b",
          9420 => x"21",
          9421 => x"00",
          9422 => x"74",
          9423 => x"69",
          9424 => x"2e",
          9425 => x"00",
          9426 => x"6c",
          9427 => x"74",
          9428 => x"6e",
          9429 => x"61",
          9430 => x"65",
          9431 => x"00",
          9432 => x"25",
          9433 => x"00",
          9434 => x"00",
          9435 => x"61",
          9436 => x"67",
          9437 => x"2e",
          9438 => x"00",
          9439 => x"79",
          9440 => x"2e",
          9441 => x"00",
          9442 => x"70",
          9443 => x"6e",
          9444 => x"2e",
          9445 => x"00",
          9446 => x"6c",
          9447 => x"30",
          9448 => x"2d",
          9449 => x"38",
          9450 => x"25",
          9451 => x"29",
          9452 => x"00",
          9453 => x"70",
          9454 => x"6d",
          9455 => x"0a",
          9456 => x"00",
          9457 => x"6d",
          9458 => x"74",
          9459 => x"00",
          9460 => x"58",
          9461 => x"32",
          9462 => x"00",
          9463 => x"0a",
          9464 => x"00",
          9465 => x"58",
          9466 => x"34",
          9467 => x"00",
          9468 => x"58",
          9469 => x"38",
          9470 => x"00",
          9471 => x"61",
          9472 => x"6e",
          9473 => x"6e",
          9474 => x"72",
          9475 => x"73",
          9476 => x"00",
          9477 => x"62",
          9478 => x"67",
          9479 => x"74",
          9480 => x"75",
          9481 => x"0a",
          9482 => x"00",
          9483 => x"61",
          9484 => x"64",
          9485 => x"72",
          9486 => x"69",
          9487 => x"00",
          9488 => x"62",
          9489 => x"67",
          9490 => x"72",
          9491 => x"69",
          9492 => x"00",
          9493 => x"63",
          9494 => x"6e",
          9495 => x"6f",
          9496 => x"40",
          9497 => x"38",
          9498 => x"2e",
          9499 => x"00",
          9500 => x"6c",
          9501 => x"20",
          9502 => x"65",
          9503 => x"25",
          9504 => x"20",
          9505 => x"0a",
          9506 => x"00",
          9507 => x"6c",
          9508 => x"74",
          9509 => x"65",
          9510 => x"6f",
          9511 => x"28",
          9512 => x"2e",
          9513 => x"00",
          9514 => x"74",
          9515 => x"69",
          9516 => x"61",
          9517 => x"69",
          9518 => x"69",
          9519 => x"2e",
          9520 => x"00",
          9521 => x"64",
          9522 => x"62",
          9523 => x"69",
          9524 => x"2e",
          9525 => x"00",
          9526 => x"00",
          9527 => x"00",
          9528 => x"5c",
          9529 => x"25",
          9530 => x"73",
          9531 => x"00",
          9532 => x"5c",
          9533 => x"25",
          9534 => x"00",
          9535 => x"5c",
          9536 => x"00",
          9537 => x"20",
          9538 => x"6d",
          9539 => x"2e",
          9540 => x"00",
          9541 => x"6e",
          9542 => x"2e",
          9543 => x"00",
          9544 => x"62",
          9545 => x"67",
          9546 => x"74",
          9547 => x"75",
          9548 => x"2e",
          9549 => x"00",
          9550 => x"25",
          9551 => x"64",
          9552 => x"3a",
          9553 => x"25",
          9554 => x"64",
          9555 => x"00",
          9556 => x"20",
          9557 => x"66",
          9558 => x"72",
          9559 => x"6f",
          9560 => x"00",
          9561 => x"72",
          9562 => x"53",
          9563 => x"63",
          9564 => x"69",
          9565 => x"00",
          9566 => x"65",
          9567 => x"65",
          9568 => x"6d",
          9569 => x"6d",
          9570 => x"65",
          9571 => x"00",
          9572 => x"20",
          9573 => x"53",
          9574 => x"4d",
          9575 => x"25",
          9576 => x"3a",
          9577 => x"58",
          9578 => x"00",
          9579 => x"20",
          9580 => x"41",
          9581 => x"20",
          9582 => x"25",
          9583 => x"3a",
          9584 => x"58",
          9585 => x"00",
          9586 => x"20",
          9587 => x"4e",
          9588 => x"41",
          9589 => x"25",
          9590 => x"3a",
          9591 => x"58",
          9592 => x"00",
          9593 => x"20",
          9594 => x"4d",
          9595 => x"20",
          9596 => x"25",
          9597 => x"3a",
          9598 => x"58",
          9599 => x"00",
          9600 => x"20",
          9601 => x"20",
          9602 => x"20",
          9603 => x"25",
          9604 => x"3a",
          9605 => x"58",
          9606 => x"00",
          9607 => x"20",
          9608 => x"43",
          9609 => x"20",
          9610 => x"44",
          9611 => x"63",
          9612 => x"3d",
          9613 => x"64",
          9614 => x"00",
          9615 => x"20",
          9616 => x"45",
          9617 => x"20",
          9618 => x"54",
          9619 => x"72",
          9620 => x"3d",
          9621 => x"64",
          9622 => x"00",
          9623 => x"20",
          9624 => x"52",
          9625 => x"52",
          9626 => x"43",
          9627 => x"6e",
          9628 => x"3d",
          9629 => x"64",
          9630 => x"00",
          9631 => x"20",
          9632 => x"48",
          9633 => x"45",
          9634 => x"53",
          9635 => x"00",
          9636 => x"20",
          9637 => x"49",
          9638 => x"00",
          9639 => x"20",
          9640 => x"54",
          9641 => x"00",
          9642 => x"20",
          9643 => x"0a",
          9644 => x"00",
          9645 => x"20",
          9646 => x"0a",
          9647 => x"00",
          9648 => x"72",
          9649 => x"65",
          9650 => x"00",
          9651 => x"20",
          9652 => x"20",
          9653 => x"65",
          9654 => x"65",
          9655 => x"72",
          9656 => x"64",
          9657 => x"73",
          9658 => x"25",
          9659 => x"0a",
          9660 => x"00",
          9661 => x"20",
          9662 => x"20",
          9663 => x"6f",
          9664 => x"53",
          9665 => x"74",
          9666 => x"64",
          9667 => x"73",
          9668 => x"25",
          9669 => x"0a",
          9670 => x"00",
          9671 => x"20",
          9672 => x"63",
          9673 => x"74",
          9674 => x"20",
          9675 => x"72",
          9676 => x"20",
          9677 => x"20",
          9678 => x"25",
          9679 => x"0a",
          9680 => x"00",
          9681 => x"63",
          9682 => x"00",
          9683 => x"20",
          9684 => x"20",
          9685 => x"20",
          9686 => x"20",
          9687 => x"20",
          9688 => x"20",
          9689 => x"20",
          9690 => x"25",
          9691 => x"0a",
          9692 => x"00",
          9693 => x"20",
          9694 => x"74",
          9695 => x"43",
          9696 => x"6b",
          9697 => x"65",
          9698 => x"20",
          9699 => x"20",
          9700 => x"25",
          9701 => x"30",
          9702 => x"48",
          9703 => x"00",
          9704 => x"20",
          9705 => x"41",
          9706 => x"6c",
          9707 => x"20",
          9708 => x"71",
          9709 => x"20",
          9710 => x"20",
          9711 => x"25",
          9712 => x"30",
          9713 => x"48",
          9714 => x"00",
          9715 => x"20",
          9716 => x"68",
          9717 => x"65",
          9718 => x"52",
          9719 => x"43",
          9720 => x"6b",
          9721 => x"65",
          9722 => x"25",
          9723 => x"30",
          9724 => x"48",
          9725 => x"00",
          9726 => x"6c",
          9727 => x"00",
          9728 => x"69",
          9729 => x"00",
          9730 => x"78",
          9731 => x"00",
          9732 => x"00",
          9733 => x"6d",
          9734 => x"00",
          9735 => x"6e",
          9736 => x"00",
          9737 => x"80",
          9738 => x"00",
          9739 => x"02",
          9740 => x"7c",
          9741 => x"00",
          9742 => x"03",
          9743 => x"78",
          9744 => x"00",
          9745 => x"04",
          9746 => x"74",
          9747 => x"00",
          9748 => x"05",
          9749 => x"70",
          9750 => x"00",
          9751 => x"06",
          9752 => x"6c",
          9753 => x"00",
          9754 => x"07",
          9755 => x"68",
          9756 => x"00",
          9757 => x"01",
          9758 => x"64",
          9759 => x"00",
          9760 => x"08",
          9761 => x"60",
          9762 => x"00",
          9763 => x"0b",
          9764 => x"5c",
          9765 => x"00",
          9766 => x"09",
          9767 => x"58",
          9768 => x"00",
          9769 => x"0a",
          9770 => x"54",
          9771 => x"00",
          9772 => x"0d",
          9773 => x"50",
          9774 => x"00",
          9775 => x"0c",
          9776 => x"4c",
          9777 => x"00",
          9778 => x"0e",
          9779 => x"48",
          9780 => x"00",
          9781 => x"0f",
          9782 => x"44",
          9783 => x"00",
          9784 => x"0f",
          9785 => x"40",
          9786 => x"00",
          9787 => x"10",
          9788 => x"3c",
          9789 => x"00",
          9790 => x"11",
          9791 => x"38",
          9792 => x"00",
          9793 => x"12",
          9794 => x"34",
          9795 => x"00",
          9796 => x"13",
          9797 => x"30",
          9798 => x"00",
          9799 => x"14",
          9800 => x"2c",
          9801 => x"00",
          9802 => x"15",
          9803 => x"00",
          9804 => x"00",
          9805 => x"00",
          9806 => x"00",
          9807 => x"7e",
          9808 => x"7e",
          9809 => x"7e",
          9810 => x"00",
          9811 => x"7e",
          9812 => x"7e",
          9813 => x"7e",
          9814 => x"00",
          9815 => x"00",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"00",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"00",
          9824 => x"00",
          9825 => x"74",
          9826 => x"00",
          9827 => x"74",
          9828 => x"00",
          9829 => x"00",
          9830 => x"64",
          9831 => x"73",
          9832 => x"00",
          9833 => x"6c",
          9834 => x"74",
          9835 => x"65",
          9836 => x"20",
          9837 => x"20",
          9838 => x"74",
          9839 => x"20",
          9840 => x"65",
          9841 => x"20",
          9842 => x"2e",
          9843 => x"00",
          9844 => x"6e",
          9845 => x"6f",
          9846 => x"2f",
          9847 => x"61",
          9848 => x"68",
          9849 => x"6f",
          9850 => x"66",
          9851 => x"2c",
          9852 => x"73",
          9853 => x"69",
          9854 => x"00",
          9855 => x"00",
          9856 => x"2c",
          9857 => x"3d",
          9858 => x"5d",
          9859 => x"00",
          9860 => x"00",
          9861 => x"33",
          9862 => x"00",
          9863 => x"4d",
          9864 => x"53",
          9865 => x"00",
          9866 => x"4e",
          9867 => x"20",
          9868 => x"46",
          9869 => x"32",
          9870 => x"00",
          9871 => x"4e",
          9872 => x"20",
          9873 => x"46",
          9874 => x"20",
          9875 => x"00",
          9876 => x"fc",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"41",
          9881 => x"80",
          9882 => x"49",
          9883 => x"8f",
          9884 => x"4f",
          9885 => x"55",
          9886 => x"9b",
          9887 => x"9f",
          9888 => x"55",
          9889 => x"a7",
          9890 => x"ab",
          9891 => x"af",
          9892 => x"b3",
          9893 => x"b7",
          9894 => x"bb",
          9895 => x"bf",
          9896 => x"c3",
          9897 => x"c7",
          9898 => x"cb",
          9899 => x"cf",
          9900 => x"d3",
          9901 => x"d7",
          9902 => x"db",
          9903 => x"df",
          9904 => x"e3",
          9905 => x"e7",
          9906 => x"eb",
          9907 => x"ef",
          9908 => x"f3",
          9909 => x"f7",
          9910 => x"fb",
          9911 => x"ff",
          9912 => x"3b",
          9913 => x"2f",
          9914 => x"3a",
          9915 => x"7c",
          9916 => x"00",
          9917 => x"04",
          9918 => x"40",
          9919 => x"00",
          9920 => x"00",
          9921 => x"02",
          9922 => x"08",
          9923 => x"20",
          9924 => x"00",
          9925 => x"00",
          9926 => x"d0",
          9927 => x"00",
          9928 => x"00",
          9929 => x"00",
          9930 => x"d8",
          9931 => x"00",
          9932 => x"00",
          9933 => x"00",
          9934 => x"e0",
          9935 => x"00",
          9936 => x"00",
          9937 => x"00",
          9938 => x"e8",
          9939 => x"00",
          9940 => x"00",
          9941 => x"00",
          9942 => x"f0",
          9943 => x"00",
          9944 => x"00",
          9945 => x"00",
          9946 => x"f8",
          9947 => x"00",
          9948 => x"00",
          9949 => x"00",
          9950 => x"00",
          9951 => x"00",
          9952 => x"00",
          9953 => x"00",
          9954 => x"08",
          9955 => x"00",
          9956 => x"00",
          9957 => x"00",
          9958 => x"10",
          9959 => x"00",
          9960 => x"00",
          9961 => x"00",
          9962 => x"18",
          9963 => x"00",
          9964 => x"00",
          9965 => x"00",
          9966 => x"1c",
          9967 => x"00",
          9968 => x"00",
          9969 => x"00",
          9970 => x"20",
          9971 => x"00",
          9972 => x"00",
          9973 => x"00",
          9974 => x"24",
          9975 => x"00",
          9976 => x"00",
          9977 => x"00",
          9978 => x"28",
          9979 => x"00",
          9980 => x"00",
          9981 => x"00",
          9982 => x"2c",
          9983 => x"00",
          9984 => x"00",
          9985 => x"00",
          9986 => x"30",
          9987 => x"00",
          9988 => x"00",
          9989 => x"00",
          9990 => x"34",
          9991 => x"00",
          9992 => x"00",
          9993 => x"00",
          9994 => x"3c",
          9995 => x"00",
          9996 => x"00",
          9997 => x"00",
          9998 => x"40",
          9999 => x"00",
         10000 => x"00",
         10001 => x"00",
         10002 => x"48",
         10003 => x"00",
         10004 => x"00",
         10005 => x"00",
         10006 => x"50",
         10007 => x"00",
         10008 => x"00",
         10009 => x"00",
         10010 => x"58",
         10011 => x"00",
         10012 => x"00",
         10013 => x"00",
         10014 => x"60",
         10015 => x"00",
         10016 => x"00",
         10017 => x"00",
         10018 => x"68",
         10019 => x"00",
         10020 => x"00",
         10021 => x"00",
         10022 => x"70",
         10023 => x"00",
         10024 => x"00",
         10025 => x"00",
         10026 => x"78",
         10027 => x"00",
         10028 => x"00",
         10029 => x"00",
         10030 => x"00",
         10031 => x"00",
         10032 => x"ff",
         10033 => x"00",
         10034 => x"ff",
         10035 => x"00",
         10036 => x"ff",
         10037 => x"00",
         10038 => x"00",
         10039 => x"00",
         10040 => x"ff",
         10041 => x"00",
         10042 => x"00",
         10043 => x"00",
         10044 => x"00",
         10045 => x"00",
         10046 => x"00",
         10047 => x"00",
         10048 => x"00",
         10049 => x"01",
         10050 => x"01",
         10051 => x"01",
         10052 => x"00",
         10053 => x"00",
         10054 => x"00",
         10055 => x"00",
         10056 => x"00",
         10057 => x"00",
         10058 => x"00",
         10059 => x"00",
         10060 => x"00",
         10061 => x"00",
         10062 => x"00",
         10063 => x"00",
         10064 => x"00",
         10065 => x"00",
         10066 => x"00",
         10067 => x"00",
         10068 => x"00",
         10069 => x"00",
         10070 => x"00",
         10071 => x"00",
         10072 => x"00",
         10073 => x"00",
         10074 => x"00",
         10075 => x"00",
         10076 => x"00",
         10077 => x"84",
         10078 => x"00",
         10079 => x"8c",
         10080 => x"00",
         10081 => x"94",
         10082 => x"00",
         10083 => x"00",
         10084 => x"00",
         10085 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"83",
             1 => x"0b",
             2 => x"b7",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"92",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"82",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"80",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"80",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a4",
           270 => x"0b",
           271 => x"0b",
           272 => x"c2",
           273 => x"0b",
           274 => x"0b",
           275 => x"e0",
           276 => x"0b",
           277 => x"0b",
           278 => x"fe",
           279 => x"0b",
           280 => x"0b",
           281 => x"9c",
           282 => x"0b",
           283 => x"0b",
           284 => x"bb",
           285 => x"0b",
           286 => x"0b",
           287 => x"db",
           288 => x"0b",
           289 => x"0b",
           290 => x"fb",
           291 => x"0b",
           292 => x"0b",
           293 => x"9b",
           294 => x"0b",
           295 => x"0b",
           296 => x"bb",
           297 => x"0b",
           298 => x"0b",
           299 => x"db",
           300 => x"0b",
           301 => x"0b",
           302 => x"fb",
           303 => x"0b",
           304 => x"0b",
           305 => x"9b",
           306 => x"0b",
           307 => x"0b",
           308 => x"bb",
           309 => x"0b",
           310 => x"0b",
           311 => x"db",
           312 => x"0b",
           313 => x"0b",
           314 => x"fb",
           315 => x"0b",
           316 => x"0b",
           317 => x"9b",
           318 => x"0b",
           319 => x"0b",
           320 => x"bb",
           321 => x"0b",
           322 => x"0b",
           323 => x"db",
           324 => x"0b",
           325 => x"0b",
           326 => x"fb",
           327 => x"0b",
           328 => x"0b",
           329 => x"9b",
           330 => x"0b",
           331 => x"0b",
           332 => x"bb",
           333 => x"0b",
           334 => x"0b",
           335 => x"db",
           336 => x"0b",
           337 => x"0b",
           338 => x"fb",
           339 => x"0b",
           340 => x"0b",
           341 => x"9b",
           342 => x"0b",
           343 => x"0b",
           344 => x"bb",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"bb",
           386 => x"f8",
           387 => x"bb",
           388 => x"e0",
           389 => x"bb",
           390 => x"d2",
           391 => x"a4",
           392 => x"90",
           393 => x"a4",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"82",
           399 => x"82",
           400 => x"82",
           401 => x"94",
           402 => x"bb",
           403 => x"e0",
           404 => x"bb",
           405 => x"e2",
           406 => x"a4",
           407 => x"90",
           408 => x"a4",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"82",
           414 => x"82",
           415 => x"82",
           416 => x"93",
           417 => x"bb",
           418 => x"e0",
           419 => x"bb",
           420 => x"be",
           421 => x"a4",
           422 => x"90",
           423 => x"a4",
           424 => x"2d",
           425 => x"08",
           426 => x"04",
           427 => x"0c",
           428 => x"2d",
           429 => x"08",
           430 => x"04",
           431 => x"0c",
           432 => x"2d",
           433 => x"08",
           434 => x"04",
           435 => x"0c",
           436 => x"2d",
           437 => x"08",
           438 => x"04",
           439 => x"0c",
           440 => x"2d",
           441 => x"08",
           442 => x"04",
           443 => x"0c",
           444 => x"2d",
           445 => x"08",
           446 => x"04",
           447 => x"0c",
           448 => x"2d",
           449 => x"08",
           450 => x"04",
           451 => x"0c",
           452 => x"2d",
           453 => x"08",
           454 => x"04",
           455 => x"0c",
           456 => x"2d",
           457 => x"08",
           458 => x"04",
           459 => x"0c",
           460 => x"2d",
           461 => x"08",
           462 => x"04",
           463 => x"0c",
           464 => x"2d",
           465 => x"08",
           466 => x"04",
           467 => x"0c",
           468 => x"2d",
           469 => x"08",
           470 => x"04",
           471 => x"0c",
           472 => x"2d",
           473 => x"08",
           474 => x"04",
           475 => x"0c",
           476 => x"2d",
           477 => x"08",
           478 => x"04",
           479 => x"0c",
           480 => x"2d",
           481 => x"08",
           482 => x"04",
           483 => x"0c",
           484 => x"2d",
           485 => x"08",
           486 => x"04",
           487 => x"0c",
           488 => x"2d",
           489 => x"08",
           490 => x"04",
           491 => x"0c",
           492 => x"2d",
           493 => x"08",
           494 => x"04",
           495 => x"0c",
           496 => x"2d",
           497 => x"08",
           498 => x"04",
           499 => x"0c",
           500 => x"2d",
           501 => x"08",
           502 => x"04",
           503 => x"0c",
           504 => x"2d",
           505 => x"08",
           506 => x"04",
           507 => x"0c",
           508 => x"2d",
           509 => x"08",
           510 => x"04",
           511 => x"0c",
           512 => x"2d",
           513 => x"08",
           514 => x"04",
           515 => x"0c",
           516 => x"2d",
           517 => x"08",
           518 => x"04",
           519 => x"0c",
           520 => x"2d",
           521 => x"08",
           522 => x"04",
           523 => x"0c",
           524 => x"2d",
           525 => x"08",
           526 => x"04",
           527 => x"0c",
           528 => x"2d",
           529 => x"08",
           530 => x"04",
           531 => x"0c",
           532 => x"2d",
           533 => x"08",
           534 => x"04",
           535 => x"0c",
           536 => x"2d",
           537 => x"08",
           538 => x"04",
           539 => x"0c",
           540 => x"2d",
           541 => x"08",
           542 => x"04",
           543 => x"0c",
           544 => x"2d",
           545 => x"08",
           546 => x"04",
           547 => x"0c",
           548 => x"2d",
           549 => x"08",
           550 => x"04",
           551 => x"0c",
           552 => x"2d",
           553 => x"08",
           554 => x"04",
           555 => x"0c",
           556 => x"2d",
           557 => x"08",
           558 => x"04",
           559 => x"0c",
           560 => x"2d",
           561 => x"08",
           562 => x"04",
           563 => x"0c",
           564 => x"2d",
           565 => x"08",
           566 => x"04",
           567 => x"0c",
           568 => x"2d",
           569 => x"08",
           570 => x"04",
           571 => x"0c",
           572 => x"2d",
           573 => x"08",
           574 => x"04",
           575 => x"0c",
           576 => x"2d",
           577 => x"08",
           578 => x"04",
           579 => x"0c",
           580 => x"2d",
           581 => x"08",
           582 => x"04",
           583 => x"0c",
           584 => x"2d",
           585 => x"08",
           586 => x"04",
           587 => x"0c",
           588 => x"2d",
           589 => x"08",
           590 => x"04",
           591 => x"0c",
           592 => x"2d",
           593 => x"08",
           594 => x"04",
           595 => x"0c",
           596 => x"2d",
           597 => x"08",
           598 => x"04",
           599 => x"00",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"53",
           608 => x"00",
           609 => x"06",
           610 => x"09",
           611 => x"05",
           612 => x"2b",
           613 => x"06",
           614 => x"04",
           615 => x"72",
           616 => x"05",
           617 => x"05",
           618 => x"72",
           619 => x"53",
           620 => x"51",
           621 => x"04",
           622 => x"70",
           623 => x"27",
           624 => x"71",
           625 => x"53",
           626 => x"0b",
           627 => x"8c",
           628 => x"f2",
           629 => x"82",
           630 => x"02",
           631 => x"0c",
           632 => x"82",
           633 => x"8c",
           634 => x"bb",
           635 => x"05",
           636 => x"a4",
           637 => x"08",
           638 => x"a4",
           639 => x"08",
           640 => x"ec",
           641 => x"84",
           642 => x"bb",
           643 => x"82",
           644 => x"f8",
           645 => x"bb",
           646 => x"05",
           647 => x"bb",
           648 => x"54",
           649 => x"82",
           650 => x"04",
           651 => x"08",
           652 => x"a4",
           653 => x"0d",
           654 => x"08",
           655 => x"85",
           656 => x"81",
           657 => x"06",
           658 => x"52",
           659 => x"80",
           660 => x"a4",
           661 => x"08",
           662 => x"8d",
           663 => x"82",
           664 => x"f4",
           665 => x"c4",
           666 => x"a4",
           667 => x"08",
           668 => x"bb",
           669 => x"05",
           670 => x"82",
           671 => x"f8",
           672 => x"bb",
           673 => x"05",
           674 => x"a4",
           675 => x"0c",
           676 => x"08",
           677 => x"8a",
           678 => x"38",
           679 => x"bb",
           680 => x"05",
           681 => x"e9",
           682 => x"a4",
           683 => x"08",
           684 => x"3f",
           685 => x"08",
           686 => x"a4",
           687 => x"0c",
           688 => x"a4",
           689 => x"08",
           690 => x"81",
           691 => x"80",
           692 => x"a4",
           693 => x"0c",
           694 => x"82",
           695 => x"fc",
           696 => x"bb",
           697 => x"05",
           698 => x"71",
           699 => x"bb",
           700 => x"05",
           701 => x"82",
           702 => x"8c",
           703 => x"bb",
           704 => x"05",
           705 => x"82",
           706 => x"fc",
           707 => x"80",
           708 => x"a4",
           709 => x"08",
           710 => x"34",
           711 => x"08",
           712 => x"70",
           713 => x"08",
           714 => x"52",
           715 => x"08",
           716 => x"82",
           717 => x"87",
           718 => x"bb",
           719 => x"82",
           720 => x"02",
           721 => x"0c",
           722 => x"86",
           723 => x"a4",
           724 => x"34",
           725 => x"08",
           726 => x"82",
           727 => x"e0",
           728 => x"0a",
           729 => x"a4",
           730 => x"0c",
           731 => x"08",
           732 => x"82",
           733 => x"fc",
           734 => x"bb",
           735 => x"05",
           736 => x"bb",
           737 => x"05",
           738 => x"bb",
           739 => x"05",
           740 => x"54",
           741 => x"82",
           742 => x"70",
           743 => x"08",
           744 => x"82",
           745 => x"ec",
           746 => x"bb",
           747 => x"05",
           748 => x"54",
           749 => x"82",
           750 => x"dc",
           751 => x"82",
           752 => x"54",
           753 => x"82",
           754 => x"04",
           755 => x"08",
           756 => x"a4",
           757 => x"0d",
           758 => x"08",
           759 => x"82",
           760 => x"fc",
           761 => x"bb",
           762 => x"05",
           763 => x"bb",
           764 => x"05",
           765 => x"bb",
           766 => x"05",
           767 => x"a3",
           768 => x"98",
           769 => x"bb",
           770 => x"05",
           771 => x"a4",
           772 => x"08",
           773 => x"98",
           774 => x"87",
           775 => x"bb",
           776 => x"82",
           777 => x"02",
           778 => x"0c",
           779 => x"80",
           780 => x"a4",
           781 => x"23",
           782 => x"08",
           783 => x"53",
           784 => x"14",
           785 => x"a4",
           786 => x"08",
           787 => x"70",
           788 => x"81",
           789 => x"06",
           790 => x"51",
           791 => x"2e",
           792 => x"0b",
           793 => x"08",
           794 => x"96",
           795 => x"bb",
           796 => x"05",
           797 => x"33",
           798 => x"bb",
           799 => x"05",
           800 => x"ff",
           801 => x"80",
           802 => x"38",
           803 => x"08",
           804 => x"81",
           805 => x"a4",
           806 => x"0c",
           807 => x"08",
           808 => x"70",
           809 => x"53",
           810 => x"95",
           811 => x"bb",
           812 => x"05",
           813 => x"73",
           814 => x"38",
           815 => x"08",
           816 => x"53",
           817 => x"81",
           818 => x"bb",
           819 => x"05",
           820 => x"b0",
           821 => x"06",
           822 => x"82",
           823 => x"e8",
           824 => x"98",
           825 => x"2c",
           826 => x"72",
           827 => x"bb",
           828 => x"05",
           829 => x"2a",
           830 => x"70",
           831 => x"51",
           832 => x"80",
           833 => x"82",
           834 => x"e4",
           835 => x"82",
           836 => x"53",
           837 => x"a4",
           838 => x"23",
           839 => x"82",
           840 => x"e8",
           841 => x"98",
           842 => x"2c",
           843 => x"2b",
           844 => x"11",
           845 => x"53",
           846 => x"72",
           847 => x"08",
           848 => x"82",
           849 => x"e8",
           850 => x"82",
           851 => x"f8",
           852 => x"15",
           853 => x"51",
           854 => x"bb",
           855 => x"05",
           856 => x"a4",
           857 => x"33",
           858 => x"70",
           859 => x"51",
           860 => x"25",
           861 => x"ff",
           862 => x"a4",
           863 => x"34",
           864 => x"08",
           865 => x"70",
           866 => x"81",
           867 => x"53",
           868 => x"38",
           869 => x"08",
           870 => x"70",
           871 => x"90",
           872 => x"2c",
           873 => x"51",
           874 => x"53",
           875 => x"a4",
           876 => x"23",
           877 => x"82",
           878 => x"e4",
           879 => x"83",
           880 => x"06",
           881 => x"72",
           882 => x"38",
           883 => x"08",
           884 => x"70",
           885 => x"98",
           886 => x"53",
           887 => x"81",
           888 => x"a4",
           889 => x"34",
           890 => x"08",
           891 => x"e0",
           892 => x"a4",
           893 => x"0c",
           894 => x"a4",
           895 => x"08",
           896 => x"92",
           897 => x"bb",
           898 => x"05",
           899 => x"2b",
           900 => x"11",
           901 => x"51",
           902 => x"04",
           903 => x"08",
           904 => x"70",
           905 => x"53",
           906 => x"a4",
           907 => x"23",
           908 => x"08",
           909 => x"70",
           910 => x"53",
           911 => x"a4",
           912 => x"23",
           913 => x"82",
           914 => x"e4",
           915 => x"81",
           916 => x"53",
           917 => x"a4",
           918 => x"23",
           919 => x"82",
           920 => x"e4",
           921 => x"80",
           922 => x"53",
           923 => x"a4",
           924 => x"23",
           925 => x"82",
           926 => x"e4",
           927 => x"88",
           928 => x"72",
           929 => x"08",
           930 => x"80",
           931 => x"a4",
           932 => x"34",
           933 => x"82",
           934 => x"e4",
           935 => x"84",
           936 => x"72",
           937 => x"08",
           938 => x"fb",
           939 => x"0b",
           940 => x"08",
           941 => x"82",
           942 => x"ec",
           943 => x"11",
           944 => x"82",
           945 => x"ec",
           946 => x"e3",
           947 => x"a4",
           948 => x"34",
           949 => x"82",
           950 => x"90",
           951 => x"bb",
           952 => x"05",
           953 => x"82",
           954 => x"90",
           955 => x"08",
           956 => x"82",
           957 => x"fc",
           958 => x"bb",
           959 => x"05",
           960 => x"51",
           961 => x"bb",
           962 => x"05",
           963 => x"39",
           964 => x"08",
           965 => x"82",
           966 => x"90",
           967 => x"05",
           968 => x"08",
           969 => x"70",
           970 => x"a4",
           971 => x"0c",
           972 => x"08",
           973 => x"70",
           974 => x"81",
           975 => x"51",
           976 => x"2e",
           977 => x"bb",
           978 => x"05",
           979 => x"2b",
           980 => x"2c",
           981 => x"a4",
           982 => x"08",
           983 => x"fa",
           984 => x"98",
           985 => x"82",
           986 => x"f4",
           987 => x"39",
           988 => x"08",
           989 => x"51",
           990 => x"82",
           991 => x"53",
           992 => x"a4",
           993 => x"23",
           994 => x"08",
           995 => x"53",
           996 => x"08",
           997 => x"73",
           998 => x"54",
           999 => x"a4",
          1000 => x"23",
          1001 => x"82",
          1002 => x"90",
          1003 => x"bb",
          1004 => x"05",
          1005 => x"82",
          1006 => x"90",
          1007 => x"08",
          1008 => x"08",
          1009 => x"82",
          1010 => x"e4",
          1011 => x"83",
          1012 => x"06",
          1013 => x"53",
          1014 => x"ab",
          1015 => x"a4",
          1016 => x"33",
          1017 => x"53",
          1018 => x"53",
          1019 => x"08",
          1020 => x"52",
          1021 => x"3f",
          1022 => x"08",
          1023 => x"bb",
          1024 => x"05",
          1025 => x"82",
          1026 => x"fc",
          1027 => x"a7",
          1028 => x"bb",
          1029 => x"72",
          1030 => x"08",
          1031 => x"82",
          1032 => x"ec",
          1033 => x"82",
          1034 => x"f4",
          1035 => x"71",
          1036 => x"72",
          1037 => x"08",
          1038 => x"8a",
          1039 => x"bb",
          1040 => x"05",
          1041 => x"2a",
          1042 => x"51",
          1043 => x"80",
          1044 => x"82",
          1045 => x"90",
          1046 => x"bb",
          1047 => x"05",
          1048 => x"82",
          1049 => x"90",
          1050 => x"08",
          1051 => x"08",
          1052 => x"53",
          1053 => x"bb",
          1054 => x"05",
          1055 => x"a4",
          1056 => x"08",
          1057 => x"bb",
          1058 => x"05",
          1059 => x"82",
          1060 => x"dc",
          1061 => x"82",
          1062 => x"dc",
          1063 => x"bb",
          1064 => x"05",
          1065 => x"a4",
          1066 => x"08",
          1067 => x"38",
          1068 => x"08",
          1069 => x"70",
          1070 => x"53",
          1071 => x"a4",
          1072 => x"23",
          1073 => x"08",
          1074 => x"30",
          1075 => x"08",
          1076 => x"82",
          1077 => x"e4",
          1078 => x"ff",
          1079 => x"53",
          1080 => x"a4",
          1081 => x"23",
          1082 => x"88",
          1083 => x"a4",
          1084 => x"23",
          1085 => x"bb",
          1086 => x"05",
          1087 => x"c0",
          1088 => x"72",
          1089 => x"08",
          1090 => x"80",
          1091 => x"bb",
          1092 => x"05",
          1093 => x"82",
          1094 => x"f4",
          1095 => x"bb",
          1096 => x"05",
          1097 => x"2a",
          1098 => x"51",
          1099 => x"80",
          1100 => x"82",
          1101 => x"90",
          1102 => x"bb",
          1103 => x"05",
          1104 => x"82",
          1105 => x"90",
          1106 => x"08",
          1107 => x"08",
          1108 => x"53",
          1109 => x"bb",
          1110 => x"05",
          1111 => x"a4",
          1112 => x"08",
          1113 => x"bb",
          1114 => x"05",
          1115 => x"82",
          1116 => x"d8",
          1117 => x"82",
          1118 => x"d8",
          1119 => x"bb",
          1120 => x"05",
          1121 => x"a4",
          1122 => x"22",
          1123 => x"51",
          1124 => x"bb",
          1125 => x"05",
          1126 => x"a8",
          1127 => x"a4",
          1128 => x"0c",
          1129 => x"08",
          1130 => x"82",
          1131 => x"f4",
          1132 => x"bb",
          1133 => x"05",
          1134 => x"70",
          1135 => x"55",
          1136 => x"82",
          1137 => x"53",
          1138 => x"82",
          1139 => x"f0",
          1140 => x"bb",
          1141 => x"05",
          1142 => x"a4",
          1143 => x"08",
          1144 => x"53",
          1145 => x"a4",
          1146 => x"a4",
          1147 => x"08",
          1148 => x"54",
          1149 => x"08",
          1150 => x"70",
          1151 => x"51",
          1152 => x"82",
          1153 => x"d0",
          1154 => x"39",
          1155 => x"08",
          1156 => x"53",
          1157 => x"11",
          1158 => x"82",
          1159 => x"d0",
          1160 => x"bb",
          1161 => x"05",
          1162 => x"bb",
          1163 => x"05",
          1164 => x"82",
          1165 => x"f0",
          1166 => x"05",
          1167 => x"08",
          1168 => x"82",
          1169 => x"f4",
          1170 => x"53",
          1171 => x"08",
          1172 => x"52",
          1173 => x"3f",
          1174 => x"08",
          1175 => x"a4",
          1176 => x"0c",
          1177 => x"a4",
          1178 => x"08",
          1179 => x"38",
          1180 => x"82",
          1181 => x"f0",
          1182 => x"bb",
          1183 => x"72",
          1184 => x"75",
          1185 => x"72",
          1186 => x"08",
          1187 => x"82",
          1188 => x"e4",
          1189 => x"b2",
          1190 => x"72",
          1191 => x"38",
          1192 => x"08",
          1193 => x"ff",
          1194 => x"72",
          1195 => x"08",
          1196 => x"82",
          1197 => x"e4",
          1198 => x"86",
          1199 => x"06",
          1200 => x"72",
          1201 => x"e7",
          1202 => x"a4",
          1203 => x"22",
          1204 => x"82",
          1205 => x"cc",
          1206 => x"bb",
          1207 => x"05",
          1208 => x"82",
          1209 => x"cc",
          1210 => x"bb",
          1211 => x"05",
          1212 => x"72",
          1213 => x"81",
          1214 => x"82",
          1215 => x"cc",
          1216 => x"05",
          1217 => x"bb",
          1218 => x"05",
          1219 => x"82",
          1220 => x"cc",
          1221 => x"05",
          1222 => x"bb",
          1223 => x"05",
          1224 => x"a4",
          1225 => x"22",
          1226 => x"08",
          1227 => x"82",
          1228 => x"e4",
          1229 => x"83",
          1230 => x"06",
          1231 => x"72",
          1232 => x"d0",
          1233 => x"a4",
          1234 => x"33",
          1235 => x"70",
          1236 => x"bb",
          1237 => x"05",
          1238 => x"51",
          1239 => x"24",
          1240 => x"bb",
          1241 => x"05",
          1242 => x"06",
          1243 => x"82",
          1244 => x"e4",
          1245 => x"39",
          1246 => x"08",
          1247 => x"53",
          1248 => x"08",
          1249 => x"73",
          1250 => x"54",
          1251 => x"a4",
          1252 => x"34",
          1253 => x"08",
          1254 => x"70",
          1255 => x"81",
          1256 => x"53",
          1257 => x"b1",
          1258 => x"a4",
          1259 => x"33",
          1260 => x"70",
          1261 => x"90",
          1262 => x"2c",
          1263 => x"51",
          1264 => x"82",
          1265 => x"ec",
          1266 => x"75",
          1267 => x"72",
          1268 => x"08",
          1269 => x"af",
          1270 => x"a4",
          1271 => x"33",
          1272 => x"70",
          1273 => x"90",
          1274 => x"2c",
          1275 => x"51",
          1276 => x"82",
          1277 => x"ec",
          1278 => x"75",
          1279 => x"72",
          1280 => x"08",
          1281 => x"82",
          1282 => x"e4",
          1283 => x"83",
          1284 => x"53",
          1285 => x"82",
          1286 => x"ec",
          1287 => x"11",
          1288 => x"82",
          1289 => x"ec",
          1290 => x"90",
          1291 => x"2c",
          1292 => x"73",
          1293 => x"82",
          1294 => x"88",
          1295 => x"a0",
          1296 => x"3f",
          1297 => x"bb",
          1298 => x"05",
          1299 => x"2a",
          1300 => x"51",
          1301 => x"80",
          1302 => x"82",
          1303 => x"88",
          1304 => x"ad",
          1305 => x"3f",
          1306 => x"82",
          1307 => x"e4",
          1308 => x"84",
          1309 => x"06",
          1310 => x"72",
          1311 => x"38",
          1312 => x"08",
          1313 => x"52",
          1314 => x"c7",
          1315 => x"82",
          1316 => x"e4",
          1317 => x"85",
          1318 => x"06",
          1319 => x"72",
          1320 => x"38",
          1321 => x"08",
          1322 => x"52",
          1323 => x"a3",
          1324 => x"a4",
          1325 => x"22",
          1326 => x"70",
          1327 => x"51",
          1328 => x"2e",
          1329 => x"bb",
          1330 => x"05",
          1331 => x"51",
          1332 => x"82",
          1333 => x"f4",
          1334 => x"72",
          1335 => x"81",
          1336 => x"82",
          1337 => x"88",
          1338 => x"82",
          1339 => x"f8",
          1340 => x"94",
          1341 => x"bb",
          1342 => x"05",
          1343 => x"2a",
          1344 => x"51",
          1345 => x"80",
          1346 => x"82",
          1347 => x"ec",
          1348 => x"11",
          1349 => x"82",
          1350 => x"ec",
          1351 => x"90",
          1352 => x"2c",
          1353 => x"73",
          1354 => x"82",
          1355 => x"88",
          1356 => x"b0",
          1357 => x"3f",
          1358 => x"bb",
          1359 => x"05",
          1360 => x"2a",
          1361 => x"51",
          1362 => x"80",
          1363 => x"82",
          1364 => x"e8",
          1365 => x"11",
          1366 => x"82",
          1367 => x"e8",
          1368 => x"98",
          1369 => x"2c",
          1370 => x"73",
          1371 => x"82",
          1372 => x"88",
          1373 => x"b0",
          1374 => x"3f",
          1375 => x"bb",
          1376 => x"05",
          1377 => x"2a",
          1378 => x"51",
          1379 => x"b0",
          1380 => x"a4",
          1381 => x"22",
          1382 => x"54",
          1383 => x"a4",
          1384 => x"23",
          1385 => x"70",
          1386 => x"53",
          1387 => x"90",
          1388 => x"a4",
          1389 => x"08",
          1390 => x"93",
          1391 => x"39",
          1392 => x"08",
          1393 => x"53",
          1394 => x"2e",
          1395 => x"97",
          1396 => x"a4",
          1397 => x"08",
          1398 => x"a4",
          1399 => x"33",
          1400 => x"3f",
          1401 => x"82",
          1402 => x"f8",
          1403 => x"72",
          1404 => x"09",
          1405 => x"cb",
          1406 => x"a4",
          1407 => x"22",
          1408 => x"53",
          1409 => x"a4",
          1410 => x"23",
          1411 => x"ff",
          1412 => x"83",
          1413 => x"81",
          1414 => x"bb",
          1415 => x"05",
          1416 => x"bb",
          1417 => x"05",
          1418 => x"52",
          1419 => x"08",
          1420 => x"81",
          1421 => x"a4",
          1422 => x"0c",
          1423 => x"3f",
          1424 => x"82",
          1425 => x"f8",
          1426 => x"72",
          1427 => x"09",
          1428 => x"cb",
          1429 => x"a4",
          1430 => x"22",
          1431 => x"53",
          1432 => x"a4",
          1433 => x"23",
          1434 => x"ff",
          1435 => x"83",
          1436 => x"80",
          1437 => x"bb",
          1438 => x"05",
          1439 => x"bb",
          1440 => x"05",
          1441 => x"52",
          1442 => x"3f",
          1443 => x"08",
          1444 => x"81",
          1445 => x"a4",
          1446 => x"0c",
          1447 => x"82",
          1448 => x"f0",
          1449 => x"bb",
          1450 => x"38",
          1451 => x"08",
          1452 => x"52",
          1453 => x"08",
          1454 => x"ff",
          1455 => x"a4",
          1456 => x"0c",
          1457 => x"08",
          1458 => x"70",
          1459 => x"91",
          1460 => x"39",
          1461 => x"08",
          1462 => x"70",
          1463 => x"81",
          1464 => x"53",
          1465 => x"80",
          1466 => x"bb",
          1467 => x"05",
          1468 => x"54",
          1469 => x"bb",
          1470 => x"05",
          1471 => x"2b",
          1472 => x"51",
          1473 => x"25",
          1474 => x"bb",
          1475 => x"05",
          1476 => x"51",
          1477 => x"d2",
          1478 => x"a4",
          1479 => x"08",
          1480 => x"a4",
          1481 => x"33",
          1482 => x"3f",
          1483 => x"bb",
          1484 => x"05",
          1485 => x"39",
          1486 => x"08",
          1487 => x"53",
          1488 => x"09",
          1489 => x"38",
          1490 => x"bb",
          1491 => x"05",
          1492 => x"82",
          1493 => x"ec",
          1494 => x"0b",
          1495 => x"08",
          1496 => x"8a",
          1497 => x"a4",
          1498 => x"23",
          1499 => x"82",
          1500 => x"88",
          1501 => x"82",
          1502 => x"f8",
          1503 => x"8f",
          1504 => x"ea",
          1505 => x"a4",
          1506 => x"08",
          1507 => x"70",
          1508 => x"08",
          1509 => x"51",
          1510 => x"a4",
          1511 => x"08",
          1512 => x"0c",
          1513 => x"82",
          1514 => x"04",
          1515 => x"08",
          1516 => x"a4",
          1517 => x"0d",
          1518 => x"bb",
          1519 => x"05",
          1520 => x"a4",
          1521 => x"08",
          1522 => x"0c",
          1523 => x"08",
          1524 => x"70",
          1525 => x"72",
          1526 => x"82",
          1527 => x"f8",
          1528 => x"81",
          1529 => x"72",
          1530 => x"81",
          1531 => x"82",
          1532 => x"88",
          1533 => x"08",
          1534 => x"0c",
          1535 => x"82",
          1536 => x"f8",
          1537 => x"72",
          1538 => x"81",
          1539 => x"81",
          1540 => x"a4",
          1541 => x"34",
          1542 => x"08",
          1543 => x"70",
          1544 => x"71",
          1545 => x"51",
          1546 => x"82",
          1547 => x"f8",
          1548 => x"bb",
          1549 => x"05",
          1550 => x"b0",
          1551 => x"06",
          1552 => x"82",
          1553 => x"88",
          1554 => x"08",
          1555 => x"0c",
          1556 => x"53",
          1557 => x"bb",
          1558 => x"05",
          1559 => x"a4",
          1560 => x"33",
          1561 => x"08",
          1562 => x"82",
          1563 => x"e8",
          1564 => x"e2",
          1565 => x"82",
          1566 => x"e8",
          1567 => x"f8",
          1568 => x"80",
          1569 => x"0b",
          1570 => x"08",
          1571 => x"82",
          1572 => x"88",
          1573 => x"08",
          1574 => x"0c",
          1575 => x"53",
          1576 => x"bb",
          1577 => x"05",
          1578 => x"39",
          1579 => x"bb",
          1580 => x"05",
          1581 => x"a4",
          1582 => x"08",
          1583 => x"05",
          1584 => x"08",
          1585 => x"33",
          1586 => x"08",
          1587 => x"80",
          1588 => x"bb",
          1589 => x"05",
          1590 => x"a0",
          1591 => x"81",
          1592 => x"a4",
          1593 => x"0c",
          1594 => x"82",
          1595 => x"f8",
          1596 => x"af",
          1597 => x"38",
          1598 => x"08",
          1599 => x"53",
          1600 => x"83",
          1601 => x"80",
          1602 => x"a4",
          1603 => x"0c",
          1604 => x"88",
          1605 => x"a4",
          1606 => x"34",
          1607 => x"bb",
          1608 => x"05",
          1609 => x"73",
          1610 => x"82",
          1611 => x"f8",
          1612 => x"72",
          1613 => x"38",
          1614 => x"0b",
          1615 => x"08",
          1616 => x"82",
          1617 => x"0b",
          1618 => x"08",
          1619 => x"80",
          1620 => x"a4",
          1621 => x"0c",
          1622 => x"08",
          1623 => x"53",
          1624 => x"81",
          1625 => x"bb",
          1626 => x"05",
          1627 => x"e0",
          1628 => x"38",
          1629 => x"08",
          1630 => x"e0",
          1631 => x"72",
          1632 => x"08",
          1633 => x"82",
          1634 => x"f8",
          1635 => x"11",
          1636 => x"82",
          1637 => x"f8",
          1638 => x"bb",
          1639 => x"05",
          1640 => x"73",
          1641 => x"82",
          1642 => x"f8",
          1643 => x"11",
          1644 => x"82",
          1645 => x"f8",
          1646 => x"bb",
          1647 => x"05",
          1648 => x"89",
          1649 => x"80",
          1650 => x"a4",
          1651 => x"0c",
          1652 => x"82",
          1653 => x"f8",
          1654 => x"bb",
          1655 => x"05",
          1656 => x"72",
          1657 => x"38",
          1658 => x"bb",
          1659 => x"05",
          1660 => x"39",
          1661 => x"08",
          1662 => x"70",
          1663 => x"08",
          1664 => x"29",
          1665 => x"08",
          1666 => x"70",
          1667 => x"a4",
          1668 => x"0c",
          1669 => x"08",
          1670 => x"70",
          1671 => x"71",
          1672 => x"51",
          1673 => x"53",
          1674 => x"bb",
          1675 => x"05",
          1676 => x"39",
          1677 => x"08",
          1678 => x"53",
          1679 => x"90",
          1680 => x"a4",
          1681 => x"08",
          1682 => x"a4",
          1683 => x"0c",
          1684 => x"08",
          1685 => x"82",
          1686 => x"fc",
          1687 => x"0c",
          1688 => x"82",
          1689 => x"ec",
          1690 => x"bb",
          1691 => x"05",
          1692 => x"98",
          1693 => x"0d",
          1694 => x"0c",
          1695 => x"a4",
          1696 => x"bb",
          1697 => x"3d",
          1698 => x"e8",
          1699 => x"bb",
          1700 => x"05",
          1701 => x"bb",
          1702 => x"05",
          1703 => x"8c",
          1704 => x"98",
          1705 => x"bb",
          1706 => x"85",
          1707 => x"bb",
          1708 => x"82",
          1709 => x"02",
          1710 => x"0c",
          1711 => x"80",
          1712 => x"a4",
          1713 => x"34",
          1714 => x"08",
          1715 => x"53",
          1716 => x"82",
          1717 => x"88",
          1718 => x"08",
          1719 => x"33",
          1720 => x"bb",
          1721 => x"05",
          1722 => x"ff",
          1723 => x"a0",
          1724 => x"06",
          1725 => x"bb",
          1726 => x"05",
          1727 => x"81",
          1728 => x"53",
          1729 => x"bb",
          1730 => x"05",
          1731 => x"ad",
          1732 => x"06",
          1733 => x"0b",
          1734 => x"08",
          1735 => x"82",
          1736 => x"88",
          1737 => x"08",
          1738 => x"0c",
          1739 => x"53",
          1740 => x"bb",
          1741 => x"05",
          1742 => x"a4",
          1743 => x"33",
          1744 => x"2e",
          1745 => x"81",
          1746 => x"bb",
          1747 => x"05",
          1748 => x"81",
          1749 => x"70",
          1750 => x"72",
          1751 => x"a4",
          1752 => x"34",
          1753 => x"08",
          1754 => x"82",
          1755 => x"e8",
          1756 => x"bb",
          1757 => x"05",
          1758 => x"2e",
          1759 => x"bb",
          1760 => x"05",
          1761 => x"2e",
          1762 => x"cd",
          1763 => x"82",
          1764 => x"f4",
          1765 => x"bb",
          1766 => x"05",
          1767 => x"81",
          1768 => x"70",
          1769 => x"72",
          1770 => x"a4",
          1771 => x"34",
          1772 => x"82",
          1773 => x"a4",
          1774 => x"34",
          1775 => x"08",
          1776 => x"70",
          1777 => x"71",
          1778 => x"51",
          1779 => x"82",
          1780 => x"f8",
          1781 => x"fe",
          1782 => x"a4",
          1783 => x"33",
          1784 => x"26",
          1785 => x"0b",
          1786 => x"08",
          1787 => x"83",
          1788 => x"bb",
          1789 => x"05",
          1790 => x"73",
          1791 => x"82",
          1792 => x"f8",
          1793 => x"72",
          1794 => x"38",
          1795 => x"0b",
          1796 => x"08",
          1797 => x"82",
          1798 => x"0b",
          1799 => x"08",
          1800 => x"b2",
          1801 => x"a4",
          1802 => x"33",
          1803 => x"27",
          1804 => x"bb",
          1805 => x"05",
          1806 => x"b9",
          1807 => x"8d",
          1808 => x"82",
          1809 => x"ec",
          1810 => x"a5",
          1811 => x"82",
          1812 => x"f4",
          1813 => x"0b",
          1814 => x"08",
          1815 => x"82",
          1816 => x"f8",
          1817 => x"a0",
          1818 => x"cf",
          1819 => x"a4",
          1820 => x"33",
          1821 => x"73",
          1822 => x"82",
          1823 => x"f8",
          1824 => x"11",
          1825 => x"82",
          1826 => x"f8",
          1827 => x"bb",
          1828 => x"05",
          1829 => x"51",
          1830 => x"bb",
          1831 => x"05",
          1832 => x"a4",
          1833 => x"33",
          1834 => x"27",
          1835 => x"bb",
          1836 => x"05",
          1837 => x"51",
          1838 => x"bb",
          1839 => x"05",
          1840 => x"a4",
          1841 => x"33",
          1842 => x"26",
          1843 => x"0b",
          1844 => x"08",
          1845 => x"81",
          1846 => x"bb",
          1847 => x"05",
          1848 => x"a4",
          1849 => x"33",
          1850 => x"74",
          1851 => x"80",
          1852 => x"a4",
          1853 => x"0c",
          1854 => x"82",
          1855 => x"f4",
          1856 => x"82",
          1857 => x"fc",
          1858 => x"82",
          1859 => x"f8",
          1860 => x"12",
          1861 => x"08",
          1862 => x"82",
          1863 => x"88",
          1864 => x"08",
          1865 => x"0c",
          1866 => x"51",
          1867 => x"72",
          1868 => x"a4",
          1869 => x"34",
          1870 => x"82",
          1871 => x"f0",
          1872 => x"72",
          1873 => x"38",
          1874 => x"08",
          1875 => x"30",
          1876 => x"08",
          1877 => x"82",
          1878 => x"8c",
          1879 => x"bb",
          1880 => x"05",
          1881 => x"53",
          1882 => x"bb",
          1883 => x"05",
          1884 => x"a4",
          1885 => x"08",
          1886 => x"0c",
          1887 => x"82",
          1888 => x"04",
          1889 => x"08",
          1890 => x"a4",
          1891 => x"0d",
          1892 => x"bb",
          1893 => x"05",
          1894 => x"ec",
          1895 => x"33",
          1896 => x"70",
          1897 => x"81",
          1898 => x"51",
          1899 => x"80",
          1900 => x"ff",
          1901 => x"a4",
          1902 => x"0c",
          1903 => x"82",
          1904 => x"88",
          1905 => x"72",
          1906 => x"a4",
          1907 => x"08",
          1908 => x"bb",
          1909 => x"05",
          1910 => x"82",
          1911 => x"fc",
          1912 => x"81",
          1913 => x"72",
          1914 => x"38",
          1915 => x"08",
          1916 => x"08",
          1917 => x"a4",
          1918 => x"33",
          1919 => x"08",
          1920 => x"2d",
          1921 => x"08",
          1922 => x"2e",
          1923 => x"ff",
          1924 => x"a4",
          1925 => x"0c",
          1926 => x"82",
          1927 => x"82",
          1928 => x"53",
          1929 => x"90",
          1930 => x"72",
          1931 => x"98",
          1932 => x"80",
          1933 => x"ff",
          1934 => x"a4",
          1935 => x"0c",
          1936 => x"08",
          1937 => x"70",
          1938 => x"08",
          1939 => x"53",
          1940 => x"08",
          1941 => x"82",
          1942 => x"87",
          1943 => x"bb",
          1944 => x"82",
          1945 => x"02",
          1946 => x"0c",
          1947 => x"80",
          1948 => x"a4",
          1949 => x"0c",
          1950 => x"08",
          1951 => x"85",
          1952 => x"81",
          1953 => x"32",
          1954 => x"51",
          1955 => x"53",
          1956 => x"8d",
          1957 => x"82",
          1958 => x"f4",
          1959 => x"f3",
          1960 => x"a4",
          1961 => x"08",
          1962 => x"82",
          1963 => x"88",
          1964 => x"05",
          1965 => x"08",
          1966 => x"53",
          1967 => x"a4",
          1968 => x"34",
          1969 => x"06",
          1970 => x"2e",
          1971 => x"bb",
          1972 => x"05",
          1973 => x"a4",
          1974 => x"08",
          1975 => x"a4",
          1976 => x"33",
          1977 => x"08",
          1978 => x"2d",
          1979 => x"08",
          1980 => x"2e",
          1981 => x"ff",
          1982 => x"a4",
          1983 => x"0c",
          1984 => x"82",
          1985 => x"f8",
          1986 => x"82",
          1987 => x"f4",
          1988 => x"82",
          1989 => x"f4",
          1990 => x"bb",
          1991 => x"3d",
          1992 => x"a4",
          1993 => x"bb",
          1994 => x"82",
          1995 => x"fe",
          1996 => x"d2",
          1997 => x"82",
          1998 => x"88",
          1999 => x"93",
          2000 => x"98",
          2001 => x"bb",
          2002 => x"84",
          2003 => x"bb",
          2004 => x"82",
          2005 => x"02",
          2006 => x"0c",
          2007 => x"82",
          2008 => x"8c",
          2009 => x"11",
          2010 => x"2a",
          2011 => x"70",
          2012 => x"51",
          2013 => x"72",
          2014 => x"38",
          2015 => x"bb",
          2016 => x"05",
          2017 => x"39",
          2018 => x"08",
          2019 => x"85",
          2020 => x"82",
          2021 => x"06",
          2022 => x"53",
          2023 => x"80",
          2024 => x"bb",
          2025 => x"05",
          2026 => x"a4",
          2027 => x"08",
          2028 => x"14",
          2029 => x"08",
          2030 => x"82",
          2031 => x"8c",
          2032 => x"08",
          2033 => x"a4",
          2034 => x"08",
          2035 => x"54",
          2036 => x"73",
          2037 => x"74",
          2038 => x"a4",
          2039 => x"08",
          2040 => x"81",
          2041 => x"0c",
          2042 => x"08",
          2043 => x"70",
          2044 => x"08",
          2045 => x"51",
          2046 => x"39",
          2047 => x"08",
          2048 => x"82",
          2049 => x"8c",
          2050 => x"82",
          2051 => x"88",
          2052 => x"81",
          2053 => x"90",
          2054 => x"54",
          2055 => x"82",
          2056 => x"53",
          2057 => x"82",
          2058 => x"8c",
          2059 => x"11",
          2060 => x"8c",
          2061 => x"bb",
          2062 => x"05",
          2063 => x"bb",
          2064 => x"05",
          2065 => x"8a",
          2066 => x"82",
          2067 => x"fc",
          2068 => x"bb",
          2069 => x"05",
          2070 => x"98",
          2071 => x"0d",
          2072 => x"0c",
          2073 => x"a4",
          2074 => x"bb",
          2075 => x"3d",
          2076 => x"a4",
          2077 => x"08",
          2078 => x"70",
          2079 => x"81",
          2080 => x"51",
          2081 => x"2e",
          2082 => x"0b",
          2083 => x"08",
          2084 => x"83",
          2085 => x"bb",
          2086 => x"05",
          2087 => x"33",
          2088 => x"70",
          2089 => x"51",
          2090 => x"80",
          2091 => x"38",
          2092 => x"08",
          2093 => x"82",
          2094 => x"88",
          2095 => x"53",
          2096 => x"70",
          2097 => x"51",
          2098 => x"14",
          2099 => x"a4",
          2100 => x"08",
          2101 => x"81",
          2102 => x"0c",
          2103 => x"08",
          2104 => x"84",
          2105 => x"82",
          2106 => x"f8",
          2107 => x"51",
          2108 => x"39",
          2109 => x"08",
          2110 => x"85",
          2111 => x"82",
          2112 => x"06",
          2113 => x"52",
          2114 => x"80",
          2115 => x"bb",
          2116 => x"05",
          2117 => x"70",
          2118 => x"a4",
          2119 => x"0c",
          2120 => x"bb",
          2121 => x"05",
          2122 => x"82",
          2123 => x"88",
          2124 => x"bb",
          2125 => x"05",
          2126 => x"85",
          2127 => x"a0",
          2128 => x"71",
          2129 => x"ff",
          2130 => x"a4",
          2131 => x"0c",
          2132 => x"82",
          2133 => x"88",
          2134 => x"08",
          2135 => x"0c",
          2136 => x"39",
          2137 => x"08",
          2138 => x"82",
          2139 => x"88",
          2140 => x"94",
          2141 => x"52",
          2142 => x"bb",
          2143 => x"82",
          2144 => x"fc",
          2145 => x"82",
          2146 => x"fc",
          2147 => x"25",
          2148 => x"82",
          2149 => x"88",
          2150 => x"bb",
          2151 => x"05",
          2152 => x"a4",
          2153 => x"08",
          2154 => x"82",
          2155 => x"f0",
          2156 => x"82",
          2157 => x"fc",
          2158 => x"2e",
          2159 => x"95",
          2160 => x"a4",
          2161 => x"08",
          2162 => x"71",
          2163 => x"08",
          2164 => x"93",
          2165 => x"a4",
          2166 => x"08",
          2167 => x"71",
          2168 => x"08",
          2169 => x"82",
          2170 => x"f4",
          2171 => x"82",
          2172 => x"ec",
          2173 => x"13",
          2174 => x"82",
          2175 => x"f8",
          2176 => x"39",
          2177 => x"08",
          2178 => x"8c",
          2179 => x"05",
          2180 => x"82",
          2181 => x"fc",
          2182 => x"81",
          2183 => x"82",
          2184 => x"f8",
          2185 => x"51",
          2186 => x"a4",
          2187 => x"08",
          2188 => x"0c",
          2189 => x"82",
          2190 => x"04",
          2191 => x"08",
          2192 => x"a4",
          2193 => x"0d",
          2194 => x"08",
          2195 => x"82",
          2196 => x"fc",
          2197 => x"bb",
          2198 => x"05",
          2199 => x"a4",
          2200 => x"0c",
          2201 => x"08",
          2202 => x"80",
          2203 => x"38",
          2204 => x"08",
          2205 => x"82",
          2206 => x"fc",
          2207 => x"81",
          2208 => x"bb",
          2209 => x"05",
          2210 => x"a4",
          2211 => x"08",
          2212 => x"bb",
          2213 => x"05",
          2214 => x"81",
          2215 => x"bb",
          2216 => x"05",
          2217 => x"a4",
          2218 => x"08",
          2219 => x"a4",
          2220 => x"0c",
          2221 => x"08",
          2222 => x"82",
          2223 => x"90",
          2224 => x"82",
          2225 => x"f8",
          2226 => x"bb",
          2227 => x"05",
          2228 => x"82",
          2229 => x"90",
          2230 => x"bb",
          2231 => x"05",
          2232 => x"82",
          2233 => x"90",
          2234 => x"bb",
          2235 => x"05",
          2236 => x"81",
          2237 => x"bb",
          2238 => x"05",
          2239 => x"82",
          2240 => x"fc",
          2241 => x"bb",
          2242 => x"05",
          2243 => x"82",
          2244 => x"f8",
          2245 => x"bb",
          2246 => x"05",
          2247 => x"a4",
          2248 => x"08",
          2249 => x"33",
          2250 => x"ae",
          2251 => x"a4",
          2252 => x"08",
          2253 => x"bb",
          2254 => x"05",
          2255 => x"a4",
          2256 => x"08",
          2257 => x"bb",
          2258 => x"05",
          2259 => x"a4",
          2260 => x"08",
          2261 => x"38",
          2262 => x"08",
          2263 => x"51",
          2264 => x"bb",
          2265 => x"05",
          2266 => x"82",
          2267 => x"f8",
          2268 => x"bb",
          2269 => x"05",
          2270 => x"71",
          2271 => x"bb",
          2272 => x"05",
          2273 => x"82",
          2274 => x"fc",
          2275 => x"ad",
          2276 => x"a4",
          2277 => x"08",
          2278 => x"98",
          2279 => x"3d",
          2280 => x"a4",
          2281 => x"bb",
          2282 => x"82",
          2283 => x"fe",
          2284 => x"bb",
          2285 => x"05",
          2286 => x"a4",
          2287 => x"0c",
          2288 => x"08",
          2289 => x"52",
          2290 => x"bb",
          2291 => x"05",
          2292 => x"82",
          2293 => x"fc",
          2294 => x"81",
          2295 => x"51",
          2296 => x"83",
          2297 => x"82",
          2298 => x"fc",
          2299 => x"05",
          2300 => x"08",
          2301 => x"82",
          2302 => x"fc",
          2303 => x"bb",
          2304 => x"05",
          2305 => x"82",
          2306 => x"51",
          2307 => x"82",
          2308 => x"04",
          2309 => x"08",
          2310 => x"a4",
          2311 => x"0d",
          2312 => x"08",
          2313 => x"82",
          2314 => x"fc",
          2315 => x"bb",
          2316 => x"05",
          2317 => x"33",
          2318 => x"08",
          2319 => x"81",
          2320 => x"a4",
          2321 => x"0c",
          2322 => x"08",
          2323 => x"53",
          2324 => x"34",
          2325 => x"08",
          2326 => x"81",
          2327 => x"a4",
          2328 => x"0c",
          2329 => x"06",
          2330 => x"2e",
          2331 => x"be",
          2332 => x"a4",
          2333 => x"08",
          2334 => x"98",
          2335 => x"3d",
          2336 => x"a4",
          2337 => x"bb",
          2338 => x"82",
          2339 => x"fd",
          2340 => x"bb",
          2341 => x"05",
          2342 => x"a4",
          2343 => x"0c",
          2344 => x"08",
          2345 => x"82",
          2346 => x"f8",
          2347 => x"bb",
          2348 => x"05",
          2349 => x"80",
          2350 => x"bb",
          2351 => x"05",
          2352 => x"82",
          2353 => x"90",
          2354 => x"bb",
          2355 => x"05",
          2356 => x"82",
          2357 => x"90",
          2358 => x"bb",
          2359 => x"05",
          2360 => x"ba",
          2361 => x"a4",
          2362 => x"08",
          2363 => x"82",
          2364 => x"f8",
          2365 => x"05",
          2366 => x"08",
          2367 => x"82",
          2368 => x"fc",
          2369 => x"52",
          2370 => x"82",
          2371 => x"fc",
          2372 => x"05",
          2373 => x"08",
          2374 => x"ff",
          2375 => x"bb",
          2376 => x"05",
          2377 => x"bb",
          2378 => x"85",
          2379 => x"bb",
          2380 => x"82",
          2381 => x"02",
          2382 => x"0c",
          2383 => x"82",
          2384 => x"90",
          2385 => x"2e",
          2386 => x"82",
          2387 => x"8c",
          2388 => x"71",
          2389 => x"a4",
          2390 => x"08",
          2391 => x"bb",
          2392 => x"05",
          2393 => x"a4",
          2394 => x"08",
          2395 => x"81",
          2396 => x"54",
          2397 => x"71",
          2398 => x"80",
          2399 => x"bb",
          2400 => x"05",
          2401 => x"33",
          2402 => x"08",
          2403 => x"81",
          2404 => x"a4",
          2405 => x"0c",
          2406 => x"06",
          2407 => x"8d",
          2408 => x"82",
          2409 => x"fc",
          2410 => x"9b",
          2411 => x"a4",
          2412 => x"08",
          2413 => x"bb",
          2414 => x"05",
          2415 => x"a4",
          2416 => x"08",
          2417 => x"38",
          2418 => x"82",
          2419 => x"90",
          2420 => x"2e",
          2421 => x"82",
          2422 => x"88",
          2423 => x"33",
          2424 => x"8d",
          2425 => x"82",
          2426 => x"fc",
          2427 => x"d7",
          2428 => x"a4",
          2429 => x"08",
          2430 => x"bb",
          2431 => x"05",
          2432 => x"a4",
          2433 => x"08",
          2434 => x"52",
          2435 => x"81",
          2436 => x"a4",
          2437 => x"0c",
          2438 => x"bb",
          2439 => x"05",
          2440 => x"82",
          2441 => x"8c",
          2442 => x"33",
          2443 => x"70",
          2444 => x"08",
          2445 => x"53",
          2446 => x"53",
          2447 => x"0b",
          2448 => x"08",
          2449 => x"82",
          2450 => x"fc",
          2451 => x"bb",
          2452 => x"3d",
          2453 => x"a4",
          2454 => x"bb",
          2455 => x"82",
          2456 => x"fd",
          2457 => x"bb",
          2458 => x"05",
          2459 => x"a4",
          2460 => x"0c",
          2461 => x"08",
          2462 => x"8d",
          2463 => x"82",
          2464 => x"fc",
          2465 => x"ec",
          2466 => x"a4",
          2467 => x"08",
          2468 => x"82",
          2469 => x"f8",
          2470 => x"05",
          2471 => x"08",
          2472 => x"70",
          2473 => x"51",
          2474 => x"2e",
          2475 => x"bb",
          2476 => x"05",
          2477 => x"82",
          2478 => x"8c",
          2479 => x"bb",
          2480 => x"05",
          2481 => x"84",
          2482 => x"39",
          2483 => x"08",
          2484 => x"ff",
          2485 => x"a4",
          2486 => x"0c",
          2487 => x"08",
          2488 => x"82",
          2489 => x"88",
          2490 => x"70",
          2491 => x"08",
          2492 => x"51",
          2493 => x"08",
          2494 => x"82",
          2495 => x"85",
          2496 => x"bb",
          2497 => x"82",
          2498 => x"02",
          2499 => x"0c",
          2500 => x"82",
          2501 => x"88",
          2502 => x"bb",
          2503 => x"05",
          2504 => x"a4",
          2505 => x"08",
          2506 => x"d4",
          2507 => x"a4",
          2508 => x"08",
          2509 => x"bb",
          2510 => x"05",
          2511 => x"a4",
          2512 => x"08",
          2513 => x"bb",
          2514 => x"05",
          2515 => x"a4",
          2516 => x"08",
          2517 => x"38",
          2518 => x"08",
          2519 => x"51",
          2520 => x"a4",
          2521 => x"08",
          2522 => x"71",
          2523 => x"a4",
          2524 => x"08",
          2525 => x"bb",
          2526 => x"05",
          2527 => x"39",
          2528 => x"08",
          2529 => x"70",
          2530 => x"0c",
          2531 => x"0d",
          2532 => x"0c",
          2533 => x"a4",
          2534 => x"bb",
          2535 => x"3d",
          2536 => x"82",
          2537 => x"fc",
          2538 => x"bb",
          2539 => x"05",
          2540 => x"b9",
          2541 => x"a4",
          2542 => x"08",
          2543 => x"a4",
          2544 => x"0c",
          2545 => x"bb",
          2546 => x"05",
          2547 => x"a4",
          2548 => x"08",
          2549 => x"0b",
          2550 => x"08",
          2551 => x"82",
          2552 => x"f4",
          2553 => x"bb",
          2554 => x"05",
          2555 => x"a4",
          2556 => x"08",
          2557 => x"38",
          2558 => x"08",
          2559 => x"30",
          2560 => x"08",
          2561 => x"80",
          2562 => x"a4",
          2563 => x"0c",
          2564 => x"08",
          2565 => x"8a",
          2566 => x"82",
          2567 => x"f0",
          2568 => x"bb",
          2569 => x"05",
          2570 => x"a4",
          2571 => x"0c",
          2572 => x"bb",
          2573 => x"05",
          2574 => x"bb",
          2575 => x"05",
          2576 => x"c5",
          2577 => x"98",
          2578 => x"bb",
          2579 => x"05",
          2580 => x"bb",
          2581 => x"05",
          2582 => x"90",
          2583 => x"a4",
          2584 => x"08",
          2585 => x"a4",
          2586 => x"0c",
          2587 => x"08",
          2588 => x"70",
          2589 => x"0c",
          2590 => x"0d",
          2591 => x"0c",
          2592 => x"a4",
          2593 => x"bb",
          2594 => x"3d",
          2595 => x"82",
          2596 => x"fc",
          2597 => x"bb",
          2598 => x"05",
          2599 => x"99",
          2600 => x"a4",
          2601 => x"08",
          2602 => x"a4",
          2603 => x"0c",
          2604 => x"bb",
          2605 => x"05",
          2606 => x"a4",
          2607 => x"08",
          2608 => x"38",
          2609 => x"08",
          2610 => x"30",
          2611 => x"08",
          2612 => x"81",
          2613 => x"a4",
          2614 => x"08",
          2615 => x"a4",
          2616 => x"08",
          2617 => x"3f",
          2618 => x"08",
          2619 => x"a4",
          2620 => x"0c",
          2621 => x"a4",
          2622 => x"08",
          2623 => x"38",
          2624 => x"08",
          2625 => x"30",
          2626 => x"08",
          2627 => x"82",
          2628 => x"f8",
          2629 => x"82",
          2630 => x"54",
          2631 => x"82",
          2632 => x"04",
          2633 => x"08",
          2634 => x"a4",
          2635 => x"0d",
          2636 => x"bb",
          2637 => x"05",
          2638 => x"bb",
          2639 => x"05",
          2640 => x"c5",
          2641 => x"98",
          2642 => x"bb",
          2643 => x"85",
          2644 => x"bb",
          2645 => x"82",
          2646 => x"02",
          2647 => x"0c",
          2648 => x"81",
          2649 => x"a4",
          2650 => x"08",
          2651 => x"a4",
          2652 => x"08",
          2653 => x"82",
          2654 => x"70",
          2655 => x"0c",
          2656 => x"0d",
          2657 => x"0c",
          2658 => x"a4",
          2659 => x"bb",
          2660 => x"3d",
          2661 => x"82",
          2662 => x"fc",
          2663 => x"0b",
          2664 => x"08",
          2665 => x"82",
          2666 => x"8c",
          2667 => x"bb",
          2668 => x"05",
          2669 => x"38",
          2670 => x"08",
          2671 => x"80",
          2672 => x"80",
          2673 => x"a4",
          2674 => x"08",
          2675 => x"82",
          2676 => x"8c",
          2677 => x"82",
          2678 => x"8c",
          2679 => x"bb",
          2680 => x"05",
          2681 => x"bb",
          2682 => x"05",
          2683 => x"39",
          2684 => x"08",
          2685 => x"80",
          2686 => x"38",
          2687 => x"08",
          2688 => x"82",
          2689 => x"88",
          2690 => x"ad",
          2691 => x"a4",
          2692 => x"08",
          2693 => x"08",
          2694 => x"31",
          2695 => x"08",
          2696 => x"82",
          2697 => x"f8",
          2698 => x"bb",
          2699 => x"05",
          2700 => x"bb",
          2701 => x"05",
          2702 => x"a4",
          2703 => x"08",
          2704 => x"bb",
          2705 => x"05",
          2706 => x"a4",
          2707 => x"08",
          2708 => x"bb",
          2709 => x"05",
          2710 => x"39",
          2711 => x"08",
          2712 => x"80",
          2713 => x"82",
          2714 => x"88",
          2715 => x"82",
          2716 => x"f4",
          2717 => x"91",
          2718 => x"a4",
          2719 => x"08",
          2720 => x"a4",
          2721 => x"0c",
          2722 => x"a4",
          2723 => x"08",
          2724 => x"0c",
          2725 => x"82",
          2726 => x"04",
          2727 => x"79",
          2728 => x"56",
          2729 => x"80",
          2730 => x"38",
          2731 => x"08",
          2732 => x"3f",
          2733 => x"08",
          2734 => x"85",
          2735 => x"80",
          2736 => x"33",
          2737 => x"2e",
          2738 => x"86",
          2739 => x"55",
          2740 => x"57",
          2741 => x"82",
          2742 => x"70",
          2743 => x"f1",
          2744 => x"bb",
          2745 => x"74",
          2746 => x"51",
          2747 => x"82",
          2748 => x"8b",
          2749 => x"33",
          2750 => x"2e",
          2751 => x"81",
          2752 => x"ff",
          2753 => x"99",
          2754 => x"38",
          2755 => x"82",
          2756 => x"89",
          2757 => x"ff",
          2758 => x"52",
          2759 => x"81",
          2760 => x"84",
          2761 => x"b0",
          2762 => x"08",
          2763 => x"fc",
          2764 => x"39",
          2765 => x"51",
          2766 => x"82",
          2767 => x"80",
          2768 => x"9f",
          2769 => x"eb",
          2770 => x"c0",
          2771 => x"39",
          2772 => x"51",
          2773 => x"82",
          2774 => x"80",
          2775 => x"9f",
          2776 => x"cf",
          2777 => x"8c",
          2778 => x"39",
          2779 => x"51",
          2780 => x"82",
          2781 => x"bb",
          2782 => x"d8",
          2783 => x"82",
          2784 => x"af",
          2785 => x"98",
          2786 => x"82",
          2787 => x"a3",
          2788 => x"cc",
          2789 => x"82",
          2790 => x"97",
          2791 => x"f8",
          2792 => x"82",
          2793 => x"8b",
          2794 => x"a8",
          2795 => x"82",
          2796 => x"e3",
          2797 => x"3d",
          2798 => x"3d",
          2799 => x"56",
          2800 => x"e7",
          2801 => x"74",
          2802 => x"e8",
          2803 => x"39",
          2804 => x"74",
          2805 => x"3f",
          2806 => x"08",
          2807 => x"fa",
          2808 => x"bb",
          2809 => x"79",
          2810 => x"82",
          2811 => x"ff",
          2812 => x"87",
          2813 => x"ec",
          2814 => x"02",
          2815 => x"e3",
          2816 => x"57",
          2817 => x"30",
          2818 => x"73",
          2819 => x"59",
          2820 => x"77",
          2821 => x"83",
          2822 => x"74",
          2823 => x"81",
          2824 => x"55",
          2825 => x"81",
          2826 => x"53",
          2827 => x"3d",
          2828 => x"81",
          2829 => x"82",
          2830 => x"57",
          2831 => x"08",
          2832 => x"bb",
          2833 => x"c0",
          2834 => x"82",
          2835 => x"59",
          2836 => x"05",
          2837 => x"53",
          2838 => x"51",
          2839 => x"3f",
          2840 => x"08",
          2841 => x"98",
          2842 => x"7a",
          2843 => x"2e",
          2844 => x"19",
          2845 => x"59",
          2846 => x"3d",
          2847 => x"81",
          2848 => x"76",
          2849 => x"07",
          2850 => x"30",
          2851 => x"72",
          2852 => x"51",
          2853 => x"2e",
          2854 => x"a2",
          2855 => x"c0",
          2856 => x"52",
          2857 => x"92",
          2858 => x"75",
          2859 => x"0c",
          2860 => x"04",
          2861 => x"7c",
          2862 => x"b7",
          2863 => x"59",
          2864 => x"53",
          2865 => x"51",
          2866 => x"82",
          2867 => x"a6",
          2868 => x"2e",
          2869 => x"81",
          2870 => x"9a",
          2871 => x"61",
          2872 => x"82",
          2873 => x"7f",
          2874 => x"78",
          2875 => x"98",
          2876 => x"39",
          2877 => x"82",
          2878 => x"8a",
          2879 => x"f3",
          2880 => x"61",
          2881 => x"05",
          2882 => x"33",
          2883 => x"68",
          2884 => x"5c",
          2885 => x"7a",
          2886 => x"f0",
          2887 => x"b7",
          2888 => x"f8",
          2889 => x"3f",
          2890 => x"79",
          2891 => x"38",
          2892 => x"89",
          2893 => x"2e",
          2894 => x"c4",
          2895 => x"53",
          2896 => x"8e",
          2897 => x"52",
          2898 => x"51",
          2899 => x"3f",
          2900 => x"a3",
          2901 => x"ac",
          2902 => x"55",
          2903 => x"74",
          2904 => x"7a",
          2905 => x"72",
          2906 => x"a2",
          2907 => x"b8",
          2908 => x"39",
          2909 => x"51",
          2910 => x"84",
          2911 => x"39",
          2912 => x"72",
          2913 => x"38",
          2914 => x"82",
          2915 => x"ff",
          2916 => x"88",
          2917 => x"98",
          2918 => x"3f",
          2919 => x"82",
          2920 => x"52",
          2921 => x"ab",
          2922 => x"39",
          2923 => x"51",
          2924 => x"80",
          2925 => x"27",
          2926 => x"74",
          2927 => x"55",
          2928 => x"72",
          2929 => x"38",
          2930 => x"53",
          2931 => x"83",
          2932 => x"75",
          2933 => x"81",
          2934 => x"53",
          2935 => x"90",
          2936 => x"fe",
          2937 => x"82",
          2938 => x"52",
          2939 => x"39",
          2940 => x"08",
          2941 => x"e2",
          2942 => x"15",
          2943 => x"39",
          2944 => x"51",
          2945 => x"78",
          2946 => x"5c",
          2947 => x"3f",
          2948 => x"08",
          2949 => x"98",
          2950 => x"76",
          2951 => x"81",
          2952 => x"a0",
          2953 => x"bb",
          2954 => x"2b",
          2955 => x"70",
          2956 => x"30",
          2957 => x"70",
          2958 => x"07",
          2959 => x"06",
          2960 => x"59",
          2961 => x"80",
          2962 => x"38",
          2963 => x"09",
          2964 => x"38",
          2965 => x"39",
          2966 => x"72",
          2967 => x"b7",
          2968 => x"72",
          2969 => x"0c",
          2970 => x"04",
          2971 => x"02",
          2972 => x"82",
          2973 => x"82",
          2974 => x"55",
          2975 => x"3f",
          2976 => x"22",
          2977 => x"3f",
          2978 => x"54",
          2979 => x"53",
          2980 => x"33",
          2981 => x"cc",
          2982 => x"bb",
          2983 => x"2e",
          2984 => x"fc",
          2985 => x"0d",
          2986 => x"0d",
          2987 => x"80",
          2988 => x"a7",
          2989 => x"9c",
          2990 => x"a3",
          2991 => x"c7",
          2992 => x"9c",
          2993 => x"81",
          2994 => x"06",
          2995 => x"80",
          2996 => x"81",
          2997 => x"3f",
          2998 => x"51",
          2999 => x"80",
          3000 => x"3f",
          3001 => x"70",
          3002 => x"52",
          3003 => x"92",
          3004 => x"9b",
          3005 => x"a4",
          3006 => x"8b",
          3007 => x"9b",
          3008 => x"83",
          3009 => x"06",
          3010 => x"80",
          3011 => x"81",
          3012 => x"3f",
          3013 => x"51",
          3014 => x"80",
          3015 => x"3f",
          3016 => x"70",
          3017 => x"52",
          3018 => x"92",
          3019 => x"9b",
          3020 => x"a4",
          3021 => x"cf",
          3022 => x"9b",
          3023 => x"85",
          3024 => x"06",
          3025 => x"80",
          3026 => x"81",
          3027 => x"3f",
          3028 => x"51",
          3029 => x"80",
          3030 => x"3f",
          3031 => x"70",
          3032 => x"52",
          3033 => x"92",
          3034 => x"9a",
          3035 => x"a4",
          3036 => x"93",
          3037 => x"9a",
          3038 => x"87",
          3039 => x"06",
          3040 => x"80",
          3041 => x"81",
          3042 => x"3f",
          3043 => x"51",
          3044 => x"80",
          3045 => x"3f",
          3046 => x"70",
          3047 => x"52",
          3048 => x"92",
          3049 => x"9a",
          3050 => x"a5",
          3051 => x"d7",
          3052 => x"9a",
          3053 => x"ab",
          3054 => x"0d",
          3055 => x"0d",
          3056 => x"05",
          3057 => x"70",
          3058 => x"80",
          3059 => x"ee",
          3060 => x"0b",
          3061 => x"33",
          3062 => x"38",
          3063 => x"a5",
          3064 => x"d2",
          3065 => x"fc",
          3066 => x"bb",
          3067 => x"70",
          3068 => x"08",
          3069 => x"82",
          3070 => x"51",
          3071 => x"0b",
          3072 => x"34",
          3073 => x"b6",
          3074 => x"73",
          3075 => x"81",
          3076 => x"82",
          3077 => x"74",
          3078 => x"81",
          3079 => x"82",
          3080 => x"80",
          3081 => x"82",
          3082 => x"51",
          3083 => x"91",
          3084 => x"98",
          3085 => x"be",
          3086 => x"0b",
          3087 => x"94",
          3088 => x"82",
          3089 => x"54",
          3090 => x"09",
          3091 => x"38",
          3092 => x"53",
          3093 => x"51",
          3094 => x"80",
          3095 => x"98",
          3096 => x"0d",
          3097 => x"0d",
          3098 => x"82",
          3099 => x"40",
          3100 => x"7d",
          3101 => x"e8",
          3102 => x"98",
          3103 => x"06",
          3104 => x"2e",
          3105 => x"a3",
          3106 => x"5a",
          3107 => x"a5",
          3108 => x"51",
          3109 => x"7d",
          3110 => x"82",
          3111 => x"80",
          3112 => x"82",
          3113 => x"7e",
          3114 => x"82",
          3115 => x"91",
          3116 => x"70",
          3117 => x"a6",
          3118 => x"c8",
          3119 => x"70",
          3120 => x"f8",
          3121 => x"fd",
          3122 => x"3d",
          3123 => x"51",
          3124 => x"82",
          3125 => x"90",
          3126 => x"2c",
          3127 => x"80",
          3128 => x"d4",
          3129 => x"c1",
          3130 => x"38",
          3131 => x"83",
          3132 => x"ab",
          3133 => x"79",
          3134 => x"b3",
          3135 => x"24",
          3136 => x"80",
          3137 => x"38",
          3138 => x"79",
          3139 => x"83",
          3140 => x"2e",
          3141 => x"8e",
          3142 => x"bd",
          3143 => x"38",
          3144 => x"90",
          3145 => x"2e",
          3146 => x"79",
          3147 => x"88",
          3148 => x"39",
          3149 => x"85",
          3150 => x"80",
          3151 => x"bd",
          3152 => x"39",
          3153 => x"2e",
          3154 => x"79",
          3155 => x"b0",
          3156 => x"d0",
          3157 => x"38",
          3158 => x"24",
          3159 => x"80",
          3160 => x"f6",
          3161 => x"c3",
          3162 => x"38",
          3163 => x"79",
          3164 => x"8c",
          3165 => x"80",
          3166 => x"c2",
          3167 => x"39",
          3168 => x"2e",
          3169 => x"79",
          3170 => x"92",
          3171 => x"f8",
          3172 => x"38",
          3173 => x"2e",
          3174 => x"8d",
          3175 => x"81",
          3176 => x"c1",
          3177 => x"85",
          3178 => x"38",
          3179 => x"b5",
          3180 => x"11",
          3181 => x"05",
          3182 => x"3f",
          3183 => x"08",
          3184 => x"a6",
          3185 => x"b1",
          3186 => x"fe",
          3187 => x"ff",
          3188 => x"d1",
          3189 => x"bb",
          3190 => x"2e",
          3191 => x"64",
          3192 => x"80",
          3193 => x"cf",
          3194 => x"02",
          3195 => x"33",
          3196 => x"ec",
          3197 => x"98",
          3198 => x"06",
          3199 => x"38",
          3200 => x"51",
          3201 => x"81",
          3202 => x"39",
          3203 => x"51",
          3204 => x"b5",
          3205 => x"11",
          3206 => x"05",
          3207 => x"3f",
          3208 => x"08",
          3209 => x"8e",
          3210 => x"80",
          3211 => x"d3",
          3212 => x"80",
          3213 => x"82",
          3214 => x"52",
          3215 => x"51",
          3216 => x"b5",
          3217 => x"11",
          3218 => x"05",
          3219 => x"3f",
          3220 => x"08",
          3221 => x"38",
          3222 => x"fc",
          3223 => x"3d",
          3224 => x"53",
          3225 => x"51",
          3226 => x"82",
          3227 => x"86",
          3228 => x"98",
          3229 => x"53",
          3230 => x"52",
          3231 => x"b1",
          3232 => x"80",
          3233 => x"53",
          3234 => x"84",
          3235 => x"bc",
          3236 => x"80",
          3237 => x"82",
          3238 => x"81",
          3239 => x"a6",
          3240 => x"e0",
          3241 => x"fc",
          3242 => x"3d",
          3243 => x"51",
          3244 => x"82",
          3245 => x"b6",
          3246 => x"05",
          3247 => x"c7",
          3248 => x"82",
          3249 => x"52",
          3250 => x"ab",
          3251 => x"39",
          3252 => x"84",
          3253 => x"8b",
          3254 => x"98",
          3255 => x"ff",
          3256 => x"5c",
          3257 => x"82",
          3258 => x"b6",
          3259 => x"05",
          3260 => x"93",
          3261 => x"98",
          3262 => x"ff",
          3263 => x"5a",
          3264 => x"82",
          3265 => x"82",
          3266 => x"82",
          3267 => x"80",
          3268 => x"82",
          3269 => x"81",
          3270 => x"79",
          3271 => x"7b",
          3272 => x"3f",
          3273 => x"08",
          3274 => x"8a",
          3275 => x"98",
          3276 => x"e3",
          3277 => x"39",
          3278 => x"80",
          3279 => x"84",
          3280 => x"ef",
          3281 => x"98",
          3282 => x"fa",
          3283 => x"3d",
          3284 => x"53",
          3285 => x"51",
          3286 => x"82",
          3287 => x"80",
          3288 => x"38",
          3289 => x"f8",
          3290 => x"84",
          3291 => x"c3",
          3292 => x"98",
          3293 => x"82",
          3294 => x"43",
          3295 => x"51",
          3296 => x"64",
          3297 => x"7a",
          3298 => x"ea",
          3299 => x"79",
          3300 => x"05",
          3301 => x"7b",
          3302 => x"81",
          3303 => x"3d",
          3304 => x"53",
          3305 => x"51",
          3306 => x"82",
          3307 => x"80",
          3308 => x"38",
          3309 => x"fc",
          3310 => x"84",
          3311 => x"f3",
          3312 => x"98",
          3313 => x"f9",
          3314 => x"3d",
          3315 => x"53",
          3316 => x"51",
          3317 => x"82",
          3318 => x"80",
          3319 => x"38",
          3320 => x"51",
          3321 => x"64",
          3322 => x"27",
          3323 => x"62",
          3324 => x"81",
          3325 => x"7a",
          3326 => x"05",
          3327 => x"b5",
          3328 => x"11",
          3329 => x"05",
          3330 => x"3f",
          3331 => x"08",
          3332 => x"a2",
          3333 => x"fe",
          3334 => x"ff",
          3335 => x"cd",
          3336 => x"bb",
          3337 => x"2e",
          3338 => x"b5",
          3339 => x"11",
          3340 => x"05",
          3341 => x"3f",
          3342 => x"08",
          3343 => x"f6",
          3344 => x"88",
          3345 => x"3f",
          3346 => x"64",
          3347 => x"62",
          3348 => x"33",
          3349 => x"79",
          3350 => x"38",
          3351 => x"54",
          3352 => x"7a",
          3353 => x"98",
          3354 => x"eb",
          3355 => x"63",
          3356 => x"5b",
          3357 => x"a7",
          3358 => x"fd",
          3359 => x"ff",
          3360 => x"ff",
          3361 => x"cc",
          3362 => x"bb",
          3363 => x"df",
          3364 => x"84",
          3365 => x"80",
          3366 => x"82",
          3367 => x"45",
          3368 => x"82",
          3369 => x"5a",
          3370 => x"88",
          3371 => x"c4",
          3372 => x"39",
          3373 => x"33",
          3374 => x"2e",
          3375 => x"b9",
          3376 => x"ab",
          3377 => x"87",
          3378 => x"80",
          3379 => x"82",
          3380 => x"45",
          3381 => x"ba",
          3382 => x"79",
          3383 => x"38",
          3384 => x"08",
          3385 => x"82",
          3386 => x"fc",
          3387 => x"b5",
          3388 => x"11",
          3389 => x"05",
          3390 => x"3f",
          3391 => x"08",
          3392 => x"82",
          3393 => x"5a",
          3394 => x"89",
          3395 => x"c0",
          3396 => x"cc",
          3397 => x"85",
          3398 => x"80",
          3399 => x"82",
          3400 => x"44",
          3401 => x"ba",
          3402 => x"79",
          3403 => x"38",
          3404 => x"08",
          3405 => x"82",
          3406 => x"5a",
          3407 => x"88",
          3408 => x"d8",
          3409 => x"39",
          3410 => x"33",
          3411 => x"2e",
          3412 => x"b9",
          3413 => x"88",
          3414 => x"ec",
          3415 => x"44",
          3416 => x"f8",
          3417 => x"84",
          3418 => x"c7",
          3419 => x"98",
          3420 => x"a7",
          3421 => x"5d",
          3422 => x"2e",
          3423 => x"5d",
          3424 => x"70",
          3425 => x"07",
          3426 => x"60",
          3427 => x"5b",
          3428 => x"2e",
          3429 => x"a0",
          3430 => x"88",
          3431 => x"b4",
          3432 => x"3f",
          3433 => x"54",
          3434 => x"52",
          3435 => x"cf",
          3436 => x"c4",
          3437 => x"39",
          3438 => x"80",
          3439 => x"84",
          3440 => x"ef",
          3441 => x"98",
          3442 => x"f5",
          3443 => x"3d",
          3444 => x"53",
          3445 => x"51",
          3446 => x"82",
          3447 => x"80",
          3448 => x"64",
          3449 => x"cf",
          3450 => x"34",
          3451 => x"45",
          3452 => x"fc",
          3453 => x"84",
          3454 => x"b7",
          3455 => x"98",
          3456 => x"f5",
          3457 => x"70",
          3458 => x"82",
          3459 => x"ff",
          3460 => x"80",
          3461 => x"51",
          3462 => x"7a",
          3463 => x"5a",
          3464 => x"f5",
          3465 => x"7a",
          3466 => x"b5",
          3467 => x"11",
          3468 => x"05",
          3469 => x"3f",
          3470 => x"08",
          3471 => x"38",
          3472 => x"80",
          3473 => x"7a",
          3474 => x"05",
          3475 => x"39",
          3476 => x"51",
          3477 => x"ff",
          3478 => x"3d",
          3479 => x"53",
          3480 => x"51",
          3481 => x"82",
          3482 => x"80",
          3483 => x"38",
          3484 => x"f0",
          3485 => x"84",
          3486 => x"b0",
          3487 => x"98",
          3488 => x"a6",
          3489 => x"02",
          3490 => x"22",
          3491 => x"05",
          3492 => x"42",
          3493 => x"f0",
          3494 => x"84",
          3495 => x"8c",
          3496 => x"98",
          3497 => x"f4",
          3498 => x"70",
          3499 => x"82",
          3500 => x"ff",
          3501 => x"80",
          3502 => x"51",
          3503 => x"7a",
          3504 => x"5a",
          3505 => x"f3",
          3506 => x"9f",
          3507 => x"61",
          3508 => x"d6",
          3509 => x"fe",
          3510 => x"ff",
          3511 => x"c1",
          3512 => x"bb",
          3513 => x"2e",
          3514 => x"5a",
          3515 => x"05",
          3516 => x"82",
          3517 => x"79",
          3518 => x"39",
          3519 => x"51",
          3520 => x"ff",
          3521 => x"3d",
          3522 => x"53",
          3523 => x"51",
          3524 => x"82",
          3525 => x"80",
          3526 => x"38",
          3527 => x"f0",
          3528 => x"84",
          3529 => x"84",
          3530 => x"98",
          3531 => x"a0",
          3532 => x"71",
          3533 => x"84",
          3534 => x"3d",
          3535 => x"53",
          3536 => x"51",
          3537 => x"82",
          3538 => x"e5",
          3539 => x"39",
          3540 => x"54",
          3541 => x"f0",
          3542 => x"fb",
          3543 => x"52",
          3544 => x"99",
          3545 => x"7a",
          3546 => x"ae",
          3547 => x"38",
          3548 => x"9b",
          3549 => x"fe",
          3550 => x"ff",
          3551 => x"c0",
          3552 => x"bb",
          3553 => x"2e",
          3554 => x"61",
          3555 => x"61",
          3556 => x"ff",
          3557 => x"a7",
          3558 => x"e8",
          3559 => x"39",
          3560 => x"51",
          3561 => x"82",
          3562 => x"3f",
          3563 => x"82",
          3564 => x"cb",
          3565 => x"51",
          3566 => x"f1",
          3567 => x"a8",
          3568 => x"c0",
          3569 => x"81",
          3570 => x"94",
          3571 => x"80",
          3572 => x"c0",
          3573 => x"f1",
          3574 => x"a8",
          3575 => x"a4",
          3576 => x"83",
          3577 => x"94",
          3578 => x"80",
          3579 => x"c0",
          3580 => x"f1",
          3581 => x"3d",
          3582 => x"53",
          3583 => x"51",
          3584 => x"82",
          3585 => x"80",
          3586 => x"38",
          3587 => x"a8",
          3588 => x"a3",
          3589 => x"5a",
          3590 => x"3d",
          3591 => x"53",
          3592 => x"51",
          3593 => x"82",
          3594 => x"80",
          3595 => x"38",
          3596 => x"a8",
          3597 => x"a3",
          3598 => x"5a",
          3599 => x"bb",
          3600 => x"2e",
          3601 => x"82",
          3602 => x"52",
          3603 => x"51",
          3604 => x"3f",
          3605 => x"82",
          3606 => x"ca",
          3607 => x"a2",
          3608 => x"d2",
          3609 => x"c4",
          3610 => x"3f",
          3611 => x"a8",
          3612 => x"3f",
          3613 => x"7a",
          3614 => x"5a",
          3615 => x"f0",
          3616 => x"7e",
          3617 => x"80",
          3618 => x"38",
          3619 => x"84",
          3620 => x"cf",
          3621 => x"98",
          3622 => x"5d",
          3623 => x"b2",
          3624 => x"24",
          3625 => x"81",
          3626 => x"80",
          3627 => x"83",
          3628 => x"80",
          3629 => x"a9",
          3630 => x"55",
          3631 => x"54",
          3632 => x"a9",
          3633 => x"3d",
          3634 => x"51",
          3635 => x"3f",
          3636 => x"aa",
          3637 => x"3d",
          3638 => x"51",
          3639 => x"3f",
          3640 => x"55",
          3641 => x"54",
          3642 => x"a9",
          3643 => x"3d",
          3644 => x"51",
          3645 => x"3f",
          3646 => x"54",
          3647 => x"a9",
          3648 => x"3d",
          3649 => x"51",
          3650 => x"3f",
          3651 => x"59",
          3652 => x"58",
          3653 => x"57",
          3654 => x"55",
          3655 => x"e0",
          3656 => x"e0",
          3657 => x"3d",
          3658 => x"51",
          3659 => x"82",
          3660 => x"82",
          3661 => x"09",
          3662 => x"72",
          3663 => x"51",
          3664 => x"80",
          3665 => x"26",
          3666 => x"5b",
          3667 => x"5a",
          3668 => x"8d",
          3669 => x"70",
          3670 => x"5e",
          3671 => x"bc",
          3672 => x"32",
          3673 => x"07",
          3674 => x"38",
          3675 => x"09",
          3676 => x"c2",
          3677 => x"84",
          3678 => x"3f",
          3679 => x"f5",
          3680 => x"0b",
          3681 => x"34",
          3682 => x"8c",
          3683 => x"55",
          3684 => x"52",
          3685 => x"8c",
          3686 => x"98",
          3687 => x"75",
          3688 => x"87",
          3689 => x"73",
          3690 => x"3f",
          3691 => x"98",
          3692 => x"0c",
          3693 => x"9c",
          3694 => x"55",
          3695 => x"52",
          3696 => x"e0",
          3697 => x"98",
          3698 => x"75",
          3699 => x"87",
          3700 => x"73",
          3701 => x"3f",
          3702 => x"98",
          3703 => x"0c",
          3704 => x"0b",
          3705 => x"84",
          3706 => x"83",
          3707 => x"94",
          3708 => x"fa",
          3709 => x"fc",
          3710 => x"02",
          3711 => x"05",
          3712 => x"82",
          3713 => x"87",
          3714 => x"13",
          3715 => x"0c",
          3716 => x"0c",
          3717 => x"3f",
          3718 => x"82",
          3719 => x"c6",
          3720 => x"aa",
          3721 => x"dc",
          3722 => x"a8",
          3723 => x"3f",
          3724 => x"b8",
          3725 => x"3f",
          3726 => x"3d",
          3727 => x"83",
          3728 => x"2b",
          3729 => x"3f",
          3730 => x"08",
          3731 => x"72",
          3732 => x"54",
          3733 => x"25",
          3734 => x"82",
          3735 => x"84",
          3736 => x"fc",
          3737 => x"70",
          3738 => x"80",
          3739 => x"72",
          3740 => x"8a",
          3741 => x"51",
          3742 => x"09",
          3743 => x"38",
          3744 => x"f1",
          3745 => x"51",
          3746 => x"09",
          3747 => x"38",
          3748 => x"81",
          3749 => x"73",
          3750 => x"81",
          3751 => x"84",
          3752 => x"52",
          3753 => x"52",
          3754 => x"2e",
          3755 => x"54",
          3756 => x"9d",
          3757 => x"38",
          3758 => x"12",
          3759 => x"33",
          3760 => x"a0",
          3761 => x"81",
          3762 => x"2e",
          3763 => x"ea",
          3764 => x"33",
          3765 => x"a0",
          3766 => x"06",
          3767 => x"54",
          3768 => x"70",
          3769 => x"25",
          3770 => x"51",
          3771 => x"2e",
          3772 => x"72",
          3773 => x"54",
          3774 => x"0c",
          3775 => x"82",
          3776 => x"86",
          3777 => x"fc",
          3778 => x"53",
          3779 => x"2e",
          3780 => x"3d",
          3781 => x"72",
          3782 => x"90",
          3783 => x"98",
          3784 => x"80",
          3785 => x"74",
          3786 => x"bb",
          3787 => x"3d",
          3788 => x"3d",
          3789 => x"11",
          3790 => x"52",
          3791 => x"70",
          3792 => x"98",
          3793 => x"33",
          3794 => x"82",
          3795 => x"26",
          3796 => x"84",
          3797 => x"83",
          3798 => x"26",
          3799 => x"85",
          3800 => x"84",
          3801 => x"26",
          3802 => x"86",
          3803 => x"85",
          3804 => x"26",
          3805 => x"88",
          3806 => x"86",
          3807 => x"e7",
          3808 => x"38",
          3809 => x"54",
          3810 => x"87",
          3811 => x"cc",
          3812 => x"87",
          3813 => x"0c",
          3814 => x"c0",
          3815 => x"82",
          3816 => x"c0",
          3817 => x"83",
          3818 => x"c0",
          3819 => x"84",
          3820 => x"c0",
          3821 => x"85",
          3822 => x"c0",
          3823 => x"86",
          3824 => x"c0",
          3825 => x"74",
          3826 => x"a4",
          3827 => x"c0",
          3828 => x"80",
          3829 => x"98",
          3830 => x"52",
          3831 => x"98",
          3832 => x"0d",
          3833 => x"0d",
          3834 => x"c0",
          3835 => x"81",
          3836 => x"c0",
          3837 => x"5e",
          3838 => x"87",
          3839 => x"08",
          3840 => x"1c",
          3841 => x"98",
          3842 => x"79",
          3843 => x"87",
          3844 => x"08",
          3845 => x"1c",
          3846 => x"98",
          3847 => x"79",
          3848 => x"87",
          3849 => x"08",
          3850 => x"1c",
          3851 => x"98",
          3852 => x"7b",
          3853 => x"87",
          3854 => x"08",
          3855 => x"1c",
          3856 => x"0c",
          3857 => x"ff",
          3858 => x"83",
          3859 => x"58",
          3860 => x"57",
          3861 => x"56",
          3862 => x"55",
          3863 => x"54",
          3864 => x"53",
          3865 => x"ff",
          3866 => x"aa",
          3867 => x"9a",
          3868 => x"3d",
          3869 => x"3d",
          3870 => x"05",
          3871 => x"b8",
          3872 => x"ff",
          3873 => x"55",
          3874 => x"84",
          3875 => x"2e",
          3876 => x"c0",
          3877 => x"70",
          3878 => x"2a",
          3879 => x"53",
          3880 => x"80",
          3881 => x"71",
          3882 => x"81",
          3883 => x"70",
          3884 => x"81",
          3885 => x"06",
          3886 => x"80",
          3887 => x"71",
          3888 => x"81",
          3889 => x"70",
          3890 => x"73",
          3891 => x"51",
          3892 => x"80",
          3893 => x"2e",
          3894 => x"c0",
          3895 => x"74",
          3896 => x"82",
          3897 => x"87",
          3898 => x"ff",
          3899 => x"8f",
          3900 => x"30",
          3901 => x"51",
          3902 => x"82",
          3903 => x"83",
          3904 => x"f9",
          3905 => x"a7",
          3906 => x"77",
          3907 => x"81",
          3908 => x"7a",
          3909 => x"eb",
          3910 => x"b8",
          3911 => x"ff",
          3912 => x"87",
          3913 => x"53",
          3914 => x"86",
          3915 => x"94",
          3916 => x"08",
          3917 => x"70",
          3918 => x"56",
          3919 => x"2e",
          3920 => x"91",
          3921 => x"06",
          3922 => x"d7",
          3923 => x"32",
          3924 => x"51",
          3925 => x"2e",
          3926 => x"93",
          3927 => x"06",
          3928 => x"ff",
          3929 => x"81",
          3930 => x"87",
          3931 => x"54",
          3932 => x"86",
          3933 => x"94",
          3934 => x"74",
          3935 => x"82",
          3936 => x"89",
          3937 => x"f9",
          3938 => x"54",
          3939 => x"70",
          3940 => x"53",
          3941 => x"77",
          3942 => x"38",
          3943 => x"06",
          3944 => x"b9",
          3945 => x"81",
          3946 => x"57",
          3947 => x"c0",
          3948 => x"75",
          3949 => x"38",
          3950 => x"94",
          3951 => x"70",
          3952 => x"81",
          3953 => x"52",
          3954 => x"8c",
          3955 => x"2a",
          3956 => x"51",
          3957 => x"38",
          3958 => x"70",
          3959 => x"51",
          3960 => x"8d",
          3961 => x"2a",
          3962 => x"51",
          3963 => x"be",
          3964 => x"ff",
          3965 => x"c0",
          3966 => x"70",
          3967 => x"38",
          3968 => x"90",
          3969 => x"0c",
          3970 => x"33",
          3971 => x"06",
          3972 => x"70",
          3973 => x"76",
          3974 => x"0c",
          3975 => x"04",
          3976 => x"82",
          3977 => x"70",
          3978 => x"54",
          3979 => x"94",
          3980 => x"80",
          3981 => x"87",
          3982 => x"51",
          3983 => x"82",
          3984 => x"06",
          3985 => x"70",
          3986 => x"38",
          3987 => x"06",
          3988 => x"94",
          3989 => x"80",
          3990 => x"87",
          3991 => x"52",
          3992 => x"81",
          3993 => x"bb",
          3994 => x"84",
          3995 => x"ff",
          3996 => x"bb",
          3997 => x"ff",
          3998 => x"98",
          3999 => x"3d",
          4000 => x"b8",
          4001 => x"ff",
          4002 => x"87",
          4003 => x"52",
          4004 => x"86",
          4005 => x"94",
          4006 => x"08",
          4007 => x"70",
          4008 => x"51",
          4009 => x"70",
          4010 => x"38",
          4011 => x"06",
          4012 => x"94",
          4013 => x"80",
          4014 => x"87",
          4015 => x"52",
          4016 => x"98",
          4017 => x"2c",
          4018 => x"71",
          4019 => x"0c",
          4020 => x"04",
          4021 => x"87",
          4022 => x"08",
          4023 => x"8a",
          4024 => x"70",
          4025 => x"b4",
          4026 => x"9e",
          4027 => x"b9",
          4028 => x"c0",
          4029 => x"82",
          4030 => x"87",
          4031 => x"08",
          4032 => x"0c",
          4033 => x"98",
          4034 => x"c8",
          4035 => x"9e",
          4036 => x"b9",
          4037 => x"c0",
          4038 => x"82",
          4039 => x"87",
          4040 => x"08",
          4041 => x"0c",
          4042 => x"b0",
          4043 => x"d8",
          4044 => x"9e",
          4045 => x"b9",
          4046 => x"c0",
          4047 => x"82",
          4048 => x"87",
          4049 => x"08",
          4050 => x"0c",
          4051 => x"c0",
          4052 => x"e8",
          4053 => x"9e",
          4054 => x"b9",
          4055 => x"c0",
          4056 => x"51",
          4057 => x"f0",
          4058 => x"9e",
          4059 => x"b9",
          4060 => x"c0",
          4061 => x"82",
          4062 => x"87",
          4063 => x"08",
          4064 => x"0c",
          4065 => x"ba",
          4066 => x"0b",
          4067 => x"90",
          4068 => x"80",
          4069 => x"52",
          4070 => x"2e",
          4071 => x"52",
          4072 => x"81",
          4073 => x"87",
          4074 => x"08",
          4075 => x"0a",
          4076 => x"52",
          4077 => x"83",
          4078 => x"71",
          4079 => x"34",
          4080 => x"c0",
          4081 => x"70",
          4082 => x"06",
          4083 => x"70",
          4084 => x"38",
          4085 => x"82",
          4086 => x"80",
          4087 => x"9e",
          4088 => x"88",
          4089 => x"51",
          4090 => x"80",
          4091 => x"81",
          4092 => x"ba",
          4093 => x"0b",
          4094 => x"90",
          4095 => x"80",
          4096 => x"52",
          4097 => x"2e",
          4098 => x"52",
          4099 => x"85",
          4100 => x"87",
          4101 => x"08",
          4102 => x"80",
          4103 => x"52",
          4104 => x"83",
          4105 => x"71",
          4106 => x"34",
          4107 => x"c0",
          4108 => x"70",
          4109 => x"06",
          4110 => x"70",
          4111 => x"38",
          4112 => x"82",
          4113 => x"80",
          4114 => x"9e",
          4115 => x"82",
          4116 => x"51",
          4117 => x"80",
          4118 => x"81",
          4119 => x"ba",
          4120 => x"0b",
          4121 => x"90",
          4122 => x"80",
          4123 => x"52",
          4124 => x"2e",
          4125 => x"52",
          4126 => x"89",
          4127 => x"87",
          4128 => x"08",
          4129 => x"80",
          4130 => x"52",
          4131 => x"83",
          4132 => x"71",
          4133 => x"34",
          4134 => x"c0",
          4135 => x"70",
          4136 => x"51",
          4137 => x"80",
          4138 => x"81",
          4139 => x"ba",
          4140 => x"c0",
          4141 => x"70",
          4142 => x"70",
          4143 => x"51",
          4144 => x"ba",
          4145 => x"0b",
          4146 => x"90",
          4147 => x"80",
          4148 => x"52",
          4149 => x"83",
          4150 => x"71",
          4151 => x"34",
          4152 => x"90",
          4153 => x"f0",
          4154 => x"2a",
          4155 => x"70",
          4156 => x"34",
          4157 => x"c0",
          4158 => x"70",
          4159 => x"52",
          4160 => x"2e",
          4161 => x"52",
          4162 => x"8f",
          4163 => x"9e",
          4164 => x"87",
          4165 => x"70",
          4166 => x"34",
          4167 => x"04",
          4168 => x"82",
          4169 => x"ff",
          4170 => x"82",
          4171 => x"54",
          4172 => x"89",
          4173 => x"e4",
          4174 => x"c8",
          4175 => x"f8",
          4176 => x"c0",
          4177 => x"82",
          4178 => x"80",
          4179 => x"82",
          4180 => x"82",
          4181 => x"11",
          4182 => x"ab",
          4183 => x"90",
          4184 => x"ba",
          4185 => x"73",
          4186 => x"38",
          4187 => x"08",
          4188 => x"08",
          4189 => x"82",
          4190 => x"ff",
          4191 => x"82",
          4192 => x"54",
          4193 => x"94",
          4194 => x"bc",
          4195 => x"c0",
          4196 => x"52",
          4197 => x"51",
          4198 => x"3f",
          4199 => x"33",
          4200 => x"2e",
          4201 => x"b9",
          4202 => x"b9",
          4203 => x"54",
          4204 => x"e4",
          4205 => x"9f",
          4206 => x"86",
          4207 => x"80",
          4208 => x"82",
          4209 => x"82",
          4210 => x"11",
          4211 => x"ac",
          4212 => x"90",
          4213 => x"ba",
          4214 => x"73",
          4215 => x"38",
          4216 => x"33",
          4217 => x"9c",
          4218 => x"eb",
          4219 => x"8f",
          4220 => x"80",
          4221 => x"82",
          4222 => x"52",
          4223 => x"51",
          4224 => x"3f",
          4225 => x"33",
          4226 => x"2e",
          4227 => x"ba",
          4228 => x"82",
          4229 => x"ff",
          4230 => x"82",
          4231 => x"54",
          4232 => x"89",
          4233 => x"fc",
          4234 => x"d8",
          4235 => x"83",
          4236 => x"80",
          4237 => x"82",
          4238 => x"ff",
          4239 => x"82",
          4240 => x"54",
          4241 => x"89",
          4242 => x"9c",
          4243 => x"b4",
          4244 => x"89",
          4245 => x"80",
          4246 => x"82",
          4247 => x"ff",
          4248 => x"82",
          4249 => x"54",
          4250 => x"89",
          4251 => x"b4",
          4252 => x"90",
          4253 => x"c0",
          4254 => x"88",
          4255 => x"e4",
          4256 => x"ad",
          4257 => x"8e",
          4258 => x"b9",
          4259 => x"82",
          4260 => x"ff",
          4261 => x"82",
          4262 => x"52",
          4263 => x"51",
          4264 => x"3f",
          4265 => x"51",
          4266 => x"3f",
          4267 => x"22",
          4268 => x"cc",
          4269 => x"9f",
          4270 => x"f4",
          4271 => x"84",
          4272 => x"51",
          4273 => x"82",
          4274 => x"bd",
          4275 => x"76",
          4276 => x"54",
          4277 => x"08",
          4278 => x"f4",
          4279 => x"f7",
          4280 => x"87",
          4281 => x"80",
          4282 => x"82",
          4283 => x"56",
          4284 => x"52",
          4285 => x"ac",
          4286 => x"98",
          4287 => x"c0",
          4288 => x"31",
          4289 => x"bb",
          4290 => x"82",
          4291 => x"ff",
          4292 => x"82",
          4293 => x"54",
          4294 => x"a9",
          4295 => x"fc",
          4296 => x"84",
          4297 => x"51",
          4298 => x"82",
          4299 => x"bd",
          4300 => x"76",
          4301 => x"54",
          4302 => x"08",
          4303 => x"cc",
          4304 => x"93",
          4305 => x"b0",
          4306 => x"b8",
          4307 => x"0d",
          4308 => x"0d",
          4309 => x"33",
          4310 => x"71",
          4311 => x"38",
          4312 => x"82",
          4313 => x"52",
          4314 => x"82",
          4315 => x"9d",
          4316 => x"80",
          4317 => x"82",
          4318 => x"91",
          4319 => x"90",
          4320 => x"82",
          4321 => x"85",
          4322 => x"9c",
          4323 => x"f4",
          4324 => x"0d",
          4325 => x"80",
          4326 => x"3d",
          4327 => x"96",
          4328 => x"52",
          4329 => x"0c",
          4330 => x"70",
          4331 => x"0c",
          4332 => x"3d",
          4333 => x"3d",
          4334 => x"96",
          4335 => x"82",
          4336 => x"52",
          4337 => x"73",
          4338 => x"ba",
          4339 => x"70",
          4340 => x"0c",
          4341 => x"83",
          4342 => x"80",
          4343 => x"96",
          4344 => x"82",
          4345 => x"87",
          4346 => x"0c",
          4347 => x"0d",
          4348 => x"70",
          4349 => x"98",
          4350 => x"2c",
          4351 => x"70",
          4352 => x"53",
          4353 => x"51",
          4354 => x"b0",
          4355 => x"55",
          4356 => x"25",
          4357 => x"b0",
          4358 => x"12",
          4359 => x"97",
          4360 => x"33",
          4361 => x"70",
          4362 => x"81",
          4363 => x"81",
          4364 => x"bb",
          4365 => x"3d",
          4366 => x"3d",
          4367 => x"84",
          4368 => x"33",
          4369 => x"55",
          4370 => x"2e",
          4371 => x"51",
          4372 => x"3f",
          4373 => x"b5",
          4374 => x"51",
          4375 => x"3f",
          4376 => x"05",
          4377 => x"34",
          4378 => x"06",
          4379 => x"76",
          4380 => x"90",
          4381 => x"34",
          4382 => x"04",
          4383 => x"7c",
          4384 => x"b7",
          4385 => x"88",
          4386 => x"33",
          4387 => x"33",
          4388 => x"82",
          4389 => x"70",
          4390 => x"59",
          4391 => x"74",
          4392 => x"38",
          4393 => x"b5",
          4394 => x"f0",
          4395 => x"29",
          4396 => x"05",
          4397 => x"54",
          4398 => x"9d",
          4399 => x"bb",
          4400 => x"0c",
          4401 => x"33",
          4402 => x"82",
          4403 => x"70",
          4404 => x"5a",
          4405 => x"a7",
          4406 => x"78",
          4407 => x"ff",
          4408 => x"82",
          4409 => x"81",
          4410 => x"82",
          4411 => x"74",
          4412 => x"55",
          4413 => x"87",
          4414 => x"82",
          4415 => x"77",
          4416 => x"38",
          4417 => x"08",
          4418 => x"2e",
          4419 => x"ba",
          4420 => x"74",
          4421 => x"3d",
          4422 => x"76",
          4423 => x"75",
          4424 => x"c3",
          4425 => x"ec",
          4426 => x"51",
          4427 => x"3f",
          4428 => x"08",
          4429 => x"a0",
          4430 => x"0d",
          4431 => x"0d",
          4432 => x"53",
          4433 => x"08",
          4434 => x"2e",
          4435 => x"51",
          4436 => x"80",
          4437 => x"14",
          4438 => x"54",
          4439 => x"e6",
          4440 => x"82",
          4441 => x"82",
          4442 => x"52",
          4443 => x"95",
          4444 => x"80",
          4445 => x"82",
          4446 => x"51",
          4447 => x"80",
          4448 => x"ec",
          4449 => x"0d",
          4450 => x"0d",
          4451 => x"52",
          4452 => x"08",
          4453 => x"ed",
          4454 => x"98",
          4455 => x"38",
          4456 => x"08",
          4457 => x"52",
          4458 => x"52",
          4459 => x"bb",
          4460 => x"98",
          4461 => x"ba",
          4462 => x"ff",
          4463 => x"82",
          4464 => x"55",
          4465 => x"bb",
          4466 => x"9d",
          4467 => x"98",
          4468 => x"70",
          4469 => x"80",
          4470 => x"53",
          4471 => x"17",
          4472 => x"52",
          4473 => x"ef",
          4474 => x"2e",
          4475 => x"ff",
          4476 => x"3d",
          4477 => x"3d",
          4478 => x"08",
          4479 => x"5a",
          4480 => x"58",
          4481 => x"82",
          4482 => x"51",
          4483 => x"3f",
          4484 => x"08",
          4485 => x"ff",
          4486 => x"ec",
          4487 => x"80",
          4488 => x"3d",
          4489 => x"81",
          4490 => x"82",
          4491 => x"80",
          4492 => x"75",
          4493 => x"ee",
          4494 => x"98",
          4495 => x"58",
          4496 => x"82",
          4497 => x"25",
          4498 => x"bb",
          4499 => x"05",
          4500 => x"55",
          4501 => x"74",
          4502 => x"70",
          4503 => x"2a",
          4504 => x"78",
          4505 => x"38",
          4506 => x"38",
          4507 => x"08",
          4508 => x"53",
          4509 => x"8d",
          4510 => x"98",
          4511 => x"89",
          4512 => x"a4",
          4513 => x"fc",
          4514 => x"2e",
          4515 => x"9b",
          4516 => x"79",
          4517 => x"fc",
          4518 => x"ff",
          4519 => x"ab",
          4520 => x"82",
          4521 => x"74",
          4522 => x"77",
          4523 => x"0c",
          4524 => x"04",
          4525 => x"7c",
          4526 => x"71",
          4527 => x"59",
          4528 => x"a0",
          4529 => x"06",
          4530 => x"33",
          4531 => x"77",
          4532 => x"38",
          4533 => x"5b",
          4534 => x"56",
          4535 => x"a0",
          4536 => x"06",
          4537 => x"75",
          4538 => x"80",
          4539 => x"29",
          4540 => x"05",
          4541 => x"55",
          4542 => x"3f",
          4543 => x"08",
          4544 => x"74",
          4545 => x"bc",
          4546 => x"bb",
          4547 => x"c6",
          4548 => x"33",
          4549 => x"2e",
          4550 => x"82",
          4551 => x"b6",
          4552 => x"3f",
          4553 => x"1a",
          4554 => x"fc",
          4555 => x"05",
          4556 => x"ff",
          4557 => x"98",
          4558 => x"9a",
          4559 => x"53",
          4560 => x"51",
          4561 => x"82",
          4562 => x"81",
          4563 => x"74",
          4564 => x"54",
          4565 => x"14",
          4566 => x"06",
          4567 => x"74",
          4568 => x"38",
          4569 => x"82",
          4570 => x"8c",
          4571 => x"d3",
          4572 => x"3d",
          4573 => x"08",
          4574 => x"59",
          4575 => x"0b",
          4576 => x"82",
          4577 => x"82",
          4578 => x"55",
          4579 => x"cb",
          4580 => x"ba",
          4581 => x"55",
          4582 => x"81",
          4583 => x"2e",
          4584 => x"81",
          4585 => x"55",
          4586 => x"2e",
          4587 => x"a8",
          4588 => x"3f",
          4589 => x"08",
          4590 => x"0c",
          4591 => x"08",
          4592 => x"92",
          4593 => x"76",
          4594 => x"98",
          4595 => x"cc",
          4596 => x"bb",
          4597 => x"2e",
          4598 => x"b3",
          4599 => x"ab",
          4600 => x"f7",
          4601 => x"98",
          4602 => x"ba",
          4603 => x"80",
          4604 => x"3d",
          4605 => x"81",
          4606 => x"82",
          4607 => x"56",
          4608 => x"08",
          4609 => x"81",
          4610 => x"38",
          4611 => x"08",
          4612 => x"92",
          4613 => x"98",
          4614 => x"0b",
          4615 => x"08",
          4616 => x"82",
          4617 => x"ff",
          4618 => x"55",
          4619 => x"34",
          4620 => x"81",
          4621 => x"75",
          4622 => x"3f",
          4623 => x"81",
          4624 => x"54",
          4625 => x"83",
          4626 => x"74",
          4627 => x"81",
          4628 => x"38",
          4629 => x"82",
          4630 => x"76",
          4631 => x"ba",
          4632 => x"2e",
          4633 => x"d5",
          4634 => x"5d",
          4635 => x"82",
          4636 => x"98",
          4637 => x"2c",
          4638 => x"ff",
          4639 => x"78",
          4640 => x"82",
          4641 => x"70",
          4642 => x"98",
          4643 => x"c0",
          4644 => x"2b",
          4645 => x"71",
          4646 => x"70",
          4647 => x"b0",
          4648 => x"08",
          4649 => x"51",
          4650 => x"59",
          4651 => x"5d",
          4652 => x"73",
          4653 => x"e9",
          4654 => x"27",
          4655 => x"81",
          4656 => x"81",
          4657 => x"70",
          4658 => x"55",
          4659 => x"80",
          4660 => x"53",
          4661 => x"51",
          4662 => x"82",
          4663 => x"81",
          4664 => x"73",
          4665 => x"38",
          4666 => x"c0",
          4667 => x"b1",
          4668 => x"80",
          4669 => x"80",
          4670 => x"98",
          4671 => x"ff",
          4672 => x"55",
          4673 => x"97",
          4674 => x"74",
          4675 => x"f5",
          4676 => x"bb",
          4677 => x"ff",
          4678 => x"cc",
          4679 => x"80",
          4680 => x"2e",
          4681 => x"81",
          4682 => x"82",
          4683 => x"74",
          4684 => x"98",
          4685 => x"c0",
          4686 => x"2b",
          4687 => x"70",
          4688 => x"82",
          4689 => x"a8",
          4690 => x"51",
          4691 => x"58",
          4692 => x"77",
          4693 => x"06",
          4694 => x"82",
          4695 => x"08",
          4696 => x"0b",
          4697 => x"34",
          4698 => x"d2",
          4699 => x"39",
          4700 => x"c4",
          4701 => x"d2",
          4702 => x"af",
          4703 => x"7d",
          4704 => x"73",
          4705 => x"e1",
          4706 => x"29",
          4707 => x"05",
          4708 => x"04",
          4709 => x"33",
          4710 => x"2e",
          4711 => x"82",
          4712 => x"55",
          4713 => x"ab",
          4714 => x"2b",
          4715 => x"51",
          4716 => x"24",
          4717 => x"1a",
          4718 => x"81",
          4719 => x"81",
          4720 => x"81",
          4721 => x"70",
          4722 => x"d2",
          4723 => x"51",
          4724 => x"82",
          4725 => x"81",
          4726 => x"74",
          4727 => x"34",
          4728 => x"ae",
          4729 => x"34",
          4730 => x"33",
          4731 => x"25",
          4732 => x"14",
          4733 => x"d2",
          4734 => x"d2",
          4735 => x"81",
          4736 => x"81",
          4737 => x"70",
          4738 => x"d2",
          4739 => x"51",
          4740 => x"77",
          4741 => x"74",
          4742 => x"52",
          4743 => x"86",
          4744 => x"80",
          4745 => x"80",
          4746 => x"98",
          4747 => x"c8",
          4748 => x"55",
          4749 => x"df",
          4750 => x"cc",
          4751 => x"2b",
          4752 => x"82",
          4753 => x"5a",
          4754 => x"74",
          4755 => x"99",
          4756 => x"ff",
          4757 => x"74",
          4758 => x"29",
          4759 => x"05",
          4760 => x"82",
          4761 => x"56",
          4762 => x"75",
          4763 => x"fb",
          4764 => x"7a",
          4765 => x"81",
          4766 => x"d2",
          4767 => x"52",
          4768 => x"51",
          4769 => x"81",
          4770 => x"d2",
          4771 => x"81",
          4772 => x"55",
          4773 => x"fb",
          4774 => x"d2",
          4775 => x"05",
          4776 => x"d2",
          4777 => x"15",
          4778 => x"d2",
          4779 => x"51",
          4780 => x"3f",
          4781 => x"33",
          4782 => x"70",
          4783 => x"d2",
          4784 => x"51",
          4785 => x"74",
          4786 => x"74",
          4787 => x"14",
          4788 => x"73",
          4789 => x"a8",
          4790 => x"81",
          4791 => x"81",
          4792 => x"70",
          4793 => x"d2",
          4794 => x"51",
          4795 => x"24",
          4796 => x"51",
          4797 => x"3f",
          4798 => x"33",
          4799 => x"70",
          4800 => x"d2",
          4801 => x"51",
          4802 => x"74",
          4803 => x"38",
          4804 => x"a8",
          4805 => x"81",
          4806 => x"81",
          4807 => x"70",
          4808 => x"d2",
          4809 => x"51",
          4810 => x"25",
          4811 => x"b9",
          4812 => x"c8",
          4813 => x"54",
          4814 => x"8a",
          4815 => x"e6",
          4816 => x"c8",
          4817 => x"f6",
          4818 => x"bb",
          4819 => x"ff",
          4820 => x"96",
          4821 => x"c8",
          4822 => x"80",
          4823 => x"81",
          4824 => x"79",
          4825 => x"3f",
          4826 => x"7a",
          4827 => x"82",
          4828 => x"80",
          4829 => x"c8",
          4830 => x"bb",
          4831 => x"3d",
          4832 => x"d2",
          4833 => x"73",
          4834 => x"dd",
          4835 => x"ff",
          4836 => x"82",
          4837 => x"ff",
          4838 => x"82",
          4839 => x"73",
          4840 => x"54",
          4841 => x"d2",
          4842 => x"d2",
          4843 => x"55",
          4844 => x"f9",
          4845 => x"14",
          4846 => x"d2",
          4847 => x"98",
          4848 => x"2c",
          4849 => x"06",
          4850 => x"74",
          4851 => x"38",
          4852 => x"81",
          4853 => x"34",
          4854 => x"ff",
          4855 => x"74",
          4856 => x"29",
          4857 => x"05",
          4858 => x"82",
          4859 => x"58",
          4860 => x"75",
          4861 => x"a0",
          4862 => x"aa",
          4863 => x"cc",
          4864 => x"2b",
          4865 => x"82",
          4866 => x"57",
          4867 => x"74",
          4868 => x"d5",
          4869 => x"ff",
          4870 => x"74",
          4871 => x"29",
          4872 => x"05",
          4873 => x"82",
          4874 => x"58",
          4875 => x"75",
          4876 => x"f8",
          4877 => x"d2",
          4878 => x"81",
          4879 => x"d2",
          4880 => x"56",
          4881 => x"27",
          4882 => x"81",
          4883 => x"82",
          4884 => x"74",
          4885 => x"52",
          4886 => x"ca",
          4887 => x"cc",
          4888 => x"ff",
          4889 => x"c8",
          4890 => x"54",
          4891 => x"db",
          4892 => x"39",
          4893 => x"53",
          4894 => x"a9",
          4895 => x"ba",
          4896 => x"82",
          4897 => x"80",
          4898 => x"c8",
          4899 => x"39",
          4900 => x"82",
          4901 => x"55",
          4902 => x"a6",
          4903 => x"ff",
          4904 => x"82",
          4905 => x"82",
          4906 => x"82",
          4907 => x"81",
          4908 => x"05",
          4909 => x"79",
          4910 => x"ca",
          4911 => x"81",
          4912 => x"84",
          4913 => x"98",
          4914 => x"08",
          4915 => x"80",
          4916 => x"74",
          4917 => x"ce",
          4918 => x"98",
          4919 => x"c8",
          4920 => x"98",
          4921 => x"06",
          4922 => x"74",
          4923 => x"ff",
          4924 => x"ff",
          4925 => x"fa",
          4926 => x"55",
          4927 => x"f6",
          4928 => x"51",
          4929 => x"3f",
          4930 => x"93",
          4931 => x"06",
          4932 => x"ba",
          4933 => x"74",
          4934 => x"38",
          4935 => x"ad",
          4936 => x"bb",
          4937 => x"d2",
          4938 => x"bb",
          4939 => x"ff",
          4940 => x"53",
          4941 => x"51",
          4942 => x"3f",
          4943 => x"7a",
          4944 => x"ba",
          4945 => x"08",
          4946 => x"80",
          4947 => x"74",
          4948 => x"d2",
          4949 => x"98",
          4950 => x"c8",
          4951 => x"98",
          4952 => x"06",
          4953 => x"74",
          4954 => x"ff",
          4955 => x"81",
          4956 => x"81",
          4957 => x"89",
          4958 => x"d2",
          4959 => x"7a",
          4960 => x"cc",
          4961 => x"c8",
          4962 => x"51",
          4963 => x"f5",
          4964 => x"d2",
          4965 => x"81",
          4966 => x"d2",
          4967 => x"56",
          4968 => x"27",
          4969 => x"81",
          4970 => x"82",
          4971 => x"74",
          4972 => x"52",
          4973 => x"ee",
          4974 => x"39",
          4975 => x"33",
          4976 => x"2e",
          4977 => x"88",
          4978 => x"da",
          4979 => x"cc",
          4980 => x"54",
          4981 => x"cc",
          4982 => x"39",
          4983 => x"83",
          4984 => x"82",
          4985 => x"84",
          4986 => x"bb",
          4987 => x"80",
          4988 => x"83",
          4989 => x"ff",
          4990 => x"82",
          4991 => x"54",
          4992 => x"74",
          4993 => x"76",
          4994 => x"82",
          4995 => x"54",
          4996 => x"34",
          4997 => x"34",
          4998 => x"08",
          4999 => x"15",
          5000 => x"15",
          5001 => x"90",
          5002 => x"8c",
          5003 => x"fe",
          5004 => x"70",
          5005 => x"06",
          5006 => x"58",
          5007 => x"74",
          5008 => x"73",
          5009 => x"82",
          5010 => x"70",
          5011 => x"bb",
          5012 => x"f8",
          5013 => x"55",
          5014 => x"34",
          5015 => x"34",
          5016 => x"04",
          5017 => x"73",
          5018 => x"84",
          5019 => x"38",
          5020 => x"2a",
          5021 => x"83",
          5022 => x"51",
          5023 => x"82",
          5024 => x"83",
          5025 => x"f9",
          5026 => x"a6",
          5027 => x"84",
          5028 => x"22",
          5029 => x"bb",
          5030 => x"83",
          5031 => x"74",
          5032 => x"11",
          5033 => x"12",
          5034 => x"2b",
          5035 => x"05",
          5036 => x"71",
          5037 => x"06",
          5038 => x"2a",
          5039 => x"59",
          5040 => x"57",
          5041 => x"71",
          5042 => x"81",
          5043 => x"bb",
          5044 => x"75",
          5045 => x"54",
          5046 => x"34",
          5047 => x"34",
          5048 => x"08",
          5049 => x"33",
          5050 => x"71",
          5051 => x"70",
          5052 => x"ff",
          5053 => x"52",
          5054 => x"05",
          5055 => x"ff",
          5056 => x"2a",
          5057 => x"71",
          5058 => x"72",
          5059 => x"53",
          5060 => x"34",
          5061 => x"08",
          5062 => x"76",
          5063 => x"17",
          5064 => x"0d",
          5065 => x"0d",
          5066 => x"08",
          5067 => x"9e",
          5068 => x"83",
          5069 => x"86",
          5070 => x"12",
          5071 => x"2b",
          5072 => x"07",
          5073 => x"52",
          5074 => x"05",
          5075 => x"85",
          5076 => x"88",
          5077 => x"88",
          5078 => x"56",
          5079 => x"13",
          5080 => x"13",
          5081 => x"90",
          5082 => x"84",
          5083 => x"12",
          5084 => x"2b",
          5085 => x"07",
          5086 => x"52",
          5087 => x"12",
          5088 => x"33",
          5089 => x"07",
          5090 => x"54",
          5091 => x"70",
          5092 => x"73",
          5093 => x"82",
          5094 => x"13",
          5095 => x"12",
          5096 => x"2b",
          5097 => x"ff",
          5098 => x"88",
          5099 => x"53",
          5100 => x"73",
          5101 => x"14",
          5102 => x"0d",
          5103 => x"0d",
          5104 => x"22",
          5105 => x"08",
          5106 => x"71",
          5107 => x"81",
          5108 => x"88",
          5109 => x"88",
          5110 => x"33",
          5111 => x"71",
          5112 => x"90",
          5113 => x"5f",
          5114 => x"5a",
          5115 => x"54",
          5116 => x"80",
          5117 => x"51",
          5118 => x"82",
          5119 => x"70",
          5120 => x"81",
          5121 => x"8b",
          5122 => x"2b",
          5123 => x"70",
          5124 => x"33",
          5125 => x"07",
          5126 => x"8f",
          5127 => x"51",
          5128 => x"53",
          5129 => x"72",
          5130 => x"2a",
          5131 => x"82",
          5132 => x"83",
          5133 => x"bb",
          5134 => x"16",
          5135 => x"12",
          5136 => x"2b",
          5137 => x"07",
          5138 => x"55",
          5139 => x"33",
          5140 => x"71",
          5141 => x"70",
          5142 => x"06",
          5143 => x"57",
          5144 => x"52",
          5145 => x"71",
          5146 => x"88",
          5147 => x"fb",
          5148 => x"bb",
          5149 => x"84",
          5150 => x"22",
          5151 => x"72",
          5152 => x"33",
          5153 => x"71",
          5154 => x"83",
          5155 => x"5b",
          5156 => x"52",
          5157 => x"33",
          5158 => x"71",
          5159 => x"02",
          5160 => x"05",
          5161 => x"70",
          5162 => x"51",
          5163 => x"71",
          5164 => x"81",
          5165 => x"bb",
          5166 => x"15",
          5167 => x"12",
          5168 => x"2b",
          5169 => x"07",
          5170 => x"52",
          5171 => x"12",
          5172 => x"33",
          5173 => x"07",
          5174 => x"54",
          5175 => x"70",
          5176 => x"72",
          5177 => x"82",
          5178 => x"14",
          5179 => x"83",
          5180 => x"88",
          5181 => x"bb",
          5182 => x"54",
          5183 => x"04",
          5184 => x"7b",
          5185 => x"08",
          5186 => x"70",
          5187 => x"06",
          5188 => x"53",
          5189 => x"82",
          5190 => x"76",
          5191 => x"11",
          5192 => x"83",
          5193 => x"8b",
          5194 => x"2b",
          5195 => x"70",
          5196 => x"33",
          5197 => x"71",
          5198 => x"53",
          5199 => x"53",
          5200 => x"59",
          5201 => x"25",
          5202 => x"80",
          5203 => x"51",
          5204 => x"81",
          5205 => x"14",
          5206 => x"33",
          5207 => x"71",
          5208 => x"76",
          5209 => x"2a",
          5210 => x"58",
          5211 => x"14",
          5212 => x"ff",
          5213 => x"87",
          5214 => x"bb",
          5215 => x"19",
          5216 => x"85",
          5217 => x"88",
          5218 => x"88",
          5219 => x"5b",
          5220 => x"84",
          5221 => x"85",
          5222 => x"bb",
          5223 => x"53",
          5224 => x"14",
          5225 => x"87",
          5226 => x"bb",
          5227 => x"76",
          5228 => x"75",
          5229 => x"82",
          5230 => x"18",
          5231 => x"12",
          5232 => x"2b",
          5233 => x"80",
          5234 => x"88",
          5235 => x"55",
          5236 => x"74",
          5237 => x"15",
          5238 => x"0d",
          5239 => x"0d",
          5240 => x"bb",
          5241 => x"38",
          5242 => x"71",
          5243 => x"38",
          5244 => x"8c",
          5245 => x"0d",
          5246 => x"0d",
          5247 => x"58",
          5248 => x"82",
          5249 => x"83",
          5250 => x"82",
          5251 => x"84",
          5252 => x"12",
          5253 => x"2b",
          5254 => x"59",
          5255 => x"81",
          5256 => x"75",
          5257 => x"cb",
          5258 => x"29",
          5259 => x"81",
          5260 => x"88",
          5261 => x"81",
          5262 => x"79",
          5263 => x"ff",
          5264 => x"7f",
          5265 => x"51",
          5266 => x"77",
          5267 => x"38",
          5268 => x"85",
          5269 => x"5a",
          5270 => x"33",
          5271 => x"71",
          5272 => x"57",
          5273 => x"38",
          5274 => x"ff",
          5275 => x"7a",
          5276 => x"80",
          5277 => x"82",
          5278 => x"11",
          5279 => x"12",
          5280 => x"2b",
          5281 => x"ff",
          5282 => x"52",
          5283 => x"55",
          5284 => x"83",
          5285 => x"80",
          5286 => x"26",
          5287 => x"74",
          5288 => x"2e",
          5289 => x"77",
          5290 => x"81",
          5291 => x"75",
          5292 => x"3f",
          5293 => x"82",
          5294 => x"79",
          5295 => x"f7",
          5296 => x"bb",
          5297 => x"1c",
          5298 => x"87",
          5299 => x"8b",
          5300 => x"2b",
          5301 => x"5e",
          5302 => x"7a",
          5303 => x"ff",
          5304 => x"88",
          5305 => x"56",
          5306 => x"15",
          5307 => x"ff",
          5308 => x"85",
          5309 => x"bb",
          5310 => x"83",
          5311 => x"72",
          5312 => x"33",
          5313 => x"71",
          5314 => x"70",
          5315 => x"5b",
          5316 => x"56",
          5317 => x"19",
          5318 => x"19",
          5319 => x"90",
          5320 => x"84",
          5321 => x"12",
          5322 => x"2b",
          5323 => x"07",
          5324 => x"55",
          5325 => x"78",
          5326 => x"76",
          5327 => x"82",
          5328 => x"70",
          5329 => x"84",
          5330 => x"12",
          5331 => x"2b",
          5332 => x"2a",
          5333 => x"52",
          5334 => x"84",
          5335 => x"85",
          5336 => x"bb",
          5337 => x"84",
          5338 => x"82",
          5339 => x"8d",
          5340 => x"fe",
          5341 => x"52",
          5342 => x"08",
          5343 => x"dc",
          5344 => x"71",
          5345 => x"38",
          5346 => x"ed",
          5347 => x"98",
          5348 => x"82",
          5349 => x"84",
          5350 => x"ee",
          5351 => x"66",
          5352 => x"70",
          5353 => x"bb",
          5354 => x"2e",
          5355 => x"84",
          5356 => x"3f",
          5357 => x"7e",
          5358 => x"3f",
          5359 => x"08",
          5360 => x"39",
          5361 => x"7b",
          5362 => x"3f",
          5363 => x"ba",
          5364 => x"f5",
          5365 => x"bb",
          5366 => x"ff",
          5367 => x"bb",
          5368 => x"71",
          5369 => x"70",
          5370 => x"06",
          5371 => x"73",
          5372 => x"81",
          5373 => x"88",
          5374 => x"75",
          5375 => x"ff",
          5376 => x"88",
          5377 => x"73",
          5378 => x"70",
          5379 => x"33",
          5380 => x"07",
          5381 => x"53",
          5382 => x"48",
          5383 => x"54",
          5384 => x"56",
          5385 => x"80",
          5386 => x"76",
          5387 => x"06",
          5388 => x"83",
          5389 => x"42",
          5390 => x"33",
          5391 => x"71",
          5392 => x"70",
          5393 => x"70",
          5394 => x"33",
          5395 => x"71",
          5396 => x"53",
          5397 => x"56",
          5398 => x"25",
          5399 => x"75",
          5400 => x"ff",
          5401 => x"54",
          5402 => x"81",
          5403 => x"18",
          5404 => x"2e",
          5405 => x"8f",
          5406 => x"f6",
          5407 => x"83",
          5408 => x"58",
          5409 => x"7f",
          5410 => x"74",
          5411 => x"78",
          5412 => x"3f",
          5413 => x"7f",
          5414 => x"75",
          5415 => x"38",
          5416 => x"11",
          5417 => x"33",
          5418 => x"07",
          5419 => x"f4",
          5420 => x"52",
          5421 => x"b7",
          5422 => x"98",
          5423 => x"ff",
          5424 => x"7c",
          5425 => x"2b",
          5426 => x"08",
          5427 => x"53",
          5428 => x"9a",
          5429 => x"bb",
          5430 => x"84",
          5431 => x"ff",
          5432 => x"5c",
          5433 => x"60",
          5434 => x"74",
          5435 => x"38",
          5436 => x"c9",
          5437 => x"90",
          5438 => x"11",
          5439 => x"33",
          5440 => x"07",
          5441 => x"f4",
          5442 => x"52",
          5443 => x"df",
          5444 => x"98",
          5445 => x"ff",
          5446 => x"7c",
          5447 => x"2b",
          5448 => x"08",
          5449 => x"53",
          5450 => x"9a",
          5451 => x"bb",
          5452 => x"84",
          5453 => x"05",
          5454 => x"73",
          5455 => x"06",
          5456 => x"7b",
          5457 => x"f9",
          5458 => x"bb",
          5459 => x"82",
          5460 => x"80",
          5461 => x"7d",
          5462 => x"82",
          5463 => x"51",
          5464 => x"3f",
          5465 => x"98",
          5466 => x"7a",
          5467 => x"38",
          5468 => x"52",
          5469 => x"8f",
          5470 => x"83",
          5471 => x"90",
          5472 => x"05",
          5473 => x"3f",
          5474 => x"82",
          5475 => x"94",
          5476 => x"fc",
          5477 => x"77",
          5478 => x"54",
          5479 => x"82",
          5480 => x"55",
          5481 => x"08",
          5482 => x"38",
          5483 => x"52",
          5484 => x"08",
          5485 => x"cf",
          5486 => x"bb",
          5487 => x"3d",
          5488 => x"3d",
          5489 => x"05",
          5490 => x"52",
          5491 => x"87",
          5492 => x"94",
          5493 => x"71",
          5494 => x"0c",
          5495 => x"04",
          5496 => x"02",
          5497 => x"02",
          5498 => x"05",
          5499 => x"83",
          5500 => x"26",
          5501 => x"72",
          5502 => x"c0",
          5503 => x"53",
          5504 => x"74",
          5505 => x"38",
          5506 => x"73",
          5507 => x"c0",
          5508 => x"51",
          5509 => x"85",
          5510 => x"98",
          5511 => x"52",
          5512 => x"82",
          5513 => x"70",
          5514 => x"38",
          5515 => x"8c",
          5516 => x"ec",
          5517 => x"fc",
          5518 => x"52",
          5519 => x"87",
          5520 => x"08",
          5521 => x"2e",
          5522 => x"82",
          5523 => x"34",
          5524 => x"13",
          5525 => x"82",
          5526 => x"86",
          5527 => x"f3",
          5528 => x"62",
          5529 => x"05",
          5530 => x"57",
          5531 => x"83",
          5532 => x"fe",
          5533 => x"bb",
          5534 => x"06",
          5535 => x"71",
          5536 => x"71",
          5537 => x"2b",
          5538 => x"80",
          5539 => x"92",
          5540 => x"c0",
          5541 => x"41",
          5542 => x"5a",
          5543 => x"87",
          5544 => x"0c",
          5545 => x"84",
          5546 => x"08",
          5547 => x"70",
          5548 => x"53",
          5549 => x"2e",
          5550 => x"08",
          5551 => x"70",
          5552 => x"34",
          5553 => x"80",
          5554 => x"53",
          5555 => x"2e",
          5556 => x"53",
          5557 => x"26",
          5558 => x"80",
          5559 => x"87",
          5560 => x"08",
          5561 => x"38",
          5562 => x"8c",
          5563 => x"80",
          5564 => x"78",
          5565 => x"99",
          5566 => x"0c",
          5567 => x"8c",
          5568 => x"08",
          5569 => x"51",
          5570 => x"38",
          5571 => x"8d",
          5572 => x"17",
          5573 => x"81",
          5574 => x"53",
          5575 => x"2e",
          5576 => x"fc",
          5577 => x"52",
          5578 => x"7d",
          5579 => x"ed",
          5580 => x"80",
          5581 => x"71",
          5582 => x"38",
          5583 => x"53",
          5584 => x"98",
          5585 => x"0d",
          5586 => x"0d",
          5587 => x"02",
          5588 => x"05",
          5589 => x"58",
          5590 => x"80",
          5591 => x"fc",
          5592 => x"bb",
          5593 => x"06",
          5594 => x"71",
          5595 => x"81",
          5596 => x"38",
          5597 => x"2b",
          5598 => x"80",
          5599 => x"92",
          5600 => x"c0",
          5601 => x"40",
          5602 => x"5a",
          5603 => x"c0",
          5604 => x"76",
          5605 => x"76",
          5606 => x"75",
          5607 => x"2a",
          5608 => x"51",
          5609 => x"80",
          5610 => x"7a",
          5611 => x"5c",
          5612 => x"81",
          5613 => x"81",
          5614 => x"06",
          5615 => x"80",
          5616 => x"87",
          5617 => x"08",
          5618 => x"38",
          5619 => x"8c",
          5620 => x"80",
          5621 => x"77",
          5622 => x"99",
          5623 => x"0c",
          5624 => x"8c",
          5625 => x"08",
          5626 => x"51",
          5627 => x"38",
          5628 => x"8d",
          5629 => x"70",
          5630 => x"84",
          5631 => x"5b",
          5632 => x"2e",
          5633 => x"fc",
          5634 => x"52",
          5635 => x"7d",
          5636 => x"f8",
          5637 => x"80",
          5638 => x"71",
          5639 => x"38",
          5640 => x"53",
          5641 => x"98",
          5642 => x"0d",
          5643 => x"0d",
          5644 => x"05",
          5645 => x"02",
          5646 => x"05",
          5647 => x"54",
          5648 => x"fe",
          5649 => x"98",
          5650 => x"53",
          5651 => x"80",
          5652 => x"0b",
          5653 => x"8c",
          5654 => x"71",
          5655 => x"dc",
          5656 => x"24",
          5657 => x"84",
          5658 => x"92",
          5659 => x"54",
          5660 => x"8d",
          5661 => x"39",
          5662 => x"80",
          5663 => x"cb",
          5664 => x"70",
          5665 => x"81",
          5666 => x"52",
          5667 => x"8a",
          5668 => x"98",
          5669 => x"71",
          5670 => x"c0",
          5671 => x"52",
          5672 => x"81",
          5673 => x"c0",
          5674 => x"53",
          5675 => x"82",
          5676 => x"71",
          5677 => x"39",
          5678 => x"39",
          5679 => x"77",
          5680 => x"81",
          5681 => x"72",
          5682 => x"84",
          5683 => x"73",
          5684 => x"0c",
          5685 => x"04",
          5686 => x"74",
          5687 => x"71",
          5688 => x"2b",
          5689 => x"98",
          5690 => x"84",
          5691 => x"fd",
          5692 => x"83",
          5693 => x"12",
          5694 => x"2b",
          5695 => x"07",
          5696 => x"70",
          5697 => x"2b",
          5698 => x"07",
          5699 => x"0c",
          5700 => x"56",
          5701 => x"3d",
          5702 => x"3d",
          5703 => x"84",
          5704 => x"22",
          5705 => x"72",
          5706 => x"54",
          5707 => x"2a",
          5708 => x"34",
          5709 => x"04",
          5710 => x"73",
          5711 => x"70",
          5712 => x"05",
          5713 => x"88",
          5714 => x"72",
          5715 => x"54",
          5716 => x"2a",
          5717 => x"70",
          5718 => x"34",
          5719 => x"51",
          5720 => x"83",
          5721 => x"fe",
          5722 => x"75",
          5723 => x"51",
          5724 => x"92",
          5725 => x"81",
          5726 => x"73",
          5727 => x"55",
          5728 => x"51",
          5729 => x"3d",
          5730 => x"3d",
          5731 => x"76",
          5732 => x"72",
          5733 => x"05",
          5734 => x"11",
          5735 => x"38",
          5736 => x"04",
          5737 => x"78",
          5738 => x"56",
          5739 => x"81",
          5740 => x"74",
          5741 => x"56",
          5742 => x"31",
          5743 => x"52",
          5744 => x"80",
          5745 => x"71",
          5746 => x"38",
          5747 => x"98",
          5748 => x"0d",
          5749 => x"0d",
          5750 => x"51",
          5751 => x"73",
          5752 => x"81",
          5753 => x"33",
          5754 => x"38",
          5755 => x"bb",
          5756 => x"3d",
          5757 => x"0b",
          5758 => x"0c",
          5759 => x"82",
          5760 => x"04",
          5761 => x"7b",
          5762 => x"83",
          5763 => x"5a",
          5764 => x"80",
          5765 => x"54",
          5766 => x"53",
          5767 => x"53",
          5768 => x"52",
          5769 => x"3f",
          5770 => x"08",
          5771 => x"81",
          5772 => x"82",
          5773 => x"83",
          5774 => x"16",
          5775 => x"18",
          5776 => x"18",
          5777 => x"58",
          5778 => x"9f",
          5779 => x"33",
          5780 => x"2e",
          5781 => x"93",
          5782 => x"76",
          5783 => x"52",
          5784 => x"51",
          5785 => x"83",
          5786 => x"79",
          5787 => x"0c",
          5788 => x"04",
          5789 => x"78",
          5790 => x"80",
          5791 => x"17",
          5792 => x"38",
          5793 => x"fc",
          5794 => x"98",
          5795 => x"bb",
          5796 => x"38",
          5797 => x"53",
          5798 => x"81",
          5799 => x"f7",
          5800 => x"bb",
          5801 => x"2e",
          5802 => x"55",
          5803 => x"b0",
          5804 => x"82",
          5805 => x"88",
          5806 => x"f8",
          5807 => x"70",
          5808 => x"c0",
          5809 => x"98",
          5810 => x"bb",
          5811 => x"91",
          5812 => x"55",
          5813 => x"09",
          5814 => x"f0",
          5815 => x"33",
          5816 => x"2e",
          5817 => x"80",
          5818 => x"80",
          5819 => x"98",
          5820 => x"17",
          5821 => x"fd",
          5822 => x"d4",
          5823 => x"b2",
          5824 => x"96",
          5825 => x"85",
          5826 => x"75",
          5827 => x"3f",
          5828 => x"e4",
          5829 => x"98",
          5830 => x"9c",
          5831 => x"08",
          5832 => x"17",
          5833 => x"3f",
          5834 => x"52",
          5835 => x"51",
          5836 => x"a0",
          5837 => x"05",
          5838 => x"0c",
          5839 => x"75",
          5840 => x"33",
          5841 => x"3f",
          5842 => x"34",
          5843 => x"52",
          5844 => x"51",
          5845 => x"82",
          5846 => x"80",
          5847 => x"81",
          5848 => x"bb",
          5849 => x"3d",
          5850 => x"3d",
          5851 => x"1a",
          5852 => x"fe",
          5853 => x"54",
          5854 => x"73",
          5855 => x"8a",
          5856 => x"71",
          5857 => x"08",
          5858 => x"75",
          5859 => x"0c",
          5860 => x"04",
          5861 => x"7a",
          5862 => x"56",
          5863 => x"77",
          5864 => x"38",
          5865 => x"08",
          5866 => x"38",
          5867 => x"54",
          5868 => x"2e",
          5869 => x"72",
          5870 => x"38",
          5871 => x"8d",
          5872 => x"39",
          5873 => x"81",
          5874 => x"b6",
          5875 => x"2a",
          5876 => x"2a",
          5877 => x"05",
          5878 => x"55",
          5879 => x"82",
          5880 => x"81",
          5881 => x"83",
          5882 => x"b4",
          5883 => x"17",
          5884 => x"a4",
          5885 => x"55",
          5886 => x"57",
          5887 => x"3f",
          5888 => x"08",
          5889 => x"74",
          5890 => x"14",
          5891 => x"70",
          5892 => x"07",
          5893 => x"71",
          5894 => x"52",
          5895 => x"72",
          5896 => x"75",
          5897 => x"58",
          5898 => x"76",
          5899 => x"15",
          5900 => x"73",
          5901 => x"3f",
          5902 => x"08",
          5903 => x"76",
          5904 => x"06",
          5905 => x"05",
          5906 => x"3f",
          5907 => x"08",
          5908 => x"06",
          5909 => x"76",
          5910 => x"15",
          5911 => x"73",
          5912 => x"3f",
          5913 => x"08",
          5914 => x"82",
          5915 => x"06",
          5916 => x"05",
          5917 => x"3f",
          5918 => x"08",
          5919 => x"58",
          5920 => x"58",
          5921 => x"98",
          5922 => x"0d",
          5923 => x"0d",
          5924 => x"5a",
          5925 => x"59",
          5926 => x"82",
          5927 => x"98",
          5928 => x"82",
          5929 => x"33",
          5930 => x"2e",
          5931 => x"72",
          5932 => x"38",
          5933 => x"8d",
          5934 => x"39",
          5935 => x"81",
          5936 => x"f7",
          5937 => x"2a",
          5938 => x"2a",
          5939 => x"05",
          5940 => x"55",
          5941 => x"82",
          5942 => x"59",
          5943 => x"08",
          5944 => x"74",
          5945 => x"16",
          5946 => x"16",
          5947 => x"59",
          5948 => x"53",
          5949 => x"8f",
          5950 => x"2b",
          5951 => x"74",
          5952 => x"71",
          5953 => x"72",
          5954 => x"0b",
          5955 => x"74",
          5956 => x"17",
          5957 => x"75",
          5958 => x"3f",
          5959 => x"08",
          5960 => x"98",
          5961 => x"38",
          5962 => x"06",
          5963 => x"78",
          5964 => x"54",
          5965 => x"77",
          5966 => x"33",
          5967 => x"71",
          5968 => x"51",
          5969 => x"34",
          5970 => x"76",
          5971 => x"17",
          5972 => x"75",
          5973 => x"3f",
          5974 => x"08",
          5975 => x"98",
          5976 => x"38",
          5977 => x"ff",
          5978 => x"10",
          5979 => x"76",
          5980 => x"51",
          5981 => x"be",
          5982 => x"2a",
          5983 => x"05",
          5984 => x"f9",
          5985 => x"bb",
          5986 => x"82",
          5987 => x"ab",
          5988 => x"0a",
          5989 => x"2b",
          5990 => x"70",
          5991 => x"70",
          5992 => x"54",
          5993 => x"82",
          5994 => x"8f",
          5995 => x"07",
          5996 => x"f7",
          5997 => x"0b",
          5998 => x"78",
          5999 => x"0c",
          6000 => x"04",
          6001 => x"7a",
          6002 => x"08",
          6003 => x"59",
          6004 => x"a4",
          6005 => x"17",
          6006 => x"38",
          6007 => x"aa",
          6008 => x"73",
          6009 => x"fd",
          6010 => x"bb",
          6011 => x"82",
          6012 => x"80",
          6013 => x"39",
          6014 => x"eb",
          6015 => x"80",
          6016 => x"bb",
          6017 => x"80",
          6018 => x"52",
          6019 => x"84",
          6020 => x"98",
          6021 => x"bb",
          6022 => x"2e",
          6023 => x"82",
          6024 => x"81",
          6025 => x"82",
          6026 => x"ff",
          6027 => x"80",
          6028 => x"75",
          6029 => x"3f",
          6030 => x"08",
          6031 => x"16",
          6032 => x"90",
          6033 => x"55",
          6034 => x"27",
          6035 => x"15",
          6036 => x"84",
          6037 => x"07",
          6038 => x"17",
          6039 => x"76",
          6040 => x"a6",
          6041 => x"73",
          6042 => x"0c",
          6043 => x"04",
          6044 => x"7c",
          6045 => x"59",
          6046 => x"95",
          6047 => x"08",
          6048 => x"2e",
          6049 => x"17",
          6050 => x"b2",
          6051 => x"ae",
          6052 => x"7a",
          6053 => x"3f",
          6054 => x"82",
          6055 => x"27",
          6056 => x"82",
          6057 => x"55",
          6058 => x"08",
          6059 => x"d2",
          6060 => x"08",
          6061 => x"08",
          6062 => x"38",
          6063 => x"17",
          6064 => x"54",
          6065 => x"82",
          6066 => x"7a",
          6067 => x"06",
          6068 => x"81",
          6069 => x"17",
          6070 => x"83",
          6071 => x"75",
          6072 => x"f9",
          6073 => x"59",
          6074 => x"08",
          6075 => x"81",
          6076 => x"82",
          6077 => x"59",
          6078 => x"08",
          6079 => x"70",
          6080 => x"25",
          6081 => x"82",
          6082 => x"54",
          6083 => x"55",
          6084 => x"38",
          6085 => x"08",
          6086 => x"38",
          6087 => x"54",
          6088 => x"90",
          6089 => x"18",
          6090 => x"38",
          6091 => x"39",
          6092 => x"38",
          6093 => x"16",
          6094 => x"08",
          6095 => x"38",
          6096 => x"78",
          6097 => x"38",
          6098 => x"51",
          6099 => x"82",
          6100 => x"80",
          6101 => x"80",
          6102 => x"98",
          6103 => x"09",
          6104 => x"38",
          6105 => x"08",
          6106 => x"98",
          6107 => x"30",
          6108 => x"80",
          6109 => x"07",
          6110 => x"55",
          6111 => x"38",
          6112 => x"09",
          6113 => x"ae",
          6114 => x"80",
          6115 => x"53",
          6116 => x"51",
          6117 => x"82",
          6118 => x"82",
          6119 => x"30",
          6120 => x"98",
          6121 => x"25",
          6122 => x"79",
          6123 => x"38",
          6124 => x"8f",
          6125 => x"79",
          6126 => x"f9",
          6127 => x"bb",
          6128 => x"74",
          6129 => x"8c",
          6130 => x"17",
          6131 => x"90",
          6132 => x"54",
          6133 => x"86",
          6134 => x"90",
          6135 => x"17",
          6136 => x"54",
          6137 => x"34",
          6138 => x"56",
          6139 => x"90",
          6140 => x"80",
          6141 => x"82",
          6142 => x"55",
          6143 => x"56",
          6144 => x"82",
          6145 => x"8c",
          6146 => x"f8",
          6147 => x"70",
          6148 => x"f0",
          6149 => x"98",
          6150 => x"56",
          6151 => x"08",
          6152 => x"7b",
          6153 => x"f6",
          6154 => x"bb",
          6155 => x"bb",
          6156 => x"17",
          6157 => x"80",
          6158 => x"b4",
          6159 => x"57",
          6160 => x"77",
          6161 => x"81",
          6162 => x"15",
          6163 => x"78",
          6164 => x"81",
          6165 => x"53",
          6166 => x"15",
          6167 => x"e9",
          6168 => x"98",
          6169 => x"df",
          6170 => x"22",
          6171 => x"30",
          6172 => x"70",
          6173 => x"51",
          6174 => x"82",
          6175 => x"8a",
          6176 => x"f8",
          6177 => x"7c",
          6178 => x"56",
          6179 => x"80",
          6180 => x"f1",
          6181 => x"06",
          6182 => x"e9",
          6183 => x"18",
          6184 => x"08",
          6185 => x"38",
          6186 => x"82",
          6187 => x"38",
          6188 => x"54",
          6189 => x"74",
          6190 => x"82",
          6191 => x"22",
          6192 => x"79",
          6193 => x"38",
          6194 => x"98",
          6195 => x"cd",
          6196 => x"22",
          6197 => x"54",
          6198 => x"26",
          6199 => x"52",
          6200 => x"b0",
          6201 => x"98",
          6202 => x"bb",
          6203 => x"2e",
          6204 => x"0b",
          6205 => x"08",
          6206 => x"98",
          6207 => x"bb",
          6208 => x"85",
          6209 => x"bd",
          6210 => x"31",
          6211 => x"73",
          6212 => x"f4",
          6213 => x"bb",
          6214 => x"18",
          6215 => x"18",
          6216 => x"08",
          6217 => x"72",
          6218 => x"38",
          6219 => x"58",
          6220 => x"89",
          6221 => x"18",
          6222 => x"ff",
          6223 => x"05",
          6224 => x"80",
          6225 => x"bb",
          6226 => x"3d",
          6227 => x"3d",
          6228 => x"08",
          6229 => x"a0",
          6230 => x"54",
          6231 => x"77",
          6232 => x"80",
          6233 => x"0c",
          6234 => x"53",
          6235 => x"80",
          6236 => x"38",
          6237 => x"06",
          6238 => x"b5",
          6239 => x"98",
          6240 => x"14",
          6241 => x"92",
          6242 => x"2a",
          6243 => x"56",
          6244 => x"26",
          6245 => x"80",
          6246 => x"16",
          6247 => x"77",
          6248 => x"53",
          6249 => x"38",
          6250 => x"51",
          6251 => x"82",
          6252 => x"53",
          6253 => x"0b",
          6254 => x"08",
          6255 => x"38",
          6256 => x"bb",
          6257 => x"2e",
          6258 => x"98",
          6259 => x"bb",
          6260 => x"80",
          6261 => x"8a",
          6262 => x"15",
          6263 => x"80",
          6264 => x"14",
          6265 => x"51",
          6266 => x"82",
          6267 => x"53",
          6268 => x"bb",
          6269 => x"2e",
          6270 => x"82",
          6271 => x"98",
          6272 => x"ba",
          6273 => x"82",
          6274 => x"ff",
          6275 => x"82",
          6276 => x"52",
          6277 => x"f3",
          6278 => x"98",
          6279 => x"72",
          6280 => x"72",
          6281 => x"f2",
          6282 => x"bb",
          6283 => x"15",
          6284 => x"15",
          6285 => x"b4",
          6286 => x"0c",
          6287 => x"82",
          6288 => x"8a",
          6289 => x"f7",
          6290 => x"7d",
          6291 => x"5b",
          6292 => x"76",
          6293 => x"3f",
          6294 => x"08",
          6295 => x"98",
          6296 => x"38",
          6297 => x"08",
          6298 => x"08",
          6299 => x"f0",
          6300 => x"bb",
          6301 => x"82",
          6302 => x"80",
          6303 => x"bb",
          6304 => x"18",
          6305 => x"51",
          6306 => x"81",
          6307 => x"81",
          6308 => x"81",
          6309 => x"98",
          6310 => x"83",
          6311 => x"77",
          6312 => x"72",
          6313 => x"38",
          6314 => x"75",
          6315 => x"81",
          6316 => x"a5",
          6317 => x"98",
          6318 => x"52",
          6319 => x"8e",
          6320 => x"98",
          6321 => x"bb",
          6322 => x"2e",
          6323 => x"73",
          6324 => x"81",
          6325 => x"87",
          6326 => x"bb",
          6327 => x"3d",
          6328 => x"3d",
          6329 => x"11",
          6330 => x"ec",
          6331 => x"98",
          6332 => x"ff",
          6333 => x"33",
          6334 => x"71",
          6335 => x"81",
          6336 => x"94",
          6337 => x"d0",
          6338 => x"98",
          6339 => x"73",
          6340 => x"82",
          6341 => x"85",
          6342 => x"fc",
          6343 => x"79",
          6344 => x"ff",
          6345 => x"12",
          6346 => x"eb",
          6347 => x"70",
          6348 => x"72",
          6349 => x"81",
          6350 => x"73",
          6351 => x"94",
          6352 => x"d6",
          6353 => x"0d",
          6354 => x"0d",
          6355 => x"55",
          6356 => x"5a",
          6357 => x"08",
          6358 => x"8a",
          6359 => x"08",
          6360 => x"ee",
          6361 => x"bb",
          6362 => x"82",
          6363 => x"80",
          6364 => x"15",
          6365 => x"55",
          6366 => x"38",
          6367 => x"e6",
          6368 => x"33",
          6369 => x"70",
          6370 => x"58",
          6371 => x"86",
          6372 => x"bb",
          6373 => x"73",
          6374 => x"83",
          6375 => x"73",
          6376 => x"38",
          6377 => x"06",
          6378 => x"80",
          6379 => x"75",
          6380 => x"38",
          6381 => x"08",
          6382 => x"54",
          6383 => x"2e",
          6384 => x"83",
          6385 => x"73",
          6386 => x"38",
          6387 => x"51",
          6388 => x"82",
          6389 => x"58",
          6390 => x"08",
          6391 => x"15",
          6392 => x"38",
          6393 => x"0b",
          6394 => x"77",
          6395 => x"0c",
          6396 => x"04",
          6397 => x"77",
          6398 => x"54",
          6399 => x"51",
          6400 => x"82",
          6401 => x"55",
          6402 => x"08",
          6403 => x"14",
          6404 => x"51",
          6405 => x"82",
          6406 => x"55",
          6407 => x"08",
          6408 => x"53",
          6409 => x"08",
          6410 => x"08",
          6411 => x"3f",
          6412 => x"14",
          6413 => x"08",
          6414 => x"3f",
          6415 => x"17",
          6416 => x"bb",
          6417 => x"3d",
          6418 => x"3d",
          6419 => x"08",
          6420 => x"54",
          6421 => x"53",
          6422 => x"82",
          6423 => x"8d",
          6424 => x"08",
          6425 => x"34",
          6426 => x"15",
          6427 => x"0d",
          6428 => x"0d",
          6429 => x"57",
          6430 => x"17",
          6431 => x"08",
          6432 => x"82",
          6433 => x"89",
          6434 => x"55",
          6435 => x"14",
          6436 => x"16",
          6437 => x"71",
          6438 => x"38",
          6439 => x"09",
          6440 => x"38",
          6441 => x"73",
          6442 => x"81",
          6443 => x"ae",
          6444 => x"05",
          6445 => x"15",
          6446 => x"70",
          6447 => x"34",
          6448 => x"8a",
          6449 => x"38",
          6450 => x"05",
          6451 => x"81",
          6452 => x"17",
          6453 => x"12",
          6454 => x"34",
          6455 => x"9c",
          6456 => x"e8",
          6457 => x"bb",
          6458 => x"0c",
          6459 => x"e7",
          6460 => x"bb",
          6461 => x"17",
          6462 => x"51",
          6463 => x"82",
          6464 => x"84",
          6465 => x"3d",
          6466 => x"3d",
          6467 => x"08",
          6468 => x"61",
          6469 => x"55",
          6470 => x"2e",
          6471 => x"55",
          6472 => x"2e",
          6473 => x"80",
          6474 => x"94",
          6475 => x"1c",
          6476 => x"81",
          6477 => x"61",
          6478 => x"56",
          6479 => x"2e",
          6480 => x"83",
          6481 => x"73",
          6482 => x"70",
          6483 => x"25",
          6484 => x"51",
          6485 => x"38",
          6486 => x"0c",
          6487 => x"51",
          6488 => x"26",
          6489 => x"80",
          6490 => x"34",
          6491 => x"51",
          6492 => x"82",
          6493 => x"55",
          6494 => x"91",
          6495 => x"1d",
          6496 => x"8b",
          6497 => x"79",
          6498 => x"3f",
          6499 => x"57",
          6500 => x"55",
          6501 => x"2e",
          6502 => x"80",
          6503 => x"18",
          6504 => x"1a",
          6505 => x"70",
          6506 => x"2a",
          6507 => x"07",
          6508 => x"5a",
          6509 => x"8c",
          6510 => x"54",
          6511 => x"81",
          6512 => x"39",
          6513 => x"70",
          6514 => x"2a",
          6515 => x"75",
          6516 => x"8c",
          6517 => x"2e",
          6518 => x"a0",
          6519 => x"38",
          6520 => x"0c",
          6521 => x"76",
          6522 => x"38",
          6523 => x"b8",
          6524 => x"70",
          6525 => x"5a",
          6526 => x"76",
          6527 => x"38",
          6528 => x"70",
          6529 => x"dc",
          6530 => x"72",
          6531 => x"80",
          6532 => x"51",
          6533 => x"73",
          6534 => x"38",
          6535 => x"18",
          6536 => x"1a",
          6537 => x"55",
          6538 => x"2e",
          6539 => x"83",
          6540 => x"73",
          6541 => x"70",
          6542 => x"25",
          6543 => x"51",
          6544 => x"38",
          6545 => x"75",
          6546 => x"81",
          6547 => x"81",
          6548 => x"27",
          6549 => x"73",
          6550 => x"38",
          6551 => x"70",
          6552 => x"32",
          6553 => x"80",
          6554 => x"2a",
          6555 => x"56",
          6556 => x"81",
          6557 => x"57",
          6558 => x"f5",
          6559 => x"2b",
          6560 => x"25",
          6561 => x"80",
          6562 => x"b4",
          6563 => x"57",
          6564 => x"e6",
          6565 => x"bb",
          6566 => x"2e",
          6567 => x"18",
          6568 => x"1a",
          6569 => x"56",
          6570 => x"3f",
          6571 => x"08",
          6572 => x"e8",
          6573 => x"54",
          6574 => x"80",
          6575 => x"17",
          6576 => x"34",
          6577 => x"11",
          6578 => x"74",
          6579 => x"75",
          6580 => x"80",
          6581 => x"3f",
          6582 => x"08",
          6583 => x"9f",
          6584 => x"99",
          6585 => x"e0",
          6586 => x"ff",
          6587 => x"79",
          6588 => x"74",
          6589 => x"57",
          6590 => x"77",
          6591 => x"76",
          6592 => x"38",
          6593 => x"73",
          6594 => x"09",
          6595 => x"38",
          6596 => x"84",
          6597 => x"27",
          6598 => x"39",
          6599 => x"f2",
          6600 => x"80",
          6601 => x"54",
          6602 => x"34",
          6603 => x"58",
          6604 => x"f2",
          6605 => x"bb",
          6606 => x"82",
          6607 => x"80",
          6608 => x"1b",
          6609 => x"51",
          6610 => x"82",
          6611 => x"56",
          6612 => x"08",
          6613 => x"9c",
          6614 => x"33",
          6615 => x"80",
          6616 => x"38",
          6617 => x"bf",
          6618 => x"86",
          6619 => x"15",
          6620 => x"2a",
          6621 => x"51",
          6622 => x"92",
          6623 => x"79",
          6624 => x"e4",
          6625 => x"bb",
          6626 => x"2e",
          6627 => x"52",
          6628 => x"ba",
          6629 => x"39",
          6630 => x"33",
          6631 => x"80",
          6632 => x"74",
          6633 => x"81",
          6634 => x"38",
          6635 => x"70",
          6636 => x"82",
          6637 => x"54",
          6638 => x"96",
          6639 => x"06",
          6640 => x"2e",
          6641 => x"ff",
          6642 => x"1c",
          6643 => x"80",
          6644 => x"81",
          6645 => x"ba",
          6646 => x"b6",
          6647 => x"2a",
          6648 => x"51",
          6649 => x"38",
          6650 => x"70",
          6651 => x"81",
          6652 => x"55",
          6653 => x"e1",
          6654 => x"08",
          6655 => x"1d",
          6656 => x"7c",
          6657 => x"3f",
          6658 => x"08",
          6659 => x"fa",
          6660 => x"82",
          6661 => x"8f",
          6662 => x"f6",
          6663 => x"5b",
          6664 => x"70",
          6665 => x"59",
          6666 => x"73",
          6667 => x"c6",
          6668 => x"81",
          6669 => x"70",
          6670 => x"52",
          6671 => x"8d",
          6672 => x"38",
          6673 => x"09",
          6674 => x"a5",
          6675 => x"d0",
          6676 => x"ff",
          6677 => x"53",
          6678 => x"91",
          6679 => x"73",
          6680 => x"d0",
          6681 => x"71",
          6682 => x"f7",
          6683 => x"82",
          6684 => x"55",
          6685 => x"55",
          6686 => x"81",
          6687 => x"74",
          6688 => x"56",
          6689 => x"12",
          6690 => x"70",
          6691 => x"38",
          6692 => x"81",
          6693 => x"51",
          6694 => x"51",
          6695 => x"89",
          6696 => x"70",
          6697 => x"53",
          6698 => x"70",
          6699 => x"51",
          6700 => x"09",
          6701 => x"38",
          6702 => x"38",
          6703 => x"77",
          6704 => x"70",
          6705 => x"2a",
          6706 => x"07",
          6707 => x"51",
          6708 => x"8f",
          6709 => x"84",
          6710 => x"83",
          6711 => x"94",
          6712 => x"74",
          6713 => x"38",
          6714 => x"0c",
          6715 => x"86",
          6716 => x"e4",
          6717 => x"82",
          6718 => x"8c",
          6719 => x"fa",
          6720 => x"56",
          6721 => x"17",
          6722 => x"b0",
          6723 => x"52",
          6724 => x"e0",
          6725 => x"82",
          6726 => x"81",
          6727 => x"b2",
          6728 => x"b4",
          6729 => x"98",
          6730 => x"ff",
          6731 => x"55",
          6732 => x"d5",
          6733 => x"06",
          6734 => x"80",
          6735 => x"33",
          6736 => x"81",
          6737 => x"81",
          6738 => x"81",
          6739 => x"eb",
          6740 => x"70",
          6741 => x"07",
          6742 => x"73",
          6743 => x"81",
          6744 => x"81",
          6745 => x"83",
          6746 => x"90",
          6747 => x"16",
          6748 => x"3f",
          6749 => x"08",
          6750 => x"98",
          6751 => x"9d",
          6752 => x"82",
          6753 => x"81",
          6754 => x"e0",
          6755 => x"bb",
          6756 => x"82",
          6757 => x"80",
          6758 => x"82",
          6759 => x"bb",
          6760 => x"3d",
          6761 => x"3d",
          6762 => x"84",
          6763 => x"05",
          6764 => x"80",
          6765 => x"51",
          6766 => x"82",
          6767 => x"58",
          6768 => x"0b",
          6769 => x"08",
          6770 => x"38",
          6771 => x"08",
          6772 => x"d2",
          6773 => x"08",
          6774 => x"56",
          6775 => x"86",
          6776 => x"75",
          6777 => x"fe",
          6778 => x"54",
          6779 => x"2e",
          6780 => x"14",
          6781 => x"ca",
          6782 => x"98",
          6783 => x"06",
          6784 => x"54",
          6785 => x"38",
          6786 => x"86",
          6787 => x"82",
          6788 => x"06",
          6789 => x"56",
          6790 => x"38",
          6791 => x"80",
          6792 => x"81",
          6793 => x"52",
          6794 => x"51",
          6795 => x"82",
          6796 => x"81",
          6797 => x"81",
          6798 => x"83",
          6799 => x"87",
          6800 => x"2e",
          6801 => x"82",
          6802 => x"06",
          6803 => x"56",
          6804 => x"38",
          6805 => x"74",
          6806 => x"a3",
          6807 => x"98",
          6808 => x"06",
          6809 => x"2e",
          6810 => x"80",
          6811 => x"3d",
          6812 => x"83",
          6813 => x"15",
          6814 => x"53",
          6815 => x"8d",
          6816 => x"15",
          6817 => x"3f",
          6818 => x"08",
          6819 => x"70",
          6820 => x"0c",
          6821 => x"16",
          6822 => x"80",
          6823 => x"80",
          6824 => x"54",
          6825 => x"84",
          6826 => x"5b",
          6827 => x"80",
          6828 => x"7a",
          6829 => x"fc",
          6830 => x"bb",
          6831 => x"ff",
          6832 => x"77",
          6833 => x"81",
          6834 => x"76",
          6835 => x"81",
          6836 => x"2e",
          6837 => x"8d",
          6838 => x"26",
          6839 => x"bf",
          6840 => x"f4",
          6841 => x"98",
          6842 => x"ff",
          6843 => x"84",
          6844 => x"81",
          6845 => x"38",
          6846 => x"51",
          6847 => x"82",
          6848 => x"83",
          6849 => x"58",
          6850 => x"80",
          6851 => x"db",
          6852 => x"bb",
          6853 => x"77",
          6854 => x"80",
          6855 => x"82",
          6856 => x"c4",
          6857 => x"11",
          6858 => x"06",
          6859 => x"8d",
          6860 => x"26",
          6861 => x"74",
          6862 => x"78",
          6863 => x"c1",
          6864 => x"59",
          6865 => x"15",
          6866 => x"2e",
          6867 => x"13",
          6868 => x"72",
          6869 => x"38",
          6870 => x"eb",
          6871 => x"14",
          6872 => x"3f",
          6873 => x"08",
          6874 => x"98",
          6875 => x"23",
          6876 => x"57",
          6877 => x"83",
          6878 => x"c7",
          6879 => x"d8",
          6880 => x"98",
          6881 => x"ff",
          6882 => x"8d",
          6883 => x"14",
          6884 => x"3f",
          6885 => x"08",
          6886 => x"14",
          6887 => x"3f",
          6888 => x"08",
          6889 => x"06",
          6890 => x"72",
          6891 => x"97",
          6892 => x"22",
          6893 => x"84",
          6894 => x"5a",
          6895 => x"83",
          6896 => x"14",
          6897 => x"79",
          6898 => x"fa",
          6899 => x"bb",
          6900 => x"82",
          6901 => x"80",
          6902 => x"38",
          6903 => x"08",
          6904 => x"ff",
          6905 => x"38",
          6906 => x"83",
          6907 => x"83",
          6908 => x"74",
          6909 => x"85",
          6910 => x"89",
          6911 => x"76",
          6912 => x"c3",
          6913 => x"70",
          6914 => x"7b",
          6915 => x"73",
          6916 => x"17",
          6917 => x"ac",
          6918 => x"55",
          6919 => x"09",
          6920 => x"38",
          6921 => x"51",
          6922 => x"82",
          6923 => x"83",
          6924 => x"53",
          6925 => x"82",
          6926 => x"82",
          6927 => x"e0",
          6928 => x"ab",
          6929 => x"98",
          6930 => x"0c",
          6931 => x"53",
          6932 => x"56",
          6933 => x"81",
          6934 => x"13",
          6935 => x"74",
          6936 => x"82",
          6937 => x"74",
          6938 => x"81",
          6939 => x"06",
          6940 => x"83",
          6941 => x"2a",
          6942 => x"72",
          6943 => x"26",
          6944 => x"ff",
          6945 => x"0c",
          6946 => x"15",
          6947 => x"0b",
          6948 => x"76",
          6949 => x"81",
          6950 => x"38",
          6951 => x"51",
          6952 => x"82",
          6953 => x"83",
          6954 => x"53",
          6955 => x"09",
          6956 => x"f9",
          6957 => x"52",
          6958 => x"b8",
          6959 => x"98",
          6960 => x"38",
          6961 => x"08",
          6962 => x"84",
          6963 => x"d8",
          6964 => x"bb",
          6965 => x"ff",
          6966 => x"72",
          6967 => x"2e",
          6968 => x"80",
          6969 => x"14",
          6970 => x"3f",
          6971 => x"08",
          6972 => x"a4",
          6973 => x"81",
          6974 => x"84",
          6975 => x"d7",
          6976 => x"bb",
          6977 => x"8a",
          6978 => x"2e",
          6979 => x"9d",
          6980 => x"14",
          6981 => x"3f",
          6982 => x"08",
          6983 => x"84",
          6984 => x"d7",
          6985 => x"bb",
          6986 => x"15",
          6987 => x"34",
          6988 => x"22",
          6989 => x"72",
          6990 => x"23",
          6991 => x"23",
          6992 => x"15",
          6993 => x"75",
          6994 => x"0c",
          6995 => x"04",
          6996 => x"77",
          6997 => x"73",
          6998 => x"38",
          6999 => x"72",
          7000 => x"38",
          7001 => x"71",
          7002 => x"38",
          7003 => x"84",
          7004 => x"52",
          7005 => x"09",
          7006 => x"38",
          7007 => x"51",
          7008 => x"82",
          7009 => x"81",
          7010 => x"88",
          7011 => x"08",
          7012 => x"39",
          7013 => x"73",
          7014 => x"74",
          7015 => x"0c",
          7016 => x"04",
          7017 => x"02",
          7018 => x"7a",
          7019 => x"fc",
          7020 => x"f4",
          7021 => x"54",
          7022 => x"bb",
          7023 => x"bc",
          7024 => x"98",
          7025 => x"82",
          7026 => x"70",
          7027 => x"73",
          7028 => x"38",
          7029 => x"78",
          7030 => x"2e",
          7031 => x"74",
          7032 => x"0c",
          7033 => x"80",
          7034 => x"80",
          7035 => x"70",
          7036 => x"51",
          7037 => x"82",
          7038 => x"54",
          7039 => x"98",
          7040 => x"0d",
          7041 => x"0d",
          7042 => x"05",
          7043 => x"33",
          7044 => x"54",
          7045 => x"84",
          7046 => x"bf",
          7047 => x"98",
          7048 => x"53",
          7049 => x"05",
          7050 => x"fa",
          7051 => x"98",
          7052 => x"bb",
          7053 => x"a4",
          7054 => x"68",
          7055 => x"70",
          7056 => x"c6",
          7057 => x"98",
          7058 => x"bb",
          7059 => x"38",
          7060 => x"05",
          7061 => x"2b",
          7062 => x"80",
          7063 => x"86",
          7064 => x"06",
          7065 => x"2e",
          7066 => x"74",
          7067 => x"38",
          7068 => x"09",
          7069 => x"38",
          7070 => x"f8",
          7071 => x"98",
          7072 => x"39",
          7073 => x"33",
          7074 => x"73",
          7075 => x"77",
          7076 => x"81",
          7077 => x"73",
          7078 => x"38",
          7079 => x"bc",
          7080 => x"07",
          7081 => x"b4",
          7082 => x"2a",
          7083 => x"51",
          7084 => x"2e",
          7085 => x"62",
          7086 => x"e8",
          7087 => x"bb",
          7088 => x"82",
          7089 => x"52",
          7090 => x"51",
          7091 => x"62",
          7092 => x"8b",
          7093 => x"53",
          7094 => x"51",
          7095 => x"80",
          7096 => x"05",
          7097 => x"3f",
          7098 => x"0b",
          7099 => x"75",
          7100 => x"f1",
          7101 => x"11",
          7102 => x"80",
          7103 => x"97",
          7104 => x"51",
          7105 => x"82",
          7106 => x"55",
          7107 => x"08",
          7108 => x"b7",
          7109 => x"c4",
          7110 => x"05",
          7111 => x"2a",
          7112 => x"51",
          7113 => x"80",
          7114 => x"84",
          7115 => x"39",
          7116 => x"70",
          7117 => x"54",
          7118 => x"a9",
          7119 => x"06",
          7120 => x"2e",
          7121 => x"55",
          7122 => x"73",
          7123 => x"d6",
          7124 => x"bb",
          7125 => x"ff",
          7126 => x"0c",
          7127 => x"bb",
          7128 => x"f8",
          7129 => x"2a",
          7130 => x"51",
          7131 => x"2e",
          7132 => x"80",
          7133 => x"7a",
          7134 => x"a0",
          7135 => x"a4",
          7136 => x"53",
          7137 => x"e6",
          7138 => x"bb",
          7139 => x"bb",
          7140 => x"1b",
          7141 => x"05",
          7142 => x"d3",
          7143 => x"98",
          7144 => x"98",
          7145 => x"0c",
          7146 => x"56",
          7147 => x"84",
          7148 => x"90",
          7149 => x"0b",
          7150 => x"80",
          7151 => x"0c",
          7152 => x"1a",
          7153 => x"2a",
          7154 => x"51",
          7155 => x"2e",
          7156 => x"82",
          7157 => x"80",
          7158 => x"38",
          7159 => x"08",
          7160 => x"8a",
          7161 => x"89",
          7162 => x"59",
          7163 => x"76",
          7164 => x"d7",
          7165 => x"bb",
          7166 => x"82",
          7167 => x"81",
          7168 => x"82",
          7169 => x"98",
          7170 => x"09",
          7171 => x"38",
          7172 => x"78",
          7173 => x"30",
          7174 => x"80",
          7175 => x"77",
          7176 => x"38",
          7177 => x"06",
          7178 => x"c3",
          7179 => x"1a",
          7180 => x"38",
          7181 => x"06",
          7182 => x"2e",
          7183 => x"52",
          7184 => x"a6",
          7185 => x"98",
          7186 => x"82",
          7187 => x"75",
          7188 => x"bb",
          7189 => x"9c",
          7190 => x"39",
          7191 => x"74",
          7192 => x"bb",
          7193 => x"3d",
          7194 => x"3d",
          7195 => x"65",
          7196 => x"5d",
          7197 => x"0c",
          7198 => x"05",
          7199 => x"f9",
          7200 => x"bb",
          7201 => x"82",
          7202 => x"8a",
          7203 => x"33",
          7204 => x"2e",
          7205 => x"56",
          7206 => x"90",
          7207 => x"06",
          7208 => x"74",
          7209 => x"b6",
          7210 => x"82",
          7211 => x"34",
          7212 => x"aa",
          7213 => x"91",
          7214 => x"56",
          7215 => x"8c",
          7216 => x"1a",
          7217 => x"74",
          7218 => x"38",
          7219 => x"80",
          7220 => x"38",
          7221 => x"70",
          7222 => x"56",
          7223 => x"b2",
          7224 => x"11",
          7225 => x"77",
          7226 => x"5b",
          7227 => x"38",
          7228 => x"88",
          7229 => x"8f",
          7230 => x"08",
          7231 => x"d5",
          7232 => x"bb",
          7233 => x"81",
          7234 => x"9f",
          7235 => x"2e",
          7236 => x"74",
          7237 => x"98",
          7238 => x"7e",
          7239 => x"3f",
          7240 => x"08",
          7241 => x"83",
          7242 => x"98",
          7243 => x"89",
          7244 => x"77",
          7245 => x"d6",
          7246 => x"7f",
          7247 => x"58",
          7248 => x"75",
          7249 => x"75",
          7250 => x"77",
          7251 => x"7c",
          7252 => x"33",
          7253 => x"3f",
          7254 => x"08",
          7255 => x"7e",
          7256 => x"56",
          7257 => x"2e",
          7258 => x"16",
          7259 => x"55",
          7260 => x"94",
          7261 => x"53",
          7262 => x"b0",
          7263 => x"31",
          7264 => x"05",
          7265 => x"3f",
          7266 => x"56",
          7267 => x"9c",
          7268 => x"19",
          7269 => x"06",
          7270 => x"31",
          7271 => x"76",
          7272 => x"7b",
          7273 => x"08",
          7274 => x"d1",
          7275 => x"bb",
          7276 => x"81",
          7277 => x"94",
          7278 => x"ff",
          7279 => x"05",
          7280 => x"cf",
          7281 => x"76",
          7282 => x"17",
          7283 => x"1e",
          7284 => x"18",
          7285 => x"5e",
          7286 => x"39",
          7287 => x"82",
          7288 => x"90",
          7289 => x"f2",
          7290 => x"63",
          7291 => x"40",
          7292 => x"7e",
          7293 => x"fc",
          7294 => x"51",
          7295 => x"82",
          7296 => x"55",
          7297 => x"08",
          7298 => x"18",
          7299 => x"80",
          7300 => x"74",
          7301 => x"39",
          7302 => x"70",
          7303 => x"81",
          7304 => x"56",
          7305 => x"80",
          7306 => x"38",
          7307 => x"0b",
          7308 => x"82",
          7309 => x"39",
          7310 => x"19",
          7311 => x"83",
          7312 => x"18",
          7313 => x"56",
          7314 => x"27",
          7315 => x"09",
          7316 => x"2e",
          7317 => x"94",
          7318 => x"83",
          7319 => x"56",
          7320 => x"38",
          7321 => x"22",
          7322 => x"89",
          7323 => x"55",
          7324 => x"75",
          7325 => x"18",
          7326 => x"9c",
          7327 => x"85",
          7328 => x"08",
          7329 => x"d7",
          7330 => x"bb",
          7331 => x"82",
          7332 => x"80",
          7333 => x"38",
          7334 => x"ff",
          7335 => x"ff",
          7336 => x"38",
          7337 => x"0c",
          7338 => x"85",
          7339 => x"19",
          7340 => x"b0",
          7341 => x"19",
          7342 => x"81",
          7343 => x"74",
          7344 => x"3f",
          7345 => x"08",
          7346 => x"98",
          7347 => x"7e",
          7348 => x"3f",
          7349 => x"08",
          7350 => x"d2",
          7351 => x"98",
          7352 => x"89",
          7353 => x"78",
          7354 => x"d5",
          7355 => x"7f",
          7356 => x"58",
          7357 => x"75",
          7358 => x"75",
          7359 => x"78",
          7360 => x"7c",
          7361 => x"33",
          7362 => x"3f",
          7363 => x"08",
          7364 => x"7e",
          7365 => x"78",
          7366 => x"74",
          7367 => x"38",
          7368 => x"b0",
          7369 => x"31",
          7370 => x"05",
          7371 => x"51",
          7372 => x"7e",
          7373 => x"83",
          7374 => x"89",
          7375 => x"db",
          7376 => x"08",
          7377 => x"26",
          7378 => x"51",
          7379 => x"82",
          7380 => x"fd",
          7381 => x"77",
          7382 => x"55",
          7383 => x"0c",
          7384 => x"83",
          7385 => x"80",
          7386 => x"55",
          7387 => x"83",
          7388 => x"9c",
          7389 => x"7e",
          7390 => x"3f",
          7391 => x"08",
          7392 => x"75",
          7393 => x"94",
          7394 => x"ff",
          7395 => x"05",
          7396 => x"3f",
          7397 => x"0b",
          7398 => x"7b",
          7399 => x"08",
          7400 => x"76",
          7401 => x"08",
          7402 => x"1c",
          7403 => x"08",
          7404 => x"5c",
          7405 => x"83",
          7406 => x"74",
          7407 => x"fd",
          7408 => x"18",
          7409 => x"07",
          7410 => x"19",
          7411 => x"75",
          7412 => x"0c",
          7413 => x"04",
          7414 => x"7a",
          7415 => x"05",
          7416 => x"56",
          7417 => x"82",
          7418 => x"57",
          7419 => x"08",
          7420 => x"90",
          7421 => x"86",
          7422 => x"06",
          7423 => x"73",
          7424 => x"e9",
          7425 => x"08",
          7426 => x"cc",
          7427 => x"bb",
          7428 => x"82",
          7429 => x"80",
          7430 => x"16",
          7431 => x"33",
          7432 => x"55",
          7433 => x"34",
          7434 => x"53",
          7435 => x"08",
          7436 => x"3f",
          7437 => x"52",
          7438 => x"c9",
          7439 => x"88",
          7440 => x"96",
          7441 => x"f0",
          7442 => x"92",
          7443 => x"ca",
          7444 => x"81",
          7445 => x"34",
          7446 => x"df",
          7447 => x"98",
          7448 => x"33",
          7449 => x"55",
          7450 => x"17",
          7451 => x"bb",
          7452 => x"3d",
          7453 => x"3d",
          7454 => x"52",
          7455 => x"3f",
          7456 => x"08",
          7457 => x"98",
          7458 => x"86",
          7459 => x"52",
          7460 => x"bc",
          7461 => x"98",
          7462 => x"bb",
          7463 => x"38",
          7464 => x"08",
          7465 => x"82",
          7466 => x"86",
          7467 => x"ff",
          7468 => x"3d",
          7469 => x"3f",
          7470 => x"0b",
          7471 => x"08",
          7472 => x"82",
          7473 => x"82",
          7474 => x"80",
          7475 => x"bb",
          7476 => x"3d",
          7477 => x"3d",
          7478 => x"93",
          7479 => x"52",
          7480 => x"e9",
          7481 => x"bb",
          7482 => x"82",
          7483 => x"80",
          7484 => x"58",
          7485 => x"3d",
          7486 => x"e0",
          7487 => x"bb",
          7488 => x"82",
          7489 => x"bc",
          7490 => x"c7",
          7491 => x"98",
          7492 => x"73",
          7493 => x"38",
          7494 => x"12",
          7495 => x"39",
          7496 => x"33",
          7497 => x"70",
          7498 => x"55",
          7499 => x"2e",
          7500 => x"7f",
          7501 => x"54",
          7502 => x"82",
          7503 => x"94",
          7504 => x"39",
          7505 => x"08",
          7506 => x"81",
          7507 => x"85",
          7508 => x"bb",
          7509 => x"3d",
          7510 => x"3d",
          7511 => x"5b",
          7512 => x"34",
          7513 => x"3d",
          7514 => x"52",
          7515 => x"e8",
          7516 => x"bb",
          7517 => x"82",
          7518 => x"82",
          7519 => x"43",
          7520 => x"11",
          7521 => x"58",
          7522 => x"80",
          7523 => x"38",
          7524 => x"3d",
          7525 => x"d5",
          7526 => x"bb",
          7527 => x"82",
          7528 => x"82",
          7529 => x"52",
          7530 => x"c8",
          7531 => x"98",
          7532 => x"bb",
          7533 => x"c1",
          7534 => x"7b",
          7535 => x"3f",
          7536 => x"08",
          7537 => x"74",
          7538 => x"3f",
          7539 => x"08",
          7540 => x"98",
          7541 => x"38",
          7542 => x"51",
          7543 => x"82",
          7544 => x"57",
          7545 => x"08",
          7546 => x"52",
          7547 => x"f2",
          7548 => x"bb",
          7549 => x"a6",
          7550 => x"74",
          7551 => x"3f",
          7552 => x"08",
          7553 => x"98",
          7554 => x"cc",
          7555 => x"2e",
          7556 => x"86",
          7557 => x"81",
          7558 => x"81",
          7559 => x"3d",
          7560 => x"52",
          7561 => x"c9",
          7562 => x"3d",
          7563 => x"11",
          7564 => x"5a",
          7565 => x"2e",
          7566 => x"b9",
          7567 => x"16",
          7568 => x"33",
          7569 => x"73",
          7570 => x"16",
          7571 => x"26",
          7572 => x"75",
          7573 => x"38",
          7574 => x"05",
          7575 => x"6f",
          7576 => x"ff",
          7577 => x"55",
          7578 => x"74",
          7579 => x"38",
          7580 => x"11",
          7581 => x"74",
          7582 => x"39",
          7583 => x"09",
          7584 => x"38",
          7585 => x"11",
          7586 => x"74",
          7587 => x"82",
          7588 => x"70",
          7589 => x"b4",
          7590 => x"08",
          7591 => x"5c",
          7592 => x"73",
          7593 => x"38",
          7594 => x"1a",
          7595 => x"55",
          7596 => x"38",
          7597 => x"73",
          7598 => x"38",
          7599 => x"76",
          7600 => x"74",
          7601 => x"33",
          7602 => x"05",
          7603 => x"15",
          7604 => x"ba",
          7605 => x"05",
          7606 => x"ff",
          7607 => x"06",
          7608 => x"57",
          7609 => x"18",
          7610 => x"54",
          7611 => x"70",
          7612 => x"34",
          7613 => x"ee",
          7614 => x"34",
          7615 => x"98",
          7616 => x"0d",
          7617 => x"0d",
          7618 => x"3d",
          7619 => x"71",
          7620 => x"ec",
          7621 => x"bb",
          7622 => x"82",
          7623 => x"82",
          7624 => x"15",
          7625 => x"82",
          7626 => x"15",
          7627 => x"76",
          7628 => x"90",
          7629 => x"81",
          7630 => x"06",
          7631 => x"72",
          7632 => x"56",
          7633 => x"54",
          7634 => x"17",
          7635 => x"78",
          7636 => x"38",
          7637 => x"22",
          7638 => x"59",
          7639 => x"78",
          7640 => x"76",
          7641 => x"51",
          7642 => x"3f",
          7643 => x"08",
          7644 => x"54",
          7645 => x"53",
          7646 => x"3f",
          7647 => x"08",
          7648 => x"38",
          7649 => x"75",
          7650 => x"18",
          7651 => x"31",
          7652 => x"57",
          7653 => x"b1",
          7654 => x"08",
          7655 => x"38",
          7656 => x"51",
          7657 => x"82",
          7658 => x"54",
          7659 => x"08",
          7660 => x"9a",
          7661 => x"98",
          7662 => x"81",
          7663 => x"bb",
          7664 => x"16",
          7665 => x"16",
          7666 => x"2e",
          7667 => x"76",
          7668 => x"dc",
          7669 => x"31",
          7670 => x"18",
          7671 => x"90",
          7672 => x"81",
          7673 => x"06",
          7674 => x"56",
          7675 => x"9a",
          7676 => x"74",
          7677 => x"3f",
          7678 => x"08",
          7679 => x"98",
          7680 => x"82",
          7681 => x"56",
          7682 => x"52",
          7683 => x"84",
          7684 => x"98",
          7685 => x"ff",
          7686 => x"81",
          7687 => x"38",
          7688 => x"98",
          7689 => x"a6",
          7690 => x"16",
          7691 => x"39",
          7692 => x"16",
          7693 => x"75",
          7694 => x"53",
          7695 => x"aa",
          7696 => x"79",
          7697 => x"3f",
          7698 => x"08",
          7699 => x"0b",
          7700 => x"82",
          7701 => x"39",
          7702 => x"16",
          7703 => x"bb",
          7704 => x"2a",
          7705 => x"08",
          7706 => x"15",
          7707 => x"15",
          7708 => x"90",
          7709 => x"16",
          7710 => x"33",
          7711 => x"53",
          7712 => x"34",
          7713 => x"06",
          7714 => x"2e",
          7715 => x"9c",
          7716 => x"85",
          7717 => x"16",
          7718 => x"72",
          7719 => x"0c",
          7720 => x"04",
          7721 => x"79",
          7722 => x"75",
          7723 => x"8a",
          7724 => x"89",
          7725 => x"52",
          7726 => x"05",
          7727 => x"3f",
          7728 => x"08",
          7729 => x"98",
          7730 => x"38",
          7731 => x"7a",
          7732 => x"d8",
          7733 => x"bb",
          7734 => x"82",
          7735 => x"80",
          7736 => x"16",
          7737 => x"2b",
          7738 => x"74",
          7739 => x"86",
          7740 => x"84",
          7741 => x"06",
          7742 => x"73",
          7743 => x"38",
          7744 => x"52",
          7745 => x"da",
          7746 => x"98",
          7747 => x"0c",
          7748 => x"14",
          7749 => x"23",
          7750 => x"51",
          7751 => x"82",
          7752 => x"55",
          7753 => x"09",
          7754 => x"38",
          7755 => x"39",
          7756 => x"84",
          7757 => x"0c",
          7758 => x"82",
          7759 => x"89",
          7760 => x"fc",
          7761 => x"87",
          7762 => x"53",
          7763 => x"e7",
          7764 => x"bb",
          7765 => x"38",
          7766 => x"08",
          7767 => x"3d",
          7768 => x"3d",
          7769 => x"89",
          7770 => x"54",
          7771 => x"54",
          7772 => x"82",
          7773 => x"53",
          7774 => x"08",
          7775 => x"74",
          7776 => x"bb",
          7777 => x"73",
          7778 => x"3f",
          7779 => x"08",
          7780 => x"39",
          7781 => x"08",
          7782 => x"d3",
          7783 => x"bb",
          7784 => x"82",
          7785 => x"84",
          7786 => x"06",
          7787 => x"53",
          7788 => x"bb",
          7789 => x"38",
          7790 => x"51",
          7791 => x"72",
          7792 => x"cf",
          7793 => x"bb",
          7794 => x"32",
          7795 => x"72",
          7796 => x"70",
          7797 => x"08",
          7798 => x"54",
          7799 => x"bb",
          7800 => x"3d",
          7801 => x"3d",
          7802 => x"80",
          7803 => x"70",
          7804 => x"52",
          7805 => x"3f",
          7806 => x"08",
          7807 => x"98",
          7808 => x"64",
          7809 => x"d6",
          7810 => x"bb",
          7811 => x"82",
          7812 => x"a0",
          7813 => x"cb",
          7814 => x"98",
          7815 => x"73",
          7816 => x"38",
          7817 => x"39",
          7818 => x"88",
          7819 => x"75",
          7820 => x"3f",
          7821 => x"98",
          7822 => x"0d",
          7823 => x"0d",
          7824 => x"5c",
          7825 => x"3d",
          7826 => x"93",
          7827 => x"d6",
          7828 => x"98",
          7829 => x"bb",
          7830 => x"80",
          7831 => x"0c",
          7832 => x"11",
          7833 => x"90",
          7834 => x"56",
          7835 => x"74",
          7836 => x"75",
          7837 => x"e4",
          7838 => x"81",
          7839 => x"5b",
          7840 => x"82",
          7841 => x"75",
          7842 => x"73",
          7843 => x"81",
          7844 => x"82",
          7845 => x"76",
          7846 => x"f0",
          7847 => x"f4",
          7848 => x"98",
          7849 => x"d1",
          7850 => x"98",
          7851 => x"ce",
          7852 => x"98",
          7853 => x"82",
          7854 => x"07",
          7855 => x"05",
          7856 => x"53",
          7857 => x"98",
          7858 => x"26",
          7859 => x"f9",
          7860 => x"08",
          7861 => x"08",
          7862 => x"98",
          7863 => x"81",
          7864 => x"58",
          7865 => x"3f",
          7866 => x"08",
          7867 => x"98",
          7868 => x"38",
          7869 => x"77",
          7870 => x"5d",
          7871 => x"74",
          7872 => x"81",
          7873 => x"b4",
          7874 => x"bb",
          7875 => x"bb",
          7876 => x"ff",
          7877 => x"30",
          7878 => x"1b",
          7879 => x"5b",
          7880 => x"39",
          7881 => x"ff",
          7882 => x"82",
          7883 => x"f0",
          7884 => x"30",
          7885 => x"1b",
          7886 => x"5b",
          7887 => x"83",
          7888 => x"58",
          7889 => x"92",
          7890 => x"0c",
          7891 => x"12",
          7892 => x"33",
          7893 => x"54",
          7894 => x"34",
          7895 => x"98",
          7896 => x"0d",
          7897 => x"0d",
          7898 => x"fc",
          7899 => x"52",
          7900 => x"3f",
          7901 => x"08",
          7902 => x"98",
          7903 => x"38",
          7904 => x"56",
          7905 => x"38",
          7906 => x"70",
          7907 => x"81",
          7908 => x"55",
          7909 => x"80",
          7910 => x"38",
          7911 => x"54",
          7912 => x"08",
          7913 => x"38",
          7914 => x"82",
          7915 => x"53",
          7916 => x"52",
          7917 => x"8c",
          7918 => x"98",
          7919 => x"19",
          7920 => x"c9",
          7921 => x"08",
          7922 => x"ff",
          7923 => x"82",
          7924 => x"ff",
          7925 => x"06",
          7926 => x"56",
          7927 => x"08",
          7928 => x"81",
          7929 => x"82",
          7930 => x"75",
          7931 => x"54",
          7932 => x"08",
          7933 => x"27",
          7934 => x"17",
          7935 => x"bb",
          7936 => x"76",
          7937 => x"3f",
          7938 => x"08",
          7939 => x"08",
          7940 => x"90",
          7941 => x"c0",
          7942 => x"90",
          7943 => x"80",
          7944 => x"75",
          7945 => x"75",
          7946 => x"bb",
          7947 => x"3d",
          7948 => x"3d",
          7949 => x"a0",
          7950 => x"05",
          7951 => x"51",
          7952 => x"82",
          7953 => x"55",
          7954 => x"08",
          7955 => x"78",
          7956 => x"08",
          7957 => x"70",
          7958 => x"ae",
          7959 => x"98",
          7960 => x"bb",
          7961 => x"db",
          7962 => x"fb",
          7963 => x"85",
          7964 => x"06",
          7965 => x"86",
          7966 => x"c7",
          7967 => x"2b",
          7968 => x"24",
          7969 => x"02",
          7970 => x"33",
          7971 => x"58",
          7972 => x"76",
          7973 => x"6b",
          7974 => x"cc",
          7975 => x"bb",
          7976 => x"84",
          7977 => x"06",
          7978 => x"73",
          7979 => x"d4",
          7980 => x"82",
          7981 => x"94",
          7982 => x"81",
          7983 => x"5a",
          7984 => x"08",
          7985 => x"8a",
          7986 => x"54",
          7987 => x"82",
          7988 => x"55",
          7989 => x"08",
          7990 => x"82",
          7991 => x"52",
          7992 => x"e5",
          7993 => x"98",
          7994 => x"bb",
          7995 => x"38",
          7996 => x"cf",
          7997 => x"98",
          7998 => x"88",
          7999 => x"98",
          8000 => x"38",
          8001 => x"c2",
          8002 => x"98",
          8003 => x"98",
          8004 => x"82",
          8005 => x"07",
          8006 => x"55",
          8007 => x"2e",
          8008 => x"80",
          8009 => x"80",
          8010 => x"77",
          8011 => x"3f",
          8012 => x"08",
          8013 => x"38",
          8014 => x"ba",
          8015 => x"bb",
          8016 => x"74",
          8017 => x"0c",
          8018 => x"04",
          8019 => x"82",
          8020 => x"c0",
          8021 => x"3d",
          8022 => x"3f",
          8023 => x"08",
          8024 => x"98",
          8025 => x"38",
          8026 => x"52",
          8027 => x"52",
          8028 => x"3f",
          8029 => x"08",
          8030 => x"98",
          8031 => x"88",
          8032 => x"39",
          8033 => x"08",
          8034 => x"81",
          8035 => x"38",
          8036 => x"05",
          8037 => x"2a",
          8038 => x"55",
          8039 => x"81",
          8040 => x"5a",
          8041 => x"3d",
          8042 => x"c1",
          8043 => x"bb",
          8044 => x"55",
          8045 => x"98",
          8046 => x"87",
          8047 => x"98",
          8048 => x"09",
          8049 => x"38",
          8050 => x"bb",
          8051 => x"2e",
          8052 => x"86",
          8053 => x"81",
          8054 => x"81",
          8055 => x"bb",
          8056 => x"78",
          8057 => x"3f",
          8058 => x"08",
          8059 => x"98",
          8060 => x"38",
          8061 => x"52",
          8062 => x"ff",
          8063 => x"78",
          8064 => x"b4",
          8065 => x"54",
          8066 => x"15",
          8067 => x"b2",
          8068 => x"ca",
          8069 => x"b6",
          8070 => x"53",
          8071 => x"53",
          8072 => x"3f",
          8073 => x"b4",
          8074 => x"d4",
          8075 => x"b6",
          8076 => x"54",
          8077 => x"d5",
          8078 => x"53",
          8079 => x"11",
          8080 => x"d7",
          8081 => x"81",
          8082 => x"34",
          8083 => x"a4",
          8084 => x"98",
          8085 => x"bb",
          8086 => x"38",
          8087 => x"0a",
          8088 => x"05",
          8089 => x"d0",
          8090 => x"64",
          8091 => x"c9",
          8092 => x"54",
          8093 => x"15",
          8094 => x"81",
          8095 => x"34",
          8096 => x"b8",
          8097 => x"bb",
          8098 => x"8b",
          8099 => x"75",
          8100 => x"ff",
          8101 => x"73",
          8102 => x"0c",
          8103 => x"04",
          8104 => x"a9",
          8105 => x"51",
          8106 => x"82",
          8107 => x"ff",
          8108 => x"a9",
          8109 => x"ee",
          8110 => x"98",
          8111 => x"bb",
          8112 => x"d3",
          8113 => x"a9",
          8114 => x"9d",
          8115 => x"58",
          8116 => x"82",
          8117 => x"55",
          8118 => x"08",
          8119 => x"02",
          8120 => x"33",
          8121 => x"54",
          8122 => x"82",
          8123 => x"53",
          8124 => x"52",
          8125 => x"88",
          8126 => x"b4",
          8127 => x"53",
          8128 => x"3d",
          8129 => x"ff",
          8130 => x"aa",
          8131 => x"73",
          8132 => x"3f",
          8133 => x"08",
          8134 => x"98",
          8135 => x"63",
          8136 => x"81",
          8137 => x"65",
          8138 => x"2e",
          8139 => x"55",
          8140 => x"82",
          8141 => x"84",
          8142 => x"06",
          8143 => x"73",
          8144 => x"3f",
          8145 => x"08",
          8146 => x"98",
          8147 => x"38",
          8148 => x"53",
          8149 => x"95",
          8150 => x"16",
          8151 => x"87",
          8152 => x"05",
          8153 => x"34",
          8154 => x"70",
          8155 => x"81",
          8156 => x"55",
          8157 => x"74",
          8158 => x"73",
          8159 => x"78",
          8160 => x"83",
          8161 => x"16",
          8162 => x"2a",
          8163 => x"51",
          8164 => x"80",
          8165 => x"38",
          8166 => x"80",
          8167 => x"52",
          8168 => x"be",
          8169 => x"98",
          8170 => x"51",
          8171 => x"3f",
          8172 => x"bb",
          8173 => x"2e",
          8174 => x"82",
          8175 => x"52",
          8176 => x"b5",
          8177 => x"bb",
          8178 => x"80",
          8179 => x"58",
          8180 => x"98",
          8181 => x"38",
          8182 => x"54",
          8183 => x"09",
          8184 => x"38",
          8185 => x"52",
          8186 => x"af",
          8187 => x"81",
          8188 => x"34",
          8189 => x"bb",
          8190 => x"38",
          8191 => x"ca",
          8192 => x"98",
          8193 => x"bb",
          8194 => x"38",
          8195 => x"b5",
          8196 => x"bb",
          8197 => x"74",
          8198 => x"0c",
          8199 => x"04",
          8200 => x"02",
          8201 => x"33",
          8202 => x"80",
          8203 => x"57",
          8204 => x"95",
          8205 => x"52",
          8206 => x"d2",
          8207 => x"bb",
          8208 => x"82",
          8209 => x"80",
          8210 => x"5a",
          8211 => x"3d",
          8212 => x"c9",
          8213 => x"bb",
          8214 => x"82",
          8215 => x"b8",
          8216 => x"cf",
          8217 => x"a0",
          8218 => x"55",
          8219 => x"75",
          8220 => x"71",
          8221 => x"33",
          8222 => x"74",
          8223 => x"57",
          8224 => x"8b",
          8225 => x"54",
          8226 => x"15",
          8227 => x"ff",
          8228 => x"82",
          8229 => x"55",
          8230 => x"98",
          8231 => x"0d",
          8232 => x"0d",
          8233 => x"53",
          8234 => x"05",
          8235 => x"51",
          8236 => x"82",
          8237 => x"55",
          8238 => x"08",
          8239 => x"76",
          8240 => x"93",
          8241 => x"51",
          8242 => x"82",
          8243 => x"55",
          8244 => x"08",
          8245 => x"80",
          8246 => x"81",
          8247 => x"86",
          8248 => x"38",
          8249 => x"86",
          8250 => x"90",
          8251 => x"54",
          8252 => x"ff",
          8253 => x"76",
          8254 => x"83",
          8255 => x"51",
          8256 => x"3f",
          8257 => x"08",
          8258 => x"bb",
          8259 => x"3d",
          8260 => x"3d",
          8261 => x"5c",
          8262 => x"98",
          8263 => x"52",
          8264 => x"d1",
          8265 => x"bb",
          8266 => x"bb",
          8267 => x"70",
          8268 => x"08",
          8269 => x"51",
          8270 => x"80",
          8271 => x"38",
          8272 => x"06",
          8273 => x"80",
          8274 => x"38",
          8275 => x"5f",
          8276 => x"3d",
          8277 => x"ff",
          8278 => x"82",
          8279 => x"57",
          8280 => x"08",
          8281 => x"74",
          8282 => x"c3",
          8283 => x"bb",
          8284 => x"82",
          8285 => x"bf",
          8286 => x"98",
          8287 => x"98",
          8288 => x"59",
          8289 => x"81",
          8290 => x"56",
          8291 => x"33",
          8292 => x"16",
          8293 => x"27",
          8294 => x"56",
          8295 => x"80",
          8296 => x"80",
          8297 => x"ff",
          8298 => x"70",
          8299 => x"56",
          8300 => x"e8",
          8301 => x"76",
          8302 => x"81",
          8303 => x"80",
          8304 => x"57",
          8305 => x"78",
          8306 => x"51",
          8307 => x"2e",
          8308 => x"73",
          8309 => x"38",
          8310 => x"08",
          8311 => x"b1",
          8312 => x"bb",
          8313 => x"82",
          8314 => x"a7",
          8315 => x"33",
          8316 => x"c3",
          8317 => x"2e",
          8318 => x"e4",
          8319 => x"2e",
          8320 => x"56",
          8321 => x"05",
          8322 => x"e3",
          8323 => x"98",
          8324 => x"76",
          8325 => x"0c",
          8326 => x"04",
          8327 => x"82",
          8328 => x"ff",
          8329 => x"9d",
          8330 => x"fa",
          8331 => x"98",
          8332 => x"98",
          8333 => x"82",
          8334 => x"83",
          8335 => x"53",
          8336 => x"3d",
          8337 => x"ff",
          8338 => x"73",
          8339 => x"70",
          8340 => x"52",
          8341 => x"9f",
          8342 => x"bc",
          8343 => x"74",
          8344 => x"6d",
          8345 => x"70",
          8346 => x"af",
          8347 => x"bb",
          8348 => x"2e",
          8349 => x"70",
          8350 => x"57",
          8351 => x"fd",
          8352 => x"98",
          8353 => x"8d",
          8354 => x"2b",
          8355 => x"81",
          8356 => x"86",
          8357 => x"98",
          8358 => x"9f",
          8359 => x"ff",
          8360 => x"54",
          8361 => x"8a",
          8362 => x"70",
          8363 => x"06",
          8364 => x"ff",
          8365 => x"38",
          8366 => x"15",
          8367 => x"80",
          8368 => x"74",
          8369 => x"e0",
          8370 => x"89",
          8371 => x"98",
          8372 => x"81",
          8373 => x"88",
          8374 => x"26",
          8375 => x"39",
          8376 => x"86",
          8377 => x"81",
          8378 => x"ff",
          8379 => x"38",
          8380 => x"54",
          8381 => x"81",
          8382 => x"81",
          8383 => x"78",
          8384 => x"5a",
          8385 => x"6d",
          8386 => x"81",
          8387 => x"57",
          8388 => x"9f",
          8389 => x"38",
          8390 => x"54",
          8391 => x"81",
          8392 => x"b1",
          8393 => x"2e",
          8394 => x"a7",
          8395 => x"15",
          8396 => x"54",
          8397 => x"09",
          8398 => x"38",
          8399 => x"76",
          8400 => x"41",
          8401 => x"52",
          8402 => x"52",
          8403 => x"b3",
          8404 => x"98",
          8405 => x"bb",
          8406 => x"f7",
          8407 => x"74",
          8408 => x"e5",
          8409 => x"98",
          8410 => x"bb",
          8411 => x"38",
          8412 => x"38",
          8413 => x"74",
          8414 => x"39",
          8415 => x"08",
          8416 => x"81",
          8417 => x"38",
          8418 => x"74",
          8419 => x"38",
          8420 => x"51",
          8421 => x"3f",
          8422 => x"08",
          8423 => x"98",
          8424 => x"a0",
          8425 => x"98",
          8426 => x"51",
          8427 => x"3f",
          8428 => x"0b",
          8429 => x"8b",
          8430 => x"67",
          8431 => x"a7",
          8432 => x"81",
          8433 => x"34",
          8434 => x"ad",
          8435 => x"bb",
          8436 => x"73",
          8437 => x"bb",
          8438 => x"3d",
          8439 => x"3d",
          8440 => x"02",
          8441 => x"cb",
          8442 => x"3d",
          8443 => x"72",
          8444 => x"5a",
          8445 => x"82",
          8446 => x"58",
          8447 => x"08",
          8448 => x"91",
          8449 => x"77",
          8450 => x"7c",
          8451 => x"38",
          8452 => x"59",
          8453 => x"90",
          8454 => x"81",
          8455 => x"06",
          8456 => x"73",
          8457 => x"54",
          8458 => x"82",
          8459 => x"39",
          8460 => x"8b",
          8461 => x"11",
          8462 => x"2b",
          8463 => x"54",
          8464 => x"fe",
          8465 => x"ff",
          8466 => x"70",
          8467 => x"07",
          8468 => x"bb",
          8469 => x"8c",
          8470 => x"40",
          8471 => x"55",
          8472 => x"88",
          8473 => x"08",
          8474 => x"38",
          8475 => x"77",
          8476 => x"56",
          8477 => x"51",
          8478 => x"3f",
          8479 => x"55",
          8480 => x"08",
          8481 => x"38",
          8482 => x"bb",
          8483 => x"2e",
          8484 => x"82",
          8485 => x"ff",
          8486 => x"38",
          8487 => x"08",
          8488 => x"16",
          8489 => x"2e",
          8490 => x"87",
          8491 => x"74",
          8492 => x"74",
          8493 => x"81",
          8494 => x"38",
          8495 => x"ff",
          8496 => x"2e",
          8497 => x"7b",
          8498 => x"80",
          8499 => x"81",
          8500 => x"81",
          8501 => x"06",
          8502 => x"56",
          8503 => x"52",
          8504 => x"af",
          8505 => x"bb",
          8506 => x"82",
          8507 => x"80",
          8508 => x"81",
          8509 => x"56",
          8510 => x"d3",
          8511 => x"ff",
          8512 => x"7c",
          8513 => x"55",
          8514 => x"b3",
          8515 => x"1b",
          8516 => x"1b",
          8517 => x"33",
          8518 => x"54",
          8519 => x"34",
          8520 => x"fe",
          8521 => x"08",
          8522 => x"74",
          8523 => x"75",
          8524 => x"16",
          8525 => x"33",
          8526 => x"73",
          8527 => x"77",
          8528 => x"bb",
          8529 => x"3d",
          8530 => x"3d",
          8531 => x"02",
          8532 => x"eb",
          8533 => x"3d",
          8534 => x"59",
          8535 => x"8b",
          8536 => x"82",
          8537 => x"24",
          8538 => x"82",
          8539 => x"84",
          8540 => x"d0",
          8541 => x"51",
          8542 => x"2e",
          8543 => x"75",
          8544 => x"98",
          8545 => x"06",
          8546 => x"7e",
          8547 => x"d0",
          8548 => x"98",
          8549 => x"06",
          8550 => x"56",
          8551 => x"74",
          8552 => x"76",
          8553 => x"81",
          8554 => x"8a",
          8555 => x"b2",
          8556 => x"fc",
          8557 => x"52",
          8558 => x"a4",
          8559 => x"bb",
          8560 => x"38",
          8561 => x"80",
          8562 => x"74",
          8563 => x"26",
          8564 => x"15",
          8565 => x"74",
          8566 => x"38",
          8567 => x"80",
          8568 => x"84",
          8569 => x"92",
          8570 => x"80",
          8571 => x"38",
          8572 => x"06",
          8573 => x"2e",
          8574 => x"56",
          8575 => x"78",
          8576 => x"89",
          8577 => x"2b",
          8578 => x"43",
          8579 => x"38",
          8580 => x"30",
          8581 => x"77",
          8582 => x"91",
          8583 => x"c2",
          8584 => x"f8",
          8585 => x"52",
          8586 => x"a4",
          8587 => x"56",
          8588 => x"08",
          8589 => x"77",
          8590 => x"77",
          8591 => x"98",
          8592 => x"45",
          8593 => x"bf",
          8594 => x"8e",
          8595 => x"26",
          8596 => x"74",
          8597 => x"48",
          8598 => x"75",
          8599 => x"38",
          8600 => x"81",
          8601 => x"fa",
          8602 => x"2a",
          8603 => x"56",
          8604 => x"2e",
          8605 => x"87",
          8606 => x"82",
          8607 => x"38",
          8608 => x"55",
          8609 => x"83",
          8610 => x"81",
          8611 => x"56",
          8612 => x"80",
          8613 => x"38",
          8614 => x"83",
          8615 => x"06",
          8616 => x"78",
          8617 => x"91",
          8618 => x"0b",
          8619 => x"22",
          8620 => x"80",
          8621 => x"74",
          8622 => x"38",
          8623 => x"56",
          8624 => x"17",
          8625 => x"57",
          8626 => x"2e",
          8627 => x"75",
          8628 => x"79",
          8629 => x"fe",
          8630 => x"82",
          8631 => x"84",
          8632 => x"05",
          8633 => x"5e",
          8634 => x"80",
          8635 => x"98",
          8636 => x"8a",
          8637 => x"fd",
          8638 => x"75",
          8639 => x"38",
          8640 => x"78",
          8641 => x"8c",
          8642 => x"0b",
          8643 => x"22",
          8644 => x"80",
          8645 => x"74",
          8646 => x"38",
          8647 => x"56",
          8648 => x"17",
          8649 => x"57",
          8650 => x"2e",
          8651 => x"75",
          8652 => x"79",
          8653 => x"fe",
          8654 => x"82",
          8655 => x"10",
          8656 => x"82",
          8657 => x"9f",
          8658 => x"38",
          8659 => x"bb",
          8660 => x"82",
          8661 => x"05",
          8662 => x"2a",
          8663 => x"56",
          8664 => x"17",
          8665 => x"81",
          8666 => x"60",
          8667 => x"65",
          8668 => x"12",
          8669 => x"30",
          8670 => x"74",
          8671 => x"59",
          8672 => x"7d",
          8673 => x"81",
          8674 => x"76",
          8675 => x"41",
          8676 => x"76",
          8677 => x"90",
          8678 => x"62",
          8679 => x"51",
          8680 => x"26",
          8681 => x"75",
          8682 => x"31",
          8683 => x"65",
          8684 => x"fe",
          8685 => x"82",
          8686 => x"58",
          8687 => x"09",
          8688 => x"38",
          8689 => x"08",
          8690 => x"26",
          8691 => x"78",
          8692 => x"79",
          8693 => x"78",
          8694 => x"86",
          8695 => x"82",
          8696 => x"06",
          8697 => x"83",
          8698 => x"82",
          8699 => x"27",
          8700 => x"8f",
          8701 => x"55",
          8702 => x"26",
          8703 => x"59",
          8704 => x"62",
          8705 => x"74",
          8706 => x"38",
          8707 => x"88",
          8708 => x"98",
          8709 => x"26",
          8710 => x"86",
          8711 => x"1a",
          8712 => x"79",
          8713 => x"38",
          8714 => x"80",
          8715 => x"2e",
          8716 => x"83",
          8717 => x"9f",
          8718 => x"8b",
          8719 => x"06",
          8720 => x"74",
          8721 => x"84",
          8722 => x"52",
          8723 => x"a2",
          8724 => x"53",
          8725 => x"52",
          8726 => x"a2",
          8727 => x"80",
          8728 => x"51",
          8729 => x"3f",
          8730 => x"34",
          8731 => x"ff",
          8732 => x"1b",
          8733 => x"a2",
          8734 => x"90",
          8735 => x"83",
          8736 => x"70",
          8737 => x"80",
          8738 => x"55",
          8739 => x"ff",
          8740 => x"66",
          8741 => x"ff",
          8742 => x"38",
          8743 => x"ff",
          8744 => x"1b",
          8745 => x"f2",
          8746 => x"74",
          8747 => x"51",
          8748 => x"3f",
          8749 => x"1c",
          8750 => x"98",
          8751 => x"a0",
          8752 => x"ff",
          8753 => x"51",
          8754 => x"3f",
          8755 => x"1b",
          8756 => x"e4",
          8757 => x"2e",
          8758 => x"80",
          8759 => x"88",
          8760 => x"80",
          8761 => x"ff",
          8762 => x"7c",
          8763 => x"51",
          8764 => x"3f",
          8765 => x"1b",
          8766 => x"bc",
          8767 => x"b0",
          8768 => x"a0",
          8769 => x"52",
          8770 => x"ff",
          8771 => x"ff",
          8772 => x"c0",
          8773 => x"0b",
          8774 => x"34",
          8775 => x"b4",
          8776 => x"c7",
          8777 => x"39",
          8778 => x"0a",
          8779 => x"51",
          8780 => x"3f",
          8781 => x"ff",
          8782 => x"1b",
          8783 => x"da",
          8784 => x"0b",
          8785 => x"a9",
          8786 => x"34",
          8787 => x"b4",
          8788 => x"1b",
          8789 => x"8f",
          8790 => x"d5",
          8791 => x"1b",
          8792 => x"ff",
          8793 => x"81",
          8794 => x"7a",
          8795 => x"ff",
          8796 => x"81",
          8797 => x"98",
          8798 => x"38",
          8799 => x"09",
          8800 => x"ee",
          8801 => x"60",
          8802 => x"7a",
          8803 => x"ff",
          8804 => x"84",
          8805 => x"52",
          8806 => x"9f",
          8807 => x"8b",
          8808 => x"52",
          8809 => x"9f",
          8810 => x"8a",
          8811 => x"52",
          8812 => x"51",
          8813 => x"3f",
          8814 => x"83",
          8815 => x"ff",
          8816 => x"82",
          8817 => x"1b",
          8818 => x"ec",
          8819 => x"d5",
          8820 => x"ff",
          8821 => x"75",
          8822 => x"05",
          8823 => x"7e",
          8824 => x"e5",
          8825 => x"60",
          8826 => x"52",
          8827 => x"9a",
          8828 => x"53",
          8829 => x"51",
          8830 => x"3f",
          8831 => x"58",
          8832 => x"09",
          8833 => x"38",
          8834 => x"51",
          8835 => x"3f",
          8836 => x"1b",
          8837 => x"a0",
          8838 => x"52",
          8839 => x"91",
          8840 => x"ff",
          8841 => x"81",
          8842 => x"f8",
          8843 => x"7a",
          8844 => x"84",
          8845 => x"61",
          8846 => x"26",
          8847 => x"57",
          8848 => x"53",
          8849 => x"51",
          8850 => x"3f",
          8851 => x"08",
          8852 => x"84",
          8853 => x"bb",
          8854 => x"7a",
          8855 => x"aa",
          8856 => x"75",
          8857 => x"56",
          8858 => x"81",
          8859 => x"80",
          8860 => x"38",
          8861 => x"83",
          8862 => x"63",
          8863 => x"74",
          8864 => x"38",
          8865 => x"54",
          8866 => x"52",
          8867 => x"99",
          8868 => x"bb",
          8869 => x"c1",
          8870 => x"75",
          8871 => x"56",
          8872 => x"8c",
          8873 => x"2e",
          8874 => x"56",
          8875 => x"ff",
          8876 => x"84",
          8877 => x"2e",
          8878 => x"56",
          8879 => x"58",
          8880 => x"38",
          8881 => x"77",
          8882 => x"ff",
          8883 => x"82",
          8884 => x"78",
          8885 => x"c2",
          8886 => x"1b",
          8887 => x"34",
          8888 => x"16",
          8889 => x"82",
          8890 => x"83",
          8891 => x"84",
          8892 => x"67",
          8893 => x"fd",
          8894 => x"51",
          8895 => x"3f",
          8896 => x"16",
          8897 => x"98",
          8898 => x"bf",
          8899 => x"86",
          8900 => x"bb",
          8901 => x"16",
          8902 => x"83",
          8903 => x"ff",
          8904 => x"66",
          8905 => x"1b",
          8906 => x"8c",
          8907 => x"77",
          8908 => x"7e",
          8909 => x"91",
          8910 => x"82",
          8911 => x"a2",
          8912 => x"80",
          8913 => x"ff",
          8914 => x"81",
          8915 => x"98",
          8916 => x"89",
          8917 => x"8a",
          8918 => x"86",
          8919 => x"98",
          8920 => x"82",
          8921 => x"99",
          8922 => x"f5",
          8923 => x"60",
          8924 => x"79",
          8925 => x"5a",
          8926 => x"78",
          8927 => x"8d",
          8928 => x"55",
          8929 => x"fc",
          8930 => x"51",
          8931 => x"7a",
          8932 => x"81",
          8933 => x"8c",
          8934 => x"74",
          8935 => x"38",
          8936 => x"81",
          8937 => x"81",
          8938 => x"8a",
          8939 => x"06",
          8940 => x"76",
          8941 => x"76",
          8942 => x"55",
          8943 => x"98",
          8944 => x"0d",
          8945 => x"0d",
          8946 => x"05",
          8947 => x"59",
          8948 => x"2e",
          8949 => x"87",
          8950 => x"76",
          8951 => x"84",
          8952 => x"80",
          8953 => x"38",
          8954 => x"77",
          8955 => x"56",
          8956 => x"34",
          8957 => x"bb",
          8958 => x"38",
          8959 => x"05",
          8960 => x"8c",
          8961 => x"08",
          8962 => x"3f",
          8963 => x"70",
          8964 => x"07",
          8965 => x"30",
          8966 => x"56",
          8967 => x"0c",
          8968 => x"18",
          8969 => x"0d",
          8970 => x"0d",
          8971 => x"08",
          8972 => x"75",
          8973 => x"89",
          8974 => x"54",
          8975 => x"16",
          8976 => x"51",
          8977 => x"82",
          8978 => x"91",
          8979 => x"08",
          8980 => x"81",
          8981 => x"88",
          8982 => x"83",
          8983 => x"74",
          8984 => x"0c",
          8985 => x"04",
          8986 => x"75",
          8987 => x"53",
          8988 => x"51",
          8989 => x"3f",
          8990 => x"85",
          8991 => x"ea",
          8992 => x"80",
          8993 => x"6a",
          8994 => x"70",
          8995 => x"d8",
          8996 => x"72",
          8997 => x"3f",
          8998 => x"8d",
          8999 => x"0d",
          9000 => x"ff",
          9001 => x"ff",
          9002 => x"00",
          9003 => x"ff",
          9004 => x"2b",
          9005 => x"2b",
          9006 => x"2b",
          9007 => x"2b",
          9008 => x"2b",
          9009 => x"2b",
          9010 => x"2b",
          9011 => x"2b",
          9012 => x"2b",
          9013 => x"2b",
          9014 => x"2b",
          9015 => x"2b",
          9016 => x"2b",
          9017 => x"2b",
          9018 => x"2b",
          9019 => x"2b",
          9020 => x"2b",
          9021 => x"2b",
          9022 => x"2b",
          9023 => x"2b",
          9024 => x"43",
          9025 => x"43",
          9026 => x"43",
          9027 => x"43",
          9028 => x"43",
          9029 => x"49",
          9030 => x"4a",
          9031 => x"4b",
          9032 => x"4d",
          9033 => x"4a",
          9034 => x"48",
          9035 => x"4c",
          9036 => x"4d",
          9037 => x"4c",
          9038 => x"4d",
          9039 => x"4c",
          9040 => x"4b",
          9041 => x"48",
          9042 => x"4b",
          9043 => x"4b",
          9044 => x"4c",
          9045 => x"48",
          9046 => x"48",
          9047 => x"4c",
          9048 => x"4d",
          9049 => x"4d",
          9050 => x"4d",
          9051 => x"0e",
          9052 => x"17",
          9053 => x"17",
          9054 => x"0e",
          9055 => x"17",
          9056 => x"17",
          9057 => x"17",
          9058 => x"17",
          9059 => x"17",
          9060 => x"17",
          9061 => x"17",
          9062 => x"0e",
          9063 => x"17",
          9064 => x"0e",
          9065 => x"0e",
          9066 => x"17",
          9067 => x"17",
          9068 => x"17",
          9069 => x"17",
          9070 => x"17",
          9071 => x"17",
          9072 => x"17",
          9073 => x"17",
          9074 => x"17",
          9075 => x"17",
          9076 => x"17",
          9077 => x"17",
          9078 => x"17",
          9079 => x"17",
          9080 => x"17",
          9081 => x"17",
          9082 => x"17",
          9083 => x"17",
          9084 => x"17",
          9085 => x"17",
          9086 => x"17",
          9087 => x"17",
          9088 => x"17",
          9089 => x"17",
          9090 => x"17",
          9091 => x"17",
          9092 => x"17",
          9093 => x"17",
          9094 => x"17",
          9095 => x"17",
          9096 => x"17",
          9097 => x"17",
          9098 => x"17",
          9099 => x"17",
          9100 => x"17",
          9101 => x"17",
          9102 => x"0f",
          9103 => x"17",
          9104 => x"17",
          9105 => x"17",
          9106 => x"17",
          9107 => x"11",
          9108 => x"17",
          9109 => x"17",
          9110 => x"17",
          9111 => x"17",
          9112 => x"17",
          9113 => x"17",
          9114 => x"17",
          9115 => x"17",
          9116 => x"17",
          9117 => x"17",
          9118 => x"0e",
          9119 => x"10",
          9120 => x"0e",
          9121 => x"0e",
          9122 => x"0e",
          9123 => x"17",
          9124 => x"10",
          9125 => x"17",
          9126 => x"17",
          9127 => x"0e",
          9128 => x"17",
          9129 => x"17",
          9130 => x"10",
          9131 => x"10",
          9132 => x"17",
          9133 => x"17",
          9134 => x"0f",
          9135 => x"17",
          9136 => x"11",
          9137 => x"17",
          9138 => x"17",
          9139 => x"11",
          9140 => x"6e",
          9141 => x"00",
          9142 => x"6f",
          9143 => x"00",
          9144 => x"6e",
          9145 => x"00",
          9146 => x"6f",
          9147 => x"00",
          9148 => x"78",
          9149 => x"00",
          9150 => x"6c",
          9151 => x"00",
          9152 => x"6f",
          9153 => x"00",
          9154 => x"69",
          9155 => x"00",
          9156 => x"75",
          9157 => x"00",
          9158 => x"62",
          9159 => x"68",
          9160 => x"77",
          9161 => x"64",
          9162 => x"65",
          9163 => x"64",
          9164 => x"65",
          9165 => x"6c",
          9166 => x"00",
          9167 => x"70",
          9168 => x"73",
          9169 => x"74",
          9170 => x"73",
          9171 => x"00",
          9172 => x"66",
          9173 => x"00",
          9174 => x"73",
          9175 => x"00",
          9176 => x"61",
          9177 => x"00",
          9178 => x"61",
          9179 => x"00",
          9180 => x"6c",
          9181 => x"00",
          9182 => x"00",
          9183 => x"73",
          9184 => x"72",
          9185 => x"0a",
          9186 => x"74",
          9187 => x"61",
          9188 => x"72",
          9189 => x"2e",
          9190 => x"00",
          9191 => x"73",
          9192 => x"6f",
          9193 => x"65",
          9194 => x"2e",
          9195 => x"00",
          9196 => x"20",
          9197 => x"65",
          9198 => x"75",
          9199 => x"0a",
          9200 => x"20",
          9201 => x"68",
          9202 => x"75",
          9203 => x"0a",
          9204 => x"76",
          9205 => x"64",
          9206 => x"6c",
          9207 => x"6d",
          9208 => x"00",
          9209 => x"63",
          9210 => x"20",
          9211 => x"69",
          9212 => x"0a",
          9213 => x"6c",
          9214 => x"6c",
          9215 => x"64",
          9216 => x"78",
          9217 => x"73",
          9218 => x"00",
          9219 => x"6c",
          9220 => x"61",
          9221 => x"65",
          9222 => x"76",
          9223 => x"64",
          9224 => x"00",
          9225 => x"20",
          9226 => x"77",
          9227 => x"65",
          9228 => x"6f",
          9229 => x"74",
          9230 => x"0a",
          9231 => x"69",
          9232 => x"6e",
          9233 => x"65",
          9234 => x"73",
          9235 => x"76",
          9236 => x"64",
          9237 => x"00",
          9238 => x"73",
          9239 => x"6f",
          9240 => x"6e",
          9241 => x"65",
          9242 => x"00",
          9243 => x"20",
          9244 => x"70",
          9245 => x"62",
          9246 => x"66",
          9247 => x"73",
          9248 => x"65",
          9249 => x"6f",
          9250 => x"20",
          9251 => x"64",
          9252 => x"2e",
          9253 => x"00",
          9254 => x"72",
          9255 => x"20",
          9256 => x"72",
          9257 => x"2e",
          9258 => x"00",
          9259 => x"6d",
          9260 => x"74",
          9261 => x"70",
          9262 => x"74",
          9263 => x"20",
          9264 => x"63",
          9265 => x"65",
          9266 => x"00",
          9267 => x"6c",
          9268 => x"73",
          9269 => x"63",
          9270 => x"2e",
          9271 => x"00",
          9272 => x"73",
          9273 => x"69",
          9274 => x"6e",
          9275 => x"65",
          9276 => x"79",
          9277 => x"00",
          9278 => x"6f",
          9279 => x"6e",
          9280 => x"70",
          9281 => x"66",
          9282 => x"73",
          9283 => x"00",
          9284 => x"72",
          9285 => x"74",
          9286 => x"20",
          9287 => x"6f",
          9288 => x"63",
          9289 => x"00",
          9290 => x"63",
          9291 => x"73",
          9292 => x"00",
          9293 => x"6b",
          9294 => x"6e",
          9295 => x"72",
          9296 => x"0a",
          9297 => x"6c",
          9298 => x"79",
          9299 => x"20",
          9300 => x"61",
          9301 => x"6c",
          9302 => x"79",
          9303 => x"2f",
          9304 => x"2e",
          9305 => x"00",
          9306 => x"61",
          9307 => x"00",
          9308 => x"38",
          9309 => x"00",
          9310 => x"20",
          9311 => x"34",
          9312 => x"00",
          9313 => x"20",
          9314 => x"20",
          9315 => x"00",
          9316 => x"32",
          9317 => x"00",
          9318 => x"00",
          9319 => x"00",
          9320 => x"0a",
          9321 => x"55",
          9322 => x"00",
          9323 => x"2a",
          9324 => x"20",
          9325 => x"00",
          9326 => x"2f",
          9327 => x"32",
          9328 => x"00",
          9329 => x"2e",
          9330 => x"00",
          9331 => x"50",
          9332 => x"72",
          9333 => x"25",
          9334 => x"29",
          9335 => x"20",
          9336 => x"2a",
          9337 => x"00",
          9338 => x"55",
          9339 => x"49",
          9340 => x"72",
          9341 => x"74",
          9342 => x"6e",
          9343 => x"72",
          9344 => x"00",
          9345 => x"6d",
          9346 => x"69",
          9347 => x"72",
          9348 => x"74",
          9349 => x"00",
          9350 => x"32",
          9351 => x"74",
          9352 => x"75",
          9353 => x"00",
          9354 => x"43",
          9355 => x"52",
          9356 => x"6e",
          9357 => x"72",
          9358 => x"0a",
          9359 => x"43",
          9360 => x"57",
          9361 => x"6e",
          9362 => x"72",
          9363 => x"0a",
          9364 => x"52",
          9365 => x"52",
          9366 => x"6e",
          9367 => x"72",
          9368 => x"0a",
          9369 => x"52",
          9370 => x"54",
          9371 => x"6e",
          9372 => x"72",
          9373 => x"0a",
          9374 => x"52",
          9375 => x"52",
          9376 => x"6e",
          9377 => x"72",
          9378 => x"0a",
          9379 => x"52",
          9380 => x"54",
          9381 => x"6e",
          9382 => x"72",
          9383 => x"0a",
          9384 => x"74",
          9385 => x"67",
          9386 => x"20",
          9387 => x"65",
          9388 => x"2e",
          9389 => x"00",
          9390 => x"61",
          9391 => x"6e",
          9392 => x"69",
          9393 => x"2e",
          9394 => x"00",
          9395 => x"74",
          9396 => x"65",
          9397 => x"61",
          9398 => x"00",
          9399 => x"75",
          9400 => x"68",
          9401 => x"00",
          9402 => x"00",
          9403 => x"69",
          9404 => x"20",
          9405 => x"69",
          9406 => x"69",
          9407 => x"73",
          9408 => x"64",
          9409 => x"72",
          9410 => x"2c",
          9411 => x"65",
          9412 => x"20",
          9413 => x"74",
          9414 => x"6e",
          9415 => x"6c",
          9416 => x"00",
          9417 => x"00",
          9418 => x"64",
          9419 => x"73",
          9420 => x"64",
          9421 => x"00",
          9422 => x"69",
          9423 => x"6c",
          9424 => x"64",
          9425 => x"00",
          9426 => x"69",
          9427 => x"20",
          9428 => x"69",
          9429 => x"69",
          9430 => x"73",
          9431 => x"00",
          9432 => x"3d",
          9433 => x"00",
          9434 => x"3a",
          9435 => x"65",
          9436 => x"6e",
          9437 => x"2e",
          9438 => x"00",
          9439 => x"70",
          9440 => x"67",
          9441 => x"00",
          9442 => x"6d",
          9443 => x"69",
          9444 => x"2e",
          9445 => x"00",
          9446 => x"38",
          9447 => x"25",
          9448 => x"29",
          9449 => x"30",
          9450 => x"28",
          9451 => x"78",
          9452 => x"00",
          9453 => x"6d",
          9454 => x"65",
          9455 => x"79",
          9456 => x"00",
          9457 => x"6f",
          9458 => x"65",
          9459 => x"0a",
          9460 => x"38",
          9461 => x"30",
          9462 => x"00",
          9463 => x"3f",
          9464 => x"00",
          9465 => x"38",
          9466 => x"30",
          9467 => x"00",
          9468 => x"38",
          9469 => x"30",
          9470 => x"00",
          9471 => x"73",
          9472 => x"69",
          9473 => x"69",
          9474 => x"72",
          9475 => x"74",
          9476 => x"00",
          9477 => x"61",
          9478 => x"6e",
          9479 => x"6e",
          9480 => x"72",
          9481 => x"73",
          9482 => x"00",
          9483 => x"73",
          9484 => x"65",
          9485 => x"61",
          9486 => x"66",
          9487 => x"0a",
          9488 => x"61",
          9489 => x"6e",
          9490 => x"61",
          9491 => x"66",
          9492 => x"0a",
          9493 => x"65",
          9494 => x"69",
          9495 => x"63",
          9496 => x"20",
          9497 => x"30",
          9498 => x"2e",
          9499 => x"00",
          9500 => x"6c",
          9501 => x"67",
          9502 => x"64",
          9503 => x"20",
          9504 => x"78",
          9505 => x"2e",
          9506 => x"00",
          9507 => x"6c",
          9508 => x"65",
          9509 => x"6e",
          9510 => x"63",
          9511 => x"20",
          9512 => x"29",
          9513 => x"00",
          9514 => x"73",
          9515 => x"74",
          9516 => x"20",
          9517 => x"6c",
          9518 => x"74",
          9519 => x"2e",
          9520 => x"00",
          9521 => x"6c",
          9522 => x"65",
          9523 => x"74",
          9524 => x"2e",
          9525 => x"00",
          9526 => x"55",
          9527 => x"6e",
          9528 => x"3a",
          9529 => x"5c",
          9530 => x"25",
          9531 => x"00",
          9532 => x"3a",
          9533 => x"5c",
          9534 => x"00",
          9535 => x"3a",
          9536 => x"00",
          9537 => x"64",
          9538 => x"6d",
          9539 => x"64",
          9540 => x"00",
          9541 => x"6e",
          9542 => x"67",
          9543 => x"0a",
          9544 => x"61",
          9545 => x"6e",
          9546 => x"6e",
          9547 => x"72",
          9548 => x"73",
          9549 => x"0a",
          9550 => x"2f",
          9551 => x"25",
          9552 => x"64",
          9553 => x"3a",
          9554 => x"25",
          9555 => x"0a",
          9556 => x"43",
          9557 => x"6e",
          9558 => x"75",
          9559 => x"69",
          9560 => x"00",
          9561 => x"66",
          9562 => x"20",
          9563 => x"20",
          9564 => x"66",
          9565 => x"00",
          9566 => x"44",
          9567 => x"63",
          9568 => x"69",
          9569 => x"65",
          9570 => x"74",
          9571 => x"0a",
          9572 => x"20",
          9573 => x"20",
          9574 => x"41",
          9575 => x"28",
          9576 => x"58",
          9577 => x"38",
          9578 => x"0a",
          9579 => x"20",
          9580 => x"52",
          9581 => x"20",
          9582 => x"28",
          9583 => x"58",
          9584 => x"38",
          9585 => x"0a",
          9586 => x"20",
          9587 => x"53",
          9588 => x"52",
          9589 => x"28",
          9590 => x"58",
          9591 => x"38",
          9592 => x"0a",
          9593 => x"20",
          9594 => x"41",
          9595 => x"20",
          9596 => x"28",
          9597 => x"58",
          9598 => x"38",
          9599 => x"0a",
          9600 => x"20",
          9601 => x"4d",
          9602 => x"20",
          9603 => x"28",
          9604 => x"58",
          9605 => x"38",
          9606 => x"0a",
          9607 => x"20",
          9608 => x"20",
          9609 => x"44",
          9610 => x"28",
          9611 => x"69",
          9612 => x"20",
          9613 => x"32",
          9614 => x"0a",
          9615 => x"20",
          9616 => x"4d",
          9617 => x"20",
          9618 => x"28",
          9619 => x"65",
          9620 => x"20",
          9621 => x"32",
          9622 => x"0a",
          9623 => x"20",
          9624 => x"54",
          9625 => x"54",
          9626 => x"28",
          9627 => x"6e",
          9628 => x"73",
          9629 => x"32",
          9630 => x"0a",
          9631 => x"20",
          9632 => x"53",
          9633 => x"4e",
          9634 => x"55",
          9635 => x"00",
          9636 => x"20",
          9637 => x"20",
          9638 => x"0a",
          9639 => x"20",
          9640 => x"43",
          9641 => x"00",
          9642 => x"20",
          9643 => x"32",
          9644 => x"00",
          9645 => x"20",
          9646 => x"49",
          9647 => x"00",
          9648 => x"64",
          9649 => x"73",
          9650 => x"0a",
          9651 => x"20",
          9652 => x"55",
          9653 => x"73",
          9654 => x"56",
          9655 => x"6f",
          9656 => x"64",
          9657 => x"73",
          9658 => x"20",
          9659 => x"58",
          9660 => x"00",
          9661 => x"20",
          9662 => x"55",
          9663 => x"6d",
          9664 => x"20",
          9665 => x"72",
          9666 => x"64",
          9667 => x"73",
          9668 => x"20",
          9669 => x"58",
          9670 => x"00",
          9671 => x"20",
          9672 => x"61",
          9673 => x"53",
          9674 => x"74",
          9675 => x"64",
          9676 => x"73",
          9677 => x"20",
          9678 => x"20",
          9679 => x"58",
          9680 => x"00",
          9681 => x"73",
          9682 => x"00",
          9683 => x"20",
          9684 => x"55",
          9685 => x"20",
          9686 => x"20",
          9687 => x"20",
          9688 => x"20",
          9689 => x"20",
          9690 => x"20",
          9691 => x"58",
          9692 => x"00",
          9693 => x"20",
          9694 => x"73",
          9695 => x"20",
          9696 => x"63",
          9697 => x"72",
          9698 => x"20",
          9699 => x"20",
          9700 => x"20",
          9701 => x"25",
          9702 => x"4d",
          9703 => x"00",
          9704 => x"20",
          9705 => x"52",
          9706 => x"43",
          9707 => x"6b",
          9708 => x"65",
          9709 => x"20",
          9710 => x"20",
          9711 => x"20",
          9712 => x"25",
          9713 => x"4d",
          9714 => x"00",
          9715 => x"20",
          9716 => x"73",
          9717 => x"6e",
          9718 => x"44",
          9719 => x"20",
          9720 => x"63",
          9721 => x"72",
          9722 => x"20",
          9723 => x"25",
          9724 => x"4d",
          9725 => x"00",
          9726 => x"61",
          9727 => x"00",
          9728 => x"64",
          9729 => x"00",
          9730 => x"65",
          9731 => x"00",
          9732 => x"4f",
          9733 => x"4f",
          9734 => x"00",
          9735 => x"6b",
          9736 => x"6e",
          9737 => x"99",
          9738 => x"00",
          9739 => x"00",
          9740 => x"99",
          9741 => x"00",
          9742 => x"00",
          9743 => x"99",
          9744 => x"00",
          9745 => x"00",
          9746 => x"99",
          9747 => x"00",
          9748 => x"00",
          9749 => x"99",
          9750 => x"00",
          9751 => x"00",
          9752 => x"99",
          9753 => x"00",
          9754 => x"00",
          9755 => x"99",
          9756 => x"00",
          9757 => x"00",
          9758 => x"99",
          9759 => x"00",
          9760 => x"00",
          9761 => x"99",
          9762 => x"00",
          9763 => x"00",
          9764 => x"99",
          9765 => x"00",
          9766 => x"00",
          9767 => x"99",
          9768 => x"00",
          9769 => x"00",
          9770 => x"99",
          9771 => x"00",
          9772 => x"00",
          9773 => x"99",
          9774 => x"00",
          9775 => x"00",
          9776 => x"99",
          9777 => x"00",
          9778 => x"00",
          9779 => x"99",
          9780 => x"00",
          9781 => x"00",
          9782 => x"99",
          9783 => x"00",
          9784 => x"00",
          9785 => x"99",
          9786 => x"00",
          9787 => x"00",
          9788 => x"99",
          9789 => x"00",
          9790 => x"00",
          9791 => x"99",
          9792 => x"00",
          9793 => x"00",
          9794 => x"99",
          9795 => x"00",
          9796 => x"00",
          9797 => x"99",
          9798 => x"00",
          9799 => x"00",
          9800 => x"99",
          9801 => x"00",
          9802 => x"00",
          9803 => x"44",
          9804 => x"43",
          9805 => x"42",
          9806 => x"41",
          9807 => x"36",
          9808 => x"35",
          9809 => x"34",
          9810 => x"46",
          9811 => x"33",
          9812 => x"32",
          9813 => x"31",
          9814 => x"00",
          9815 => x"00",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"00",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"00",
          9824 => x"00",
          9825 => x"73",
          9826 => x"79",
          9827 => x"73",
          9828 => x"00",
          9829 => x"00",
          9830 => x"34",
          9831 => x"25",
          9832 => x"00",
          9833 => x"69",
          9834 => x"20",
          9835 => x"72",
          9836 => x"74",
          9837 => x"65",
          9838 => x"73",
          9839 => x"79",
          9840 => x"6c",
          9841 => x"6f",
          9842 => x"46",
          9843 => x"00",
          9844 => x"6e",
          9845 => x"20",
          9846 => x"6e",
          9847 => x"65",
          9848 => x"20",
          9849 => x"74",
          9850 => x"20",
          9851 => x"65",
          9852 => x"69",
          9853 => x"6c",
          9854 => x"2e",
          9855 => x"00",
          9856 => x"2b",
          9857 => x"3c",
          9858 => x"5b",
          9859 => x"00",
          9860 => x"54",
          9861 => x"54",
          9862 => x"00",
          9863 => x"90",
          9864 => x"4f",
          9865 => x"30",
          9866 => x"20",
          9867 => x"45",
          9868 => x"20",
          9869 => x"33",
          9870 => x"20",
          9871 => x"20",
          9872 => x"45",
          9873 => x"20",
          9874 => x"20",
          9875 => x"20",
          9876 => x"99",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"45",
          9881 => x"8f",
          9882 => x"45",
          9883 => x"8e",
          9884 => x"92",
          9885 => x"55",
          9886 => x"9a",
          9887 => x"9e",
          9888 => x"4f",
          9889 => x"a6",
          9890 => x"aa",
          9891 => x"ae",
          9892 => x"b2",
          9893 => x"b6",
          9894 => x"ba",
          9895 => x"be",
          9896 => x"c2",
          9897 => x"c6",
          9898 => x"ca",
          9899 => x"ce",
          9900 => x"d2",
          9901 => x"d6",
          9902 => x"da",
          9903 => x"de",
          9904 => x"e2",
          9905 => x"e6",
          9906 => x"ea",
          9907 => x"ee",
          9908 => x"f2",
          9909 => x"f6",
          9910 => x"fa",
          9911 => x"fe",
          9912 => x"2c",
          9913 => x"5d",
          9914 => x"2a",
          9915 => x"3f",
          9916 => x"00",
          9917 => x"00",
          9918 => x"00",
          9919 => x"02",
          9920 => x"00",
          9921 => x"00",
          9922 => x"00",
          9923 => x"00",
          9924 => x"00",
          9925 => x"00",
          9926 => x"8e",
          9927 => x"01",
          9928 => x"00",
          9929 => x"00",
          9930 => x"8e",
          9931 => x"01",
          9932 => x"00",
          9933 => x"00",
          9934 => x"8e",
          9935 => x"03",
          9936 => x"00",
          9937 => x"00",
          9938 => x"8e",
          9939 => x"03",
          9940 => x"00",
          9941 => x"00",
          9942 => x"8e",
          9943 => x"03",
          9944 => x"00",
          9945 => x"00",
          9946 => x"8e",
          9947 => x"04",
          9948 => x"00",
          9949 => x"00",
          9950 => x"8f",
          9951 => x"04",
          9952 => x"00",
          9953 => x"00",
          9954 => x"8f",
          9955 => x"04",
          9956 => x"00",
          9957 => x"00",
          9958 => x"8f",
          9959 => x"04",
          9960 => x"00",
          9961 => x"00",
          9962 => x"8f",
          9963 => x"04",
          9964 => x"00",
          9965 => x"00",
          9966 => x"8f",
          9967 => x"04",
          9968 => x"00",
          9969 => x"00",
          9970 => x"8f",
          9971 => x"04",
          9972 => x"00",
          9973 => x"00",
          9974 => x"8f",
          9975 => x"05",
          9976 => x"00",
          9977 => x"00",
          9978 => x"8f",
          9979 => x"05",
          9980 => x"00",
          9981 => x"00",
          9982 => x"8f",
          9983 => x"05",
          9984 => x"00",
          9985 => x"00",
          9986 => x"8f",
          9987 => x"05",
          9988 => x"00",
          9989 => x"00",
          9990 => x"8f",
          9991 => x"07",
          9992 => x"00",
          9993 => x"00",
          9994 => x"8f",
          9995 => x"07",
          9996 => x"00",
          9997 => x"00",
          9998 => x"8f",
          9999 => x"08",
         10000 => x"00",
         10001 => x"00",
         10002 => x"8f",
         10003 => x"08",
         10004 => x"00",
         10005 => x"00",
         10006 => x"8f",
         10007 => x"08",
         10008 => x"00",
         10009 => x"00",
         10010 => x"8f",
         10011 => x"08",
         10012 => x"00",
         10013 => x"00",
         10014 => x"8f",
         10015 => x"09",
         10016 => x"00",
         10017 => x"00",
         10018 => x"8f",
         10019 => x"09",
         10020 => x"00",
         10021 => x"00",
         10022 => x"8f",
         10023 => x"09",
         10024 => x"00",
         10025 => x"00",
         10026 => x"8f",
         10027 => x"09",
         10028 => x"00",
         10029 => x"00",
         10030 => x"00",
         10031 => x"00",
         10032 => x"7f",
         10033 => x"00",
         10034 => x"7f",
         10035 => x"00",
         10036 => x"7f",
         10037 => x"00",
         10038 => x"00",
         10039 => x"00",
         10040 => x"ff",
         10041 => x"00",
         10042 => x"00",
         10043 => x"78",
         10044 => x"00",
         10045 => x"e1",
         10046 => x"e1",
         10047 => x"e1",
         10048 => x"00",
         10049 => x"01",
         10050 => x"01",
         10051 => x"10",
         10052 => x"00",
         10053 => x"00",
         10054 => x"00",
         10055 => x"00",
         10056 => x"00",
         10057 => x"00",
         10058 => x"00",
         10059 => x"00",
         10060 => x"00",
         10061 => x"00",
         10062 => x"00",
         10063 => x"00",
         10064 => x"00",
         10065 => x"00",
         10066 => x"00",
         10067 => x"00",
         10068 => x"00",
         10069 => x"00",
         10070 => x"00",
         10071 => x"00",
         10072 => x"00",
         10073 => x"00",
         10074 => x"00",
         10075 => x"00",
         10076 => x"00",
         10077 => x"99",
         10078 => x"00",
         10079 => x"99",
         10080 => x"00",
         10081 => x"99",
         10082 => x"00",
         10083 => x"00",
         10084 => x"00",
         10085 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"83",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8c",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"80",
           387 => x"82",
           388 => x"82",
           389 => x"82",
           390 => x"be",
           391 => x"bb",
           392 => x"e0",
           393 => x"bb",
           394 => x"83",
           395 => x"a4",
           396 => x"90",
           397 => x"a4",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"82",
           403 => x"82",
           404 => x"82",
           405 => x"bc",
           406 => x"bb",
           407 => x"e0",
           408 => x"bb",
           409 => x"b2",
           410 => x"a4",
           411 => x"90",
           412 => x"a4",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"82",
           418 => x"82",
           419 => x"82",
           420 => x"96",
           421 => x"bb",
           422 => x"e0",
           423 => x"bb",
           424 => x"cb",
           425 => x"a4",
           426 => x"90",
           427 => x"a4",
           428 => x"9f",
           429 => x"a4",
           430 => x"90",
           431 => x"a4",
           432 => x"fd",
           433 => x"a4",
           434 => x"90",
           435 => x"a4",
           436 => x"b9",
           437 => x"a4",
           438 => x"90",
           439 => x"a4",
           440 => x"b1",
           441 => x"a4",
           442 => x"90",
           443 => x"a4",
           444 => x"e4",
           445 => x"a4",
           446 => x"90",
           447 => x"a4",
           448 => x"84",
           449 => x"a4",
           450 => x"90",
           451 => x"a4",
           452 => x"f5",
           453 => x"a4",
           454 => x"90",
           455 => x"a4",
           456 => x"e9",
           457 => x"a4",
           458 => x"90",
           459 => x"a4",
           460 => x"e6",
           461 => x"a4",
           462 => x"90",
           463 => x"a4",
           464 => x"84",
           465 => x"a4",
           466 => x"90",
           467 => x"a4",
           468 => x"e4",
           469 => x"a4",
           470 => x"90",
           471 => x"a4",
           472 => x"d7",
           473 => x"a4",
           474 => x"90",
           475 => x"a4",
           476 => x"a3",
           477 => x"a4",
           478 => x"90",
           479 => x"a4",
           480 => x"c2",
           481 => x"a4",
           482 => x"90",
           483 => x"a4",
           484 => x"e1",
           485 => x"a4",
           486 => x"90",
           487 => x"a4",
           488 => x"cb",
           489 => x"a4",
           490 => x"90",
           491 => x"a4",
           492 => x"b1",
           493 => x"a4",
           494 => x"90",
           495 => x"a4",
           496 => x"9f",
           497 => x"a4",
           498 => x"90",
           499 => x"a4",
           500 => x"e5",
           501 => x"a4",
           502 => x"90",
           503 => x"a4",
           504 => x"9f",
           505 => x"a4",
           506 => x"90",
           507 => x"a4",
           508 => x"a0",
           509 => x"a4",
           510 => x"90",
           511 => x"a4",
           512 => x"d5",
           513 => x"a4",
           514 => x"90",
           515 => x"a4",
           516 => x"ae",
           517 => x"a4",
           518 => x"90",
           519 => x"a4",
           520 => x"d9",
           521 => x"a4",
           522 => x"90",
           523 => x"a4",
           524 => x"bc",
           525 => x"a4",
           526 => x"90",
           527 => x"a4",
           528 => x"91",
           529 => x"a4",
           530 => x"90",
           531 => x"a4",
           532 => x"9b",
           533 => x"a4",
           534 => x"90",
           535 => x"a4",
           536 => x"dd",
           537 => x"a4",
           538 => x"90",
           539 => x"a4",
           540 => x"a3",
           541 => x"a4",
           542 => x"90",
           543 => x"a4",
           544 => x"c9",
           545 => x"a4",
           546 => x"90",
           547 => x"a4",
           548 => x"fe",
           549 => x"a4",
           550 => x"90",
           551 => x"a4",
           552 => x"ea",
           553 => x"a4",
           554 => x"90",
           555 => x"a4",
           556 => x"de",
           557 => x"a4",
           558 => x"90",
           559 => x"a4",
           560 => x"c8",
           561 => x"a4",
           562 => x"90",
           563 => x"a4",
           564 => x"ac",
           565 => x"a4",
           566 => x"90",
           567 => x"a4",
           568 => x"e2",
           569 => x"a4",
           570 => x"90",
           571 => x"a4",
           572 => x"86",
           573 => x"a4",
           574 => x"90",
           575 => x"a4",
           576 => x"ea",
           577 => x"a4",
           578 => x"90",
           579 => x"a4",
           580 => x"96",
           581 => x"a4",
           582 => x"90",
           583 => x"a4",
           584 => x"f2",
           585 => x"a4",
           586 => x"90",
           587 => x"a4",
           588 => x"9a",
           589 => x"a4",
           590 => x"90",
           591 => x"a4",
           592 => x"92",
           593 => x"a4",
           594 => x"90",
           595 => x"a4",
           596 => x"dc",
           597 => x"a4",
           598 => x"90",
           599 => x"00",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"00",
           609 => x"ff",
           610 => x"06",
           611 => x"83",
           612 => x"10",
           613 => x"fc",
           614 => x"51",
           615 => x"80",
           616 => x"ff",
           617 => x"06",
           618 => x"52",
           619 => x"0a",
           620 => x"38",
           621 => x"51",
           622 => x"98",
           623 => x"f4",
           624 => x"80",
           625 => x"05",
           626 => x"0b",
           627 => x"04",
           628 => x"80",
           629 => x"00",
           630 => x"08",
           631 => x"a4",
           632 => x"0d",
           633 => x"08",
           634 => x"82",
           635 => x"fc",
           636 => x"bb",
           637 => x"05",
           638 => x"bb",
           639 => x"05",
           640 => x"d2",
           641 => x"54",
           642 => x"82",
           643 => x"70",
           644 => x"08",
           645 => x"82",
           646 => x"f8",
           647 => x"82",
           648 => x"51",
           649 => x"0d",
           650 => x"0c",
           651 => x"a4",
           652 => x"bb",
           653 => x"3d",
           654 => x"a4",
           655 => x"08",
           656 => x"70",
           657 => x"81",
           658 => x"51",
           659 => x"38",
           660 => x"bb",
           661 => x"05",
           662 => x"38",
           663 => x"0b",
           664 => x"08",
           665 => x"81",
           666 => x"bb",
           667 => x"05",
           668 => x"82",
           669 => x"8c",
           670 => x"0b",
           671 => x"08",
           672 => x"82",
           673 => x"88",
           674 => x"bb",
           675 => x"05",
           676 => x"a4",
           677 => x"08",
           678 => x"f6",
           679 => x"82",
           680 => x"8c",
           681 => x"80",
           682 => x"bb",
           683 => x"05",
           684 => x"b2",
           685 => x"98",
           686 => x"bb",
           687 => x"05",
           688 => x"bb",
           689 => x"05",
           690 => x"09",
           691 => x"38",
           692 => x"bb",
           693 => x"05",
           694 => x"39",
           695 => x"08",
           696 => x"82",
           697 => x"f8",
           698 => x"53",
           699 => x"82",
           700 => x"8c",
           701 => x"05",
           702 => x"08",
           703 => x"82",
           704 => x"fc",
           705 => x"05",
           706 => x"08",
           707 => x"ff",
           708 => x"bb",
           709 => x"05",
           710 => x"72",
           711 => x"a4",
           712 => x"08",
           713 => x"a4",
           714 => x"0c",
           715 => x"a4",
           716 => x"08",
           717 => x"0c",
           718 => x"82",
           719 => x"04",
           720 => x"08",
           721 => x"a4",
           722 => x"0d",
           723 => x"bb",
           724 => x"05",
           725 => x"a4",
           726 => x"08",
           727 => x"08",
           728 => x"fe",
           729 => x"bb",
           730 => x"05",
           731 => x"a4",
           732 => x"70",
           733 => x"08",
           734 => x"82",
           735 => x"fc",
           736 => x"82",
           737 => x"8c",
           738 => x"82",
           739 => x"e0",
           740 => x"51",
           741 => x"3f",
           742 => x"08",
           743 => x"a4",
           744 => x"0c",
           745 => x"08",
           746 => x"82",
           747 => x"88",
           748 => x"51",
           749 => x"34",
           750 => x"08",
           751 => x"70",
           752 => x"0c",
           753 => x"0d",
           754 => x"0c",
           755 => x"a4",
           756 => x"bb",
           757 => x"3d",
           758 => x"a4",
           759 => x"70",
           760 => x"08",
           761 => x"82",
           762 => x"fc",
           763 => x"82",
           764 => x"8c",
           765 => x"82",
           766 => x"88",
           767 => x"54",
           768 => x"bb",
           769 => x"82",
           770 => x"f8",
           771 => x"bb",
           772 => x"05",
           773 => x"bb",
           774 => x"54",
           775 => x"82",
           776 => x"04",
           777 => x"08",
           778 => x"a4",
           779 => x"0d",
           780 => x"bb",
           781 => x"05",
           782 => x"a4",
           783 => x"08",
           784 => x"8c",
           785 => x"bb",
           786 => x"05",
           787 => x"33",
           788 => x"70",
           789 => x"81",
           790 => x"51",
           791 => x"80",
           792 => x"ff",
           793 => x"a4",
           794 => x"0c",
           795 => x"82",
           796 => x"8c",
           797 => x"72",
           798 => x"82",
           799 => x"f8",
           800 => x"81",
           801 => x"72",
           802 => x"fa",
           803 => x"a4",
           804 => x"08",
           805 => x"bb",
           806 => x"05",
           807 => x"a4",
           808 => x"22",
           809 => x"51",
           810 => x"2e",
           811 => x"82",
           812 => x"f8",
           813 => x"af",
           814 => x"fc",
           815 => x"a4",
           816 => x"33",
           817 => x"26",
           818 => x"82",
           819 => x"f8",
           820 => x"72",
           821 => x"81",
           822 => x"38",
           823 => x"08",
           824 => x"70",
           825 => x"98",
           826 => x"53",
           827 => x"82",
           828 => x"e4",
           829 => x"83",
           830 => x"32",
           831 => x"51",
           832 => x"72",
           833 => x"38",
           834 => x"08",
           835 => x"70",
           836 => x"51",
           837 => x"bb",
           838 => x"05",
           839 => x"39",
           840 => x"08",
           841 => x"70",
           842 => x"98",
           843 => x"83",
           844 => x"73",
           845 => x"51",
           846 => x"53",
           847 => x"a4",
           848 => x"34",
           849 => x"08",
           850 => x"54",
           851 => x"08",
           852 => x"70",
           853 => x"51",
           854 => x"82",
           855 => x"e8",
           856 => x"bb",
           857 => x"05",
           858 => x"2b",
           859 => x"51",
           860 => x"80",
           861 => x"80",
           862 => x"bb",
           863 => x"05",
           864 => x"a4",
           865 => x"22",
           866 => x"70",
           867 => x"51",
           868 => x"db",
           869 => x"a4",
           870 => x"33",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"bb",
           876 => x"05",
           877 => x"39",
           878 => x"08",
           879 => x"70",
           880 => x"81",
           881 => x"53",
           882 => x"9d",
           883 => x"a4",
           884 => x"33",
           885 => x"70",
           886 => x"51",
           887 => x"38",
           888 => x"bb",
           889 => x"05",
           890 => x"a4",
           891 => x"33",
           892 => x"bb",
           893 => x"05",
           894 => x"bb",
           895 => x"05",
           896 => x"26",
           897 => x"82",
           898 => x"c4",
           899 => x"82",
           900 => x"ec",
           901 => x"51",
           902 => x"72",
           903 => x"a4",
           904 => x"22",
           905 => x"51",
           906 => x"bb",
           907 => x"05",
           908 => x"a4",
           909 => x"22",
           910 => x"51",
           911 => x"bb",
           912 => x"05",
           913 => x"39",
           914 => x"08",
           915 => x"70",
           916 => x"51",
           917 => x"bb",
           918 => x"05",
           919 => x"39",
           920 => x"08",
           921 => x"70",
           922 => x"51",
           923 => x"bb",
           924 => x"05",
           925 => x"39",
           926 => x"08",
           927 => x"70",
           928 => x"53",
           929 => x"a4",
           930 => x"23",
           931 => x"bb",
           932 => x"05",
           933 => x"39",
           934 => x"08",
           935 => x"70",
           936 => x"53",
           937 => x"a4",
           938 => x"23",
           939 => x"bf",
           940 => x"a4",
           941 => x"34",
           942 => x"08",
           943 => x"ff",
           944 => x"72",
           945 => x"08",
           946 => x"80",
           947 => x"bb",
           948 => x"05",
           949 => x"39",
           950 => x"08",
           951 => x"82",
           952 => x"90",
           953 => x"05",
           954 => x"08",
           955 => x"70",
           956 => x"72",
           957 => x"08",
           958 => x"82",
           959 => x"ec",
           960 => x"11",
           961 => x"82",
           962 => x"ec",
           963 => x"ef",
           964 => x"a4",
           965 => x"08",
           966 => x"08",
           967 => x"84",
           968 => x"a4",
           969 => x"0c",
           970 => x"bb",
           971 => x"05",
           972 => x"a4",
           973 => x"22",
           974 => x"70",
           975 => x"51",
           976 => x"80",
           977 => x"82",
           978 => x"e8",
           979 => x"98",
           980 => x"98",
           981 => x"bb",
           982 => x"05",
           983 => x"ad",
           984 => x"bb",
           985 => x"72",
           986 => x"08",
           987 => x"99",
           988 => x"a4",
           989 => x"08",
           990 => x"3f",
           991 => x"08",
           992 => x"bb",
           993 => x"05",
           994 => x"a4",
           995 => x"22",
           996 => x"a4",
           997 => x"22",
           998 => x"54",
           999 => x"bb",
          1000 => x"05",
          1001 => x"39",
          1002 => x"08",
          1003 => x"82",
          1004 => x"90",
          1005 => x"05",
          1006 => x"08",
          1007 => x"70",
          1008 => x"a4",
          1009 => x"0c",
          1010 => x"08",
          1011 => x"70",
          1012 => x"81",
          1013 => x"51",
          1014 => x"2e",
          1015 => x"bb",
          1016 => x"05",
          1017 => x"2b",
          1018 => x"2c",
          1019 => x"a4",
          1020 => x"08",
          1021 => x"e3",
          1022 => x"98",
          1023 => x"82",
          1024 => x"f4",
          1025 => x"39",
          1026 => x"08",
          1027 => x"51",
          1028 => x"82",
          1029 => x"53",
          1030 => x"a4",
          1031 => x"23",
          1032 => x"08",
          1033 => x"53",
          1034 => x"08",
          1035 => x"73",
          1036 => x"54",
          1037 => x"a4",
          1038 => x"23",
          1039 => x"82",
          1040 => x"e4",
          1041 => x"82",
          1042 => x"06",
          1043 => x"72",
          1044 => x"38",
          1045 => x"08",
          1046 => x"82",
          1047 => x"90",
          1048 => x"05",
          1049 => x"08",
          1050 => x"70",
          1051 => x"a4",
          1052 => x"0c",
          1053 => x"82",
          1054 => x"90",
          1055 => x"bb",
          1056 => x"05",
          1057 => x"82",
          1058 => x"90",
          1059 => x"08",
          1060 => x"08",
          1061 => x"53",
          1062 => x"08",
          1063 => x"82",
          1064 => x"fc",
          1065 => x"bb",
          1066 => x"05",
          1067 => x"a4",
          1068 => x"a4",
          1069 => x"22",
          1070 => x"51",
          1071 => x"bb",
          1072 => x"05",
          1073 => x"a4",
          1074 => x"08",
          1075 => x"a4",
          1076 => x"0c",
          1077 => x"08",
          1078 => x"70",
          1079 => x"51",
          1080 => x"bb",
          1081 => x"05",
          1082 => x"39",
          1083 => x"bb",
          1084 => x"05",
          1085 => x"82",
          1086 => x"e4",
          1087 => x"80",
          1088 => x"53",
          1089 => x"a4",
          1090 => x"23",
          1091 => x"82",
          1092 => x"f8",
          1093 => x"0b",
          1094 => x"08",
          1095 => x"82",
          1096 => x"e4",
          1097 => x"82",
          1098 => x"06",
          1099 => x"72",
          1100 => x"38",
          1101 => x"08",
          1102 => x"82",
          1103 => x"90",
          1104 => x"05",
          1105 => x"08",
          1106 => x"70",
          1107 => x"a4",
          1108 => x"0c",
          1109 => x"82",
          1110 => x"90",
          1111 => x"bb",
          1112 => x"05",
          1113 => x"82",
          1114 => x"90",
          1115 => x"08",
          1116 => x"08",
          1117 => x"53",
          1118 => x"08",
          1119 => x"82",
          1120 => x"fc",
          1121 => x"bb",
          1122 => x"05",
          1123 => x"06",
          1124 => x"82",
          1125 => x"e4",
          1126 => x"bb",
          1127 => x"bb",
          1128 => x"05",
          1129 => x"a4",
          1130 => x"08",
          1131 => x"08",
          1132 => x"82",
          1133 => x"fc",
          1134 => x"55",
          1135 => x"54",
          1136 => x"3f",
          1137 => x"08",
          1138 => x"34",
          1139 => x"08",
          1140 => x"82",
          1141 => x"d4",
          1142 => x"bb",
          1143 => x"05",
          1144 => x"51",
          1145 => x"27",
          1146 => x"bb",
          1147 => x"05",
          1148 => x"33",
          1149 => x"a4",
          1150 => x"33",
          1151 => x"11",
          1152 => x"72",
          1153 => x"08",
          1154 => x"97",
          1155 => x"a4",
          1156 => x"08",
          1157 => x"b0",
          1158 => x"72",
          1159 => x"08",
          1160 => x"82",
          1161 => x"d4",
          1162 => x"82",
          1163 => x"d0",
          1164 => x"34",
          1165 => x"08",
          1166 => x"81",
          1167 => x"a4",
          1168 => x"0c",
          1169 => x"08",
          1170 => x"70",
          1171 => x"a4",
          1172 => x"08",
          1173 => x"cd",
          1174 => x"98",
          1175 => x"bb",
          1176 => x"05",
          1177 => x"bb",
          1178 => x"05",
          1179 => x"84",
          1180 => x"39",
          1181 => x"08",
          1182 => x"82",
          1183 => x"55",
          1184 => x"70",
          1185 => x"53",
          1186 => x"a4",
          1187 => x"34",
          1188 => x"08",
          1189 => x"70",
          1190 => x"53",
          1191 => x"94",
          1192 => x"a4",
          1193 => x"22",
          1194 => x"53",
          1195 => x"a4",
          1196 => x"23",
          1197 => x"08",
          1198 => x"70",
          1199 => x"81",
          1200 => x"53",
          1201 => x"80",
          1202 => x"bb",
          1203 => x"05",
          1204 => x"2b",
          1205 => x"08",
          1206 => x"82",
          1207 => x"cc",
          1208 => x"2c",
          1209 => x"08",
          1210 => x"82",
          1211 => x"f4",
          1212 => x"53",
          1213 => x"09",
          1214 => x"38",
          1215 => x"08",
          1216 => x"fe",
          1217 => x"82",
          1218 => x"c8",
          1219 => x"39",
          1220 => x"08",
          1221 => x"ff",
          1222 => x"82",
          1223 => x"c8",
          1224 => x"bb",
          1225 => x"05",
          1226 => x"a4",
          1227 => x"23",
          1228 => x"08",
          1229 => x"70",
          1230 => x"81",
          1231 => x"53",
          1232 => x"80",
          1233 => x"bb",
          1234 => x"05",
          1235 => x"2b",
          1236 => x"82",
          1237 => x"fc",
          1238 => x"51",
          1239 => x"74",
          1240 => x"82",
          1241 => x"e4",
          1242 => x"f7",
          1243 => x"72",
          1244 => x"08",
          1245 => x"9d",
          1246 => x"a4",
          1247 => x"33",
          1248 => x"a4",
          1249 => x"33",
          1250 => x"54",
          1251 => x"bb",
          1252 => x"05",
          1253 => x"a4",
          1254 => x"22",
          1255 => x"70",
          1256 => x"51",
          1257 => x"2e",
          1258 => x"bb",
          1259 => x"05",
          1260 => x"2b",
          1261 => x"70",
          1262 => x"88",
          1263 => x"51",
          1264 => x"54",
          1265 => x"08",
          1266 => x"70",
          1267 => x"53",
          1268 => x"a4",
          1269 => x"23",
          1270 => x"bb",
          1271 => x"05",
          1272 => x"2b",
          1273 => x"70",
          1274 => x"88",
          1275 => x"51",
          1276 => x"54",
          1277 => x"08",
          1278 => x"70",
          1279 => x"53",
          1280 => x"a4",
          1281 => x"23",
          1282 => x"08",
          1283 => x"70",
          1284 => x"51",
          1285 => x"38",
          1286 => x"08",
          1287 => x"ff",
          1288 => x"72",
          1289 => x"08",
          1290 => x"73",
          1291 => x"90",
          1292 => x"80",
          1293 => x"38",
          1294 => x"08",
          1295 => x"52",
          1296 => x"90",
          1297 => x"82",
          1298 => x"e4",
          1299 => x"81",
          1300 => x"06",
          1301 => x"72",
          1302 => x"38",
          1303 => x"08",
          1304 => x"52",
          1305 => x"ec",
          1306 => x"39",
          1307 => x"08",
          1308 => x"70",
          1309 => x"81",
          1310 => x"53",
          1311 => x"90",
          1312 => x"a4",
          1313 => x"08",
          1314 => x"95",
          1315 => x"39",
          1316 => x"08",
          1317 => x"70",
          1318 => x"81",
          1319 => x"53",
          1320 => x"8e",
          1321 => x"a4",
          1322 => x"08",
          1323 => x"95",
          1324 => x"bb",
          1325 => x"05",
          1326 => x"2a",
          1327 => x"51",
          1328 => x"80",
          1329 => x"82",
          1330 => x"88",
          1331 => x"b0",
          1332 => x"3f",
          1333 => x"08",
          1334 => x"53",
          1335 => x"09",
          1336 => x"38",
          1337 => x"08",
          1338 => x"52",
          1339 => x"08",
          1340 => x"51",
          1341 => x"82",
          1342 => x"e4",
          1343 => x"88",
          1344 => x"06",
          1345 => x"72",
          1346 => x"38",
          1347 => x"08",
          1348 => x"ff",
          1349 => x"72",
          1350 => x"08",
          1351 => x"73",
          1352 => x"90",
          1353 => x"80",
          1354 => x"38",
          1355 => x"08",
          1356 => x"52",
          1357 => x"9c",
          1358 => x"82",
          1359 => x"e4",
          1360 => x"83",
          1361 => x"06",
          1362 => x"72",
          1363 => x"38",
          1364 => x"08",
          1365 => x"ff",
          1366 => x"72",
          1367 => x"08",
          1368 => x"73",
          1369 => x"98",
          1370 => x"80",
          1371 => x"38",
          1372 => x"08",
          1373 => x"52",
          1374 => x"d8",
          1375 => x"82",
          1376 => x"e4",
          1377 => x"87",
          1378 => x"06",
          1379 => x"72",
          1380 => x"bb",
          1381 => x"05",
          1382 => x"54",
          1383 => x"bb",
          1384 => x"05",
          1385 => x"2b",
          1386 => x"51",
          1387 => x"25",
          1388 => x"bb",
          1389 => x"05",
          1390 => x"51",
          1391 => x"d2",
          1392 => x"a4",
          1393 => x"33",
          1394 => x"e3",
          1395 => x"06",
          1396 => x"bb",
          1397 => x"05",
          1398 => x"bb",
          1399 => x"05",
          1400 => x"f0",
          1401 => x"39",
          1402 => x"08",
          1403 => x"53",
          1404 => x"2e",
          1405 => x"80",
          1406 => x"bb",
          1407 => x"05",
          1408 => x"51",
          1409 => x"bb",
          1410 => x"05",
          1411 => x"ff",
          1412 => x"72",
          1413 => x"2e",
          1414 => x"82",
          1415 => x"88",
          1416 => x"82",
          1417 => x"fc",
          1418 => x"33",
          1419 => x"a4",
          1420 => x"08",
          1421 => x"bb",
          1422 => x"05",
          1423 => x"94",
          1424 => x"39",
          1425 => x"08",
          1426 => x"53",
          1427 => x"2e",
          1428 => x"80",
          1429 => x"bb",
          1430 => x"05",
          1431 => x"51",
          1432 => x"bb",
          1433 => x"05",
          1434 => x"ff",
          1435 => x"72",
          1436 => x"2e",
          1437 => x"82",
          1438 => x"88",
          1439 => x"82",
          1440 => x"fc",
          1441 => x"33",
          1442 => x"c8",
          1443 => x"a4",
          1444 => x"08",
          1445 => x"bb",
          1446 => x"05",
          1447 => x"39",
          1448 => x"08",
          1449 => x"82",
          1450 => x"a9",
          1451 => x"a4",
          1452 => x"08",
          1453 => x"a4",
          1454 => x"08",
          1455 => x"bb",
          1456 => x"05",
          1457 => x"a4",
          1458 => x"08",
          1459 => x"53",
          1460 => x"cc",
          1461 => x"a4",
          1462 => x"22",
          1463 => x"70",
          1464 => x"51",
          1465 => x"2e",
          1466 => x"82",
          1467 => x"ec",
          1468 => x"11",
          1469 => x"82",
          1470 => x"ec",
          1471 => x"90",
          1472 => x"2c",
          1473 => x"73",
          1474 => x"82",
          1475 => x"88",
          1476 => x"a0",
          1477 => x"3f",
          1478 => x"bb",
          1479 => x"05",
          1480 => x"bb",
          1481 => x"05",
          1482 => x"a8",
          1483 => x"82",
          1484 => x"e4",
          1485 => x"b7",
          1486 => x"a4",
          1487 => x"33",
          1488 => x"2e",
          1489 => x"a8",
          1490 => x"82",
          1491 => x"e4",
          1492 => x"0b",
          1493 => x"08",
          1494 => x"80",
          1495 => x"a4",
          1496 => x"34",
          1497 => x"bb",
          1498 => x"05",
          1499 => x"39",
          1500 => x"08",
          1501 => x"52",
          1502 => x"08",
          1503 => x"51",
          1504 => x"e9",
          1505 => x"bb",
          1506 => x"05",
          1507 => x"08",
          1508 => x"a4",
          1509 => x"0c",
          1510 => x"bb",
          1511 => x"05",
          1512 => x"98",
          1513 => x"0d",
          1514 => x"0c",
          1515 => x"a4",
          1516 => x"bb",
          1517 => x"3d",
          1518 => x"82",
          1519 => x"f0",
          1520 => x"bb",
          1521 => x"05",
          1522 => x"73",
          1523 => x"a4",
          1524 => x"08",
          1525 => x"53",
          1526 => x"72",
          1527 => x"08",
          1528 => x"72",
          1529 => x"53",
          1530 => x"09",
          1531 => x"38",
          1532 => x"08",
          1533 => x"70",
          1534 => x"71",
          1535 => x"39",
          1536 => x"08",
          1537 => x"53",
          1538 => x"09",
          1539 => x"38",
          1540 => x"bb",
          1541 => x"05",
          1542 => x"a4",
          1543 => x"08",
          1544 => x"05",
          1545 => x"08",
          1546 => x"33",
          1547 => x"08",
          1548 => x"82",
          1549 => x"f8",
          1550 => x"72",
          1551 => x"81",
          1552 => x"38",
          1553 => x"08",
          1554 => x"70",
          1555 => x"71",
          1556 => x"51",
          1557 => x"82",
          1558 => x"f8",
          1559 => x"bb",
          1560 => x"05",
          1561 => x"a4",
          1562 => x"0c",
          1563 => x"08",
          1564 => x"80",
          1565 => x"38",
          1566 => x"08",
          1567 => x"80",
          1568 => x"38",
          1569 => x"90",
          1570 => x"a4",
          1571 => x"34",
          1572 => x"08",
          1573 => x"70",
          1574 => x"71",
          1575 => x"51",
          1576 => x"82",
          1577 => x"f8",
          1578 => x"a4",
          1579 => x"82",
          1580 => x"f4",
          1581 => x"bb",
          1582 => x"05",
          1583 => x"81",
          1584 => x"70",
          1585 => x"72",
          1586 => x"a4",
          1587 => x"34",
          1588 => x"82",
          1589 => x"f8",
          1590 => x"72",
          1591 => x"38",
          1592 => x"bb",
          1593 => x"05",
          1594 => x"39",
          1595 => x"08",
          1596 => x"53",
          1597 => x"90",
          1598 => x"a4",
          1599 => x"33",
          1600 => x"26",
          1601 => x"39",
          1602 => x"bb",
          1603 => x"05",
          1604 => x"39",
          1605 => x"bb",
          1606 => x"05",
          1607 => x"82",
          1608 => x"f8",
          1609 => x"af",
          1610 => x"38",
          1611 => x"08",
          1612 => x"53",
          1613 => x"83",
          1614 => x"80",
          1615 => x"a4",
          1616 => x"0c",
          1617 => x"8a",
          1618 => x"a4",
          1619 => x"34",
          1620 => x"bb",
          1621 => x"05",
          1622 => x"a4",
          1623 => x"33",
          1624 => x"27",
          1625 => x"82",
          1626 => x"f8",
          1627 => x"80",
          1628 => x"94",
          1629 => x"a4",
          1630 => x"33",
          1631 => x"53",
          1632 => x"a4",
          1633 => x"34",
          1634 => x"08",
          1635 => x"d0",
          1636 => x"72",
          1637 => x"08",
          1638 => x"82",
          1639 => x"f8",
          1640 => x"90",
          1641 => x"38",
          1642 => x"08",
          1643 => x"f9",
          1644 => x"72",
          1645 => x"08",
          1646 => x"82",
          1647 => x"f8",
          1648 => x"72",
          1649 => x"38",
          1650 => x"bb",
          1651 => x"05",
          1652 => x"39",
          1653 => x"08",
          1654 => x"82",
          1655 => x"f4",
          1656 => x"54",
          1657 => x"8d",
          1658 => x"82",
          1659 => x"ec",
          1660 => x"f7",
          1661 => x"a4",
          1662 => x"33",
          1663 => x"a4",
          1664 => x"08",
          1665 => x"a4",
          1666 => x"33",
          1667 => x"bb",
          1668 => x"05",
          1669 => x"a4",
          1670 => x"08",
          1671 => x"05",
          1672 => x"08",
          1673 => x"55",
          1674 => x"82",
          1675 => x"f8",
          1676 => x"a5",
          1677 => x"a4",
          1678 => x"33",
          1679 => x"2e",
          1680 => x"bb",
          1681 => x"05",
          1682 => x"bb",
          1683 => x"05",
          1684 => x"a4",
          1685 => x"08",
          1686 => x"08",
          1687 => x"71",
          1688 => x"0b",
          1689 => x"08",
          1690 => x"82",
          1691 => x"ec",
          1692 => x"bb",
          1693 => x"3d",
          1694 => x"a4",
          1695 => x"bb",
          1696 => x"82",
          1697 => x"fd",
          1698 => x"d2",
          1699 => x"82",
          1700 => x"8c",
          1701 => x"82",
          1702 => x"88",
          1703 => x"df",
          1704 => x"bb",
          1705 => x"82",
          1706 => x"54",
          1707 => x"82",
          1708 => x"04",
          1709 => x"08",
          1710 => x"a4",
          1711 => x"0d",
          1712 => x"bb",
          1713 => x"05",
          1714 => x"a4",
          1715 => x"08",
          1716 => x"0c",
          1717 => x"08",
          1718 => x"70",
          1719 => x"72",
          1720 => x"82",
          1721 => x"f8",
          1722 => x"81",
          1723 => x"72",
          1724 => x"81",
          1725 => x"82",
          1726 => x"88",
          1727 => x"08",
          1728 => x"0c",
          1729 => x"82",
          1730 => x"f8",
          1731 => x"72",
          1732 => x"81",
          1733 => x"81",
          1734 => x"a4",
          1735 => x"34",
          1736 => x"08",
          1737 => x"70",
          1738 => x"71",
          1739 => x"51",
          1740 => x"82",
          1741 => x"f8",
          1742 => x"bb",
          1743 => x"05",
          1744 => x"b0",
          1745 => x"06",
          1746 => x"82",
          1747 => x"88",
          1748 => x"08",
          1749 => x"0c",
          1750 => x"53",
          1751 => x"bb",
          1752 => x"05",
          1753 => x"a4",
          1754 => x"33",
          1755 => x"08",
          1756 => x"82",
          1757 => x"e8",
          1758 => x"e2",
          1759 => x"82",
          1760 => x"e8",
          1761 => x"f8",
          1762 => x"80",
          1763 => x"0b",
          1764 => x"08",
          1765 => x"82",
          1766 => x"88",
          1767 => x"08",
          1768 => x"0c",
          1769 => x"53",
          1770 => x"bb",
          1771 => x"05",
          1772 => x"39",
          1773 => x"bb",
          1774 => x"05",
          1775 => x"a4",
          1776 => x"08",
          1777 => x"05",
          1778 => x"08",
          1779 => x"33",
          1780 => x"08",
          1781 => x"80",
          1782 => x"bb",
          1783 => x"05",
          1784 => x"a0",
          1785 => x"81",
          1786 => x"a4",
          1787 => x"0c",
          1788 => x"82",
          1789 => x"f8",
          1790 => x"af",
          1791 => x"38",
          1792 => x"08",
          1793 => x"53",
          1794 => x"83",
          1795 => x"80",
          1796 => x"a4",
          1797 => x"0c",
          1798 => x"88",
          1799 => x"a4",
          1800 => x"34",
          1801 => x"bb",
          1802 => x"05",
          1803 => x"73",
          1804 => x"82",
          1805 => x"f8",
          1806 => x"72",
          1807 => x"38",
          1808 => x"0b",
          1809 => x"08",
          1810 => x"82",
          1811 => x"0b",
          1812 => x"08",
          1813 => x"80",
          1814 => x"a4",
          1815 => x"0c",
          1816 => x"08",
          1817 => x"53",
          1818 => x"81",
          1819 => x"bb",
          1820 => x"05",
          1821 => x"e0",
          1822 => x"38",
          1823 => x"08",
          1824 => x"e0",
          1825 => x"72",
          1826 => x"08",
          1827 => x"82",
          1828 => x"f8",
          1829 => x"11",
          1830 => x"82",
          1831 => x"f8",
          1832 => x"bb",
          1833 => x"05",
          1834 => x"73",
          1835 => x"82",
          1836 => x"f8",
          1837 => x"11",
          1838 => x"82",
          1839 => x"f8",
          1840 => x"bb",
          1841 => x"05",
          1842 => x"89",
          1843 => x"80",
          1844 => x"a4",
          1845 => x"0c",
          1846 => x"82",
          1847 => x"f8",
          1848 => x"bb",
          1849 => x"05",
          1850 => x"72",
          1851 => x"38",
          1852 => x"bb",
          1853 => x"05",
          1854 => x"39",
          1855 => x"08",
          1856 => x"70",
          1857 => x"08",
          1858 => x"29",
          1859 => x"08",
          1860 => x"70",
          1861 => x"a4",
          1862 => x"0c",
          1863 => x"08",
          1864 => x"70",
          1865 => x"71",
          1866 => x"51",
          1867 => x"53",
          1868 => x"bb",
          1869 => x"05",
          1870 => x"39",
          1871 => x"08",
          1872 => x"53",
          1873 => x"90",
          1874 => x"a4",
          1875 => x"08",
          1876 => x"a4",
          1877 => x"0c",
          1878 => x"08",
          1879 => x"82",
          1880 => x"fc",
          1881 => x"0c",
          1882 => x"82",
          1883 => x"ec",
          1884 => x"bb",
          1885 => x"05",
          1886 => x"98",
          1887 => x"0d",
          1888 => x"0c",
          1889 => x"a4",
          1890 => x"bb",
          1891 => x"3d",
          1892 => x"82",
          1893 => x"f8",
          1894 => x"d2",
          1895 => x"11",
          1896 => x"2a",
          1897 => x"70",
          1898 => x"51",
          1899 => x"72",
          1900 => x"38",
          1901 => x"bb",
          1902 => x"05",
          1903 => x"39",
          1904 => x"08",
          1905 => x"53",
          1906 => x"bb",
          1907 => x"05",
          1908 => x"82",
          1909 => x"88",
          1910 => x"72",
          1911 => x"08",
          1912 => x"72",
          1913 => x"53",
          1914 => x"b0",
          1915 => x"ec",
          1916 => x"ec",
          1917 => x"bb",
          1918 => x"05",
          1919 => x"11",
          1920 => x"72",
          1921 => x"98",
          1922 => x"80",
          1923 => x"38",
          1924 => x"bb",
          1925 => x"05",
          1926 => x"39",
          1927 => x"08",
          1928 => x"08",
          1929 => x"51",
          1930 => x"53",
          1931 => x"bb",
          1932 => x"72",
          1933 => x"38",
          1934 => x"bb",
          1935 => x"05",
          1936 => x"a4",
          1937 => x"08",
          1938 => x"a4",
          1939 => x"0c",
          1940 => x"a4",
          1941 => x"08",
          1942 => x"0c",
          1943 => x"82",
          1944 => x"04",
          1945 => x"08",
          1946 => x"a4",
          1947 => x"0d",
          1948 => x"bb",
          1949 => x"05",
          1950 => x"a4",
          1951 => x"08",
          1952 => x"70",
          1953 => x"81",
          1954 => x"06",
          1955 => x"51",
          1956 => x"2e",
          1957 => x"0b",
          1958 => x"08",
          1959 => x"80",
          1960 => x"bb",
          1961 => x"05",
          1962 => x"33",
          1963 => x"08",
          1964 => x"81",
          1965 => x"a4",
          1966 => x"0c",
          1967 => x"bb",
          1968 => x"05",
          1969 => x"ff",
          1970 => x"80",
          1971 => x"82",
          1972 => x"8c",
          1973 => x"bb",
          1974 => x"05",
          1975 => x"bb",
          1976 => x"05",
          1977 => x"11",
          1978 => x"72",
          1979 => x"98",
          1980 => x"80",
          1981 => x"38",
          1982 => x"bb",
          1983 => x"05",
          1984 => x"39",
          1985 => x"08",
          1986 => x"70",
          1987 => x"08",
          1988 => x"53",
          1989 => x"08",
          1990 => x"82",
          1991 => x"87",
          1992 => x"bb",
          1993 => x"82",
          1994 => x"02",
          1995 => x"0c",
          1996 => x"82",
          1997 => x"52",
          1998 => x"08",
          1999 => x"51",
          2000 => x"bb",
          2001 => x"82",
          2002 => x"53",
          2003 => x"82",
          2004 => x"04",
          2005 => x"08",
          2006 => x"a4",
          2007 => x"0d",
          2008 => x"08",
          2009 => x"85",
          2010 => x"81",
          2011 => x"32",
          2012 => x"51",
          2013 => x"53",
          2014 => x"8d",
          2015 => x"82",
          2016 => x"fc",
          2017 => x"cb",
          2018 => x"a4",
          2019 => x"08",
          2020 => x"70",
          2021 => x"81",
          2022 => x"51",
          2023 => x"2e",
          2024 => x"82",
          2025 => x"8c",
          2026 => x"bb",
          2027 => x"05",
          2028 => x"8c",
          2029 => x"14",
          2030 => x"38",
          2031 => x"08",
          2032 => x"70",
          2033 => x"bb",
          2034 => x"05",
          2035 => x"54",
          2036 => x"34",
          2037 => x"05",
          2038 => x"bb",
          2039 => x"05",
          2040 => x"08",
          2041 => x"12",
          2042 => x"a4",
          2043 => x"08",
          2044 => x"a4",
          2045 => x"0c",
          2046 => x"d7",
          2047 => x"a4",
          2048 => x"08",
          2049 => x"08",
          2050 => x"53",
          2051 => x"08",
          2052 => x"70",
          2053 => x"53",
          2054 => x"51",
          2055 => x"2d",
          2056 => x"08",
          2057 => x"38",
          2058 => x"08",
          2059 => x"8c",
          2060 => x"05",
          2061 => x"82",
          2062 => x"88",
          2063 => x"82",
          2064 => x"fc",
          2065 => x"53",
          2066 => x"0b",
          2067 => x"08",
          2068 => x"82",
          2069 => x"fc",
          2070 => x"bb",
          2071 => x"3d",
          2072 => x"a4",
          2073 => x"bb",
          2074 => x"82",
          2075 => x"f9",
          2076 => x"bb",
          2077 => x"05",
          2078 => x"33",
          2079 => x"70",
          2080 => x"51",
          2081 => x"80",
          2082 => x"ff",
          2083 => x"a4",
          2084 => x"0c",
          2085 => x"82",
          2086 => x"88",
          2087 => x"11",
          2088 => x"2a",
          2089 => x"51",
          2090 => x"71",
          2091 => x"c5",
          2092 => x"a4",
          2093 => x"08",
          2094 => x"08",
          2095 => x"53",
          2096 => x"33",
          2097 => x"06",
          2098 => x"85",
          2099 => x"bb",
          2100 => x"05",
          2101 => x"08",
          2102 => x"12",
          2103 => x"a4",
          2104 => x"08",
          2105 => x"70",
          2106 => x"08",
          2107 => x"51",
          2108 => x"b6",
          2109 => x"a4",
          2110 => x"08",
          2111 => x"70",
          2112 => x"81",
          2113 => x"51",
          2114 => x"2e",
          2115 => x"82",
          2116 => x"88",
          2117 => x"08",
          2118 => x"bb",
          2119 => x"05",
          2120 => x"82",
          2121 => x"fc",
          2122 => x"38",
          2123 => x"08",
          2124 => x"82",
          2125 => x"88",
          2126 => x"53",
          2127 => x"70",
          2128 => x"52",
          2129 => x"34",
          2130 => x"bb",
          2131 => x"05",
          2132 => x"39",
          2133 => x"08",
          2134 => x"70",
          2135 => x"71",
          2136 => x"a1",
          2137 => x"a4",
          2138 => x"08",
          2139 => x"08",
          2140 => x"52",
          2141 => x"51",
          2142 => x"82",
          2143 => x"70",
          2144 => x"08",
          2145 => x"52",
          2146 => x"08",
          2147 => x"80",
          2148 => x"38",
          2149 => x"08",
          2150 => x"82",
          2151 => x"f4",
          2152 => x"bb",
          2153 => x"05",
          2154 => x"33",
          2155 => x"08",
          2156 => x"52",
          2157 => x"08",
          2158 => x"ff",
          2159 => x"06",
          2160 => x"bb",
          2161 => x"05",
          2162 => x"52",
          2163 => x"a4",
          2164 => x"34",
          2165 => x"bb",
          2166 => x"05",
          2167 => x"52",
          2168 => x"a4",
          2169 => x"34",
          2170 => x"08",
          2171 => x"52",
          2172 => x"08",
          2173 => x"85",
          2174 => x"0b",
          2175 => x"08",
          2176 => x"a6",
          2177 => x"a4",
          2178 => x"08",
          2179 => x"81",
          2180 => x"0c",
          2181 => x"08",
          2182 => x"70",
          2183 => x"70",
          2184 => x"08",
          2185 => x"51",
          2186 => x"bb",
          2187 => x"05",
          2188 => x"98",
          2189 => x"0d",
          2190 => x"0c",
          2191 => x"a4",
          2192 => x"bb",
          2193 => x"3d",
          2194 => x"a4",
          2195 => x"08",
          2196 => x"08",
          2197 => x"82",
          2198 => x"8c",
          2199 => x"bb",
          2200 => x"05",
          2201 => x"a4",
          2202 => x"08",
          2203 => x"a2",
          2204 => x"a4",
          2205 => x"08",
          2206 => x"08",
          2207 => x"26",
          2208 => x"82",
          2209 => x"f8",
          2210 => x"bb",
          2211 => x"05",
          2212 => x"82",
          2213 => x"fc",
          2214 => x"27",
          2215 => x"82",
          2216 => x"fc",
          2217 => x"bb",
          2218 => x"05",
          2219 => x"bb",
          2220 => x"05",
          2221 => x"a4",
          2222 => x"08",
          2223 => x"08",
          2224 => x"05",
          2225 => x"08",
          2226 => x"82",
          2227 => x"90",
          2228 => x"05",
          2229 => x"08",
          2230 => x"82",
          2231 => x"90",
          2232 => x"05",
          2233 => x"08",
          2234 => x"82",
          2235 => x"90",
          2236 => x"2e",
          2237 => x"82",
          2238 => x"fc",
          2239 => x"05",
          2240 => x"08",
          2241 => x"82",
          2242 => x"f8",
          2243 => x"05",
          2244 => x"08",
          2245 => x"82",
          2246 => x"fc",
          2247 => x"bb",
          2248 => x"05",
          2249 => x"71",
          2250 => x"ff",
          2251 => x"bb",
          2252 => x"05",
          2253 => x"82",
          2254 => x"90",
          2255 => x"bb",
          2256 => x"05",
          2257 => x"82",
          2258 => x"90",
          2259 => x"bb",
          2260 => x"05",
          2261 => x"ba",
          2262 => x"a4",
          2263 => x"08",
          2264 => x"82",
          2265 => x"f8",
          2266 => x"05",
          2267 => x"08",
          2268 => x"82",
          2269 => x"fc",
          2270 => x"52",
          2271 => x"82",
          2272 => x"fc",
          2273 => x"05",
          2274 => x"08",
          2275 => x"ff",
          2276 => x"bb",
          2277 => x"05",
          2278 => x"bb",
          2279 => x"85",
          2280 => x"bb",
          2281 => x"82",
          2282 => x"02",
          2283 => x"0c",
          2284 => x"82",
          2285 => x"88",
          2286 => x"bb",
          2287 => x"05",
          2288 => x"a4",
          2289 => x"08",
          2290 => x"82",
          2291 => x"fc",
          2292 => x"05",
          2293 => x"08",
          2294 => x"70",
          2295 => x"51",
          2296 => x"2e",
          2297 => x"39",
          2298 => x"08",
          2299 => x"ff",
          2300 => x"a4",
          2301 => x"0c",
          2302 => x"08",
          2303 => x"82",
          2304 => x"88",
          2305 => x"70",
          2306 => x"0c",
          2307 => x"0d",
          2308 => x"0c",
          2309 => x"a4",
          2310 => x"bb",
          2311 => x"3d",
          2312 => x"a4",
          2313 => x"08",
          2314 => x"08",
          2315 => x"82",
          2316 => x"8c",
          2317 => x"71",
          2318 => x"a4",
          2319 => x"08",
          2320 => x"bb",
          2321 => x"05",
          2322 => x"a4",
          2323 => x"08",
          2324 => x"72",
          2325 => x"a4",
          2326 => x"08",
          2327 => x"bb",
          2328 => x"05",
          2329 => x"ff",
          2330 => x"80",
          2331 => x"ff",
          2332 => x"bb",
          2333 => x"05",
          2334 => x"bb",
          2335 => x"84",
          2336 => x"bb",
          2337 => x"82",
          2338 => x"02",
          2339 => x"0c",
          2340 => x"82",
          2341 => x"88",
          2342 => x"bb",
          2343 => x"05",
          2344 => x"a4",
          2345 => x"08",
          2346 => x"08",
          2347 => x"82",
          2348 => x"90",
          2349 => x"2e",
          2350 => x"82",
          2351 => x"90",
          2352 => x"05",
          2353 => x"08",
          2354 => x"82",
          2355 => x"90",
          2356 => x"05",
          2357 => x"08",
          2358 => x"82",
          2359 => x"90",
          2360 => x"2e",
          2361 => x"bb",
          2362 => x"05",
          2363 => x"33",
          2364 => x"08",
          2365 => x"81",
          2366 => x"a4",
          2367 => x"0c",
          2368 => x"08",
          2369 => x"52",
          2370 => x"34",
          2371 => x"08",
          2372 => x"81",
          2373 => x"a4",
          2374 => x"0c",
          2375 => x"82",
          2376 => x"88",
          2377 => x"82",
          2378 => x"51",
          2379 => x"82",
          2380 => x"04",
          2381 => x"08",
          2382 => x"a4",
          2383 => x"0d",
          2384 => x"08",
          2385 => x"80",
          2386 => x"38",
          2387 => x"08",
          2388 => x"52",
          2389 => x"bb",
          2390 => x"05",
          2391 => x"82",
          2392 => x"8c",
          2393 => x"bb",
          2394 => x"05",
          2395 => x"72",
          2396 => x"53",
          2397 => x"71",
          2398 => x"38",
          2399 => x"82",
          2400 => x"88",
          2401 => x"71",
          2402 => x"a4",
          2403 => x"08",
          2404 => x"bb",
          2405 => x"05",
          2406 => x"ff",
          2407 => x"70",
          2408 => x"0b",
          2409 => x"08",
          2410 => x"81",
          2411 => x"bb",
          2412 => x"05",
          2413 => x"82",
          2414 => x"90",
          2415 => x"bb",
          2416 => x"05",
          2417 => x"84",
          2418 => x"39",
          2419 => x"08",
          2420 => x"80",
          2421 => x"38",
          2422 => x"08",
          2423 => x"70",
          2424 => x"70",
          2425 => x"0b",
          2426 => x"08",
          2427 => x"80",
          2428 => x"bb",
          2429 => x"05",
          2430 => x"82",
          2431 => x"8c",
          2432 => x"bb",
          2433 => x"05",
          2434 => x"52",
          2435 => x"38",
          2436 => x"bb",
          2437 => x"05",
          2438 => x"82",
          2439 => x"88",
          2440 => x"33",
          2441 => x"08",
          2442 => x"70",
          2443 => x"31",
          2444 => x"a4",
          2445 => x"0c",
          2446 => x"52",
          2447 => x"80",
          2448 => x"a4",
          2449 => x"0c",
          2450 => x"08",
          2451 => x"82",
          2452 => x"85",
          2453 => x"bb",
          2454 => x"82",
          2455 => x"02",
          2456 => x"0c",
          2457 => x"82",
          2458 => x"88",
          2459 => x"bb",
          2460 => x"05",
          2461 => x"a4",
          2462 => x"08",
          2463 => x"0b",
          2464 => x"08",
          2465 => x"80",
          2466 => x"bb",
          2467 => x"05",
          2468 => x"33",
          2469 => x"08",
          2470 => x"81",
          2471 => x"a4",
          2472 => x"0c",
          2473 => x"06",
          2474 => x"80",
          2475 => x"82",
          2476 => x"8c",
          2477 => x"05",
          2478 => x"08",
          2479 => x"82",
          2480 => x"8c",
          2481 => x"2e",
          2482 => x"be",
          2483 => x"a4",
          2484 => x"08",
          2485 => x"bb",
          2486 => x"05",
          2487 => x"a4",
          2488 => x"08",
          2489 => x"08",
          2490 => x"31",
          2491 => x"a4",
          2492 => x"0c",
          2493 => x"a4",
          2494 => x"08",
          2495 => x"0c",
          2496 => x"82",
          2497 => x"04",
          2498 => x"08",
          2499 => x"a4",
          2500 => x"0d",
          2501 => x"08",
          2502 => x"82",
          2503 => x"fc",
          2504 => x"bb",
          2505 => x"05",
          2506 => x"80",
          2507 => x"bb",
          2508 => x"05",
          2509 => x"82",
          2510 => x"90",
          2511 => x"bb",
          2512 => x"05",
          2513 => x"82",
          2514 => x"90",
          2515 => x"bb",
          2516 => x"05",
          2517 => x"a9",
          2518 => x"a4",
          2519 => x"08",
          2520 => x"bb",
          2521 => x"05",
          2522 => x"71",
          2523 => x"bb",
          2524 => x"05",
          2525 => x"82",
          2526 => x"fc",
          2527 => x"be",
          2528 => x"a4",
          2529 => x"08",
          2530 => x"98",
          2531 => x"3d",
          2532 => x"a4",
          2533 => x"bb",
          2534 => x"82",
          2535 => x"f9",
          2536 => x"0b",
          2537 => x"08",
          2538 => x"82",
          2539 => x"88",
          2540 => x"25",
          2541 => x"bb",
          2542 => x"05",
          2543 => x"bb",
          2544 => x"05",
          2545 => x"82",
          2546 => x"f4",
          2547 => x"bb",
          2548 => x"05",
          2549 => x"81",
          2550 => x"a4",
          2551 => x"0c",
          2552 => x"08",
          2553 => x"82",
          2554 => x"fc",
          2555 => x"bb",
          2556 => x"05",
          2557 => x"b9",
          2558 => x"a4",
          2559 => x"08",
          2560 => x"a4",
          2561 => x"0c",
          2562 => x"bb",
          2563 => x"05",
          2564 => x"a4",
          2565 => x"08",
          2566 => x"0b",
          2567 => x"08",
          2568 => x"82",
          2569 => x"f0",
          2570 => x"bb",
          2571 => x"05",
          2572 => x"82",
          2573 => x"8c",
          2574 => x"82",
          2575 => x"88",
          2576 => x"82",
          2577 => x"bb",
          2578 => x"82",
          2579 => x"f8",
          2580 => x"82",
          2581 => x"fc",
          2582 => x"2e",
          2583 => x"bb",
          2584 => x"05",
          2585 => x"bb",
          2586 => x"05",
          2587 => x"a4",
          2588 => x"08",
          2589 => x"98",
          2590 => x"3d",
          2591 => x"a4",
          2592 => x"bb",
          2593 => x"82",
          2594 => x"fb",
          2595 => x"0b",
          2596 => x"08",
          2597 => x"82",
          2598 => x"88",
          2599 => x"25",
          2600 => x"bb",
          2601 => x"05",
          2602 => x"bb",
          2603 => x"05",
          2604 => x"82",
          2605 => x"fc",
          2606 => x"bb",
          2607 => x"05",
          2608 => x"90",
          2609 => x"a4",
          2610 => x"08",
          2611 => x"a4",
          2612 => x"0c",
          2613 => x"bb",
          2614 => x"05",
          2615 => x"bb",
          2616 => x"05",
          2617 => x"a2",
          2618 => x"98",
          2619 => x"bb",
          2620 => x"05",
          2621 => x"bb",
          2622 => x"05",
          2623 => x"90",
          2624 => x"a4",
          2625 => x"08",
          2626 => x"a4",
          2627 => x"0c",
          2628 => x"08",
          2629 => x"70",
          2630 => x"0c",
          2631 => x"0d",
          2632 => x"0c",
          2633 => x"a4",
          2634 => x"bb",
          2635 => x"3d",
          2636 => x"82",
          2637 => x"8c",
          2638 => x"82",
          2639 => x"88",
          2640 => x"80",
          2641 => x"bb",
          2642 => x"82",
          2643 => x"54",
          2644 => x"82",
          2645 => x"04",
          2646 => x"08",
          2647 => x"a4",
          2648 => x"0d",
          2649 => x"bb",
          2650 => x"05",
          2651 => x"bb",
          2652 => x"05",
          2653 => x"3f",
          2654 => x"08",
          2655 => x"98",
          2656 => x"3d",
          2657 => x"a4",
          2658 => x"bb",
          2659 => x"82",
          2660 => x"fd",
          2661 => x"0b",
          2662 => x"08",
          2663 => x"80",
          2664 => x"a4",
          2665 => x"0c",
          2666 => x"08",
          2667 => x"82",
          2668 => x"88",
          2669 => x"b9",
          2670 => x"a4",
          2671 => x"08",
          2672 => x"38",
          2673 => x"bb",
          2674 => x"05",
          2675 => x"38",
          2676 => x"08",
          2677 => x"10",
          2678 => x"08",
          2679 => x"82",
          2680 => x"fc",
          2681 => x"82",
          2682 => x"fc",
          2683 => x"b8",
          2684 => x"a4",
          2685 => x"08",
          2686 => x"e1",
          2687 => x"a4",
          2688 => x"08",
          2689 => x"08",
          2690 => x"26",
          2691 => x"bb",
          2692 => x"05",
          2693 => x"a4",
          2694 => x"08",
          2695 => x"a4",
          2696 => x"0c",
          2697 => x"08",
          2698 => x"82",
          2699 => x"fc",
          2700 => x"82",
          2701 => x"f8",
          2702 => x"bb",
          2703 => x"05",
          2704 => x"82",
          2705 => x"fc",
          2706 => x"bb",
          2707 => x"05",
          2708 => x"82",
          2709 => x"8c",
          2710 => x"95",
          2711 => x"a4",
          2712 => x"08",
          2713 => x"38",
          2714 => x"08",
          2715 => x"70",
          2716 => x"08",
          2717 => x"51",
          2718 => x"bb",
          2719 => x"05",
          2720 => x"bb",
          2721 => x"05",
          2722 => x"bb",
          2723 => x"05",
          2724 => x"98",
          2725 => x"0d",
          2726 => x"0c",
          2727 => x"0d",
          2728 => x"70",
          2729 => x"74",
          2730 => x"e3",
          2731 => x"75",
          2732 => x"f3",
          2733 => x"98",
          2734 => x"0c",
          2735 => x"54",
          2736 => x"74",
          2737 => x"a0",
          2738 => x"06",
          2739 => x"15",
          2740 => x"80",
          2741 => x"29",
          2742 => x"05",
          2743 => x"56",
          2744 => x"82",
          2745 => x"53",
          2746 => x"08",
          2747 => x"3f",
          2748 => x"08",
          2749 => x"16",
          2750 => x"81",
          2751 => x"38",
          2752 => x"81",
          2753 => x"54",
          2754 => x"c9",
          2755 => x"73",
          2756 => x"0c",
          2757 => x"04",
          2758 => x"73",
          2759 => x"26",
          2760 => x"71",
          2761 => x"99",
          2762 => x"71",
          2763 => x"9e",
          2764 => x"80",
          2765 => x"88",
          2766 => x"39",
          2767 => x"51",
          2768 => x"82",
          2769 => x"80",
          2770 => x"9f",
          2771 => x"e4",
          2772 => x"d0",
          2773 => x"39",
          2774 => x"51",
          2775 => x"82",
          2776 => x"80",
          2777 => x"a0",
          2778 => x"c8",
          2779 => x"a4",
          2780 => x"39",
          2781 => x"51",
          2782 => x"a0",
          2783 => x"39",
          2784 => x"51",
          2785 => x"a1",
          2786 => x"39",
          2787 => x"51",
          2788 => x"a1",
          2789 => x"39",
          2790 => x"51",
          2791 => x"a1",
          2792 => x"39",
          2793 => x"51",
          2794 => x"a2",
          2795 => x"39",
          2796 => x"51",
          2797 => x"83",
          2798 => x"fb",
          2799 => x"79",
          2800 => x"87",
          2801 => x"38",
          2802 => x"87",
          2803 => x"90",
          2804 => x"52",
          2805 => x"cd",
          2806 => x"98",
          2807 => x"51",
          2808 => x"82",
          2809 => x"54",
          2810 => x"52",
          2811 => x"51",
          2812 => x"3f",
          2813 => x"04",
          2814 => x"66",
          2815 => x"80",
          2816 => x"5b",
          2817 => x"78",
          2818 => x"07",
          2819 => x"57",
          2820 => x"56",
          2821 => x"26",
          2822 => x"56",
          2823 => x"70",
          2824 => x"51",
          2825 => x"74",
          2826 => x"81",
          2827 => x"8c",
          2828 => x"56",
          2829 => x"3f",
          2830 => x"08",
          2831 => x"98",
          2832 => x"82",
          2833 => x"87",
          2834 => x"0c",
          2835 => x"08",
          2836 => x"d4",
          2837 => x"80",
          2838 => x"75",
          2839 => x"8b",
          2840 => x"98",
          2841 => x"bb",
          2842 => x"38",
          2843 => x"80",
          2844 => x"74",
          2845 => x"59",
          2846 => x"96",
          2847 => x"51",
          2848 => x"3f",
          2849 => x"78",
          2850 => x"7b",
          2851 => x"2a",
          2852 => x"57",
          2853 => x"80",
          2854 => x"82",
          2855 => x"87",
          2856 => x"08",
          2857 => x"fe",
          2858 => x"56",
          2859 => x"98",
          2860 => x"0d",
          2861 => x"0d",
          2862 => x"05",
          2863 => x"58",
          2864 => x"80",
          2865 => x"7a",
          2866 => x"3f",
          2867 => x"08",
          2868 => x"80",
          2869 => x"76",
          2870 => x"38",
          2871 => x"56",
          2872 => x"54",
          2873 => x"53",
          2874 => x"51",
          2875 => x"bb",
          2876 => x"83",
          2877 => x"77",
          2878 => x"0c",
          2879 => x"04",
          2880 => x"7f",
          2881 => x"8c",
          2882 => x"05",
          2883 => x"15",
          2884 => x"5c",
          2885 => x"5e",
          2886 => x"a2",
          2887 => x"b9",
          2888 => x"a2",
          2889 => x"dd",
          2890 => x"74",
          2891 => x"fd",
          2892 => x"2e",
          2893 => x"a0",
          2894 => x"80",
          2895 => x"18",
          2896 => x"27",
          2897 => x"22",
          2898 => x"fc",
          2899 => x"88",
          2900 => x"82",
          2901 => x"e0",
          2902 => x"15",
          2903 => x"39",
          2904 => x"72",
          2905 => x"38",
          2906 => x"82",
          2907 => x"ff",
          2908 => x"88",
          2909 => x"84",
          2910 => x"3f",
          2911 => x"a0",
          2912 => x"53",
          2913 => x"8e",
          2914 => x"52",
          2915 => x"51",
          2916 => x"3f",
          2917 => x"a3",
          2918 => x"e9",
          2919 => x"55",
          2920 => x"08",
          2921 => x"e3",
          2922 => x"ff",
          2923 => x"9c",
          2924 => x"3f",
          2925 => x"79",
          2926 => x"38",
          2927 => x"33",
          2928 => x"56",
          2929 => x"83",
          2930 => x"80",
          2931 => x"27",
          2932 => x"53",
          2933 => x"70",
          2934 => x"51",
          2935 => x"2e",
          2936 => x"80",
          2937 => x"38",
          2938 => x"08",
          2939 => x"88",
          2940 => x"ec",
          2941 => x"51",
          2942 => x"81",
          2943 => x"b6",
          2944 => x"a0",
          2945 => x"3f",
          2946 => x"1c",
          2947 => x"ef",
          2948 => x"98",
          2949 => x"70",
          2950 => x"57",
          2951 => x"09",
          2952 => x"38",
          2953 => x"82",
          2954 => x"98",
          2955 => x"2c",
          2956 => x"70",
          2957 => x"32",
          2958 => x"72",
          2959 => x"07",
          2960 => x"58",
          2961 => x"57",
          2962 => x"d8",
          2963 => x"2e",
          2964 => x"85",
          2965 => x"8c",
          2966 => x"53",
          2967 => x"fd",
          2968 => x"53",
          2969 => x"98",
          2970 => x"0d",
          2971 => x"0d",
          2972 => x"33",
          2973 => x"53",
          2974 => x"52",
          2975 => x"d8",
          2976 => x"f0",
          2977 => x"ca",
          2978 => x"b8",
          2979 => x"c4",
          2980 => x"f1",
          2981 => x"a3",
          2982 => x"b6",
          2983 => x"80",
          2984 => x"a4",
          2985 => x"3d",
          2986 => x"3d",
          2987 => x"96",
          2988 => x"aa",
          2989 => x"51",
          2990 => x"82",
          2991 => x"9d",
          2992 => x"51",
          2993 => x"72",
          2994 => x"81",
          2995 => x"71",
          2996 => x"38",
          2997 => x"94",
          2998 => x"84",
          2999 => x"3f",
          3000 => x"88",
          3001 => x"2a",
          3002 => x"51",
          3003 => x"2e",
          3004 => x"51",
          3005 => x"82",
          3006 => x"9d",
          3007 => x"51",
          3008 => x"72",
          3009 => x"81",
          3010 => x"71",
          3011 => x"38",
          3012 => x"d8",
          3013 => x"a8",
          3014 => x"3f",
          3015 => x"cc",
          3016 => x"2a",
          3017 => x"51",
          3018 => x"2e",
          3019 => x"51",
          3020 => x"82",
          3021 => x"9c",
          3022 => x"51",
          3023 => x"72",
          3024 => x"81",
          3025 => x"71",
          3026 => x"38",
          3027 => x"9c",
          3028 => x"d0",
          3029 => x"3f",
          3030 => x"90",
          3031 => x"2a",
          3032 => x"51",
          3033 => x"2e",
          3034 => x"51",
          3035 => x"82",
          3036 => x"9c",
          3037 => x"51",
          3038 => x"72",
          3039 => x"81",
          3040 => x"71",
          3041 => x"38",
          3042 => x"e0",
          3043 => x"f8",
          3044 => x"3f",
          3045 => x"d4",
          3046 => x"2a",
          3047 => x"51",
          3048 => x"2e",
          3049 => x"51",
          3050 => x"82",
          3051 => x"9b",
          3052 => x"51",
          3053 => x"a8",
          3054 => x"3d",
          3055 => x"3d",
          3056 => x"84",
          3057 => x"33",
          3058 => x"56",
          3059 => x"51",
          3060 => x"0b",
          3061 => x"94",
          3062 => x"a9",
          3063 => x"82",
          3064 => x"82",
          3065 => x"80",
          3066 => x"82",
          3067 => x"30",
          3068 => x"98",
          3069 => x"25",
          3070 => x"51",
          3071 => x"0b",
          3072 => x"94",
          3073 => x"82",
          3074 => x"54",
          3075 => x"09",
          3076 => x"38",
          3077 => x"53",
          3078 => x"51",
          3079 => x"3f",
          3080 => x"08",
          3081 => x"38",
          3082 => x"08",
          3083 => x"3f",
          3084 => x"d2",
          3085 => x"88",
          3086 => x"0b",
          3087 => x"b6",
          3088 => x"0b",
          3089 => x"33",
          3090 => x"2e",
          3091 => x"8c",
          3092 => x"dc",
          3093 => x"75",
          3094 => x"3f",
          3095 => x"bb",
          3096 => x"3d",
          3097 => x"3d",
          3098 => x"71",
          3099 => x"0c",
          3100 => x"52",
          3101 => x"ca",
          3102 => x"bb",
          3103 => x"ff",
          3104 => x"7e",
          3105 => x"06",
          3106 => x"3d",
          3107 => x"82",
          3108 => x"79",
          3109 => x"3f",
          3110 => x"52",
          3111 => x"51",
          3112 => x"3f",
          3113 => x"08",
          3114 => x"38",
          3115 => x"51",
          3116 => x"81",
          3117 => x"82",
          3118 => x"d9",
          3119 => x"3d",
          3120 => x"80",
          3121 => x"51",
          3122 => x"b5",
          3123 => x"05",
          3124 => x"3f",
          3125 => x"08",
          3126 => x"90",
          3127 => x"79",
          3128 => x"89",
          3129 => x"80",
          3130 => x"d9",
          3131 => x"2e",
          3132 => x"79",
          3133 => x"38",
          3134 => x"81",
          3135 => x"82",
          3136 => x"79",
          3137 => x"af",
          3138 => x"39",
          3139 => x"82",
          3140 => x"94",
          3141 => x"38",
          3142 => x"79",
          3143 => x"ff",
          3144 => x"24",
          3145 => x"b0",
          3146 => x"38",
          3147 => x"84",
          3148 => x"c4",
          3149 => x"2e",
          3150 => x"79",
          3151 => x"86",
          3152 => x"b4",
          3153 => x"d5",
          3154 => x"38",
          3155 => x"24",
          3156 => x"80",
          3157 => x"c9",
          3158 => x"d0",
          3159 => x"79",
          3160 => x"89",
          3161 => x"80",
          3162 => x"9b",
          3163 => x"39",
          3164 => x"2e",
          3165 => x"79",
          3166 => x"8c",
          3167 => x"f8",
          3168 => x"82",
          3169 => x"38",
          3170 => x"24",
          3171 => x"80",
          3172 => x"e3",
          3173 => x"f9",
          3174 => x"38",
          3175 => x"79",
          3176 => x"8d",
          3177 => x"81",
          3178 => x"c6",
          3179 => x"39",
          3180 => x"80",
          3181 => x"84",
          3182 => x"f8",
          3183 => x"98",
          3184 => x"82",
          3185 => x"8f",
          3186 => x"3d",
          3187 => x"53",
          3188 => x"51",
          3189 => x"82",
          3190 => x"80",
          3191 => x"81",
          3192 => x"38",
          3193 => x"80",
          3194 => x"52",
          3195 => x"05",
          3196 => x"c7",
          3197 => x"bb",
          3198 => x"ff",
          3199 => x"8d",
          3200 => x"b8",
          3201 => x"3f",
          3202 => x"ab",
          3203 => x"c8",
          3204 => x"39",
          3205 => x"80",
          3206 => x"84",
          3207 => x"94",
          3208 => x"98",
          3209 => x"fd",
          3210 => x"53",
          3211 => x"80",
          3212 => x"51",
          3213 => x"3f",
          3214 => x"08",
          3215 => x"e0",
          3216 => x"39",
          3217 => x"80",
          3218 => x"84",
          3219 => x"e4",
          3220 => x"98",
          3221 => x"87",
          3222 => x"26",
          3223 => x"b5",
          3224 => x"11",
          3225 => x"05",
          3226 => x"3f",
          3227 => x"08",
          3228 => x"bb",
          3229 => x"64",
          3230 => x"e8",
          3231 => x"ff",
          3232 => x"02",
          3233 => x"33",
          3234 => x"64",
          3235 => x"82",
          3236 => x"51",
          3237 => x"3f",
          3238 => x"08",
          3239 => x"82",
          3240 => x"d5",
          3241 => x"5e",
          3242 => x"b5",
          3243 => x"05",
          3244 => x"3f",
          3245 => x"08",
          3246 => x"84",
          3247 => x"90",
          3248 => x"53",
          3249 => x"08",
          3250 => x"f2",
          3251 => x"d5",
          3252 => x"ff",
          3253 => x"8f",
          3254 => x"bb",
          3255 => x"3d",
          3256 => x"52",
          3257 => x"3f",
          3258 => x"08",
          3259 => x"84",
          3260 => x"90",
          3261 => x"bb",
          3262 => x"3d",
          3263 => x"52",
          3264 => x"3f",
          3265 => x"59",
          3266 => x"58",
          3267 => x"57",
          3268 => x"55",
          3269 => x"08",
          3270 => x"54",
          3271 => x"52",
          3272 => x"91",
          3273 => x"98",
          3274 => x"fb",
          3275 => x"bb",
          3276 => x"ef",
          3277 => x"ff",
          3278 => x"ff",
          3279 => x"ff",
          3280 => x"ce",
          3281 => x"bb",
          3282 => x"2e",
          3283 => x"b5",
          3284 => x"11",
          3285 => x"05",
          3286 => x"3f",
          3287 => x"08",
          3288 => x"d3",
          3289 => x"fe",
          3290 => x"ff",
          3291 => x"ce",
          3292 => x"bb",
          3293 => x"38",
          3294 => x"08",
          3295 => x"ec",
          3296 => x"3f",
          3297 => x"5b",
          3298 => x"81",
          3299 => x"5a",
          3300 => x"84",
          3301 => x"7b",
          3302 => x"38",
          3303 => x"b5",
          3304 => x"11",
          3305 => x"05",
          3306 => x"3f",
          3307 => x"08",
          3308 => x"83",
          3309 => x"fe",
          3310 => x"ff",
          3311 => x"cd",
          3312 => x"bb",
          3313 => x"2e",
          3314 => x"b5",
          3315 => x"11",
          3316 => x"05",
          3317 => x"3f",
          3318 => x"08",
          3319 => x"d7",
          3320 => x"fc",
          3321 => x"3f",
          3322 => x"64",
          3323 => x"38",
          3324 => x"70",
          3325 => x"33",
          3326 => x"81",
          3327 => x"39",
          3328 => x"80",
          3329 => x"84",
          3330 => x"a8",
          3331 => x"98",
          3332 => x"f9",
          3333 => x"3d",
          3334 => x"53",
          3335 => x"51",
          3336 => x"82",
          3337 => x"80",
          3338 => x"38",
          3339 => x"f8",
          3340 => x"84",
          3341 => x"fc",
          3342 => x"98",
          3343 => x"f8",
          3344 => x"a7",
          3345 => x"bd",
          3346 => x"7a",
          3347 => x"38",
          3348 => x"7c",
          3349 => x"5c",
          3350 => x"92",
          3351 => x"7b",
          3352 => x"53",
          3353 => x"a7",
          3354 => x"aa",
          3355 => x"1b",
          3356 => x"44",
          3357 => x"82",
          3358 => x"89",
          3359 => x"3d",
          3360 => x"53",
          3361 => x"51",
          3362 => x"82",
          3363 => x"80",
          3364 => x"ba",
          3365 => x"79",
          3366 => x"38",
          3367 => x"08",
          3368 => x"39",
          3369 => x"33",
          3370 => x"2e",
          3371 => x"b9",
          3372 => x"bc",
          3373 => x"86",
          3374 => x"80",
          3375 => x"82",
          3376 => x"45",
          3377 => x"ba",
          3378 => x"79",
          3379 => x"38",
          3380 => x"08",
          3381 => x"82",
          3382 => x"5a",
          3383 => x"88",
          3384 => x"dc",
          3385 => x"39",
          3386 => x"08",
          3387 => x"45",
          3388 => x"fc",
          3389 => x"84",
          3390 => x"b8",
          3391 => x"98",
          3392 => x"38",
          3393 => x"33",
          3394 => x"2e",
          3395 => x"b9",
          3396 => x"80",
          3397 => x"ba",
          3398 => x"79",
          3399 => x"38",
          3400 => x"08",
          3401 => x"82",
          3402 => x"5a",
          3403 => x"88",
          3404 => x"d0",
          3405 => x"39",
          3406 => x"33",
          3407 => x"2e",
          3408 => x"b9",
          3409 => x"99",
          3410 => x"82",
          3411 => x"80",
          3412 => x"82",
          3413 => x"44",
          3414 => x"b9",
          3415 => x"05",
          3416 => x"fe",
          3417 => x"ff",
          3418 => x"ca",
          3419 => x"bb",
          3420 => x"2e",
          3421 => x"63",
          3422 => x"88",
          3423 => x"81",
          3424 => x"32",
          3425 => x"72",
          3426 => x"70",
          3427 => x"51",
          3428 => x"80",
          3429 => x"7b",
          3430 => x"38",
          3431 => x"a7",
          3432 => x"e1",
          3433 => x"64",
          3434 => x"63",
          3435 => x"ee",
          3436 => x"a7",
          3437 => x"c2",
          3438 => x"ff",
          3439 => x"ff",
          3440 => x"c9",
          3441 => x"bb",
          3442 => x"2e",
          3443 => x"b5",
          3444 => x"11",
          3445 => x"05",
          3446 => x"3f",
          3447 => x"08",
          3448 => x"38",
          3449 => x"80",
          3450 => x"7a",
          3451 => x"05",
          3452 => x"fe",
          3453 => x"ff",
          3454 => x"c9",
          3455 => x"bb",
          3456 => x"38",
          3457 => x"64",
          3458 => x"52",
          3459 => x"51",
          3460 => x"3f",
          3461 => x"7a",
          3462 => x"3f",
          3463 => x"33",
          3464 => x"2e",
          3465 => x"9f",
          3466 => x"38",
          3467 => x"fc",
          3468 => x"84",
          3469 => x"fc",
          3470 => x"98",
          3471 => x"91",
          3472 => x"02",
          3473 => x"33",
          3474 => x"81",
          3475 => x"b7",
          3476 => x"dc",
          3477 => x"3f",
          3478 => x"b5",
          3479 => x"11",
          3480 => x"05",
          3481 => x"3f",
          3482 => x"08",
          3483 => x"c7",
          3484 => x"fe",
          3485 => x"ff",
          3486 => x"c2",
          3487 => x"bb",
          3488 => x"2e",
          3489 => x"5a",
          3490 => x"05",
          3491 => x"82",
          3492 => x"79",
          3493 => x"fe",
          3494 => x"ff",
          3495 => x"c2",
          3496 => x"bb",
          3497 => x"38",
          3498 => x"61",
          3499 => x"52",
          3500 => x"51",
          3501 => x"3f",
          3502 => x"7a",
          3503 => x"3f",
          3504 => x"33",
          3505 => x"2e",
          3506 => x"79",
          3507 => x"38",
          3508 => x"42",
          3509 => x"3d",
          3510 => x"53",
          3511 => x"51",
          3512 => x"82",
          3513 => x"80",
          3514 => x"61",
          3515 => x"c2",
          3516 => x"70",
          3517 => x"23",
          3518 => x"af",
          3519 => x"dc",
          3520 => x"3f",
          3521 => x"b5",
          3522 => x"11",
          3523 => x"05",
          3524 => x"3f",
          3525 => x"08",
          3526 => x"9b",
          3527 => x"fe",
          3528 => x"ff",
          3529 => x"c1",
          3530 => x"bb",
          3531 => x"2e",
          3532 => x"61",
          3533 => x"61",
          3534 => x"b5",
          3535 => x"11",
          3536 => x"05",
          3537 => x"3f",
          3538 => x"08",
          3539 => x"e7",
          3540 => x"08",
          3541 => x"a7",
          3542 => x"a4",
          3543 => x"f8",
          3544 => x"c6",
          3545 => x"46",
          3546 => x"79",
          3547 => x"c7",
          3548 => x"27",
          3549 => x"3d",
          3550 => x"53",
          3551 => x"51",
          3552 => x"82",
          3553 => x"80",
          3554 => x"61",
          3555 => x"5a",
          3556 => x"42",
          3557 => x"82",
          3558 => x"cb",
          3559 => x"b1",
          3560 => x"fc",
          3561 => x"3f",
          3562 => x"8b",
          3563 => x"39",
          3564 => x"51",
          3565 => x"a2",
          3566 => x"3f",
          3567 => x"82",
          3568 => x"cb",
          3569 => x"80",
          3570 => x"c0",
          3571 => x"84",
          3572 => x"87",
          3573 => x"0c",
          3574 => x"82",
          3575 => x"cb",
          3576 => x"80",
          3577 => x"c0",
          3578 => x"8c",
          3579 => x"87",
          3580 => x"0c",
          3581 => x"b5",
          3582 => x"11",
          3583 => x"05",
          3584 => x"3f",
          3585 => x"08",
          3586 => x"ab",
          3587 => x"82",
          3588 => x"ff",
          3589 => x"64",
          3590 => x"b5",
          3591 => x"11",
          3592 => x"05",
          3593 => x"3f",
          3594 => x"08",
          3595 => x"87",
          3596 => x"82",
          3597 => x"ff",
          3598 => x"64",
          3599 => x"82",
          3600 => x"80",
          3601 => x"38",
          3602 => x"08",
          3603 => x"8c",
          3604 => x"84",
          3605 => x"39",
          3606 => x"51",
          3607 => x"ff",
          3608 => x"f0",
          3609 => x"a9",
          3610 => x"99",
          3611 => x"ff",
          3612 => x"ad",
          3613 => x"39",
          3614 => x"33",
          3615 => x"2e",
          3616 => x"7e",
          3617 => x"79",
          3618 => x"d6",
          3619 => x"ff",
          3620 => x"83",
          3621 => x"bb",
          3622 => x"81",
          3623 => x"2e",
          3624 => x"82",
          3625 => x"7c",
          3626 => x"38",
          3627 => x"7c",
          3628 => x"38",
          3629 => x"82",
          3630 => x"7b",
          3631 => x"dc",
          3632 => x"82",
          3633 => x"b5",
          3634 => x"05",
          3635 => x"f0",
          3636 => x"82",
          3637 => x"b5",
          3638 => x"05",
          3639 => x"e0",
          3640 => x"7b",
          3641 => x"dc",
          3642 => x"82",
          3643 => x"b5",
          3644 => x"05",
          3645 => x"c8",
          3646 => x"7b",
          3647 => x"82",
          3648 => x"b5",
          3649 => x"05",
          3650 => x"b4",
          3651 => x"e8",
          3652 => x"bc",
          3653 => x"c8",
          3654 => x"65",
          3655 => x"82",
          3656 => x"82",
          3657 => x"b5",
          3658 => x"05",
          3659 => x"3f",
          3660 => x"08",
          3661 => x"08",
          3662 => x"70",
          3663 => x"25",
          3664 => x"40",
          3665 => x"83",
          3666 => x"81",
          3667 => x"06",
          3668 => x"2e",
          3669 => x"1d",
          3670 => x"06",
          3671 => x"fe",
          3672 => x"81",
          3673 => x"32",
          3674 => x"8a",
          3675 => x"2e",
          3676 => x"ee",
          3677 => x"aa",
          3678 => x"89",
          3679 => x"39",
          3680 => x"80",
          3681 => x"c8",
          3682 => x"94",
          3683 => x"54",
          3684 => x"80",
          3685 => x"df",
          3686 => x"bb",
          3687 => x"2b",
          3688 => x"53",
          3689 => x"52",
          3690 => x"f9",
          3691 => x"bb",
          3692 => x"75",
          3693 => x"94",
          3694 => x"54",
          3695 => x"80",
          3696 => x"de",
          3697 => x"bb",
          3698 => x"2b",
          3699 => x"53",
          3700 => x"52",
          3701 => x"cd",
          3702 => x"bb",
          3703 => x"75",
          3704 => x"83",
          3705 => x"94",
          3706 => x"80",
          3707 => x"c0",
          3708 => x"80",
          3709 => x"80",
          3710 => x"83",
          3711 => x"99",
          3712 => x"5c",
          3713 => x"0b",
          3714 => x"88",
          3715 => x"72",
          3716 => x"ec",
          3717 => x"bd",
          3718 => x"3f",
          3719 => x"51",
          3720 => x"82",
          3721 => x"c6",
          3722 => x"dd",
          3723 => x"e6",
          3724 => x"e8",
          3725 => x"ae",
          3726 => x"fe",
          3727 => x"52",
          3728 => x"88",
          3729 => x"d9",
          3730 => x"98",
          3731 => x"06",
          3732 => x"14",
          3733 => x"80",
          3734 => x"71",
          3735 => x"0c",
          3736 => x"04",
          3737 => x"76",
          3738 => x"55",
          3739 => x"54",
          3740 => x"81",
          3741 => x"33",
          3742 => x"2e",
          3743 => x"86",
          3744 => x"53",
          3745 => x"33",
          3746 => x"2e",
          3747 => x"86",
          3748 => x"53",
          3749 => x"52",
          3750 => x"09",
          3751 => x"38",
          3752 => x"12",
          3753 => x"33",
          3754 => x"a2",
          3755 => x"81",
          3756 => x"2e",
          3757 => x"ea",
          3758 => x"81",
          3759 => x"72",
          3760 => x"70",
          3761 => x"38",
          3762 => x"80",
          3763 => x"73",
          3764 => x"72",
          3765 => x"70",
          3766 => x"81",
          3767 => x"81",
          3768 => x"32",
          3769 => x"80",
          3770 => x"51",
          3771 => x"80",
          3772 => x"80",
          3773 => x"05",
          3774 => x"75",
          3775 => x"70",
          3776 => x"0c",
          3777 => x"04",
          3778 => x"76",
          3779 => x"80",
          3780 => x"86",
          3781 => x"52",
          3782 => x"b9",
          3783 => x"bb",
          3784 => x"38",
          3785 => x"39",
          3786 => x"82",
          3787 => x"86",
          3788 => x"fc",
          3789 => x"82",
          3790 => x"05",
          3791 => x"52",
          3792 => x"81",
          3793 => x"13",
          3794 => x"51",
          3795 => x"9e",
          3796 => x"38",
          3797 => x"51",
          3798 => x"97",
          3799 => x"38",
          3800 => x"51",
          3801 => x"bb",
          3802 => x"38",
          3803 => x"51",
          3804 => x"bb",
          3805 => x"38",
          3806 => x"55",
          3807 => x"87",
          3808 => x"d9",
          3809 => x"22",
          3810 => x"73",
          3811 => x"80",
          3812 => x"0b",
          3813 => x"9c",
          3814 => x"87",
          3815 => x"0c",
          3816 => x"87",
          3817 => x"0c",
          3818 => x"87",
          3819 => x"0c",
          3820 => x"87",
          3821 => x"0c",
          3822 => x"87",
          3823 => x"0c",
          3824 => x"87",
          3825 => x"0c",
          3826 => x"98",
          3827 => x"87",
          3828 => x"0c",
          3829 => x"c0",
          3830 => x"80",
          3831 => x"bb",
          3832 => x"3d",
          3833 => x"3d",
          3834 => x"87",
          3835 => x"5d",
          3836 => x"87",
          3837 => x"08",
          3838 => x"23",
          3839 => x"b8",
          3840 => x"82",
          3841 => x"c0",
          3842 => x"5a",
          3843 => x"34",
          3844 => x"b0",
          3845 => x"84",
          3846 => x"c0",
          3847 => x"5a",
          3848 => x"34",
          3849 => x"a8",
          3850 => x"86",
          3851 => x"c0",
          3852 => x"5c",
          3853 => x"23",
          3854 => x"a0",
          3855 => x"8a",
          3856 => x"7d",
          3857 => x"ff",
          3858 => x"7b",
          3859 => x"06",
          3860 => x"33",
          3861 => x"33",
          3862 => x"33",
          3863 => x"33",
          3864 => x"33",
          3865 => x"ff",
          3866 => x"82",
          3867 => x"ff",
          3868 => x"8f",
          3869 => x"fb",
          3870 => x"9f",
          3871 => x"b9",
          3872 => x"81",
          3873 => x"55",
          3874 => x"94",
          3875 => x"80",
          3876 => x"87",
          3877 => x"51",
          3878 => x"96",
          3879 => x"06",
          3880 => x"70",
          3881 => x"38",
          3882 => x"70",
          3883 => x"51",
          3884 => x"72",
          3885 => x"81",
          3886 => x"70",
          3887 => x"38",
          3888 => x"70",
          3889 => x"51",
          3890 => x"38",
          3891 => x"06",
          3892 => x"94",
          3893 => x"80",
          3894 => x"87",
          3895 => x"52",
          3896 => x"74",
          3897 => x"0c",
          3898 => x"04",
          3899 => x"02",
          3900 => x"70",
          3901 => x"2a",
          3902 => x"70",
          3903 => x"34",
          3904 => x"04",
          3905 => x"02",
          3906 => x"58",
          3907 => x"09",
          3908 => x"38",
          3909 => x"51",
          3910 => x"b9",
          3911 => x"81",
          3912 => x"56",
          3913 => x"84",
          3914 => x"2e",
          3915 => x"c0",
          3916 => x"72",
          3917 => x"2a",
          3918 => x"55",
          3919 => x"80",
          3920 => x"73",
          3921 => x"81",
          3922 => x"72",
          3923 => x"81",
          3924 => x"06",
          3925 => x"80",
          3926 => x"73",
          3927 => x"81",
          3928 => x"72",
          3929 => x"75",
          3930 => x"53",
          3931 => x"80",
          3932 => x"2e",
          3933 => x"c0",
          3934 => x"77",
          3935 => x"0b",
          3936 => x"0c",
          3937 => x"04",
          3938 => x"79",
          3939 => x"33",
          3940 => x"06",
          3941 => x"70",
          3942 => x"fc",
          3943 => x"ff",
          3944 => x"82",
          3945 => x"70",
          3946 => x"59",
          3947 => x"87",
          3948 => x"51",
          3949 => x"86",
          3950 => x"94",
          3951 => x"08",
          3952 => x"70",
          3953 => x"54",
          3954 => x"2e",
          3955 => x"91",
          3956 => x"06",
          3957 => x"d7",
          3958 => x"32",
          3959 => x"51",
          3960 => x"2e",
          3961 => x"93",
          3962 => x"06",
          3963 => x"ff",
          3964 => x"81",
          3965 => x"87",
          3966 => x"52",
          3967 => x"86",
          3968 => x"94",
          3969 => x"72",
          3970 => x"74",
          3971 => x"ff",
          3972 => x"57",
          3973 => x"38",
          3974 => x"98",
          3975 => x"0d",
          3976 => x"0d",
          3977 => x"33",
          3978 => x"06",
          3979 => x"c0",
          3980 => x"72",
          3981 => x"38",
          3982 => x"94",
          3983 => x"70",
          3984 => x"81",
          3985 => x"51",
          3986 => x"e2",
          3987 => x"ff",
          3988 => x"c0",
          3989 => x"70",
          3990 => x"38",
          3991 => x"90",
          3992 => x"70",
          3993 => x"82",
          3994 => x"51",
          3995 => x"04",
          3996 => x"82",
          3997 => x"81",
          3998 => x"bb",
          3999 => x"fe",
          4000 => x"b9",
          4001 => x"81",
          4002 => x"53",
          4003 => x"84",
          4004 => x"2e",
          4005 => x"c0",
          4006 => x"71",
          4007 => x"2a",
          4008 => x"51",
          4009 => x"52",
          4010 => x"a0",
          4011 => x"ff",
          4012 => x"c0",
          4013 => x"70",
          4014 => x"38",
          4015 => x"90",
          4016 => x"70",
          4017 => x"98",
          4018 => x"51",
          4019 => x"98",
          4020 => x"0d",
          4021 => x"0d",
          4022 => x"80",
          4023 => x"2a",
          4024 => x"51",
          4025 => x"84",
          4026 => x"c0",
          4027 => x"82",
          4028 => x"87",
          4029 => x"08",
          4030 => x"0c",
          4031 => x"94",
          4032 => x"c4",
          4033 => x"9e",
          4034 => x"b9",
          4035 => x"c0",
          4036 => x"82",
          4037 => x"87",
          4038 => x"08",
          4039 => x"0c",
          4040 => x"ac",
          4041 => x"d4",
          4042 => x"9e",
          4043 => x"b9",
          4044 => x"c0",
          4045 => x"82",
          4046 => x"87",
          4047 => x"08",
          4048 => x"0c",
          4049 => x"bc",
          4050 => x"e4",
          4051 => x"9e",
          4052 => x"b9",
          4053 => x"c0",
          4054 => x"82",
          4055 => x"87",
          4056 => x"08",
          4057 => x"b9",
          4058 => x"c0",
          4059 => x"82",
          4060 => x"87",
          4061 => x"08",
          4062 => x"0c",
          4063 => x"8c",
          4064 => x"fc",
          4065 => x"82",
          4066 => x"80",
          4067 => x"9e",
          4068 => x"84",
          4069 => x"51",
          4070 => x"80",
          4071 => x"81",
          4072 => x"ba",
          4073 => x"0b",
          4074 => x"90",
          4075 => x"80",
          4076 => x"52",
          4077 => x"2e",
          4078 => x"52",
          4079 => x"82",
          4080 => x"87",
          4081 => x"08",
          4082 => x"0a",
          4083 => x"52",
          4084 => x"83",
          4085 => x"71",
          4086 => x"34",
          4087 => x"c0",
          4088 => x"70",
          4089 => x"06",
          4090 => x"70",
          4091 => x"38",
          4092 => x"82",
          4093 => x"80",
          4094 => x"9e",
          4095 => x"a0",
          4096 => x"51",
          4097 => x"80",
          4098 => x"81",
          4099 => x"ba",
          4100 => x"0b",
          4101 => x"90",
          4102 => x"80",
          4103 => x"52",
          4104 => x"2e",
          4105 => x"52",
          4106 => x"86",
          4107 => x"87",
          4108 => x"08",
          4109 => x"80",
          4110 => x"52",
          4111 => x"83",
          4112 => x"71",
          4113 => x"34",
          4114 => x"c0",
          4115 => x"70",
          4116 => x"06",
          4117 => x"70",
          4118 => x"38",
          4119 => x"82",
          4120 => x"80",
          4121 => x"9e",
          4122 => x"81",
          4123 => x"51",
          4124 => x"80",
          4125 => x"81",
          4126 => x"ba",
          4127 => x"0b",
          4128 => x"90",
          4129 => x"c0",
          4130 => x"52",
          4131 => x"2e",
          4132 => x"52",
          4133 => x"8a",
          4134 => x"87",
          4135 => x"08",
          4136 => x"06",
          4137 => x"70",
          4138 => x"38",
          4139 => x"82",
          4140 => x"87",
          4141 => x"08",
          4142 => x"06",
          4143 => x"51",
          4144 => x"82",
          4145 => x"80",
          4146 => x"9e",
          4147 => x"84",
          4148 => x"52",
          4149 => x"2e",
          4150 => x"52",
          4151 => x"8d",
          4152 => x"9e",
          4153 => x"83",
          4154 => x"84",
          4155 => x"51",
          4156 => x"8e",
          4157 => x"87",
          4158 => x"08",
          4159 => x"51",
          4160 => x"80",
          4161 => x"81",
          4162 => x"ba",
          4163 => x"c0",
          4164 => x"70",
          4165 => x"51",
          4166 => x"90",
          4167 => x"0d",
          4168 => x"0d",
          4169 => x"51",
          4170 => x"3f",
          4171 => x"33",
          4172 => x"2e",
          4173 => x"aa",
          4174 => x"b8",
          4175 => x"aa",
          4176 => x"b8",
          4177 => x"ba",
          4178 => x"73",
          4179 => x"38",
          4180 => x"08",
          4181 => x"08",
          4182 => x"82",
          4183 => x"ff",
          4184 => x"82",
          4185 => x"54",
          4186 => x"94",
          4187 => x"d4",
          4188 => x"d8",
          4189 => x"52",
          4190 => x"51",
          4191 => x"3f",
          4192 => x"33",
          4193 => x"2e",
          4194 => x"b9",
          4195 => x"b9",
          4196 => x"54",
          4197 => x"c8",
          4198 => x"bc",
          4199 => x"85",
          4200 => x"80",
          4201 => x"82",
          4202 => x"82",
          4203 => x"11",
          4204 => x"ab",
          4205 => x"90",
          4206 => x"ba",
          4207 => x"73",
          4208 => x"38",
          4209 => x"08",
          4210 => x"08",
          4211 => x"82",
          4212 => x"ff",
          4213 => x"82",
          4214 => x"54",
          4215 => x"8e",
          4216 => x"8c",
          4217 => x"ac",
          4218 => x"8f",
          4219 => x"ba",
          4220 => x"73",
          4221 => x"38",
          4222 => x"33",
          4223 => x"bc",
          4224 => x"d4",
          4225 => x"8d",
          4226 => x"80",
          4227 => x"82",
          4228 => x"52",
          4229 => x"51",
          4230 => x"3f",
          4231 => x"33",
          4232 => x"2e",
          4233 => x"ac",
          4234 => x"b6",
          4235 => x"ba",
          4236 => x"73",
          4237 => x"38",
          4238 => x"51",
          4239 => x"3f",
          4240 => x"33",
          4241 => x"2e",
          4242 => x"ad",
          4243 => x"b6",
          4244 => x"ba",
          4245 => x"73",
          4246 => x"38",
          4247 => x"51",
          4248 => x"3f",
          4249 => x"33",
          4250 => x"2e",
          4251 => x"ad",
          4252 => x"b6",
          4253 => x"ad",
          4254 => x"b6",
          4255 => x"b9",
          4256 => x"82",
          4257 => x"ff",
          4258 => x"82",
          4259 => x"52",
          4260 => x"51",
          4261 => x"3f",
          4262 => x"08",
          4263 => x"9c",
          4264 => x"b4",
          4265 => x"c4",
          4266 => x"d9",
          4267 => x"f0",
          4268 => x"ae",
          4269 => x"8e",
          4270 => x"b9",
          4271 => x"bd",
          4272 => x"75",
          4273 => x"3f",
          4274 => x"08",
          4275 => x"29",
          4276 => x"54",
          4277 => x"98",
          4278 => x"ae",
          4279 => x"8d",
          4280 => x"ba",
          4281 => x"73",
          4282 => x"38",
          4283 => x"08",
          4284 => x"c0",
          4285 => x"cc",
          4286 => x"bb",
          4287 => x"84",
          4288 => x"71",
          4289 => x"82",
          4290 => x"52",
          4291 => x"51",
          4292 => x"3f",
          4293 => x"33",
          4294 => x"2e",
          4295 => x"b9",
          4296 => x"bd",
          4297 => x"75",
          4298 => x"3f",
          4299 => x"08",
          4300 => x"29",
          4301 => x"54",
          4302 => x"98",
          4303 => x"af",
          4304 => x"8d",
          4305 => x"a7",
          4306 => x"b4",
          4307 => x"3d",
          4308 => x"3d",
          4309 => x"05",
          4310 => x"52",
          4311 => x"aa",
          4312 => x"29",
          4313 => x"05",
          4314 => x"04",
          4315 => x"51",
          4316 => x"b0",
          4317 => x"39",
          4318 => x"51",
          4319 => x"b0",
          4320 => x"39",
          4321 => x"51",
          4322 => x"b0",
          4323 => x"b3",
          4324 => x"3d",
          4325 => x"88",
          4326 => x"ff",
          4327 => x"c0",
          4328 => x"08",
          4329 => x"72",
          4330 => x"07",
          4331 => x"94",
          4332 => x"83",
          4333 => x"ff",
          4334 => x"c0",
          4335 => x"08",
          4336 => x"0c",
          4337 => x"0c",
          4338 => x"82",
          4339 => x"06",
          4340 => x"94",
          4341 => x"51",
          4342 => x"04",
          4343 => x"c0",
          4344 => x"04",
          4345 => x"08",
          4346 => x"84",
          4347 => x"3d",
          4348 => x"2b",
          4349 => x"79",
          4350 => x"98",
          4351 => x"13",
          4352 => x"51",
          4353 => x"51",
          4354 => x"82",
          4355 => x"33",
          4356 => x"74",
          4357 => x"82",
          4358 => x"08",
          4359 => x"05",
          4360 => x"71",
          4361 => x"52",
          4362 => x"09",
          4363 => x"38",
          4364 => x"82",
          4365 => x"85",
          4366 => x"fc",
          4367 => x"02",
          4368 => x"05",
          4369 => x"54",
          4370 => x"80",
          4371 => x"88",
          4372 => x"d3",
          4373 => x"ff",
          4374 => x"88",
          4375 => x"c7",
          4376 => x"ff",
          4377 => x"73",
          4378 => x"ff",
          4379 => x"39",
          4380 => x"b2",
          4381 => x"73",
          4382 => x"0d",
          4383 => x"0d",
          4384 => x"05",
          4385 => x"02",
          4386 => x"05",
          4387 => x"f0",
          4388 => x"29",
          4389 => x"05",
          4390 => x"59",
          4391 => x"59",
          4392 => x"86",
          4393 => x"9a",
          4394 => x"ba",
          4395 => x"84",
          4396 => x"98",
          4397 => x"70",
          4398 => x"5a",
          4399 => x"82",
          4400 => x"75",
          4401 => x"f0",
          4402 => x"29",
          4403 => x"05",
          4404 => x"56",
          4405 => x"2e",
          4406 => x"53",
          4407 => x"51",
          4408 => x"3f",
          4409 => x"33",
          4410 => x"74",
          4411 => x"34",
          4412 => x"06",
          4413 => x"27",
          4414 => x"0b",
          4415 => x"34",
          4416 => x"b6",
          4417 => x"ec",
          4418 => x"80",
          4419 => x"82",
          4420 => x"55",
          4421 => x"8c",
          4422 => x"54",
          4423 => x"52",
          4424 => x"d9",
          4425 => x"ba",
          4426 => x"8a",
          4427 => x"d0",
          4428 => x"ec",
          4429 => x"dd",
          4430 => x"3d",
          4431 => x"3d",
          4432 => x"98",
          4433 => x"72",
          4434 => x"80",
          4435 => x"71",
          4436 => x"3f",
          4437 => x"ff",
          4438 => x"54",
          4439 => x"25",
          4440 => x"0b",
          4441 => x"34",
          4442 => x"08",
          4443 => x"2e",
          4444 => x"51",
          4445 => x"3f",
          4446 => x"08",
          4447 => x"3f",
          4448 => x"ba",
          4449 => x"3d",
          4450 => x"3d",
          4451 => x"80",
          4452 => x"ec",
          4453 => x"e2",
          4454 => x"bb",
          4455 => x"d3",
          4456 => x"ec",
          4457 => x"f8",
          4458 => x"70",
          4459 => x"8b",
          4460 => x"bb",
          4461 => x"2e",
          4462 => x"51",
          4463 => x"3f",
          4464 => x"08",
          4465 => x"82",
          4466 => x"25",
          4467 => x"bb",
          4468 => x"05",
          4469 => x"55",
          4470 => x"75",
          4471 => x"81",
          4472 => x"98",
          4473 => x"87",
          4474 => x"ff",
          4475 => x"06",
          4476 => x"a6",
          4477 => x"d9",
          4478 => x"3d",
          4479 => x"08",
          4480 => x"70",
          4481 => x"52",
          4482 => x"08",
          4483 => x"f6",
          4484 => x"98",
          4485 => x"38",
          4486 => x"ba",
          4487 => x"55",
          4488 => x"8b",
          4489 => x"56",
          4490 => x"3f",
          4491 => x"08",
          4492 => x"38",
          4493 => x"ba",
          4494 => x"bb",
          4495 => x"18",
          4496 => x"0b",
          4497 => x"08",
          4498 => x"82",
          4499 => x"ff",
          4500 => x"55",
          4501 => x"34",
          4502 => x"30",
          4503 => x"9f",
          4504 => x"55",
          4505 => x"85",
          4506 => x"ac",
          4507 => x"ec",
          4508 => x"08",
          4509 => x"e1",
          4510 => x"bb",
          4511 => x"2e",
          4512 => x"b3",
          4513 => x"ad",
          4514 => x"77",
          4515 => x"06",
          4516 => x"52",
          4517 => x"ba",
          4518 => x"51",
          4519 => x"3f",
          4520 => x"54",
          4521 => x"08",
          4522 => x"58",
          4523 => x"98",
          4524 => x"0d",
          4525 => x"0d",
          4526 => x"5c",
          4527 => x"57",
          4528 => x"73",
          4529 => x"81",
          4530 => x"78",
          4531 => x"56",
          4532 => x"98",
          4533 => x"70",
          4534 => x"33",
          4535 => x"73",
          4536 => x"81",
          4537 => x"75",
          4538 => x"38",
          4539 => x"88",
          4540 => x"f4",
          4541 => x"52",
          4542 => x"ab",
          4543 => x"98",
          4544 => x"52",
          4545 => x"ff",
          4546 => x"82",
          4547 => x"80",
          4548 => x"15",
          4549 => x"81",
          4550 => x"74",
          4551 => x"38",
          4552 => x"e6",
          4553 => x"81",
          4554 => x"3d",
          4555 => x"f8",
          4556 => x"a6",
          4557 => x"bb",
          4558 => x"2e",
          4559 => x"1b",
          4560 => x"77",
          4561 => x"3f",
          4562 => x"08",
          4563 => x"55",
          4564 => x"74",
          4565 => x"81",
          4566 => x"ff",
          4567 => x"82",
          4568 => x"8a",
          4569 => x"73",
          4570 => x"0c",
          4571 => x"04",
          4572 => x"b0",
          4573 => x"3d",
          4574 => x"08",
          4575 => x"80",
          4576 => x"34",
          4577 => x"33",
          4578 => x"08",
          4579 => x"81",
          4580 => x"82",
          4581 => x"55",
          4582 => x"38",
          4583 => x"80",
          4584 => x"38",
          4585 => x"06",
          4586 => x"80",
          4587 => x"38",
          4588 => x"c0",
          4589 => x"98",
          4590 => x"ec",
          4591 => x"98",
          4592 => x"81",
          4593 => x"53",
          4594 => x"bb",
          4595 => x"80",
          4596 => x"82",
          4597 => x"80",
          4598 => x"82",
          4599 => x"ff",
          4600 => x"80",
          4601 => x"bb",
          4602 => x"82",
          4603 => x"53",
          4604 => x"90",
          4605 => x"54",
          4606 => x"3f",
          4607 => x"08",
          4608 => x"98",
          4609 => x"09",
          4610 => x"d0",
          4611 => x"98",
          4612 => x"b7",
          4613 => x"bb",
          4614 => x"80",
          4615 => x"98",
          4616 => x"38",
          4617 => x"08",
          4618 => x"17",
          4619 => x"74",
          4620 => x"74",
          4621 => x"52",
          4622 => x"c1",
          4623 => x"70",
          4624 => x"5c",
          4625 => x"27",
          4626 => x"5b",
          4627 => x"09",
          4628 => x"97",
          4629 => x"75",
          4630 => x"34",
          4631 => x"82",
          4632 => x"80",
          4633 => x"f9",
          4634 => x"3d",
          4635 => x"3f",
          4636 => x"08",
          4637 => x"98",
          4638 => x"78",
          4639 => x"38",
          4640 => x"06",
          4641 => x"33",
          4642 => x"70",
          4643 => x"d2",
          4644 => x"98",
          4645 => x"2c",
          4646 => x"05",
          4647 => x"82",
          4648 => x"70",
          4649 => x"33",
          4650 => x"51",
          4651 => x"59",
          4652 => x"56",
          4653 => x"80",
          4654 => x"74",
          4655 => x"74",
          4656 => x"29",
          4657 => x"05",
          4658 => x"51",
          4659 => x"24",
          4660 => x"76",
          4661 => x"77",
          4662 => x"3f",
          4663 => x"08",
          4664 => x"54",
          4665 => x"d7",
          4666 => x"d2",
          4667 => x"56",
          4668 => x"81",
          4669 => x"81",
          4670 => x"70",
          4671 => x"81",
          4672 => x"51",
          4673 => x"26",
          4674 => x"53",
          4675 => x"51",
          4676 => x"82",
          4677 => x"81",
          4678 => x"73",
          4679 => x"39",
          4680 => x"80",
          4681 => x"38",
          4682 => x"74",
          4683 => x"34",
          4684 => x"70",
          4685 => x"d2",
          4686 => x"98",
          4687 => x"2c",
          4688 => x"70",
          4689 => x"b0",
          4690 => x"5e",
          4691 => x"57",
          4692 => x"74",
          4693 => x"81",
          4694 => x"38",
          4695 => x"14",
          4696 => x"80",
          4697 => x"c4",
          4698 => x"82",
          4699 => x"92",
          4700 => x"d2",
          4701 => x"82",
          4702 => x"78",
          4703 => x"75",
          4704 => x"54",
          4705 => x"fd",
          4706 => x"84",
          4707 => x"94",
          4708 => x"08",
          4709 => x"cc",
          4710 => x"7e",
          4711 => x"38",
          4712 => x"33",
          4713 => x"27",
          4714 => x"98",
          4715 => x"2c",
          4716 => x"75",
          4717 => x"74",
          4718 => x"33",
          4719 => x"74",
          4720 => x"29",
          4721 => x"05",
          4722 => x"82",
          4723 => x"56",
          4724 => x"39",
          4725 => x"33",
          4726 => x"54",
          4727 => x"cc",
          4728 => x"54",
          4729 => x"74",
          4730 => x"c8",
          4731 => x"7e",
          4732 => x"81",
          4733 => x"82",
          4734 => x"82",
          4735 => x"70",
          4736 => x"29",
          4737 => x"05",
          4738 => x"82",
          4739 => x"5a",
          4740 => x"74",
          4741 => x"38",
          4742 => x"33",
          4743 => x"aa",
          4744 => x"81",
          4745 => x"81",
          4746 => x"70",
          4747 => x"d2",
          4748 => x"51",
          4749 => x"24",
          4750 => x"d2",
          4751 => x"98",
          4752 => x"2c",
          4753 => x"33",
          4754 => x"56",
          4755 => x"fc",
          4756 => x"51",
          4757 => x"3f",
          4758 => x"0a",
          4759 => x"0a",
          4760 => x"2c",
          4761 => x"33",
          4762 => x"73",
          4763 => x"38",
          4764 => x"83",
          4765 => x"0b",
          4766 => x"82",
          4767 => x"80",
          4768 => x"88",
          4769 => x"3f",
          4770 => x"82",
          4771 => x"70",
          4772 => x"55",
          4773 => x"2e",
          4774 => x"82",
          4775 => x"ff",
          4776 => x"82",
          4777 => x"ff",
          4778 => x"82",
          4779 => x"88",
          4780 => x"f3",
          4781 => x"cc",
          4782 => x"2b",
          4783 => x"82",
          4784 => x"57",
          4785 => x"74",
          4786 => x"38",
          4787 => x"81",
          4788 => x"34",
          4789 => x"ff",
          4790 => x"74",
          4791 => x"29",
          4792 => x"05",
          4793 => x"82",
          4794 => x"58",
          4795 => x"75",
          4796 => x"a0",
          4797 => x"af",
          4798 => x"cc",
          4799 => x"2b",
          4800 => x"82",
          4801 => x"57",
          4802 => x"74",
          4803 => x"da",
          4804 => x"ff",
          4805 => x"74",
          4806 => x"29",
          4807 => x"05",
          4808 => x"82",
          4809 => x"58",
          4810 => x"75",
          4811 => x"fa",
          4812 => x"d2",
          4813 => x"05",
          4814 => x"34",
          4815 => x"a7",
          4816 => x"d2",
          4817 => x"51",
          4818 => x"82",
          4819 => x"81",
          4820 => x"73",
          4821 => x"d2",
          4822 => x"73",
          4823 => x"38",
          4824 => x"52",
          4825 => x"95",
          4826 => x"80",
          4827 => x"0b",
          4828 => x"34",
          4829 => x"d2",
          4830 => x"82",
          4831 => x"af",
          4832 => x"82",
          4833 => x"54",
          4834 => x"f9",
          4835 => x"51",
          4836 => x"3f",
          4837 => x"33",
          4838 => x"73",
          4839 => x"34",
          4840 => x"06",
          4841 => x"82",
          4842 => x"82",
          4843 => x"55",
          4844 => x"2e",
          4845 => x"ff",
          4846 => x"82",
          4847 => x"74",
          4848 => x"98",
          4849 => x"ff",
          4850 => x"55",
          4851 => x"a8",
          4852 => x"54",
          4853 => x"74",
          4854 => x"51",
          4855 => x"3f",
          4856 => x"0a",
          4857 => x"0a",
          4858 => x"2c",
          4859 => x"33",
          4860 => x"75",
          4861 => x"38",
          4862 => x"a6",
          4863 => x"d2",
          4864 => x"98",
          4865 => x"2c",
          4866 => x"33",
          4867 => x"57",
          4868 => x"f8",
          4869 => x"51",
          4870 => x"3f",
          4871 => x"0a",
          4872 => x"0a",
          4873 => x"2c",
          4874 => x"33",
          4875 => x"75",
          4876 => x"38",
          4877 => x"82",
          4878 => x"70",
          4879 => x"82",
          4880 => x"59",
          4881 => x"77",
          4882 => x"38",
          4883 => x"73",
          4884 => x"34",
          4885 => x"33",
          4886 => x"a5",
          4887 => x"d2",
          4888 => x"81",
          4889 => x"d2",
          4890 => x"56",
          4891 => x"26",
          4892 => x"f6",
          4893 => x"cc",
          4894 => x"82",
          4895 => x"ef",
          4896 => x"0b",
          4897 => x"34",
          4898 => x"d2",
          4899 => x"da",
          4900 => x"38",
          4901 => x"08",
          4902 => x"2e",
          4903 => x"51",
          4904 => x"3f",
          4905 => x"08",
          4906 => x"34",
          4907 => x"08",
          4908 => x"81",
          4909 => x"52",
          4910 => x"af",
          4911 => x"5b",
          4912 => x"7a",
          4913 => x"ba",
          4914 => x"11",
          4915 => x"74",
          4916 => x"38",
          4917 => x"ad",
          4918 => x"bb",
          4919 => x"d2",
          4920 => x"bb",
          4921 => x"ff",
          4922 => x"53",
          4923 => x"51",
          4924 => x"3f",
          4925 => x"80",
          4926 => x"08",
          4927 => x"2e",
          4928 => x"74",
          4929 => x"9f",
          4930 => x"7a",
          4931 => x"81",
          4932 => x"82",
          4933 => x"55",
          4934 => x"a4",
          4935 => x"ff",
          4936 => x"82",
          4937 => x"82",
          4938 => x"82",
          4939 => x"81",
          4940 => x"05",
          4941 => x"79",
          4942 => x"cb",
          4943 => x"39",
          4944 => x"82",
          4945 => x"70",
          4946 => x"74",
          4947 => x"38",
          4948 => x"ac",
          4949 => x"bb",
          4950 => x"d2",
          4951 => x"bb",
          4952 => x"ff",
          4953 => x"53",
          4954 => x"51",
          4955 => x"3f",
          4956 => x"73",
          4957 => x"5b",
          4958 => x"82",
          4959 => x"74",
          4960 => x"d2",
          4961 => x"d2",
          4962 => x"79",
          4963 => x"3f",
          4964 => x"82",
          4965 => x"70",
          4966 => x"82",
          4967 => x"59",
          4968 => x"77",
          4969 => x"38",
          4970 => x"73",
          4971 => x"34",
          4972 => x"33",
          4973 => x"a2",
          4974 => x"ae",
          4975 => x"cc",
          4976 => x"80",
          4977 => x"38",
          4978 => x"a2",
          4979 => x"d2",
          4980 => x"05",
          4981 => x"d2",
          4982 => x"8e",
          4983 => x"0d",
          4984 => x"0b",
          4985 => x"0c",
          4986 => x"82",
          4987 => x"a0",
          4988 => x"52",
          4989 => x"51",
          4990 => x"3f",
          4991 => x"08",
          4992 => x"77",
          4993 => x"57",
          4994 => x"34",
          4995 => x"08",
          4996 => x"15",
          4997 => x"15",
          4998 => x"90",
          4999 => x"86",
          5000 => x"87",
          5001 => x"bb",
          5002 => x"bb",
          5003 => x"05",
          5004 => x"07",
          5005 => x"ff",
          5006 => x"2a",
          5007 => x"56",
          5008 => x"34",
          5009 => x"34",
          5010 => x"22",
          5011 => x"82",
          5012 => x"05",
          5013 => x"55",
          5014 => x"15",
          5015 => x"15",
          5016 => x"0d",
          5017 => x"0d",
          5018 => x"51",
          5019 => x"8f",
          5020 => x"83",
          5021 => x"70",
          5022 => x"06",
          5023 => x"70",
          5024 => x"0c",
          5025 => x"04",
          5026 => x"02",
          5027 => x"02",
          5028 => x"05",
          5029 => x"82",
          5030 => x"71",
          5031 => x"11",
          5032 => x"73",
          5033 => x"81",
          5034 => x"88",
          5035 => x"a4",
          5036 => x"22",
          5037 => x"ff",
          5038 => x"88",
          5039 => x"52",
          5040 => x"5b",
          5041 => x"55",
          5042 => x"70",
          5043 => x"82",
          5044 => x"14",
          5045 => x"52",
          5046 => x"15",
          5047 => x"15",
          5048 => x"90",
          5049 => x"70",
          5050 => x"33",
          5051 => x"07",
          5052 => x"8f",
          5053 => x"51",
          5054 => x"71",
          5055 => x"ff",
          5056 => x"88",
          5057 => x"51",
          5058 => x"34",
          5059 => x"06",
          5060 => x"12",
          5061 => x"90",
          5062 => x"71",
          5063 => x"81",
          5064 => x"3d",
          5065 => x"3d",
          5066 => x"90",
          5067 => x"05",
          5068 => x"70",
          5069 => x"11",
          5070 => x"87",
          5071 => x"8b",
          5072 => x"2b",
          5073 => x"59",
          5074 => x"72",
          5075 => x"33",
          5076 => x"71",
          5077 => x"70",
          5078 => x"56",
          5079 => x"84",
          5080 => x"85",
          5081 => x"bb",
          5082 => x"14",
          5083 => x"85",
          5084 => x"8b",
          5085 => x"2b",
          5086 => x"57",
          5087 => x"86",
          5088 => x"13",
          5089 => x"2b",
          5090 => x"2a",
          5091 => x"52",
          5092 => x"34",
          5093 => x"34",
          5094 => x"08",
          5095 => x"81",
          5096 => x"88",
          5097 => x"81",
          5098 => x"70",
          5099 => x"51",
          5100 => x"71",
          5101 => x"81",
          5102 => x"3d",
          5103 => x"3d",
          5104 => x"05",
          5105 => x"90",
          5106 => x"2b",
          5107 => x"33",
          5108 => x"71",
          5109 => x"70",
          5110 => x"70",
          5111 => x"33",
          5112 => x"71",
          5113 => x"53",
          5114 => x"52",
          5115 => x"53",
          5116 => x"25",
          5117 => x"72",
          5118 => x"3f",
          5119 => x"08",
          5120 => x"33",
          5121 => x"71",
          5122 => x"83",
          5123 => x"11",
          5124 => x"12",
          5125 => x"2b",
          5126 => x"2b",
          5127 => x"06",
          5128 => x"51",
          5129 => x"53",
          5130 => x"88",
          5131 => x"72",
          5132 => x"73",
          5133 => x"82",
          5134 => x"70",
          5135 => x"81",
          5136 => x"8b",
          5137 => x"2b",
          5138 => x"57",
          5139 => x"70",
          5140 => x"33",
          5141 => x"07",
          5142 => x"ff",
          5143 => x"2a",
          5144 => x"58",
          5145 => x"34",
          5146 => x"34",
          5147 => x"04",
          5148 => x"82",
          5149 => x"02",
          5150 => x"05",
          5151 => x"2b",
          5152 => x"11",
          5153 => x"33",
          5154 => x"71",
          5155 => x"59",
          5156 => x"56",
          5157 => x"71",
          5158 => x"33",
          5159 => x"07",
          5160 => x"a2",
          5161 => x"07",
          5162 => x"53",
          5163 => x"53",
          5164 => x"70",
          5165 => x"82",
          5166 => x"70",
          5167 => x"81",
          5168 => x"8b",
          5169 => x"2b",
          5170 => x"57",
          5171 => x"82",
          5172 => x"13",
          5173 => x"2b",
          5174 => x"2a",
          5175 => x"52",
          5176 => x"34",
          5177 => x"34",
          5178 => x"08",
          5179 => x"33",
          5180 => x"71",
          5181 => x"82",
          5182 => x"52",
          5183 => x"0d",
          5184 => x"0d",
          5185 => x"90",
          5186 => x"2a",
          5187 => x"ff",
          5188 => x"57",
          5189 => x"3f",
          5190 => x"08",
          5191 => x"71",
          5192 => x"33",
          5193 => x"71",
          5194 => x"83",
          5195 => x"11",
          5196 => x"12",
          5197 => x"2b",
          5198 => x"07",
          5199 => x"51",
          5200 => x"55",
          5201 => x"80",
          5202 => x"82",
          5203 => x"75",
          5204 => x"3f",
          5205 => x"84",
          5206 => x"15",
          5207 => x"2b",
          5208 => x"07",
          5209 => x"88",
          5210 => x"55",
          5211 => x"86",
          5212 => x"81",
          5213 => x"75",
          5214 => x"82",
          5215 => x"70",
          5216 => x"33",
          5217 => x"71",
          5218 => x"70",
          5219 => x"57",
          5220 => x"72",
          5221 => x"73",
          5222 => x"82",
          5223 => x"18",
          5224 => x"86",
          5225 => x"0b",
          5226 => x"82",
          5227 => x"53",
          5228 => x"34",
          5229 => x"34",
          5230 => x"08",
          5231 => x"81",
          5232 => x"88",
          5233 => x"82",
          5234 => x"70",
          5235 => x"51",
          5236 => x"74",
          5237 => x"81",
          5238 => x"3d",
          5239 => x"3d",
          5240 => x"82",
          5241 => x"84",
          5242 => x"3f",
          5243 => x"86",
          5244 => x"fe",
          5245 => x"3d",
          5246 => x"3d",
          5247 => x"52",
          5248 => x"3f",
          5249 => x"08",
          5250 => x"06",
          5251 => x"08",
          5252 => x"85",
          5253 => x"88",
          5254 => x"5f",
          5255 => x"5a",
          5256 => x"59",
          5257 => x"80",
          5258 => x"88",
          5259 => x"33",
          5260 => x"71",
          5261 => x"70",
          5262 => x"06",
          5263 => x"83",
          5264 => x"70",
          5265 => x"53",
          5266 => x"55",
          5267 => x"8a",
          5268 => x"2e",
          5269 => x"78",
          5270 => x"15",
          5271 => x"33",
          5272 => x"07",
          5273 => x"c2",
          5274 => x"ff",
          5275 => x"38",
          5276 => x"56",
          5277 => x"2b",
          5278 => x"08",
          5279 => x"81",
          5280 => x"88",
          5281 => x"81",
          5282 => x"51",
          5283 => x"5c",
          5284 => x"2e",
          5285 => x"55",
          5286 => x"78",
          5287 => x"38",
          5288 => x"80",
          5289 => x"38",
          5290 => x"09",
          5291 => x"38",
          5292 => x"f2",
          5293 => x"39",
          5294 => x"53",
          5295 => x"51",
          5296 => x"82",
          5297 => x"70",
          5298 => x"33",
          5299 => x"71",
          5300 => x"83",
          5301 => x"5a",
          5302 => x"05",
          5303 => x"83",
          5304 => x"70",
          5305 => x"59",
          5306 => x"84",
          5307 => x"81",
          5308 => x"76",
          5309 => x"82",
          5310 => x"75",
          5311 => x"11",
          5312 => x"11",
          5313 => x"33",
          5314 => x"07",
          5315 => x"53",
          5316 => x"5a",
          5317 => x"86",
          5318 => x"87",
          5319 => x"bb",
          5320 => x"1c",
          5321 => x"85",
          5322 => x"8b",
          5323 => x"2b",
          5324 => x"5a",
          5325 => x"54",
          5326 => x"34",
          5327 => x"34",
          5328 => x"08",
          5329 => x"1d",
          5330 => x"85",
          5331 => x"88",
          5332 => x"88",
          5333 => x"5f",
          5334 => x"73",
          5335 => x"75",
          5336 => x"82",
          5337 => x"1b",
          5338 => x"73",
          5339 => x"0c",
          5340 => x"04",
          5341 => x"74",
          5342 => x"90",
          5343 => x"f4",
          5344 => x"53",
          5345 => x"8b",
          5346 => x"fc",
          5347 => x"bb",
          5348 => x"72",
          5349 => x"0c",
          5350 => x"04",
          5351 => x"64",
          5352 => x"80",
          5353 => x"82",
          5354 => x"60",
          5355 => x"06",
          5356 => x"a9",
          5357 => x"38",
          5358 => x"b8",
          5359 => x"98",
          5360 => x"c7",
          5361 => x"38",
          5362 => x"92",
          5363 => x"83",
          5364 => x"51",
          5365 => x"82",
          5366 => x"83",
          5367 => x"82",
          5368 => x"7d",
          5369 => x"2a",
          5370 => x"ff",
          5371 => x"2b",
          5372 => x"33",
          5373 => x"71",
          5374 => x"70",
          5375 => x"83",
          5376 => x"70",
          5377 => x"05",
          5378 => x"1a",
          5379 => x"12",
          5380 => x"2b",
          5381 => x"2b",
          5382 => x"53",
          5383 => x"5c",
          5384 => x"5c",
          5385 => x"73",
          5386 => x"38",
          5387 => x"ff",
          5388 => x"70",
          5389 => x"06",
          5390 => x"16",
          5391 => x"33",
          5392 => x"07",
          5393 => x"1c",
          5394 => x"12",
          5395 => x"2b",
          5396 => x"07",
          5397 => x"52",
          5398 => x"80",
          5399 => x"78",
          5400 => x"83",
          5401 => x"41",
          5402 => x"27",
          5403 => x"60",
          5404 => x"7b",
          5405 => x"06",
          5406 => x"51",
          5407 => x"7a",
          5408 => x"06",
          5409 => x"39",
          5410 => x"7a",
          5411 => x"38",
          5412 => x"aa",
          5413 => x"39",
          5414 => x"7a",
          5415 => x"c8",
          5416 => x"82",
          5417 => x"12",
          5418 => x"2b",
          5419 => x"54",
          5420 => x"80",
          5421 => x"f7",
          5422 => x"bb",
          5423 => x"ff",
          5424 => x"54",
          5425 => x"83",
          5426 => x"90",
          5427 => x"05",
          5428 => x"ff",
          5429 => x"82",
          5430 => x"14",
          5431 => x"83",
          5432 => x"59",
          5433 => x"39",
          5434 => x"7a",
          5435 => x"d4",
          5436 => x"f5",
          5437 => x"bb",
          5438 => x"82",
          5439 => x"12",
          5440 => x"2b",
          5441 => x"54",
          5442 => x"80",
          5443 => x"f6",
          5444 => x"bb",
          5445 => x"ff",
          5446 => x"54",
          5447 => x"83",
          5448 => x"90",
          5449 => x"05",
          5450 => x"ff",
          5451 => x"82",
          5452 => x"14",
          5453 => x"62",
          5454 => x"5c",
          5455 => x"ff",
          5456 => x"39",
          5457 => x"54",
          5458 => x"82",
          5459 => x"5c",
          5460 => x"08",
          5461 => x"38",
          5462 => x"52",
          5463 => x"08",
          5464 => x"a3",
          5465 => x"f7",
          5466 => x"58",
          5467 => x"99",
          5468 => x"7a",
          5469 => x"f2",
          5470 => x"19",
          5471 => x"bb",
          5472 => x"84",
          5473 => x"f9",
          5474 => x"73",
          5475 => x"0c",
          5476 => x"04",
          5477 => x"77",
          5478 => x"52",
          5479 => x"3f",
          5480 => x"08",
          5481 => x"98",
          5482 => x"8e",
          5483 => x"80",
          5484 => x"98",
          5485 => x"a2",
          5486 => x"82",
          5487 => x"86",
          5488 => x"ff",
          5489 => x"8f",
          5490 => x"81",
          5491 => x"26",
          5492 => x"bb",
          5493 => x"52",
          5494 => x"98",
          5495 => x"0d",
          5496 => x"0d",
          5497 => x"33",
          5498 => x"9f",
          5499 => x"53",
          5500 => x"81",
          5501 => x"38",
          5502 => x"87",
          5503 => x"11",
          5504 => x"54",
          5505 => x"84",
          5506 => x"54",
          5507 => x"87",
          5508 => x"11",
          5509 => x"0c",
          5510 => x"c0",
          5511 => x"70",
          5512 => x"70",
          5513 => x"51",
          5514 => x"8a",
          5515 => x"98",
          5516 => x"70",
          5517 => x"08",
          5518 => x"06",
          5519 => x"38",
          5520 => x"8c",
          5521 => x"80",
          5522 => x"71",
          5523 => x"14",
          5524 => x"94",
          5525 => x"70",
          5526 => x"0c",
          5527 => x"04",
          5528 => x"60",
          5529 => x"8c",
          5530 => x"33",
          5531 => x"5b",
          5532 => x"5a",
          5533 => x"82",
          5534 => x"81",
          5535 => x"52",
          5536 => x"38",
          5537 => x"84",
          5538 => x"92",
          5539 => x"c0",
          5540 => x"87",
          5541 => x"13",
          5542 => x"57",
          5543 => x"0b",
          5544 => x"8c",
          5545 => x"0c",
          5546 => x"75",
          5547 => x"2a",
          5548 => x"51",
          5549 => x"80",
          5550 => x"7b",
          5551 => x"7b",
          5552 => x"5d",
          5553 => x"59",
          5554 => x"06",
          5555 => x"73",
          5556 => x"81",
          5557 => x"ff",
          5558 => x"72",
          5559 => x"38",
          5560 => x"8c",
          5561 => x"c3",
          5562 => x"98",
          5563 => x"71",
          5564 => x"38",
          5565 => x"2e",
          5566 => x"76",
          5567 => x"92",
          5568 => x"72",
          5569 => x"06",
          5570 => x"f7",
          5571 => x"5a",
          5572 => x"80",
          5573 => x"70",
          5574 => x"5a",
          5575 => x"80",
          5576 => x"73",
          5577 => x"06",
          5578 => x"38",
          5579 => x"fe",
          5580 => x"fc",
          5581 => x"52",
          5582 => x"83",
          5583 => x"71",
          5584 => x"bb",
          5585 => x"3d",
          5586 => x"3d",
          5587 => x"64",
          5588 => x"bf",
          5589 => x"40",
          5590 => x"59",
          5591 => x"58",
          5592 => x"82",
          5593 => x"81",
          5594 => x"52",
          5595 => x"09",
          5596 => x"b1",
          5597 => x"84",
          5598 => x"92",
          5599 => x"c0",
          5600 => x"87",
          5601 => x"13",
          5602 => x"56",
          5603 => x"87",
          5604 => x"0c",
          5605 => x"82",
          5606 => x"58",
          5607 => x"84",
          5608 => x"06",
          5609 => x"71",
          5610 => x"38",
          5611 => x"05",
          5612 => x"0c",
          5613 => x"73",
          5614 => x"81",
          5615 => x"71",
          5616 => x"38",
          5617 => x"8c",
          5618 => x"d0",
          5619 => x"98",
          5620 => x"71",
          5621 => x"38",
          5622 => x"2e",
          5623 => x"76",
          5624 => x"92",
          5625 => x"72",
          5626 => x"06",
          5627 => x"f7",
          5628 => x"59",
          5629 => x"1a",
          5630 => x"06",
          5631 => x"59",
          5632 => x"80",
          5633 => x"73",
          5634 => x"06",
          5635 => x"38",
          5636 => x"fe",
          5637 => x"fc",
          5638 => x"52",
          5639 => x"83",
          5640 => x"71",
          5641 => x"bb",
          5642 => x"3d",
          5643 => x"3d",
          5644 => x"84",
          5645 => x"33",
          5646 => x"a7",
          5647 => x"54",
          5648 => x"fa",
          5649 => x"bb",
          5650 => x"06",
          5651 => x"72",
          5652 => x"85",
          5653 => x"98",
          5654 => x"56",
          5655 => x"80",
          5656 => x"76",
          5657 => x"74",
          5658 => x"c0",
          5659 => x"54",
          5660 => x"2e",
          5661 => x"d4",
          5662 => x"2e",
          5663 => x"80",
          5664 => x"08",
          5665 => x"70",
          5666 => x"51",
          5667 => x"2e",
          5668 => x"c0",
          5669 => x"52",
          5670 => x"87",
          5671 => x"08",
          5672 => x"38",
          5673 => x"87",
          5674 => x"14",
          5675 => x"70",
          5676 => x"52",
          5677 => x"96",
          5678 => x"92",
          5679 => x"0a",
          5680 => x"39",
          5681 => x"0c",
          5682 => x"39",
          5683 => x"54",
          5684 => x"98",
          5685 => x"0d",
          5686 => x"0d",
          5687 => x"33",
          5688 => x"88",
          5689 => x"bb",
          5690 => x"51",
          5691 => x"04",
          5692 => x"75",
          5693 => x"82",
          5694 => x"90",
          5695 => x"2b",
          5696 => x"33",
          5697 => x"88",
          5698 => x"71",
          5699 => x"98",
          5700 => x"54",
          5701 => x"85",
          5702 => x"ff",
          5703 => x"02",
          5704 => x"05",
          5705 => x"70",
          5706 => x"05",
          5707 => x"88",
          5708 => x"72",
          5709 => x"0d",
          5710 => x"0d",
          5711 => x"52",
          5712 => x"81",
          5713 => x"70",
          5714 => x"70",
          5715 => x"05",
          5716 => x"88",
          5717 => x"72",
          5718 => x"54",
          5719 => x"2a",
          5720 => x"34",
          5721 => x"04",
          5722 => x"76",
          5723 => x"54",
          5724 => x"2e",
          5725 => x"70",
          5726 => x"33",
          5727 => x"05",
          5728 => x"11",
          5729 => x"84",
          5730 => x"fe",
          5731 => x"77",
          5732 => x"53",
          5733 => x"81",
          5734 => x"ff",
          5735 => x"f4",
          5736 => x"0d",
          5737 => x"0d",
          5738 => x"56",
          5739 => x"70",
          5740 => x"33",
          5741 => x"05",
          5742 => x"71",
          5743 => x"56",
          5744 => x"72",
          5745 => x"38",
          5746 => x"e2",
          5747 => x"bb",
          5748 => x"3d",
          5749 => x"3d",
          5750 => x"54",
          5751 => x"71",
          5752 => x"38",
          5753 => x"70",
          5754 => x"f3",
          5755 => x"82",
          5756 => x"84",
          5757 => x"80",
          5758 => x"98",
          5759 => x"0b",
          5760 => x"0c",
          5761 => x"0d",
          5762 => x"0b",
          5763 => x"56",
          5764 => x"2e",
          5765 => x"81",
          5766 => x"08",
          5767 => x"70",
          5768 => x"33",
          5769 => x"a2",
          5770 => x"98",
          5771 => x"09",
          5772 => x"38",
          5773 => x"08",
          5774 => x"b0",
          5775 => x"a4",
          5776 => x"9c",
          5777 => x"56",
          5778 => x"27",
          5779 => x"16",
          5780 => x"82",
          5781 => x"06",
          5782 => x"54",
          5783 => x"78",
          5784 => x"33",
          5785 => x"3f",
          5786 => x"5a",
          5787 => x"98",
          5788 => x"0d",
          5789 => x"0d",
          5790 => x"56",
          5791 => x"b0",
          5792 => x"af",
          5793 => x"fe",
          5794 => x"bb",
          5795 => x"82",
          5796 => x"9f",
          5797 => x"74",
          5798 => x"52",
          5799 => x"51",
          5800 => x"82",
          5801 => x"80",
          5802 => x"ff",
          5803 => x"74",
          5804 => x"76",
          5805 => x"0c",
          5806 => x"04",
          5807 => x"7a",
          5808 => x"fe",
          5809 => x"bb",
          5810 => x"82",
          5811 => x"81",
          5812 => x"33",
          5813 => x"2e",
          5814 => x"80",
          5815 => x"17",
          5816 => x"81",
          5817 => x"06",
          5818 => x"84",
          5819 => x"bb",
          5820 => x"b4",
          5821 => x"56",
          5822 => x"82",
          5823 => x"84",
          5824 => x"fc",
          5825 => x"8b",
          5826 => x"52",
          5827 => x"a9",
          5828 => x"85",
          5829 => x"84",
          5830 => x"fc",
          5831 => x"17",
          5832 => x"9c",
          5833 => x"91",
          5834 => x"08",
          5835 => x"17",
          5836 => x"3f",
          5837 => x"81",
          5838 => x"19",
          5839 => x"53",
          5840 => x"17",
          5841 => x"82",
          5842 => x"18",
          5843 => x"80",
          5844 => x"33",
          5845 => x"3f",
          5846 => x"08",
          5847 => x"38",
          5848 => x"82",
          5849 => x"8a",
          5850 => x"fb",
          5851 => x"fe",
          5852 => x"08",
          5853 => x"56",
          5854 => x"74",
          5855 => x"38",
          5856 => x"75",
          5857 => x"16",
          5858 => x"53",
          5859 => x"98",
          5860 => x"0d",
          5861 => x"0d",
          5862 => x"08",
          5863 => x"81",
          5864 => x"df",
          5865 => x"15",
          5866 => x"d7",
          5867 => x"33",
          5868 => x"82",
          5869 => x"38",
          5870 => x"89",
          5871 => x"2e",
          5872 => x"bf",
          5873 => x"2e",
          5874 => x"81",
          5875 => x"81",
          5876 => x"89",
          5877 => x"08",
          5878 => x"52",
          5879 => x"3f",
          5880 => x"08",
          5881 => x"74",
          5882 => x"14",
          5883 => x"81",
          5884 => x"2a",
          5885 => x"05",
          5886 => x"57",
          5887 => x"f5",
          5888 => x"98",
          5889 => x"38",
          5890 => x"06",
          5891 => x"33",
          5892 => x"78",
          5893 => x"06",
          5894 => x"5c",
          5895 => x"53",
          5896 => x"38",
          5897 => x"06",
          5898 => x"39",
          5899 => x"a4",
          5900 => x"52",
          5901 => x"bd",
          5902 => x"98",
          5903 => x"38",
          5904 => x"fe",
          5905 => x"b4",
          5906 => x"8d",
          5907 => x"98",
          5908 => x"ff",
          5909 => x"39",
          5910 => x"a4",
          5911 => x"52",
          5912 => x"91",
          5913 => x"98",
          5914 => x"76",
          5915 => x"fc",
          5916 => x"b4",
          5917 => x"f8",
          5918 => x"98",
          5919 => x"06",
          5920 => x"81",
          5921 => x"bb",
          5922 => x"3d",
          5923 => x"3d",
          5924 => x"7e",
          5925 => x"82",
          5926 => x"27",
          5927 => x"76",
          5928 => x"27",
          5929 => x"75",
          5930 => x"79",
          5931 => x"38",
          5932 => x"89",
          5933 => x"2e",
          5934 => x"80",
          5935 => x"2e",
          5936 => x"81",
          5937 => x"81",
          5938 => x"89",
          5939 => x"08",
          5940 => x"52",
          5941 => x"3f",
          5942 => x"08",
          5943 => x"98",
          5944 => x"38",
          5945 => x"06",
          5946 => x"81",
          5947 => x"06",
          5948 => x"77",
          5949 => x"2e",
          5950 => x"84",
          5951 => x"06",
          5952 => x"06",
          5953 => x"53",
          5954 => x"81",
          5955 => x"34",
          5956 => x"a4",
          5957 => x"52",
          5958 => x"d9",
          5959 => x"98",
          5960 => x"bb",
          5961 => x"94",
          5962 => x"ff",
          5963 => x"05",
          5964 => x"54",
          5965 => x"38",
          5966 => x"74",
          5967 => x"06",
          5968 => x"07",
          5969 => x"74",
          5970 => x"39",
          5971 => x"a4",
          5972 => x"52",
          5973 => x"9d",
          5974 => x"98",
          5975 => x"bb",
          5976 => x"d8",
          5977 => x"ff",
          5978 => x"76",
          5979 => x"06",
          5980 => x"05",
          5981 => x"3f",
          5982 => x"87",
          5983 => x"08",
          5984 => x"51",
          5985 => x"82",
          5986 => x"59",
          5987 => x"08",
          5988 => x"f0",
          5989 => x"82",
          5990 => x"06",
          5991 => x"05",
          5992 => x"54",
          5993 => x"3f",
          5994 => x"08",
          5995 => x"74",
          5996 => x"51",
          5997 => x"81",
          5998 => x"34",
          5999 => x"98",
          6000 => x"0d",
          6001 => x"0d",
          6002 => x"72",
          6003 => x"56",
          6004 => x"27",
          6005 => x"98",
          6006 => x"9d",
          6007 => x"2e",
          6008 => x"53",
          6009 => x"51",
          6010 => x"82",
          6011 => x"54",
          6012 => x"08",
          6013 => x"93",
          6014 => x"80",
          6015 => x"54",
          6016 => x"82",
          6017 => x"54",
          6018 => x"74",
          6019 => x"fb",
          6020 => x"bb",
          6021 => x"82",
          6022 => x"80",
          6023 => x"38",
          6024 => x"08",
          6025 => x"38",
          6026 => x"08",
          6027 => x"38",
          6028 => x"52",
          6029 => x"d6",
          6030 => x"98",
          6031 => x"98",
          6032 => x"11",
          6033 => x"57",
          6034 => x"74",
          6035 => x"81",
          6036 => x"0c",
          6037 => x"81",
          6038 => x"84",
          6039 => x"55",
          6040 => x"ff",
          6041 => x"54",
          6042 => x"98",
          6043 => x"0d",
          6044 => x"0d",
          6045 => x"08",
          6046 => x"79",
          6047 => x"17",
          6048 => x"80",
          6049 => x"98",
          6050 => x"26",
          6051 => x"58",
          6052 => x"52",
          6053 => x"fd",
          6054 => x"74",
          6055 => x"08",
          6056 => x"38",
          6057 => x"08",
          6058 => x"98",
          6059 => x"82",
          6060 => x"17",
          6061 => x"98",
          6062 => x"c7",
          6063 => x"90",
          6064 => x"56",
          6065 => x"2e",
          6066 => x"77",
          6067 => x"81",
          6068 => x"38",
          6069 => x"98",
          6070 => x"26",
          6071 => x"56",
          6072 => x"51",
          6073 => x"80",
          6074 => x"98",
          6075 => x"09",
          6076 => x"38",
          6077 => x"08",
          6078 => x"98",
          6079 => x"30",
          6080 => x"80",
          6081 => x"07",
          6082 => x"08",
          6083 => x"55",
          6084 => x"ef",
          6085 => x"98",
          6086 => x"95",
          6087 => x"08",
          6088 => x"27",
          6089 => x"98",
          6090 => x"89",
          6091 => x"85",
          6092 => x"db",
          6093 => x"81",
          6094 => x"17",
          6095 => x"89",
          6096 => x"75",
          6097 => x"ac",
          6098 => x"7a",
          6099 => x"3f",
          6100 => x"08",
          6101 => x"38",
          6102 => x"bb",
          6103 => x"2e",
          6104 => x"86",
          6105 => x"98",
          6106 => x"bb",
          6107 => x"70",
          6108 => x"07",
          6109 => x"7c",
          6110 => x"55",
          6111 => x"f8",
          6112 => x"2e",
          6113 => x"ff",
          6114 => x"55",
          6115 => x"ff",
          6116 => x"76",
          6117 => x"3f",
          6118 => x"08",
          6119 => x"08",
          6120 => x"bb",
          6121 => x"80",
          6122 => x"55",
          6123 => x"94",
          6124 => x"2e",
          6125 => x"53",
          6126 => x"51",
          6127 => x"82",
          6128 => x"55",
          6129 => x"75",
          6130 => x"98",
          6131 => x"05",
          6132 => x"56",
          6133 => x"26",
          6134 => x"15",
          6135 => x"84",
          6136 => x"07",
          6137 => x"18",
          6138 => x"ff",
          6139 => x"2e",
          6140 => x"39",
          6141 => x"39",
          6142 => x"08",
          6143 => x"81",
          6144 => x"74",
          6145 => x"0c",
          6146 => x"04",
          6147 => x"7a",
          6148 => x"f3",
          6149 => x"bb",
          6150 => x"81",
          6151 => x"98",
          6152 => x"38",
          6153 => x"51",
          6154 => x"82",
          6155 => x"82",
          6156 => x"b0",
          6157 => x"84",
          6158 => x"52",
          6159 => x"52",
          6160 => x"3f",
          6161 => x"39",
          6162 => x"8a",
          6163 => x"75",
          6164 => x"38",
          6165 => x"19",
          6166 => x"81",
          6167 => x"ed",
          6168 => x"bb",
          6169 => x"2e",
          6170 => x"15",
          6171 => x"70",
          6172 => x"07",
          6173 => x"53",
          6174 => x"75",
          6175 => x"0c",
          6176 => x"04",
          6177 => x"7a",
          6178 => x"58",
          6179 => x"f0",
          6180 => x"80",
          6181 => x"9f",
          6182 => x"80",
          6183 => x"90",
          6184 => x"17",
          6185 => x"aa",
          6186 => x"53",
          6187 => x"88",
          6188 => x"08",
          6189 => x"38",
          6190 => x"53",
          6191 => x"17",
          6192 => x"72",
          6193 => x"fe",
          6194 => x"08",
          6195 => x"80",
          6196 => x"16",
          6197 => x"2b",
          6198 => x"75",
          6199 => x"73",
          6200 => x"f5",
          6201 => x"bb",
          6202 => x"82",
          6203 => x"ff",
          6204 => x"81",
          6205 => x"98",
          6206 => x"38",
          6207 => x"82",
          6208 => x"26",
          6209 => x"58",
          6210 => x"73",
          6211 => x"39",
          6212 => x"51",
          6213 => x"82",
          6214 => x"98",
          6215 => x"94",
          6216 => x"17",
          6217 => x"58",
          6218 => x"9a",
          6219 => x"81",
          6220 => x"74",
          6221 => x"98",
          6222 => x"83",
          6223 => x"b4",
          6224 => x"0c",
          6225 => x"82",
          6226 => x"8a",
          6227 => x"f8",
          6228 => x"70",
          6229 => x"08",
          6230 => x"57",
          6231 => x"0a",
          6232 => x"38",
          6233 => x"15",
          6234 => x"08",
          6235 => x"72",
          6236 => x"cb",
          6237 => x"ff",
          6238 => x"81",
          6239 => x"13",
          6240 => x"94",
          6241 => x"74",
          6242 => x"85",
          6243 => x"22",
          6244 => x"73",
          6245 => x"38",
          6246 => x"8a",
          6247 => x"05",
          6248 => x"06",
          6249 => x"8a",
          6250 => x"73",
          6251 => x"3f",
          6252 => x"08",
          6253 => x"81",
          6254 => x"98",
          6255 => x"ff",
          6256 => x"82",
          6257 => x"ff",
          6258 => x"38",
          6259 => x"82",
          6260 => x"26",
          6261 => x"7b",
          6262 => x"98",
          6263 => x"55",
          6264 => x"94",
          6265 => x"73",
          6266 => x"3f",
          6267 => x"08",
          6268 => x"82",
          6269 => x"80",
          6270 => x"38",
          6271 => x"bb",
          6272 => x"2e",
          6273 => x"55",
          6274 => x"08",
          6275 => x"38",
          6276 => x"08",
          6277 => x"fb",
          6278 => x"bb",
          6279 => x"38",
          6280 => x"0c",
          6281 => x"51",
          6282 => x"82",
          6283 => x"98",
          6284 => x"90",
          6285 => x"16",
          6286 => x"15",
          6287 => x"74",
          6288 => x"0c",
          6289 => x"04",
          6290 => x"7b",
          6291 => x"5b",
          6292 => x"52",
          6293 => x"ac",
          6294 => x"98",
          6295 => x"bb",
          6296 => x"ec",
          6297 => x"98",
          6298 => x"17",
          6299 => x"51",
          6300 => x"82",
          6301 => x"54",
          6302 => x"08",
          6303 => x"82",
          6304 => x"9c",
          6305 => x"33",
          6306 => x"72",
          6307 => x"09",
          6308 => x"38",
          6309 => x"bb",
          6310 => x"72",
          6311 => x"55",
          6312 => x"53",
          6313 => x"8e",
          6314 => x"56",
          6315 => x"09",
          6316 => x"38",
          6317 => x"bb",
          6318 => x"81",
          6319 => x"fd",
          6320 => x"bb",
          6321 => x"82",
          6322 => x"80",
          6323 => x"38",
          6324 => x"09",
          6325 => x"38",
          6326 => x"82",
          6327 => x"8b",
          6328 => x"fd",
          6329 => x"9a",
          6330 => x"eb",
          6331 => x"bb",
          6332 => x"ff",
          6333 => x"70",
          6334 => x"53",
          6335 => x"09",
          6336 => x"38",
          6337 => x"eb",
          6338 => x"bb",
          6339 => x"2b",
          6340 => x"72",
          6341 => x"0c",
          6342 => x"04",
          6343 => x"77",
          6344 => x"ff",
          6345 => x"9a",
          6346 => x"55",
          6347 => x"76",
          6348 => x"53",
          6349 => x"09",
          6350 => x"38",
          6351 => x"52",
          6352 => x"eb",
          6353 => x"3d",
          6354 => x"3d",
          6355 => x"5b",
          6356 => x"08",
          6357 => x"15",
          6358 => x"81",
          6359 => x"15",
          6360 => x"51",
          6361 => x"82",
          6362 => x"58",
          6363 => x"08",
          6364 => x"9c",
          6365 => x"33",
          6366 => x"86",
          6367 => x"80",
          6368 => x"13",
          6369 => x"06",
          6370 => x"06",
          6371 => x"72",
          6372 => x"82",
          6373 => x"53",
          6374 => x"2e",
          6375 => x"53",
          6376 => x"a9",
          6377 => x"74",
          6378 => x"72",
          6379 => x"38",
          6380 => x"99",
          6381 => x"98",
          6382 => x"06",
          6383 => x"88",
          6384 => x"06",
          6385 => x"54",
          6386 => x"a0",
          6387 => x"74",
          6388 => x"3f",
          6389 => x"08",
          6390 => x"98",
          6391 => x"98",
          6392 => x"fa",
          6393 => x"80",
          6394 => x"0c",
          6395 => x"98",
          6396 => x"0d",
          6397 => x"0d",
          6398 => x"57",
          6399 => x"73",
          6400 => x"3f",
          6401 => x"08",
          6402 => x"98",
          6403 => x"98",
          6404 => x"75",
          6405 => x"3f",
          6406 => x"08",
          6407 => x"98",
          6408 => x"a0",
          6409 => x"98",
          6410 => x"14",
          6411 => x"db",
          6412 => x"a0",
          6413 => x"14",
          6414 => x"ac",
          6415 => x"83",
          6416 => x"82",
          6417 => x"87",
          6418 => x"fd",
          6419 => x"70",
          6420 => x"08",
          6421 => x"55",
          6422 => x"3f",
          6423 => x"08",
          6424 => x"13",
          6425 => x"73",
          6426 => x"83",
          6427 => x"3d",
          6428 => x"3d",
          6429 => x"57",
          6430 => x"89",
          6431 => x"17",
          6432 => x"81",
          6433 => x"70",
          6434 => x"55",
          6435 => x"08",
          6436 => x"81",
          6437 => x"52",
          6438 => x"a8",
          6439 => x"2e",
          6440 => x"84",
          6441 => x"52",
          6442 => x"09",
          6443 => x"38",
          6444 => x"81",
          6445 => x"81",
          6446 => x"73",
          6447 => x"55",
          6448 => x"55",
          6449 => x"c5",
          6450 => x"88",
          6451 => x"0b",
          6452 => x"9c",
          6453 => x"8b",
          6454 => x"17",
          6455 => x"08",
          6456 => x"52",
          6457 => x"82",
          6458 => x"76",
          6459 => x"51",
          6460 => x"82",
          6461 => x"86",
          6462 => x"12",
          6463 => x"3f",
          6464 => x"08",
          6465 => x"88",
          6466 => x"f3",
          6467 => x"70",
          6468 => x"80",
          6469 => x"51",
          6470 => x"af",
          6471 => x"81",
          6472 => x"dc",
          6473 => x"74",
          6474 => x"38",
          6475 => x"88",
          6476 => x"39",
          6477 => x"80",
          6478 => x"56",
          6479 => x"af",
          6480 => x"06",
          6481 => x"56",
          6482 => x"32",
          6483 => x"80",
          6484 => x"51",
          6485 => x"dc",
          6486 => x"1c",
          6487 => x"33",
          6488 => x"9f",
          6489 => x"ff",
          6490 => x"1c",
          6491 => x"7a",
          6492 => x"3f",
          6493 => x"08",
          6494 => x"39",
          6495 => x"a0",
          6496 => x"5e",
          6497 => x"52",
          6498 => x"ff",
          6499 => x"59",
          6500 => x"33",
          6501 => x"ae",
          6502 => x"06",
          6503 => x"78",
          6504 => x"81",
          6505 => x"32",
          6506 => x"9f",
          6507 => x"26",
          6508 => x"53",
          6509 => x"73",
          6510 => x"17",
          6511 => x"34",
          6512 => x"db",
          6513 => x"32",
          6514 => x"9f",
          6515 => x"54",
          6516 => x"2e",
          6517 => x"80",
          6518 => x"75",
          6519 => x"bd",
          6520 => x"7e",
          6521 => x"a0",
          6522 => x"bd",
          6523 => x"82",
          6524 => x"18",
          6525 => x"1a",
          6526 => x"a0",
          6527 => x"fc",
          6528 => x"32",
          6529 => x"80",
          6530 => x"30",
          6531 => x"71",
          6532 => x"51",
          6533 => x"55",
          6534 => x"ac",
          6535 => x"81",
          6536 => x"78",
          6537 => x"51",
          6538 => x"af",
          6539 => x"06",
          6540 => x"55",
          6541 => x"32",
          6542 => x"80",
          6543 => x"51",
          6544 => x"db",
          6545 => x"39",
          6546 => x"09",
          6547 => x"38",
          6548 => x"7c",
          6549 => x"54",
          6550 => x"a2",
          6551 => x"32",
          6552 => x"ae",
          6553 => x"72",
          6554 => x"9f",
          6555 => x"51",
          6556 => x"74",
          6557 => x"88",
          6558 => x"fe",
          6559 => x"98",
          6560 => x"80",
          6561 => x"75",
          6562 => x"82",
          6563 => x"33",
          6564 => x"51",
          6565 => x"82",
          6566 => x"80",
          6567 => x"78",
          6568 => x"81",
          6569 => x"5a",
          6570 => x"d2",
          6571 => x"98",
          6572 => x"80",
          6573 => x"1c",
          6574 => x"27",
          6575 => x"79",
          6576 => x"74",
          6577 => x"7a",
          6578 => x"74",
          6579 => x"39",
          6580 => x"b4",
          6581 => x"fe",
          6582 => x"98",
          6583 => x"ff",
          6584 => x"73",
          6585 => x"38",
          6586 => x"81",
          6587 => x"54",
          6588 => x"75",
          6589 => x"17",
          6590 => x"39",
          6591 => x"0c",
          6592 => x"99",
          6593 => x"54",
          6594 => x"2e",
          6595 => x"84",
          6596 => x"34",
          6597 => x"76",
          6598 => x"8b",
          6599 => x"81",
          6600 => x"56",
          6601 => x"80",
          6602 => x"1b",
          6603 => x"08",
          6604 => x"51",
          6605 => x"82",
          6606 => x"56",
          6607 => x"08",
          6608 => x"98",
          6609 => x"76",
          6610 => x"3f",
          6611 => x"08",
          6612 => x"98",
          6613 => x"38",
          6614 => x"70",
          6615 => x"73",
          6616 => x"be",
          6617 => x"33",
          6618 => x"73",
          6619 => x"8b",
          6620 => x"83",
          6621 => x"06",
          6622 => x"73",
          6623 => x"53",
          6624 => x"51",
          6625 => x"82",
          6626 => x"80",
          6627 => x"75",
          6628 => x"f3",
          6629 => x"9f",
          6630 => x"1c",
          6631 => x"74",
          6632 => x"38",
          6633 => x"09",
          6634 => x"e7",
          6635 => x"2a",
          6636 => x"77",
          6637 => x"51",
          6638 => x"2e",
          6639 => x"81",
          6640 => x"80",
          6641 => x"38",
          6642 => x"ab",
          6643 => x"55",
          6644 => x"75",
          6645 => x"73",
          6646 => x"55",
          6647 => x"82",
          6648 => x"06",
          6649 => x"ab",
          6650 => x"33",
          6651 => x"70",
          6652 => x"55",
          6653 => x"2e",
          6654 => x"1b",
          6655 => x"06",
          6656 => x"52",
          6657 => x"db",
          6658 => x"98",
          6659 => x"0c",
          6660 => x"74",
          6661 => x"0c",
          6662 => x"04",
          6663 => x"7c",
          6664 => x"08",
          6665 => x"55",
          6666 => x"59",
          6667 => x"81",
          6668 => x"70",
          6669 => x"33",
          6670 => x"52",
          6671 => x"2e",
          6672 => x"ee",
          6673 => x"2e",
          6674 => x"81",
          6675 => x"33",
          6676 => x"81",
          6677 => x"52",
          6678 => x"26",
          6679 => x"14",
          6680 => x"06",
          6681 => x"52",
          6682 => x"80",
          6683 => x"0b",
          6684 => x"59",
          6685 => x"7a",
          6686 => x"70",
          6687 => x"33",
          6688 => x"05",
          6689 => x"9f",
          6690 => x"53",
          6691 => x"89",
          6692 => x"70",
          6693 => x"54",
          6694 => x"12",
          6695 => x"26",
          6696 => x"12",
          6697 => x"06",
          6698 => x"30",
          6699 => x"51",
          6700 => x"2e",
          6701 => x"85",
          6702 => x"be",
          6703 => x"74",
          6704 => x"30",
          6705 => x"9f",
          6706 => x"2a",
          6707 => x"54",
          6708 => x"2e",
          6709 => x"15",
          6710 => x"55",
          6711 => x"ff",
          6712 => x"39",
          6713 => x"86",
          6714 => x"7c",
          6715 => x"51",
          6716 => x"d2",
          6717 => x"70",
          6718 => x"0c",
          6719 => x"04",
          6720 => x"78",
          6721 => x"83",
          6722 => x"0b",
          6723 => x"79",
          6724 => x"e2",
          6725 => x"55",
          6726 => x"08",
          6727 => x"84",
          6728 => x"df",
          6729 => x"bb",
          6730 => x"ff",
          6731 => x"83",
          6732 => x"d4",
          6733 => x"81",
          6734 => x"38",
          6735 => x"17",
          6736 => x"74",
          6737 => x"09",
          6738 => x"38",
          6739 => x"81",
          6740 => x"30",
          6741 => x"79",
          6742 => x"54",
          6743 => x"74",
          6744 => x"09",
          6745 => x"38",
          6746 => x"b4",
          6747 => x"ea",
          6748 => x"b1",
          6749 => x"98",
          6750 => x"bb",
          6751 => x"2e",
          6752 => x"53",
          6753 => x"52",
          6754 => x"51",
          6755 => x"82",
          6756 => x"55",
          6757 => x"08",
          6758 => x"38",
          6759 => x"82",
          6760 => x"88",
          6761 => x"f2",
          6762 => x"02",
          6763 => x"cb",
          6764 => x"55",
          6765 => x"60",
          6766 => x"3f",
          6767 => x"08",
          6768 => x"80",
          6769 => x"98",
          6770 => x"fc",
          6771 => x"98",
          6772 => x"82",
          6773 => x"70",
          6774 => x"8c",
          6775 => x"2e",
          6776 => x"73",
          6777 => x"81",
          6778 => x"33",
          6779 => x"80",
          6780 => x"81",
          6781 => x"d7",
          6782 => x"bb",
          6783 => x"ff",
          6784 => x"06",
          6785 => x"98",
          6786 => x"2e",
          6787 => x"74",
          6788 => x"81",
          6789 => x"8a",
          6790 => x"ac",
          6791 => x"39",
          6792 => x"77",
          6793 => x"81",
          6794 => x"33",
          6795 => x"3f",
          6796 => x"08",
          6797 => x"70",
          6798 => x"55",
          6799 => x"86",
          6800 => x"80",
          6801 => x"74",
          6802 => x"81",
          6803 => x"8a",
          6804 => x"f4",
          6805 => x"53",
          6806 => x"fd",
          6807 => x"bb",
          6808 => x"ff",
          6809 => x"82",
          6810 => x"06",
          6811 => x"8c",
          6812 => x"58",
          6813 => x"f6",
          6814 => x"58",
          6815 => x"2e",
          6816 => x"fa",
          6817 => x"e8",
          6818 => x"98",
          6819 => x"78",
          6820 => x"5a",
          6821 => x"90",
          6822 => x"75",
          6823 => x"38",
          6824 => x"3d",
          6825 => x"70",
          6826 => x"08",
          6827 => x"7a",
          6828 => x"38",
          6829 => x"51",
          6830 => x"82",
          6831 => x"81",
          6832 => x"81",
          6833 => x"38",
          6834 => x"83",
          6835 => x"38",
          6836 => x"84",
          6837 => x"38",
          6838 => x"81",
          6839 => x"38",
          6840 => x"db",
          6841 => x"bb",
          6842 => x"ff",
          6843 => x"72",
          6844 => x"09",
          6845 => x"d0",
          6846 => x"14",
          6847 => x"3f",
          6848 => x"08",
          6849 => x"06",
          6850 => x"38",
          6851 => x"51",
          6852 => x"82",
          6853 => x"58",
          6854 => x"0c",
          6855 => x"33",
          6856 => x"80",
          6857 => x"ff",
          6858 => x"ff",
          6859 => x"55",
          6860 => x"81",
          6861 => x"38",
          6862 => x"06",
          6863 => x"80",
          6864 => x"52",
          6865 => x"8a",
          6866 => x"80",
          6867 => x"ff",
          6868 => x"53",
          6869 => x"86",
          6870 => x"83",
          6871 => x"c5",
          6872 => x"f5",
          6873 => x"98",
          6874 => x"bb",
          6875 => x"15",
          6876 => x"06",
          6877 => x"76",
          6878 => x"80",
          6879 => x"da",
          6880 => x"bb",
          6881 => x"ff",
          6882 => x"74",
          6883 => x"d4",
          6884 => x"dc",
          6885 => x"98",
          6886 => x"c2",
          6887 => x"b9",
          6888 => x"98",
          6889 => x"ff",
          6890 => x"56",
          6891 => x"83",
          6892 => x"14",
          6893 => x"71",
          6894 => x"5a",
          6895 => x"26",
          6896 => x"8a",
          6897 => x"74",
          6898 => x"fe",
          6899 => x"82",
          6900 => x"55",
          6901 => x"08",
          6902 => x"ec",
          6903 => x"98",
          6904 => x"ff",
          6905 => x"83",
          6906 => x"74",
          6907 => x"26",
          6908 => x"57",
          6909 => x"26",
          6910 => x"57",
          6911 => x"56",
          6912 => x"82",
          6913 => x"15",
          6914 => x"0c",
          6915 => x"0c",
          6916 => x"a4",
          6917 => x"1d",
          6918 => x"54",
          6919 => x"2e",
          6920 => x"af",
          6921 => x"14",
          6922 => x"3f",
          6923 => x"08",
          6924 => x"06",
          6925 => x"72",
          6926 => x"79",
          6927 => x"80",
          6928 => x"d9",
          6929 => x"bb",
          6930 => x"15",
          6931 => x"2b",
          6932 => x"8d",
          6933 => x"2e",
          6934 => x"77",
          6935 => x"0c",
          6936 => x"76",
          6937 => x"38",
          6938 => x"70",
          6939 => x"81",
          6940 => x"53",
          6941 => x"89",
          6942 => x"56",
          6943 => x"08",
          6944 => x"38",
          6945 => x"15",
          6946 => x"8c",
          6947 => x"80",
          6948 => x"34",
          6949 => x"09",
          6950 => x"92",
          6951 => x"14",
          6952 => x"3f",
          6953 => x"08",
          6954 => x"06",
          6955 => x"2e",
          6956 => x"80",
          6957 => x"1b",
          6958 => x"db",
          6959 => x"bb",
          6960 => x"ea",
          6961 => x"98",
          6962 => x"34",
          6963 => x"51",
          6964 => x"82",
          6965 => x"83",
          6966 => x"53",
          6967 => x"d5",
          6968 => x"06",
          6969 => x"b4",
          6970 => x"84",
          6971 => x"98",
          6972 => x"85",
          6973 => x"09",
          6974 => x"38",
          6975 => x"51",
          6976 => x"82",
          6977 => x"86",
          6978 => x"f2",
          6979 => x"06",
          6980 => x"9c",
          6981 => x"d8",
          6982 => x"98",
          6983 => x"0c",
          6984 => x"51",
          6985 => x"82",
          6986 => x"8c",
          6987 => x"74",
          6988 => x"e0",
          6989 => x"53",
          6990 => x"e0",
          6991 => x"15",
          6992 => x"94",
          6993 => x"56",
          6994 => x"98",
          6995 => x"0d",
          6996 => x"0d",
          6997 => x"55",
          6998 => x"b9",
          6999 => x"53",
          7000 => x"b1",
          7001 => x"52",
          7002 => x"a9",
          7003 => x"22",
          7004 => x"57",
          7005 => x"2e",
          7006 => x"99",
          7007 => x"33",
          7008 => x"3f",
          7009 => x"08",
          7010 => x"71",
          7011 => x"74",
          7012 => x"83",
          7013 => x"78",
          7014 => x"52",
          7015 => x"98",
          7016 => x"0d",
          7017 => x"0d",
          7018 => x"33",
          7019 => x"3d",
          7020 => x"56",
          7021 => x"8b",
          7022 => x"82",
          7023 => x"24",
          7024 => x"bb",
          7025 => x"29",
          7026 => x"05",
          7027 => x"55",
          7028 => x"84",
          7029 => x"34",
          7030 => x"80",
          7031 => x"80",
          7032 => x"75",
          7033 => x"75",
          7034 => x"38",
          7035 => x"3d",
          7036 => x"05",
          7037 => x"3f",
          7038 => x"08",
          7039 => x"bb",
          7040 => x"3d",
          7041 => x"3d",
          7042 => x"84",
          7043 => x"05",
          7044 => x"89",
          7045 => x"2e",
          7046 => x"77",
          7047 => x"54",
          7048 => x"05",
          7049 => x"84",
          7050 => x"f6",
          7051 => x"bb",
          7052 => x"82",
          7053 => x"84",
          7054 => x"5c",
          7055 => x"3d",
          7056 => x"ed",
          7057 => x"bb",
          7058 => x"82",
          7059 => x"92",
          7060 => x"d7",
          7061 => x"98",
          7062 => x"73",
          7063 => x"38",
          7064 => x"9c",
          7065 => x"80",
          7066 => x"38",
          7067 => x"95",
          7068 => x"2e",
          7069 => x"aa",
          7070 => x"ea",
          7071 => x"bb",
          7072 => x"9e",
          7073 => x"05",
          7074 => x"54",
          7075 => x"38",
          7076 => x"70",
          7077 => x"54",
          7078 => x"8e",
          7079 => x"83",
          7080 => x"88",
          7081 => x"83",
          7082 => x"83",
          7083 => x"06",
          7084 => x"80",
          7085 => x"38",
          7086 => x"51",
          7087 => x"82",
          7088 => x"56",
          7089 => x"0a",
          7090 => x"05",
          7091 => x"3f",
          7092 => x"0b",
          7093 => x"80",
          7094 => x"7a",
          7095 => x"3f",
          7096 => x"9c",
          7097 => x"d1",
          7098 => x"81",
          7099 => x"34",
          7100 => x"80",
          7101 => x"b0",
          7102 => x"54",
          7103 => x"52",
          7104 => x"05",
          7105 => x"3f",
          7106 => x"08",
          7107 => x"98",
          7108 => x"38",
          7109 => x"82",
          7110 => x"b2",
          7111 => x"84",
          7112 => x"06",
          7113 => x"73",
          7114 => x"38",
          7115 => x"ad",
          7116 => x"2a",
          7117 => x"51",
          7118 => x"2e",
          7119 => x"81",
          7120 => x"80",
          7121 => x"87",
          7122 => x"39",
          7123 => x"51",
          7124 => x"82",
          7125 => x"7b",
          7126 => x"12",
          7127 => x"82",
          7128 => x"81",
          7129 => x"83",
          7130 => x"06",
          7131 => x"80",
          7132 => x"77",
          7133 => x"58",
          7134 => x"08",
          7135 => x"63",
          7136 => x"63",
          7137 => x"57",
          7138 => x"82",
          7139 => x"82",
          7140 => x"88",
          7141 => x"9c",
          7142 => x"d2",
          7143 => x"bb",
          7144 => x"bb",
          7145 => x"1b",
          7146 => x"0c",
          7147 => x"22",
          7148 => x"77",
          7149 => x"80",
          7150 => x"34",
          7151 => x"1a",
          7152 => x"94",
          7153 => x"85",
          7154 => x"06",
          7155 => x"80",
          7156 => x"38",
          7157 => x"08",
          7158 => x"84",
          7159 => x"98",
          7160 => x"0c",
          7161 => x"70",
          7162 => x"52",
          7163 => x"39",
          7164 => x"51",
          7165 => x"82",
          7166 => x"57",
          7167 => x"08",
          7168 => x"38",
          7169 => x"bb",
          7170 => x"2e",
          7171 => x"83",
          7172 => x"75",
          7173 => x"74",
          7174 => x"07",
          7175 => x"54",
          7176 => x"8a",
          7177 => x"75",
          7178 => x"73",
          7179 => x"98",
          7180 => x"a9",
          7181 => x"ff",
          7182 => x"80",
          7183 => x"76",
          7184 => x"d6",
          7185 => x"bb",
          7186 => x"38",
          7187 => x"39",
          7188 => x"82",
          7189 => x"05",
          7190 => x"84",
          7191 => x"0c",
          7192 => x"82",
          7193 => x"97",
          7194 => x"f2",
          7195 => x"63",
          7196 => x"40",
          7197 => x"7e",
          7198 => x"fc",
          7199 => x"51",
          7200 => x"82",
          7201 => x"55",
          7202 => x"08",
          7203 => x"19",
          7204 => x"80",
          7205 => x"74",
          7206 => x"39",
          7207 => x"81",
          7208 => x"56",
          7209 => x"82",
          7210 => x"39",
          7211 => x"1a",
          7212 => x"82",
          7213 => x"0b",
          7214 => x"81",
          7215 => x"39",
          7216 => x"94",
          7217 => x"55",
          7218 => x"83",
          7219 => x"7b",
          7220 => x"89",
          7221 => x"08",
          7222 => x"06",
          7223 => x"81",
          7224 => x"8a",
          7225 => x"05",
          7226 => x"06",
          7227 => x"a8",
          7228 => x"38",
          7229 => x"55",
          7230 => x"19",
          7231 => x"51",
          7232 => x"82",
          7233 => x"55",
          7234 => x"ff",
          7235 => x"ff",
          7236 => x"38",
          7237 => x"0c",
          7238 => x"52",
          7239 => x"cb",
          7240 => x"98",
          7241 => x"ff",
          7242 => x"bb",
          7243 => x"7c",
          7244 => x"57",
          7245 => x"80",
          7246 => x"1a",
          7247 => x"22",
          7248 => x"75",
          7249 => x"38",
          7250 => x"58",
          7251 => x"53",
          7252 => x"1b",
          7253 => x"88",
          7254 => x"98",
          7255 => x"38",
          7256 => x"33",
          7257 => x"80",
          7258 => x"b0",
          7259 => x"31",
          7260 => x"27",
          7261 => x"80",
          7262 => x"52",
          7263 => x"77",
          7264 => x"7d",
          7265 => x"e0",
          7266 => x"2b",
          7267 => x"76",
          7268 => x"94",
          7269 => x"ff",
          7270 => x"71",
          7271 => x"7b",
          7272 => x"38",
          7273 => x"19",
          7274 => x"51",
          7275 => x"82",
          7276 => x"fe",
          7277 => x"53",
          7278 => x"83",
          7279 => x"b4",
          7280 => x"51",
          7281 => x"7b",
          7282 => x"08",
          7283 => x"76",
          7284 => x"08",
          7285 => x"0c",
          7286 => x"f3",
          7287 => x"75",
          7288 => x"0c",
          7289 => x"04",
          7290 => x"60",
          7291 => x"40",
          7292 => x"80",
          7293 => x"3d",
          7294 => x"77",
          7295 => x"3f",
          7296 => x"08",
          7297 => x"98",
          7298 => x"91",
          7299 => x"74",
          7300 => x"38",
          7301 => x"b8",
          7302 => x"33",
          7303 => x"70",
          7304 => x"56",
          7305 => x"74",
          7306 => x"a4",
          7307 => x"82",
          7308 => x"34",
          7309 => x"98",
          7310 => x"91",
          7311 => x"56",
          7312 => x"94",
          7313 => x"11",
          7314 => x"76",
          7315 => x"75",
          7316 => x"80",
          7317 => x"38",
          7318 => x"70",
          7319 => x"56",
          7320 => x"fd",
          7321 => x"11",
          7322 => x"77",
          7323 => x"5c",
          7324 => x"38",
          7325 => x"88",
          7326 => x"74",
          7327 => x"52",
          7328 => x"18",
          7329 => x"51",
          7330 => x"82",
          7331 => x"55",
          7332 => x"08",
          7333 => x"ab",
          7334 => x"2e",
          7335 => x"74",
          7336 => x"95",
          7337 => x"19",
          7338 => x"08",
          7339 => x"88",
          7340 => x"55",
          7341 => x"9c",
          7342 => x"09",
          7343 => x"38",
          7344 => x"c1",
          7345 => x"98",
          7346 => x"38",
          7347 => x"52",
          7348 => x"97",
          7349 => x"98",
          7350 => x"fe",
          7351 => x"bb",
          7352 => x"7c",
          7353 => x"57",
          7354 => x"80",
          7355 => x"1b",
          7356 => x"22",
          7357 => x"75",
          7358 => x"38",
          7359 => x"59",
          7360 => x"53",
          7361 => x"1a",
          7362 => x"be",
          7363 => x"98",
          7364 => x"38",
          7365 => x"08",
          7366 => x"56",
          7367 => x"9b",
          7368 => x"53",
          7369 => x"77",
          7370 => x"7d",
          7371 => x"16",
          7372 => x"3f",
          7373 => x"0b",
          7374 => x"78",
          7375 => x"80",
          7376 => x"18",
          7377 => x"08",
          7378 => x"7e",
          7379 => x"3f",
          7380 => x"08",
          7381 => x"7e",
          7382 => x"0c",
          7383 => x"19",
          7384 => x"08",
          7385 => x"84",
          7386 => x"57",
          7387 => x"27",
          7388 => x"56",
          7389 => x"52",
          7390 => x"f9",
          7391 => x"98",
          7392 => x"38",
          7393 => x"52",
          7394 => x"83",
          7395 => x"b4",
          7396 => x"d4",
          7397 => x"81",
          7398 => x"34",
          7399 => x"7e",
          7400 => x"0c",
          7401 => x"1a",
          7402 => x"94",
          7403 => x"1b",
          7404 => x"5e",
          7405 => x"27",
          7406 => x"55",
          7407 => x"0c",
          7408 => x"90",
          7409 => x"c0",
          7410 => x"90",
          7411 => x"56",
          7412 => x"98",
          7413 => x"0d",
          7414 => x"0d",
          7415 => x"fc",
          7416 => x"52",
          7417 => x"3f",
          7418 => x"08",
          7419 => x"98",
          7420 => x"38",
          7421 => x"70",
          7422 => x"81",
          7423 => x"55",
          7424 => x"80",
          7425 => x"16",
          7426 => x"51",
          7427 => x"82",
          7428 => x"57",
          7429 => x"08",
          7430 => x"a4",
          7431 => x"11",
          7432 => x"55",
          7433 => x"16",
          7434 => x"08",
          7435 => x"75",
          7436 => x"e8",
          7437 => x"08",
          7438 => x"51",
          7439 => x"82",
          7440 => x"52",
          7441 => x"c9",
          7442 => x"52",
          7443 => x"c9",
          7444 => x"54",
          7445 => x"15",
          7446 => x"cc",
          7447 => x"bb",
          7448 => x"17",
          7449 => x"06",
          7450 => x"90",
          7451 => x"82",
          7452 => x"8a",
          7453 => x"fc",
          7454 => x"70",
          7455 => x"d9",
          7456 => x"98",
          7457 => x"bb",
          7458 => x"38",
          7459 => x"05",
          7460 => x"f1",
          7461 => x"bb",
          7462 => x"82",
          7463 => x"87",
          7464 => x"98",
          7465 => x"72",
          7466 => x"0c",
          7467 => x"04",
          7468 => x"84",
          7469 => x"e4",
          7470 => x"80",
          7471 => x"98",
          7472 => x"38",
          7473 => x"08",
          7474 => x"34",
          7475 => x"82",
          7476 => x"83",
          7477 => x"ef",
          7478 => x"53",
          7479 => x"05",
          7480 => x"51",
          7481 => x"82",
          7482 => x"55",
          7483 => x"08",
          7484 => x"76",
          7485 => x"93",
          7486 => x"51",
          7487 => x"82",
          7488 => x"55",
          7489 => x"08",
          7490 => x"80",
          7491 => x"70",
          7492 => x"56",
          7493 => x"89",
          7494 => x"94",
          7495 => x"b2",
          7496 => x"05",
          7497 => x"2a",
          7498 => x"51",
          7499 => x"80",
          7500 => x"76",
          7501 => x"52",
          7502 => x"3f",
          7503 => x"08",
          7504 => x"8e",
          7505 => x"98",
          7506 => x"09",
          7507 => x"38",
          7508 => x"82",
          7509 => x"93",
          7510 => x"e4",
          7511 => x"6f",
          7512 => x"7a",
          7513 => x"9e",
          7514 => x"05",
          7515 => x"51",
          7516 => x"82",
          7517 => x"57",
          7518 => x"08",
          7519 => x"7b",
          7520 => x"94",
          7521 => x"55",
          7522 => x"73",
          7523 => x"ed",
          7524 => x"93",
          7525 => x"55",
          7526 => x"82",
          7527 => x"57",
          7528 => x"08",
          7529 => x"68",
          7530 => x"c9",
          7531 => x"bb",
          7532 => x"82",
          7533 => x"82",
          7534 => x"52",
          7535 => x"a3",
          7536 => x"98",
          7537 => x"52",
          7538 => x"b8",
          7539 => x"98",
          7540 => x"bb",
          7541 => x"a2",
          7542 => x"74",
          7543 => x"3f",
          7544 => x"08",
          7545 => x"98",
          7546 => x"69",
          7547 => x"d9",
          7548 => x"82",
          7549 => x"2e",
          7550 => x"52",
          7551 => x"cf",
          7552 => x"98",
          7553 => x"bb",
          7554 => x"2e",
          7555 => x"84",
          7556 => x"06",
          7557 => x"57",
          7558 => x"76",
          7559 => x"9e",
          7560 => x"05",
          7561 => x"dc",
          7562 => x"90",
          7563 => x"81",
          7564 => x"56",
          7565 => x"80",
          7566 => x"02",
          7567 => x"81",
          7568 => x"70",
          7569 => x"56",
          7570 => x"81",
          7571 => x"78",
          7572 => x"38",
          7573 => x"99",
          7574 => x"81",
          7575 => x"18",
          7576 => x"18",
          7577 => x"58",
          7578 => x"33",
          7579 => x"ee",
          7580 => x"6f",
          7581 => x"af",
          7582 => x"8d",
          7583 => x"2e",
          7584 => x"8a",
          7585 => x"6f",
          7586 => x"af",
          7587 => x"0b",
          7588 => x"33",
          7589 => x"82",
          7590 => x"70",
          7591 => x"52",
          7592 => x"56",
          7593 => x"8d",
          7594 => x"70",
          7595 => x"51",
          7596 => x"f5",
          7597 => x"54",
          7598 => x"a7",
          7599 => x"74",
          7600 => x"38",
          7601 => x"73",
          7602 => x"81",
          7603 => x"81",
          7604 => x"39",
          7605 => x"81",
          7606 => x"74",
          7607 => x"81",
          7608 => x"91",
          7609 => x"6e",
          7610 => x"59",
          7611 => x"7a",
          7612 => x"5c",
          7613 => x"26",
          7614 => x"7a",
          7615 => x"bb",
          7616 => x"3d",
          7617 => x"3d",
          7618 => x"8d",
          7619 => x"54",
          7620 => x"55",
          7621 => x"82",
          7622 => x"53",
          7623 => x"08",
          7624 => x"91",
          7625 => x"72",
          7626 => x"8c",
          7627 => x"73",
          7628 => x"38",
          7629 => x"70",
          7630 => x"81",
          7631 => x"57",
          7632 => x"73",
          7633 => x"08",
          7634 => x"94",
          7635 => x"75",
          7636 => x"97",
          7637 => x"11",
          7638 => x"2b",
          7639 => x"73",
          7640 => x"38",
          7641 => x"16",
          7642 => x"b9",
          7643 => x"98",
          7644 => x"78",
          7645 => x"55",
          7646 => x"a9",
          7647 => x"98",
          7648 => x"96",
          7649 => x"70",
          7650 => x"94",
          7651 => x"71",
          7652 => x"08",
          7653 => x"53",
          7654 => x"15",
          7655 => x"a6",
          7656 => x"74",
          7657 => x"3f",
          7658 => x"08",
          7659 => x"98",
          7660 => x"81",
          7661 => x"bb",
          7662 => x"2e",
          7663 => x"82",
          7664 => x"88",
          7665 => x"98",
          7666 => x"80",
          7667 => x"38",
          7668 => x"80",
          7669 => x"77",
          7670 => x"08",
          7671 => x"0c",
          7672 => x"70",
          7673 => x"81",
          7674 => x"5a",
          7675 => x"2e",
          7676 => x"52",
          7677 => x"f9",
          7678 => x"98",
          7679 => x"bb",
          7680 => x"38",
          7681 => x"08",
          7682 => x"73",
          7683 => x"c7",
          7684 => x"bb",
          7685 => x"73",
          7686 => x"38",
          7687 => x"af",
          7688 => x"73",
          7689 => x"27",
          7690 => x"98",
          7691 => x"a0",
          7692 => x"08",
          7693 => x"0c",
          7694 => x"06",
          7695 => x"2e",
          7696 => x"52",
          7697 => x"a3",
          7698 => x"98",
          7699 => x"82",
          7700 => x"34",
          7701 => x"c4",
          7702 => x"91",
          7703 => x"53",
          7704 => x"89",
          7705 => x"98",
          7706 => x"94",
          7707 => x"8c",
          7708 => x"27",
          7709 => x"8c",
          7710 => x"15",
          7711 => x"07",
          7712 => x"16",
          7713 => x"ff",
          7714 => x"80",
          7715 => x"77",
          7716 => x"2e",
          7717 => x"9c",
          7718 => x"53",
          7719 => x"98",
          7720 => x"0d",
          7721 => x"0d",
          7722 => x"54",
          7723 => x"81",
          7724 => x"53",
          7725 => x"05",
          7726 => x"84",
          7727 => x"e7",
          7728 => x"98",
          7729 => x"bb",
          7730 => x"ea",
          7731 => x"0c",
          7732 => x"51",
          7733 => x"82",
          7734 => x"55",
          7735 => x"08",
          7736 => x"ab",
          7737 => x"98",
          7738 => x"80",
          7739 => x"38",
          7740 => x"70",
          7741 => x"81",
          7742 => x"57",
          7743 => x"ad",
          7744 => x"08",
          7745 => x"d3",
          7746 => x"bb",
          7747 => x"17",
          7748 => x"86",
          7749 => x"17",
          7750 => x"75",
          7751 => x"3f",
          7752 => x"08",
          7753 => x"2e",
          7754 => x"85",
          7755 => x"86",
          7756 => x"2e",
          7757 => x"76",
          7758 => x"73",
          7759 => x"0c",
          7760 => x"04",
          7761 => x"76",
          7762 => x"05",
          7763 => x"53",
          7764 => x"82",
          7765 => x"87",
          7766 => x"98",
          7767 => x"86",
          7768 => x"fb",
          7769 => x"79",
          7770 => x"05",
          7771 => x"56",
          7772 => x"3f",
          7773 => x"08",
          7774 => x"98",
          7775 => x"38",
          7776 => x"82",
          7777 => x"52",
          7778 => x"f8",
          7779 => x"98",
          7780 => x"ca",
          7781 => x"98",
          7782 => x"51",
          7783 => x"82",
          7784 => x"53",
          7785 => x"08",
          7786 => x"81",
          7787 => x"80",
          7788 => x"82",
          7789 => x"a6",
          7790 => x"73",
          7791 => x"3f",
          7792 => x"51",
          7793 => x"82",
          7794 => x"84",
          7795 => x"70",
          7796 => x"2c",
          7797 => x"98",
          7798 => x"51",
          7799 => x"82",
          7800 => x"87",
          7801 => x"ee",
          7802 => x"57",
          7803 => x"3d",
          7804 => x"3d",
          7805 => x"af",
          7806 => x"98",
          7807 => x"bb",
          7808 => x"38",
          7809 => x"51",
          7810 => x"82",
          7811 => x"55",
          7812 => x"08",
          7813 => x"80",
          7814 => x"70",
          7815 => x"58",
          7816 => x"85",
          7817 => x"8d",
          7818 => x"2e",
          7819 => x"52",
          7820 => x"be",
          7821 => x"bb",
          7822 => x"3d",
          7823 => x"3d",
          7824 => x"55",
          7825 => x"92",
          7826 => x"52",
          7827 => x"de",
          7828 => x"bb",
          7829 => x"82",
          7830 => x"82",
          7831 => x"74",
          7832 => x"98",
          7833 => x"11",
          7834 => x"59",
          7835 => x"75",
          7836 => x"38",
          7837 => x"81",
          7838 => x"5b",
          7839 => x"82",
          7840 => x"39",
          7841 => x"08",
          7842 => x"59",
          7843 => x"09",
          7844 => x"38",
          7845 => x"57",
          7846 => x"3d",
          7847 => x"c1",
          7848 => x"bb",
          7849 => x"2e",
          7850 => x"bb",
          7851 => x"2e",
          7852 => x"bb",
          7853 => x"70",
          7854 => x"08",
          7855 => x"7a",
          7856 => x"7f",
          7857 => x"54",
          7858 => x"77",
          7859 => x"80",
          7860 => x"15",
          7861 => x"98",
          7862 => x"75",
          7863 => x"52",
          7864 => x"52",
          7865 => x"8d",
          7866 => x"98",
          7867 => x"bb",
          7868 => x"d6",
          7869 => x"33",
          7870 => x"1a",
          7871 => x"54",
          7872 => x"09",
          7873 => x"38",
          7874 => x"ff",
          7875 => x"82",
          7876 => x"83",
          7877 => x"70",
          7878 => x"25",
          7879 => x"59",
          7880 => x"9b",
          7881 => x"51",
          7882 => x"3f",
          7883 => x"08",
          7884 => x"70",
          7885 => x"25",
          7886 => x"59",
          7887 => x"75",
          7888 => x"7a",
          7889 => x"ff",
          7890 => x"7c",
          7891 => x"90",
          7892 => x"11",
          7893 => x"56",
          7894 => x"15",
          7895 => x"bb",
          7896 => x"3d",
          7897 => x"3d",
          7898 => x"3d",
          7899 => x"70",
          7900 => x"dd",
          7901 => x"98",
          7902 => x"bb",
          7903 => x"a8",
          7904 => x"33",
          7905 => x"a0",
          7906 => x"33",
          7907 => x"70",
          7908 => x"55",
          7909 => x"73",
          7910 => x"8e",
          7911 => x"08",
          7912 => x"18",
          7913 => x"80",
          7914 => x"38",
          7915 => x"08",
          7916 => x"08",
          7917 => x"c4",
          7918 => x"bb",
          7919 => x"88",
          7920 => x"80",
          7921 => x"17",
          7922 => x"51",
          7923 => x"3f",
          7924 => x"08",
          7925 => x"81",
          7926 => x"81",
          7927 => x"98",
          7928 => x"09",
          7929 => x"38",
          7930 => x"39",
          7931 => x"77",
          7932 => x"98",
          7933 => x"08",
          7934 => x"98",
          7935 => x"82",
          7936 => x"52",
          7937 => x"bd",
          7938 => x"98",
          7939 => x"17",
          7940 => x"0c",
          7941 => x"80",
          7942 => x"73",
          7943 => x"75",
          7944 => x"38",
          7945 => x"34",
          7946 => x"82",
          7947 => x"89",
          7948 => x"e2",
          7949 => x"53",
          7950 => x"a4",
          7951 => x"3d",
          7952 => x"3f",
          7953 => x"08",
          7954 => x"98",
          7955 => x"38",
          7956 => x"3d",
          7957 => x"3d",
          7958 => x"d1",
          7959 => x"bb",
          7960 => x"82",
          7961 => x"81",
          7962 => x"80",
          7963 => x"70",
          7964 => x"81",
          7965 => x"56",
          7966 => x"81",
          7967 => x"98",
          7968 => x"74",
          7969 => x"38",
          7970 => x"05",
          7971 => x"06",
          7972 => x"55",
          7973 => x"38",
          7974 => x"51",
          7975 => x"82",
          7976 => x"74",
          7977 => x"81",
          7978 => x"56",
          7979 => x"80",
          7980 => x"54",
          7981 => x"08",
          7982 => x"2e",
          7983 => x"73",
          7984 => x"98",
          7985 => x"52",
          7986 => x"52",
          7987 => x"3f",
          7988 => x"08",
          7989 => x"98",
          7990 => x"38",
          7991 => x"08",
          7992 => x"cc",
          7993 => x"bb",
          7994 => x"82",
          7995 => x"86",
          7996 => x"80",
          7997 => x"bb",
          7998 => x"2e",
          7999 => x"bb",
          8000 => x"c0",
          8001 => x"ce",
          8002 => x"bb",
          8003 => x"bb",
          8004 => x"70",
          8005 => x"08",
          8006 => x"51",
          8007 => x"80",
          8008 => x"73",
          8009 => x"38",
          8010 => x"52",
          8011 => x"95",
          8012 => x"98",
          8013 => x"8c",
          8014 => x"ff",
          8015 => x"82",
          8016 => x"55",
          8017 => x"98",
          8018 => x"0d",
          8019 => x"0d",
          8020 => x"3d",
          8021 => x"9a",
          8022 => x"cb",
          8023 => x"98",
          8024 => x"bb",
          8025 => x"b0",
          8026 => x"69",
          8027 => x"70",
          8028 => x"97",
          8029 => x"98",
          8030 => x"bb",
          8031 => x"38",
          8032 => x"94",
          8033 => x"98",
          8034 => x"09",
          8035 => x"88",
          8036 => x"df",
          8037 => x"85",
          8038 => x"51",
          8039 => x"74",
          8040 => x"78",
          8041 => x"8a",
          8042 => x"57",
          8043 => x"82",
          8044 => x"75",
          8045 => x"bb",
          8046 => x"38",
          8047 => x"bb",
          8048 => x"2e",
          8049 => x"83",
          8050 => x"82",
          8051 => x"ff",
          8052 => x"06",
          8053 => x"54",
          8054 => x"73",
          8055 => x"82",
          8056 => x"52",
          8057 => x"a4",
          8058 => x"98",
          8059 => x"bb",
          8060 => x"9a",
          8061 => x"a0",
          8062 => x"51",
          8063 => x"3f",
          8064 => x"0b",
          8065 => x"78",
          8066 => x"bf",
          8067 => x"88",
          8068 => x"80",
          8069 => x"ff",
          8070 => x"75",
          8071 => x"11",
          8072 => x"f8",
          8073 => x"78",
          8074 => x"80",
          8075 => x"ff",
          8076 => x"78",
          8077 => x"80",
          8078 => x"7f",
          8079 => x"d4",
          8080 => x"c9",
          8081 => x"54",
          8082 => x"15",
          8083 => x"cb",
          8084 => x"bb",
          8085 => x"82",
          8086 => x"b2",
          8087 => x"b2",
          8088 => x"96",
          8089 => x"b5",
          8090 => x"53",
          8091 => x"51",
          8092 => x"64",
          8093 => x"8b",
          8094 => x"54",
          8095 => x"15",
          8096 => x"ff",
          8097 => x"82",
          8098 => x"54",
          8099 => x"53",
          8100 => x"51",
          8101 => x"3f",
          8102 => x"98",
          8103 => x"0d",
          8104 => x"0d",
          8105 => x"05",
          8106 => x"3f",
          8107 => x"3d",
          8108 => x"52",
          8109 => x"d5",
          8110 => x"bb",
          8111 => x"82",
          8112 => x"82",
          8113 => x"4d",
          8114 => x"52",
          8115 => x"52",
          8116 => x"3f",
          8117 => x"08",
          8118 => x"98",
          8119 => x"38",
          8120 => x"05",
          8121 => x"06",
          8122 => x"73",
          8123 => x"a0",
          8124 => x"08",
          8125 => x"ff",
          8126 => x"ff",
          8127 => x"ac",
          8128 => x"92",
          8129 => x"54",
          8130 => x"3f",
          8131 => x"52",
          8132 => x"f7",
          8133 => x"98",
          8134 => x"bb",
          8135 => x"38",
          8136 => x"09",
          8137 => x"38",
          8138 => x"08",
          8139 => x"88",
          8140 => x"39",
          8141 => x"08",
          8142 => x"81",
          8143 => x"38",
          8144 => x"b1",
          8145 => x"98",
          8146 => x"bb",
          8147 => x"c8",
          8148 => x"93",
          8149 => x"ff",
          8150 => x"8d",
          8151 => x"b4",
          8152 => x"af",
          8153 => x"17",
          8154 => x"33",
          8155 => x"70",
          8156 => x"55",
          8157 => x"38",
          8158 => x"54",
          8159 => x"34",
          8160 => x"0b",
          8161 => x"8b",
          8162 => x"84",
          8163 => x"06",
          8164 => x"73",
          8165 => x"e5",
          8166 => x"2e",
          8167 => x"75",
          8168 => x"c6",
          8169 => x"bb",
          8170 => x"78",
          8171 => x"bb",
          8172 => x"82",
          8173 => x"80",
          8174 => x"38",
          8175 => x"08",
          8176 => x"ff",
          8177 => x"82",
          8178 => x"79",
          8179 => x"58",
          8180 => x"bb",
          8181 => x"c0",
          8182 => x"33",
          8183 => x"2e",
          8184 => x"99",
          8185 => x"75",
          8186 => x"c6",
          8187 => x"54",
          8188 => x"15",
          8189 => x"82",
          8190 => x"9c",
          8191 => x"c8",
          8192 => x"bb",
          8193 => x"82",
          8194 => x"8c",
          8195 => x"ff",
          8196 => x"82",
          8197 => x"55",
          8198 => x"98",
          8199 => x"0d",
          8200 => x"0d",
          8201 => x"05",
          8202 => x"05",
          8203 => x"33",
          8204 => x"53",
          8205 => x"05",
          8206 => x"51",
          8207 => x"82",
          8208 => x"55",
          8209 => x"08",
          8210 => x"78",
          8211 => x"95",
          8212 => x"51",
          8213 => x"82",
          8214 => x"55",
          8215 => x"08",
          8216 => x"80",
          8217 => x"81",
          8218 => x"86",
          8219 => x"38",
          8220 => x"61",
          8221 => x"12",
          8222 => x"7a",
          8223 => x"51",
          8224 => x"74",
          8225 => x"78",
          8226 => x"83",
          8227 => x"51",
          8228 => x"3f",
          8229 => x"08",
          8230 => x"bb",
          8231 => x"3d",
          8232 => x"3d",
          8233 => x"82",
          8234 => x"d0",
          8235 => x"3d",
          8236 => x"3f",
          8237 => x"08",
          8238 => x"98",
          8239 => x"38",
          8240 => x"52",
          8241 => x"05",
          8242 => x"3f",
          8243 => x"08",
          8244 => x"98",
          8245 => x"02",
          8246 => x"33",
          8247 => x"54",
          8248 => x"a6",
          8249 => x"22",
          8250 => x"71",
          8251 => x"53",
          8252 => x"51",
          8253 => x"3f",
          8254 => x"0b",
          8255 => x"76",
          8256 => x"b8",
          8257 => x"98",
          8258 => x"82",
          8259 => x"93",
          8260 => x"ea",
          8261 => x"6b",
          8262 => x"53",
          8263 => x"05",
          8264 => x"51",
          8265 => x"82",
          8266 => x"82",
          8267 => x"30",
          8268 => x"98",
          8269 => x"25",
          8270 => x"79",
          8271 => x"85",
          8272 => x"75",
          8273 => x"73",
          8274 => x"f9",
          8275 => x"80",
          8276 => x"8d",
          8277 => x"54",
          8278 => x"3f",
          8279 => x"08",
          8280 => x"98",
          8281 => x"38",
          8282 => x"51",
          8283 => x"82",
          8284 => x"57",
          8285 => x"08",
          8286 => x"bb",
          8287 => x"bb",
          8288 => x"5b",
          8289 => x"18",
          8290 => x"18",
          8291 => x"74",
          8292 => x"81",
          8293 => x"78",
          8294 => x"8b",
          8295 => x"54",
          8296 => x"75",
          8297 => x"38",
          8298 => x"1b",
          8299 => x"55",
          8300 => x"2e",
          8301 => x"39",
          8302 => x"09",
          8303 => x"38",
          8304 => x"80",
          8305 => x"70",
          8306 => x"25",
          8307 => x"80",
          8308 => x"38",
          8309 => x"bc",
          8310 => x"11",
          8311 => x"ff",
          8312 => x"82",
          8313 => x"57",
          8314 => x"08",
          8315 => x"70",
          8316 => x"80",
          8317 => x"83",
          8318 => x"80",
          8319 => x"84",
          8320 => x"a7",
          8321 => x"b4",
          8322 => x"ad",
          8323 => x"bb",
          8324 => x"0c",
          8325 => x"98",
          8326 => x"0d",
          8327 => x"0d",
          8328 => x"3d",
          8329 => x"52",
          8330 => x"ce",
          8331 => x"bb",
          8332 => x"bb",
          8333 => x"54",
          8334 => x"08",
          8335 => x"8b",
          8336 => x"8b",
          8337 => x"59",
          8338 => x"3f",
          8339 => x"33",
          8340 => x"06",
          8341 => x"57",
          8342 => x"81",
          8343 => x"58",
          8344 => x"06",
          8345 => x"4e",
          8346 => x"ff",
          8347 => x"82",
          8348 => x"80",
          8349 => x"6c",
          8350 => x"53",
          8351 => x"ae",
          8352 => x"bb",
          8353 => x"2e",
          8354 => x"88",
          8355 => x"6d",
          8356 => x"55",
          8357 => x"bb",
          8358 => x"ff",
          8359 => x"83",
          8360 => x"51",
          8361 => x"26",
          8362 => x"15",
          8363 => x"ff",
          8364 => x"80",
          8365 => x"87",
          8366 => x"e0",
          8367 => x"74",
          8368 => x"38",
          8369 => x"b5",
          8370 => x"ae",
          8371 => x"bb",
          8372 => x"38",
          8373 => x"27",
          8374 => x"89",
          8375 => x"8b",
          8376 => x"27",
          8377 => x"55",
          8378 => x"81",
          8379 => x"8f",
          8380 => x"2a",
          8381 => x"70",
          8382 => x"34",
          8383 => x"74",
          8384 => x"05",
          8385 => x"17",
          8386 => x"70",
          8387 => x"52",
          8388 => x"73",
          8389 => x"c8",
          8390 => x"33",
          8391 => x"73",
          8392 => x"81",
          8393 => x"80",
          8394 => x"02",
          8395 => x"76",
          8396 => x"51",
          8397 => x"2e",
          8398 => x"87",
          8399 => x"57",
          8400 => x"79",
          8401 => x"80",
          8402 => x"70",
          8403 => x"ba",
          8404 => x"bb",
          8405 => x"82",
          8406 => x"80",
          8407 => x"52",
          8408 => x"bf",
          8409 => x"bb",
          8410 => x"82",
          8411 => x"8d",
          8412 => x"c4",
          8413 => x"e5",
          8414 => x"c6",
          8415 => x"98",
          8416 => x"09",
          8417 => x"cc",
          8418 => x"76",
          8419 => x"c4",
          8420 => x"74",
          8421 => x"b0",
          8422 => x"98",
          8423 => x"bb",
          8424 => x"38",
          8425 => x"bb",
          8426 => x"67",
          8427 => x"db",
          8428 => x"88",
          8429 => x"34",
          8430 => x"52",
          8431 => x"ab",
          8432 => x"54",
          8433 => x"15",
          8434 => x"ff",
          8435 => x"82",
          8436 => x"54",
          8437 => x"82",
          8438 => x"9c",
          8439 => x"f2",
          8440 => x"62",
          8441 => x"80",
          8442 => x"93",
          8443 => x"55",
          8444 => x"5e",
          8445 => x"3f",
          8446 => x"08",
          8447 => x"98",
          8448 => x"38",
          8449 => x"58",
          8450 => x"38",
          8451 => x"97",
          8452 => x"08",
          8453 => x"38",
          8454 => x"70",
          8455 => x"81",
          8456 => x"55",
          8457 => x"87",
          8458 => x"39",
          8459 => x"90",
          8460 => x"82",
          8461 => x"8a",
          8462 => x"89",
          8463 => x"7f",
          8464 => x"56",
          8465 => x"3f",
          8466 => x"06",
          8467 => x"72",
          8468 => x"82",
          8469 => x"05",
          8470 => x"7c",
          8471 => x"55",
          8472 => x"27",
          8473 => x"16",
          8474 => x"83",
          8475 => x"76",
          8476 => x"80",
          8477 => x"79",
          8478 => x"99",
          8479 => x"7f",
          8480 => x"14",
          8481 => x"83",
          8482 => x"82",
          8483 => x"81",
          8484 => x"38",
          8485 => x"08",
          8486 => x"95",
          8487 => x"98",
          8488 => x"81",
          8489 => x"7b",
          8490 => x"06",
          8491 => x"39",
          8492 => x"56",
          8493 => x"09",
          8494 => x"b9",
          8495 => x"80",
          8496 => x"80",
          8497 => x"78",
          8498 => x"7a",
          8499 => x"38",
          8500 => x"73",
          8501 => x"81",
          8502 => x"ff",
          8503 => x"74",
          8504 => x"ff",
          8505 => x"82",
          8506 => x"58",
          8507 => x"08",
          8508 => x"74",
          8509 => x"16",
          8510 => x"73",
          8511 => x"39",
          8512 => x"7e",
          8513 => x"0c",
          8514 => x"2e",
          8515 => x"88",
          8516 => x"8c",
          8517 => x"1a",
          8518 => x"07",
          8519 => x"1b",
          8520 => x"08",
          8521 => x"16",
          8522 => x"75",
          8523 => x"38",
          8524 => x"90",
          8525 => x"15",
          8526 => x"54",
          8527 => x"34",
          8528 => x"82",
          8529 => x"90",
          8530 => x"e9",
          8531 => x"6d",
          8532 => x"80",
          8533 => x"9d",
          8534 => x"5c",
          8535 => x"3f",
          8536 => x"0b",
          8537 => x"08",
          8538 => x"38",
          8539 => x"08",
          8540 => x"d2",
          8541 => x"08",
          8542 => x"80",
          8543 => x"80",
          8544 => x"bb",
          8545 => x"ff",
          8546 => x"52",
          8547 => x"a0",
          8548 => x"bb",
          8549 => x"ff",
          8550 => x"06",
          8551 => x"56",
          8552 => x"38",
          8553 => x"70",
          8554 => x"55",
          8555 => x"8b",
          8556 => x"3d",
          8557 => x"83",
          8558 => x"ff",
          8559 => x"82",
          8560 => x"99",
          8561 => x"74",
          8562 => x"38",
          8563 => x"80",
          8564 => x"ff",
          8565 => x"55",
          8566 => x"83",
          8567 => x"78",
          8568 => x"38",
          8569 => x"26",
          8570 => x"81",
          8571 => x"8b",
          8572 => x"79",
          8573 => x"80",
          8574 => x"93",
          8575 => x"39",
          8576 => x"6e",
          8577 => x"89",
          8578 => x"48",
          8579 => x"83",
          8580 => x"61",
          8581 => x"25",
          8582 => x"55",
          8583 => x"8a",
          8584 => x"3d",
          8585 => x"81",
          8586 => x"ff",
          8587 => x"81",
          8588 => x"98",
          8589 => x"38",
          8590 => x"70",
          8591 => x"bb",
          8592 => x"56",
          8593 => x"38",
          8594 => x"55",
          8595 => x"75",
          8596 => x"38",
          8597 => x"70",
          8598 => x"ff",
          8599 => x"83",
          8600 => x"78",
          8601 => x"89",
          8602 => x"81",
          8603 => x"06",
          8604 => x"80",
          8605 => x"77",
          8606 => x"74",
          8607 => x"8d",
          8608 => x"06",
          8609 => x"2e",
          8610 => x"77",
          8611 => x"93",
          8612 => x"74",
          8613 => x"cb",
          8614 => x"7d",
          8615 => x"81",
          8616 => x"38",
          8617 => x"66",
          8618 => x"81",
          8619 => x"84",
          8620 => x"74",
          8621 => x"38",
          8622 => x"98",
          8623 => x"84",
          8624 => x"82",
          8625 => x"57",
          8626 => x"80",
          8627 => x"76",
          8628 => x"38",
          8629 => x"51",
          8630 => x"3f",
          8631 => x"08",
          8632 => x"87",
          8633 => x"2a",
          8634 => x"5c",
          8635 => x"bb",
          8636 => x"80",
          8637 => x"44",
          8638 => x"0a",
          8639 => x"ec",
          8640 => x"39",
          8641 => x"66",
          8642 => x"81",
          8643 => x"f4",
          8644 => x"74",
          8645 => x"38",
          8646 => x"98",
          8647 => x"f4",
          8648 => x"82",
          8649 => x"57",
          8650 => x"80",
          8651 => x"76",
          8652 => x"38",
          8653 => x"51",
          8654 => x"3f",
          8655 => x"08",
          8656 => x"57",
          8657 => x"08",
          8658 => x"96",
          8659 => x"82",
          8660 => x"10",
          8661 => x"08",
          8662 => x"72",
          8663 => x"59",
          8664 => x"ff",
          8665 => x"5d",
          8666 => x"44",
          8667 => x"11",
          8668 => x"70",
          8669 => x"71",
          8670 => x"06",
          8671 => x"52",
          8672 => x"40",
          8673 => x"09",
          8674 => x"38",
          8675 => x"18",
          8676 => x"39",
          8677 => x"79",
          8678 => x"70",
          8679 => x"58",
          8680 => x"76",
          8681 => x"38",
          8682 => x"7d",
          8683 => x"70",
          8684 => x"55",
          8685 => x"3f",
          8686 => x"08",
          8687 => x"2e",
          8688 => x"9b",
          8689 => x"98",
          8690 => x"f5",
          8691 => x"38",
          8692 => x"38",
          8693 => x"59",
          8694 => x"38",
          8695 => x"7d",
          8696 => x"81",
          8697 => x"38",
          8698 => x"0b",
          8699 => x"08",
          8700 => x"78",
          8701 => x"1a",
          8702 => x"c0",
          8703 => x"74",
          8704 => x"39",
          8705 => x"55",
          8706 => x"8f",
          8707 => x"fd",
          8708 => x"bb",
          8709 => x"f5",
          8710 => x"78",
          8711 => x"79",
          8712 => x"80",
          8713 => x"f1",
          8714 => x"39",
          8715 => x"81",
          8716 => x"06",
          8717 => x"55",
          8718 => x"27",
          8719 => x"81",
          8720 => x"56",
          8721 => x"38",
          8722 => x"80",
          8723 => x"ff",
          8724 => x"8b",
          8725 => x"9c",
          8726 => x"ff",
          8727 => x"84",
          8728 => x"1b",
          8729 => x"b3",
          8730 => x"1c",
          8731 => x"ff",
          8732 => x"8e",
          8733 => x"a1",
          8734 => x"0b",
          8735 => x"7d",
          8736 => x"30",
          8737 => x"84",
          8738 => x"51",
          8739 => x"51",
          8740 => x"3f",
          8741 => x"83",
          8742 => x"90",
          8743 => x"ff",
          8744 => x"93",
          8745 => x"a0",
          8746 => x"39",
          8747 => x"1b",
          8748 => x"85",
          8749 => x"95",
          8750 => x"52",
          8751 => x"ff",
          8752 => x"81",
          8753 => x"1b",
          8754 => x"cf",
          8755 => x"9c",
          8756 => x"a0",
          8757 => x"83",
          8758 => x"06",
          8759 => x"82",
          8760 => x"52",
          8761 => x"51",
          8762 => x"3f",
          8763 => x"1b",
          8764 => x"c5",
          8765 => x"ac",
          8766 => x"a0",
          8767 => x"52",
          8768 => x"ff",
          8769 => x"86",
          8770 => x"51",
          8771 => x"3f",
          8772 => x"80",
          8773 => x"a9",
          8774 => x"1c",
          8775 => x"82",
          8776 => x"80",
          8777 => x"ae",
          8778 => x"b2",
          8779 => x"1b",
          8780 => x"85",
          8781 => x"ff",
          8782 => x"96",
          8783 => x"9f",
          8784 => x"80",
          8785 => x"34",
          8786 => x"1c",
          8787 => x"82",
          8788 => x"ab",
          8789 => x"a0",
          8790 => x"d4",
          8791 => x"fe",
          8792 => x"59",
          8793 => x"3f",
          8794 => x"53",
          8795 => x"51",
          8796 => x"3f",
          8797 => x"bb",
          8798 => x"e7",
          8799 => x"2e",
          8800 => x"80",
          8801 => x"54",
          8802 => x"53",
          8803 => x"51",
          8804 => x"3f",
          8805 => x"80",
          8806 => x"ff",
          8807 => x"84",
          8808 => x"d2",
          8809 => x"ff",
          8810 => x"86",
          8811 => x"f2",
          8812 => x"1b",
          8813 => x"81",
          8814 => x"52",
          8815 => x"51",
          8816 => x"3f",
          8817 => x"ec",
          8818 => x"9e",
          8819 => x"d4",
          8820 => x"51",
          8821 => x"3f",
          8822 => x"87",
          8823 => x"52",
          8824 => x"9a",
          8825 => x"54",
          8826 => x"7a",
          8827 => x"ff",
          8828 => x"65",
          8829 => x"7a",
          8830 => x"8f",
          8831 => x"80",
          8832 => x"2e",
          8833 => x"9a",
          8834 => x"7a",
          8835 => x"a9",
          8836 => x"84",
          8837 => x"9e",
          8838 => x"0a",
          8839 => x"51",
          8840 => x"ff",
          8841 => x"7d",
          8842 => x"38",
          8843 => x"52",
          8844 => x"9e",
          8845 => x"55",
          8846 => x"62",
          8847 => x"74",
          8848 => x"75",
          8849 => x"7e",
          8850 => x"fe",
          8851 => x"98",
          8852 => x"38",
          8853 => x"82",
          8854 => x"52",
          8855 => x"9e",
          8856 => x"16",
          8857 => x"56",
          8858 => x"38",
          8859 => x"77",
          8860 => x"8d",
          8861 => x"7d",
          8862 => x"38",
          8863 => x"57",
          8864 => x"83",
          8865 => x"76",
          8866 => x"7a",
          8867 => x"ff",
          8868 => x"82",
          8869 => x"81",
          8870 => x"16",
          8871 => x"56",
          8872 => x"38",
          8873 => x"83",
          8874 => x"86",
          8875 => x"ff",
          8876 => x"38",
          8877 => x"82",
          8878 => x"81",
          8879 => x"06",
          8880 => x"fe",
          8881 => x"53",
          8882 => x"51",
          8883 => x"3f",
          8884 => x"52",
          8885 => x"9c",
          8886 => x"be",
          8887 => x"75",
          8888 => x"81",
          8889 => x"0b",
          8890 => x"77",
          8891 => x"75",
          8892 => x"60",
          8893 => x"80",
          8894 => x"75",
          8895 => x"a5",
          8896 => x"85",
          8897 => x"bb",
          8898 => x"2a",
          8899 => x"75",
          8900 => x"82",
          8901 => x"87",
          8902 => x"52",
          8903 => x"51",
          8904 => x"3f",
          8905 => x"ca",
          8906 => x"9c",
          8907 => x"54",
          8908 => x"52",
          8909 => x"98",
          8910 => x"56",
          8911 => x"08",
          8912 => x"53",
          8913 => x"51",
          8914 => x"3f",
          8915 => x"bb",
          8916 => x"38",
          8917 => x"56",
          8918 => x"56",
          8919 => x"bb",
          8920 => x"75",
          8921 => x"0c",
          8922 => x"04",
          8923 => x"7d",
          8924 => x"80",
          8925 => x"05",
          8926 => x"76",
          8927 => x"38",
          8928 => x"11",
          8929 => x"53",
          8930 => x"79",
          8931 => x"3f",
          8932 => x"09",
          8933 => x"38",
          8934 => x"55",
          8935 => x"db",
          8936 => x"70",
          8937 => x"34",
          8938 => x"74",
          8939 => x"81",
          8940 => x"80",
          8941 => x"55",
          8942 => x"76",
          8943 => x"bb",
          8944 => x"3d",
          8945 => x"3d",
          8946 => x"84",
          8947 => x"33",
          8948 => x"8a",
          8949 => x"06",
          8950 => x"52",
          8951 => x"3f",
          8952 => x"56",
          8953 => x"be",
          8954 => x"08",
          8955 => x"05",
          8956 => x"75",
          8957 => x"56",
          8958 => x"a1",
          8959 => x"fc",
          8960 => x"53",
          8961 => x"76",
          8962 => x"dc",
          8963 => x"32",
          8964 => x"72",
          8965 => x"70",
          8966 => x"56",
          8967 => x"18",
          8968 => x"88",
          8969 => x"3d",
          8970 => x"3d",
          8971 => x"11",
          8972 => x"80",
          8973 => x"38",
          8974 => x"05",
          8975 => x"8c",
          8976 => x"08",
          8977 => x"3f",
          8978 => x"08",
          8979 => x"16",
          8980 => x"09",
          8981 => x"38",
          8982 => x"55",
          8983 => x"55",
          8984 => x"98",
          8985 => x"0d",
          8986 => x"0d",
          8987 => x"cc",
          8988 => x"73",
          8989 => x"93",
          8990 => x"0c",
          8991 => x"04",
          8992 => x"02",
          8993 => x"33",
          8994 => x"3d",
          8995 => x"54",
          8996 => x"52",
          8997 => x"ae",
          8998 => x"ff",
          8999 => x"3d",
          9000 => x"ff",
          9001 => x"00",
          9002 => x"ff",
          9003 => x"ff",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"00",
          9136 => x"00",
          9137 => x"00",
          9138 => x"00",
          9139 => x"00",
          9140 => x"69",
          9141 => x"00",
          9142 => x"69",
          9143 => x"6c",
          9144 => x"69",
          9145 => x"00",
          9146 => x"6c",
          9147 => x"00",
          9148 => x"65",
          9149 => x"00",
          9150 => x"63",
          9151 => x"72",
          9152 => x"63",
          9153 => x"00",
          9154 => x"64",
          9155 => x"00",
          9156 => x"64",
          9157 => x"00",
          9158 => x"65",
          9159 => x"65",
          9160 => x"65",
          9161 => x"69",
          9162 => x"69",
          9163 => x"66",
          9164 => x"66",
          9165 => x"61",
          9166 => x"00",
          9167 => x"6d",
          9168 => x"65",
          9169 => x"72",
          9170 => x"65",
          9171 => x"00",
          9172 => x"6e",
          9173 => x"00",
          9174 => x"65",
          9175 => x"00",
          9176 => x"62",
          9177 => x"63",
          9178 => x"62",
          9179 => x"63",
          9180 => x"69",
          9181 => x"00",
          9182 => x"64",
          9183 => x"69",
          9184 => x"45",
          9185 => x"72",
          9186 => x"6e",
          9187 => x"6e",
          9188 => x"65",
          9189 => x"72",
          9190 => x"00",
          9191 => x"69",
          9192 => x"6e",
          9193 => x"72",
          9194 => x"79",
          9195 => x"00",
          9196 => x"6f",
          9197 => x"6c",
          9198 => x"6f",
          9199 => x"2e",
          9200 => x"6f",
          9201 => x"74",
          9202 => x"6f",
          9203 => x"2e",
          9204 => x"6e",
          9205 => x"69",
          9206 => x"69",
          9207 => x"61",
          9208 => x"0a",
          9209 => x"63",
          9210 => x"73",
          9211 => x"6e",
          9212 => x"2e",
          9213 => x"69",
          9214 => x"61",
          9215 => x"61",
          9216 => x"65",
          9217 => x"74",
          9218 => x"00",
          9219 => x"69",
          9220 => x"68",
          9221 => x"6c",
          9222 => x"6e",
          9223 => x"69",
          9224 => x"00",
          9225 => x"44",
          9226 => x"20",
          9227 => x"74",
          9228 => x"72",
          9229 => x"63",
          9230 => x"2e",
          9231 => x"72",
          9232 => x"20",
          9233 => x"62",
          9234 => x"69",
          9235 => x"6e",
          9236 => x"69",
          9237 => x"00",
          9238 => x"69",
          9239 => x"6e",
          9240 => x"65",
          9241 => x"6c",
          9242 => x"0a",
          9243 => x"6f",
          9244 => x"6d",
          9245 => x"69",
          9246 => x"20",
          9247 => x"65",
          9248 => x"74",
          9249 => x"66",
          9250 => x"64",
          9251 => x"20",
          9252 => x"6b",
          9253 => x"00",
          9254 => x"6f",
          9255 => x"74",
          9256 => x"6f",
          9257 => x"64",
          9258 => x"00",
          9259 => x"69",
          9260 => x"75",
          9261 => x"6f",
          9262 => x"61",
          9263 => x"6e",
          9264 => x"6e",
          9265 => x"6c",
          9266 => x"0a",
          9267 => x"69",
          9268 => x"69",
          9269 => x"6f",
          9270 => x"64",
          9271 => x"00",
          9272 => x"6e",
          9273 => x"66",
          9274 => x"65",
          9275 => x"6d",
          9276 => x"72",
          9277 => x"00",
          9278 => x"6f",
          9279 => x"61",
          9280 => x"6f",
          9281 => x"20",
          9282 => x"65",
          9283 => x"00",
          9284 => x"61",
          9285 => x"65",
          9286 => x"73",
          9287 => x"63",
          9288 => x"65",
          9289 => x"0a",
          9290 => x"75",
          9291 => x"73",
          9292 => x"00",
          9293 => x"6e",
          9294 => x"77",
          9295 => x"72",
          9296 => x"2e",
          9297 => x"25",
          9298 => x"62",
          9299 => x"73",
          9300 => x"20",
          9301 => x"25",
          9302 => x"62",
          9303 => x"73",
          9304 => x"63",
          9305 => x"00",
          9306 => x"65",
          9307 => x"00",
          9308 => x"30",
          9309 => x"00",
          9310 => x"20",
          9311 => x"30",
          9312 => x"00",
          9313 => x"20",
          9314 => x"20",
          9315 => x"00",
          9316 => x"30",
          9317 => x"00",
          9318 => x"20",
          9319 => x"7c",
          9320 => x"0d",
          9321 => x"50",
          9322 => x"00",
          9323 => x"2a",
          9324 => x"73",
          9325 => x"00",
          9326 => x"32",
          9327 => x"2f",
          9328 => x"30",
          9329 => x"31",
          9330 => x"00",
          9331 => x"5a",
          9332 => x"20",
          9333 => x"20",
          9334 => x"78",
          9335 => x"73",
          9336 => x"20",
          9337 => x"0a",
          9338 => x"50",
          9339 => x"20",
          9340 => x"65",
          9341 => x"70",
          9342 => x"61",
          9343 => x"65",
          9344 => x"00",
          9345 => x"69",
          9346 => x"20",
          9347 => x"65",
          9348 => x"70",
          9349 => x"00",
          9350 => x"53",
          9351 => x"6e",
          9352 => x"72",
          9353 => x"0a",
          9354 => x"4f",
          9355 => x"20",
          9356 => x"69",
          9357 => x"72",
          9358 => x"74",
          9359 => x"4f",
          9360 => x"20",
          9361 => x"69",
          9362 => x"72",
          9363 => x"74",
          9364 => x"41",
          9365 => x"20",
          9366 => x"69",
          9367 => x"72",
          9368 => x"74",
          9369 => x"41",
          9370 => x"20",
          9371 => x"69",
          9372 => x"72",
          9373 => x"74",
          9374 => x"41",
          9375 => x"20",
          9376 => x"69",
          9377 => x"72",
          9378 => x"74",
          9379 => x"41",
          9380 => x"20",
          9381 => x"69",
          9382 => x"72",
          9383 => x"74",
          9384 => x"65",
          9385 => x"6e",
          9386 => x"70",
          9387 => x"6d",
          9388 => x"2e",
          9389 => x"00",
          9390 => x"6e",
          9391 => x"69",
          9392 => x"74",
          9393 => x"72",
          9394 => x"0a",
          9395 => x"75",
          9396 => x"78",
          9397 => x"62",
          9398 => x"00",
          9399 => x"70",
          9400 => x"2e",
          9401 => x"00",
          9402 => x"3a",
          9403 => x"61",
          9404 => x"64",
          9405 => x"20",
          9406 => x"74",
          9407 => x"69",
          9408 => x"73",
          9409 => x"61",
          9410 => x"30",
          9411 => x"6c",
          9412 => x"65",
          9413 => x"69",
          9414 => x"61",
          9415 => x"6c",
          9416 => x"00",
          9417 => x"20",
          9418 => x"61",
          9419 => x"69",
          9420 => x"69",
          9421 => x"00",
          9422 => x"6e",
          9423 => x"61",
          9424 => x"65",
          9425 => x"00",
          9426 => x"61",
          9427 => x"64",
          9428 => x"20",
          9429 => x"74",
          9430 => x"69",
          9431 => x"0a",
          9432 => x"63",
          9433 => x"0a",
          9434 => x"75",
          9435 => x"6c",
          9436 => x"69",
          9437 => x"2e",
          9438 => x"00",
          9439 => x"6f",
          9440 => x"6e",
          9441 => x"2e",
          9442 => x"6f",
          9443 => x"72",
          9444 => x"2e",
          9445 => x"00",
          9446 => x"30",
          9447 => x"28",
          9448 => x"78",
          9449 => x"25",
          9450 => x"78",
          9451 => x"38",
          9452 => x"00",
          9453 => x"75",
          9454 => x"4d",
          9455 => x"72",
          9456 => x"00",
          9457 => x"43",
          9458 => x"6c",
          9459 => x"2e",
          9460 => x"30",
          9461 => x"25",
          9462 => x"2d",
          9463 => x"3f",
          9464 => x"00",
          9465 => x"30",
          9466 => x"25",
          9467 => x"2d",
          9468 => x"30",
          9469 => x"25",
          9470 => x"2d",
          9471 => x"69",
          9472 => x"6c",
          9473 => x"20",
          9474 => x"65",
          9475 => x"70",
          9476 => x"00",
          9477 => x"6e",
          9478 => x"69",
          9479 => x"69",
          9480 => x"72",
          9481 => x"74",
          9482 => x"00",
          9483 => x"69",
          9484 => x"6c",
          9485 => x"75",
          9486 => x"20",
          9487 => x"6f",
          9488 => x"6e",
          9489 => x"69",
          9490 => x"75",
          9491 => x"20",
          9492 => x"6f",
          9493 => x"78",
          9494 => x"74",
          9495 => x"20",
          9496 => x"65",
          9497 => x"25",
          9498 => x"20",
          9499 => x"0a",
          9500 => x"61",
          9501 => x"6e",
          9502 => x"6f",
          9503 => x"40",
          9504 => x"38",
          9505 => x"2e",
          9506 => x"00",
          9507 => x"61",
          9508 => x"72",
          9509 => x"72",
          9510 => x"20",
          9511 => x"65",
          9512 => x"64",
          9513 => x"00",
          9514 => x"65",
          9515 => x"72",
          9516 => x"67",
          9517 => x"70",
          9518 => x"61",
          9519 => x"6e",
          9520 => x"0a",
          9521 => x"6f",
          9522 => x"72",
          9523 => x"6f",
          9524 => x"67",
          9525 => x"0a",
          9526 => x"50",
          9527 => x"69",
          9528 => x"64",
          9529 => x"73",
          9530 => x"2e",
          9531 => x"00",
          9532 => x"64",
          9533 => x"73",
          9534 => x"00",
          9535 => x"64",
          9536 => x"73",
          9537 => x"61",
          9538 => x"6f",
          9539 => x"6e",
          9540 => x"00",
          9541 => x"75",
          9542 => x"6e",
          9543 => x"2e",
          9544 => x"6e",
          9545 => x"69",
          9546 => x"69",
          9547 => x"72",
          9548 => x"74",
          9549 => x"2e",
          9550 => x"64",
          9551 => x"2f",
          9552 => x"25",
          9553 => x"64",
          9554 => x"2e",
          9555 => x"64",
          9556 => x"6f",
          9557 => x"6f",
          9558 => x"67",
          9559 => x"74",
          9560 => x"00",
          9561 => x"28",
          9562 => x"6d",
          9563 => x"43",
          9564 => x"6e",
          9565 => x"29",
          9566 => x"0a",
          9567 => x"69",
          9568 => x"20",
          9569 => x"6c",
          9570 => x"6e",
          9571 => x"3a",
          9572 => x"20",
          9573 => x"42",
          9574 => x"52",
          9575 => x"20",
          9576 => x"38",
          9577 => x"30",
          9578 => x"2e",
          9579 => x"20",
          9580 => x"44",
          9581 => x"20",
          9582 => x"20",
          9583 => x"38",
          9584 => x"30",
          9585 => x"2e",
          9586 => x"20",
          9587 => x"4e",
          9588 => x"42",
          9589 => x"20",
          9590 => x"38",
          9591 => x"30",
          9592 => x"2e",
          9593 => x"20",
          9594 => x"52",
          9595 => x"20",
          9596 => x"20",
          9597 => x"38",
          9598 => x"30",
          9599 => x"2e",
          9600 => x"20",
          9601 => x"41",
          9602 => x"20",
          9603 => x"20",
          9604 => x"38",
          9605 => x"30",
          9606 => x"2e",
          9607 => x"20",
          9608 => x"44",
          9609 => x"52",
          9610 => x"20",
          9611 => x"76",
          9612 => x"73",
          9613 => x"30",
          9614 => x"2e",
          9615 => x"20",
          9616 => x"49",
          9617 => x"31",
          9618 => x"20",
          9619 => x"6d",
          9620 => x"20",
          9621 => x"30",
          9622 => x"2e",
          9623 => x"20",
          9624 => x"4e",
          9625 => x"43",
          9626 => x"20",
          9627 => x"61",
          9628 => x"6c",
          9629 => x"30",
          9630 => x"2e",
          9631 => x"20",
          9632 => x"49",
          9633 => x"4f",
          9634 => x"42",
          9635 => x"00",
          9636 => x"20",
          9637 => x"42",
          9638 => x"43",
          9639 => x"20",
          9640 => x"4f",
          9641 => x"0a",
          9642 => x"20",
          9643 => x"53",
          9644 => x"00",
          9645 => x"20",
          9646 => x"50",
          9647 => x"00",
          9648 => x"64",
          9649 => x"73",
          9650 => x"3a",
          9651 => x"20",
          9652 => x"50",
          9653 => x"65",
          9654 => x"20",
          9655 => x"74",
          9656 => x"41",
          9657 => x"65",
          9658 => x"3d",
          9659 => x"38",
          9660 => x"00",
          9661 => x"20",
          9662 => x"50",
          9663 => x"65",
          9664 => x"79",
          9665 => x"61",
          9666 => x"41",
          9667 => x"65",
          9668 => x"3d",
          9669 => x"38",
          9670 => x"00",
          9671 => x"20",
          9672 => x"74",
          9673 => x"20",
          9674 => x"72",
          9675 => x"64",
          9676 => x"73",
          9677 => x"20",
          9678 => x"3d",
          9679 => x"38",
          9680 => x"00",
          9681 => x"69",
          9682 => x"0a",
          9683 => x"20",
          9684 => x"50",
          9685 => x"64",
          9686 => x"20",
          9687 => x"20",
          9688 => x"20",
          9689 => x"20",
          9690 => x"3d",
          9691 => x"34",
          9692 => x"00",
          9693 => x"20",
          9694 => x"79",
          9695 => x"6d",
          9696 => x"6f",
          9697 => x"46",
          9698 => x"20",
          9699 => x"20",
          9700 => x"3d",
          9701 => x"2e",
          9702 => x"64",
          9703 => x"0a",
          9704 => x"20",
          9705 => x"44",
          9706 => x"20",
          9707 => x"63",
          9708 => x"72",
          9709 => x"20",
          9710 => x"20",
          9711 => x"3d",
          9712 => x"2e",
          9713 => x"64",
          9714 => x"0a",
          9715 => x"20",
          9716 => x"69",
          9717 => x"6f",
          9718 => x"53",
          9719 => x"4d",
          9720 => x"6f",
          9721 => x"46",
          9722 => x"3d",
          9723 => x"2e",
          9724 => x"64",
          9725 => x"0a",
          9726 => x"6d",
          9727 => x"00",
          9728 => x"65",
          9729 => x"6d",
          9730 => x"6c",
          9731 => x"00",
          9732 => x"56",
          9733 => x"56",
          9734 => x"6e",
          9735 => x"6e",
          9736 => x"77",
          9737 => x"00",
          9738 => x"00",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"00",
          9752 => x"00",
          9753 => x"00",
          9754 => x"00",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"00",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"00",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"00",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"00",
          9788 => x"00",
          9789 => x"00",
          9790 => x"00",
          9791 => x"00",
          9792 => x"00",
          9793 => x"00",
          9794 => x"00",
          9795 => x"00",
          9796 => x"00",
          9797 => x"00",
          9798 => x"00",
          9799 => x"00",
          9800 => x"00",
          9801 => x"00",
          9802 => x"00",
          9803 => x"5b",
          9804 => x"5b",
          9805 => x"5b",
          9806 => x"5b",
          9807 => x"5b",
          9808 => x"5b",
          9809 => x"5b",
          9810 => x"30",
          9811 => x"5b",
          9812 => x"5b",
          9813 => x"5b",
          9814 => x"00",
          9815 => x"00",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"00",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"00",
          9824 => x"00",
          9825 => x"69",
          9826 => x"72",
          9827 => x"69",
          9828 => x"00",
          9829 => x"00",
          9830 => x"30",
          9831 => x"20",
          9832 => x"00",
          9833 => x"61",
          9834 => x"64",
          9835 => x"20",
          9836 => x"65",
          9837 => x"68",
          9838 => x"69",
          9839 => x"72",
          9840 => x"69",
          9841 => x"74",
          9842 => x"4f",
          9843 => x"00",
          9844 => x"61",
          9845 => x"74",
          9846 => x"65",
          9847 => x"72",
          9848 => x"65",
          9849 => x"73",
          9850 => x"79",
          9851 => x"6c",
          9852 => x"64",
          9853 => x"62",
          9854 => x"67",
          9855 => x"44",
          9856 => x"2a",
          9857 => x"3b",
          9858 => x"3f",
          9859 => x"7f",
          9860 => x"41",
          9861 => x"41",
          9862 => x"00",
          9863 => x"fe",
          9864 => x"44",
          9865 => x"2e",
          9866 => x"4f",
          9867 => x"4d",
          9868 => x"20",
          9869 => x"54",
          9870 => x"20",
          9871 => x"4f",
          9872 => x"4d",
          9873 => x"20",
          9874 => x"54",
          9875 => x"20",
          9876 => x"00",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"9a",
          9881 => x"41",
          9882 => x"45",
          9883 => x"49",
          9884 => x"92",
          9885 => x"4f",
          9886 => x"99",
          9887 => x"9d",
          9888 => x"49",
          9889 => x"a5",
          9890 => x"a9",
          9891 => x"ad",
          9892 => x"b1",
          9893 => x"b5",
          9894 => x"b9",
          9895 => x"bd",
          9896 => x"c1",
          9897 => x"c5",
          9898 => x"c9",
          9899 => x"cd",
          9900 => x"d1",
          9901 => x"d5",
          9902 => x"d9",
          9903 => x"dd",
          9904 => x"e1",
          9905 => x"e5",
          9906 => x"e9",
          9907 => x"ed",
          9908 => x"f1",
          9909 => x"f5",
          9910 => x"f9",
          9911 => x"fd",
          9912 => x"2e",
          9913 => x"5b",
          9914 => x"22",
          9915 => x"3e",
          9916 => x"00",
          9917 => x"01",
          9918 => x"10",
          9919 => x"00",
          9920 => x"00",
          9921 => x"01",
          9922 => x"04",
          9923 => x"10",
          9924 => x"00",
          9925 => x"00",
          9926 => x"00",
          9927 => x"02",
          9928 => x"00",
          9929 => x"00",
          9930 => x"00",
          9931 => x"04",
          9932 => x"00",
          9933 => x"00",
          9934 => x"00",
          9935 => x"14",
          9936 => x"00",
          9937 => x"00",
          9938 => x"00",
          9939 => x"2b",
          9940 => x"00",
          9941 => x"00",
          9942 => x"00",
          9943 => x"30",
          9944 => x"00",
          9945 => x"00",
          9946 => x"00",
          9947 => x"3c",
          9948 => x"00",
          9949 => x"00",
          9950 => x"00",
          9951 => x"3d",
          9952 => x"00",
          9953 => x"00",
          9954 => x"00",
          9955 => x"3f",
          9956 => x"00",
          9957 => x"00",
          9958 => x"00",
          9959 => x"40",
          9960 => x"00",
          9961 => x"00",
          9962 => x"00",
          9963 => x"41",
          9964 => x"00",
          9965 => x"00",
          9966 => x"00",
          9967 => x"42",
          9968 => x"00",
          9969 => x"00",
          9970 => x"00",
          9971 => x"43",
          9972 => x"00",
          9973 => x"00",
          9974 => x"00",
          9975 => x"50",
          9976 => x"00",
          9977 => x"00",
          9978 => x"00",
          9979 => x"51",
          9980 => x"00",
          9981 => x"00",
          9982 => x"00",
          9983 => x"54",
          9984 => x"00",
          9985 => x"00",
          9986 => x"00",
          9987 => x"55",
          9988 => x"00",
          9989 => x"00",
          9990 => x"00",
          9991 => x"79",
          9992 => x"00",
          9993 => x"00",
          9994 => x"00",
          9995 => x"78",
          9996 => x"00",
          9997 => x"00",
          9998 => x"00",
          9999 => x"82",
         10000 => x"00",
         10001 => x"00",
         10002 => x"00",
         10003 => x"83",
         10004 => x"00",
         10005 => x"00",
         10006 => x"00",
         10007 => x"85",
         10008 => x"00",
         10009 => x"00",
         10010 => x"00",
         10011 => x"87",
         10012 => x"00",
         10013 => x"00",
         10014 => x"00",
         10015 => x"8c",
         10016 => x"00",
         10017 => x"00",
         10018 => x"00",
         10019 => x"8d",
         10020 => x"00",
         10021 => x"00",
         10022 => x"00",
         10023 => x"8e",
         10024 => x"00",
         10025 => x"00",
         10026 => x"00",
         10027 => x"8f",
         10028 => x"00",
         10029 => x"00",
         10030 => x"00",
         10031 => x"00",
         10032 => x"00",
         10033 => x"00",
         10034 => x"00",
         10035 => x"01",
         10036 => x"00",
         10037 => x"01",
         10038 => x"81",
         10039 => x"00",
         10040 => x"7f",
         10041 => x"00",
         10042 => x"00",
         10043 => x"00",
         10044 => x"00",
         10045 => x"f5",
         10046 => x"f5",
         10047 => x"f5",
         10048 => x"00",
         10049 => x"01",
         10050 => x"01",
         10051 => x"01",
         10052 => x"00",
         10053 => x"00",
         10054 => x"00",
         10055 => x"00",
         10056 => x"00",
         10057 => x"00",
         10058 => x"00",
         10059 => x"00",
         10060 => x"00",
         10061 => x"00",
         10062 => x"00",
         10063 => x"00",
         10064 => x"00",
         10065 => x"00",
         10066 => x"00",
         10067 => x"00",
         10068 => x"00",
         10069 => x"00",
         10070 => x"00",
         10071 => x"00",
         10072 => x"00",
         10073 => x"00",
         10074 => x"00",
         10075 => x"00",
         10076 => x"00",
         10077 => x"00",
         10078 => x"00",
         10079 => x"00",
         10080 => x"00",
         10081 => x"00",
         10082 => x"00",
         10083 => x"00",
         10084 => x"00",
         10085 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"9b",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"a0",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"94",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"80",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"95",
           269 => x"0b",
           270 => x"0b",
           271 => x"b3",
           272 => x"0b",
           273 => x"0b",
           274 => x"d1",
           275 => x"0b",
           276 => x"0b",
           277 => x"ef",
           278 => x"0b",
           279 => x"0b",
           280 => x"8d",
           281 => x"0b",
           282 => x"0b",
           283 => x"ab",
           284 => x"0b",
           285 => x"0b",
           286 => x"cb",
           287 => x"0b",
           288 => x"0b",
           289 => x"eb",
           290 => x"0b",
           291 => x"0b",
           292 => x"8b",
           293 => x"0b",
           294 => x"0b",
           295 => x"ab",
           296 => x"0b",
           297 => x"0b",
           298 => x"cb",
           299 => x"0b",
           300 => x"0b",
           301 => x"eb",
           302 => x"0b",
           303 => x"0b",
           304 => x"8b",
           305 => x"0b",
           306 => x"0b",
           307 => x"ab",
           308 => x"0b",
           309 => x"0b",
           310 => x"cb",
           311 => x"0b",
           312 => x"0b",
           313 => x"eb",
           314 => x"0b",
           315 => x"0b",
           316 => x"8b",
           317 => x"0b",
           318 => x"0b",
           319 => x"ab",
           320 => x"0b",
           321 => x"0b",
           322 => x"cb",
           323 => x"0b",
           324 => x"0b",
           325 => x"eb",
           326 => x"0b",
           327 => x"0b",
           328 => x"8b",
           329 => x"0b",
           330 => x"0b",
           331 => x"ab",
           332 => x"0b",
           333 => x"0b",
           334 => x"cb",
           335 => x"0b",
           336 => x"0b",
           337 => x"eb",
           338 => x"0b",
           339 => x"0b",
           340 => x"8b",
           341 => x"0b",
           342 => x"0b",
           343 => x"ab",
           344 => x"0b",
           345 => x"0b",
           346 => x"cb",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"04",
           390 => x"0c",
           391 => x"82",
           392 => x"82",
           393 => x"82",
           394 => x"bb",
           395 => x"bb",
           396 => x"e0",
           397 => x"bb",
           398 => x"fc",
           399 => x"a4",
           400 => x"90",
           401 => x"a4",
           402 => x"2d",
           403 => x"08",
           404 => x"04",
           405 => x"0c",
           406 => x"82",
           407 => x"82",
           408 => x"82",
           409 => x"b5",
           410 => x"bb",
           411 => x"e0",
           412 => x"bb",
           413 => x"ab",
           414 => x"a4",
           415 => x"90",
           416 => x"a4",
           417 => x"2d",
           418 => x"08",
           419 => x"04",
           420 => x"0c",
           421 => x"82",
           422 => x"82",
           423 => x"82",
           424 => x"97",
           425 => x"bb",
           426 => x"e0",
           427 => x"bb",
           428 => x"fc",
           429 => x"bb",
           430 => x"e0",
           431 => x"bb",
           432 => x"fc",
           433 => x"bb",
           434 => x"e0",
           435 => x"bb",
           436 => x"f4",
           437 => x"bb",
           438 => x"e0",
           439 => x"bb",
           440 => x"f6",
           441 => x"bb",
           442 => x"e0",
           443 => x"bb",
           444 => x"f7",
           445 => x"bb",
           446 => x"e0",
           447 => x"bb",
           448 => x"dc",
           449 => x"bb",
           450 => x"e0",
           451 => x"bb",
           452 => x"e8",
           453 => x"bb",
           454 => x"e0",
           455 => x"bb",
           456 => x"e0",
           457 => x"bb",
           458 => x"e0",
           459 => x"bb",
           460 => x"e3",
           461 => x"bb",
           462 => x"e0",
           463 => x"bb",
           464 => x"ee",
           465 => x"bb",
           466 => x"e0",
           467 => x"bb",
           468 => x"f6",
           469 => x"bb",
           470 => x"e0",
           471 => x"bb",
           472 => x"e7",
           473 => x"bb",
           474 => x"e0",
           475 => x"bb",
           476 => x"f1",
           477 => x"bb",
           478 => x"e0",
           479 => x"bb",
           480 => x"f2",
           481 => x"bb",
           482 => x"e0",
           483 => x"bb",
           484 => x"f2",
           485 => x"bb",
           486 => x"e0",
           487 => x"bb",
           488 => x"fa",
           489 => x"bb",
           490 => x"e0",
           491 => x"bb",
           492 => x"f8",
           493 => x"bb",
           494 => x"e0",
           495 => x"bb",
           496 => x"fd",
           497 => x"bb",
           498 => x"e0",
           499 => x"bb",
           500 => x"f3",
           501 => x"bb",
           502 => x"e0",
           503 => x"bb",
           504 => x"80",
           505 => x"bb",
           506 => x"e0",
           507 => x"bb",
           508 => x"81",
           509 => x"bb",
           510 => x"e0",
           511 => x"bb",
           512 => x"e9",
           513 => x"bb",
           514 => x"e0",
           515 => x"bb",
           516 => x"e9",
           517 => x"bb",
           518 => x"e0",
           519 => x"bb",
           520 => x"ea",
           521 => x"bb",
           522 => x"e0",
           523 => x"bb",
           524 => x"f4",
           525 => x"bb",
           526 => x"e0",
           527 => x"bb",
           528 => x"82",
           529 => x"bb",
           530 => x"e0",
           531 => x"bb",
           532 => x"84",
           533 => x"bb",
           534 => x"e0",
           535 => x"bb",
           536 => x"87",
           537 => x"bb",
           538 => x"e0",
           539 => x"bb",
           540 => x"db",
           541 => x"bb",
           542 => x"e0",
           543 => x"bb",
           544 => x"8a",
           545 => x"bb",
           546 => x"e0",
           547 => x"bb",
           548 => x"98",
           549 => x"bb",
           550 => x"e0",
           551 => x"bb",
           552 => x"96",
           553 => x"bb",
           554 => x"e0",
           555 => x"bb",
           556 => x"ac",
           557 => x"bb",
           558 => x"e0",
           559 => x"bb",
           560 => x"ae",
           561 => x"bb",
           562 => x"e0",
           563 => x"bb",
           564 => x"b0",
           565 => x"bb",
           566 => x"e0",
           567 => x"bb",
           568 => x"f4",
           569 => x"bb",
           570 => x"e0",
           571 => x"bb",
           572 => x"f6",
           573 => x"bb",
           574 => x"e0",
           575 => x"bb",
           576 => x"f9",
           577 => x"bb",
           578 => x"e0",
           579 => x"bb",
           580 => x"d6",
           581 => x"bb",
           582 => x"e0",
           583 => x"bb",
           584 => x"a6",
           585 => x"bb",
           586 => x"e0",
           587 => x"bb",
           588 => x"a7",
           589 => x"bb",
           590 => x"e0",
           591 => x"bb",
           592 => x"ab",
           593 => x"bb",
           594 => x"e0",
           595 => x"bb",
           596 => x"a3",
           597 => x"bb",
           598 => x"e0",
           599 => x"04",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"04",
           609 => x"81",
           610 => x"83",
           611 => x"05",
           612 => x"10",
           613 => x"72",
           614 => x"51",
           615 => x"72",
           616 => x"06",
           617 => x"72",
           618 => x"10",
           619 => x"10",
           620 => x"ed",
           621 => x"53",
           622 => x"bb",
           623 => x"d2",
           624 => x"38",
           625 => x"84",
           626 => x"0b",
           627 => x"ba",
           628 => x"51",
           629 => x"04",
           630 => x"a4",
           631 => x"bb",
           632 => x"3d",
           633 => x"a4",
           634 => x"70",
           635 => x"08",
           636 => x"82",
           637 => x"fc",
           638 => x"82",
           639 => x"88",
           640 => x"82",
           641 => x"52",
           642 => x"3f",
           643 => x"08",
           644 => x"a4",
           645 => x"0c",
           646 => x"08",
           647 => x"70",
           648 => x"0c",
           649 => x"3d",
           650 => x"a4",
           651 => x"bb",
           652 => x"82",
           653 => x"fb",
           654 => x"bb",
           655 => x"05",
           656 => x"33",
           657 => x"70",
           658 => x"51",
           659 => x"8f",
           660 => x"82",
           661 => x"8c",
           662 => x"83",
           663 => x"80",
           664 => x"a4",
           665 => x"0c",
           666 => x"82",
           667 => x"8c",
           668 => x"05",
           669 => x"08",
           670 => x"80",
           671 => x"a4",
           672 => x"0c",
           673 => x"08",
           674 => x"82",
           675 => x"fc",
           676 => x"bb",
           677 => x"05",
           678 => x"80",
           679 => x"0b",
           680 => x"08",
           681 => x"25",
           682 => x"82",
           683 => x"90",
           684 => x"ab",
           685 => x"bb",
           686 => x"82",
           687 => x"f8",
           688 => x"82",
           689 => x"f8",
           690 => x"2e",
           691 => x"8d",
           692 => x"82",
           693 => x"f4",
           694 => x"d2",
           695 => x"a4",
           696 => x"08",
           697 => x"08",
           698 => x"53",
           699 => x"34",
           700 => x"08",
           701 => x"ff",
           702 => x"a4",
           703 => x"0c",
           704 => x"08",
           705 => x"81",
           706 => x"a4",
           707 => x"0c",
           708 => x"82",
           709 => x"fc",
           710 => x"80",
           711 => x"bb",
           712 => x"05",
           713 => x"bb",
           714 => x"05",
           715 => x"bb",
           716 => x"05",
           717 => x"98",
           718 => x"0d",
           719 => x"0c",
           720 => x"a4",
           721 => x"bb",
           722 => x"3d",
           723 => x"82",
           724 => x"e5",
           725 => x"bb",
           726 => x"05",
           727 => x"a4",
           728 => x"0c",
           729 => x"82",
           730 => x"e8",
           731 => x"bb",
           732 => x"05",
           733 => x"a4",
           734 => x"0c",
           735 => x"08",
           736 => x"54",
           737 => x"08",
           738 => x"53",
           739 => x"08",
           740 => x"53",
           741 => x"8d",
           742 => x"98",
           743 => x"bb",
           744 => x"05",
           745 => x"a4",
           746 => x"08",
           747 => x"08",
           748 => x"05",
           749 => x"74",
           750 => x"a4",
           751 => x"08",
           752 => x"98",
           753 => x"3d",
           754 => x"a4",
           755 => x"bb",
           756 => x"82",
           757 => x"fb",
           758 => x"bb",
           759 => x"05",
           760 => x"a4",
           761 => x"0c",
           762 => x"08",
           763 => x"54",
           764 => x"08",
           765 => x"53",
           766 => x"08",
           767 => x"52",
           768 => x"82",
           769 => x"70",
           770 => x"08",
           771 => x"82",
           772 => x"f8",
           773 => x"82",
           774 => x"51",
           775 => x"0d",
           776 => x"0c",
           777 => x"a4",
           778 => x"bb",
           779 => x"3d",
           780 => x"82",
           781 => x"e4",
           782 => x"bb",
           783 => x"05",
           784 => x"0b",
           785 => x"82",
           786 => x"88",
           787 => x"11",
           788 => x"2a",
           789 => x"70",
           790 => x"51",
           791 => x"72",
           792 => x"38",
           793 => x"bb",
           794 => x"05",
           795 => x"39",
           796 => x"08",
           797 => x"53",
           798 => x"72",
           799 => x"08",
           800 => x"72",
           801 => x"53",
           802 => x"95",
           803 => x"bb",
           804 => x"05",
           805 => x"82",
           806 => x"8c",
           807 => x"bb",
           808 => x"05",
           809 => x"06",
           810 => x"80",
           811 => x"38",
           812 => x"08",
           813 => x"53",
           814 => x"81",
           815 => x"bb",
           816 => x"05",
           817 => x"b9",
           818 => x"38",
           819 => x"08",
           820 => x"53",
           821 => x"09",
           822 => x"c5",
           823 => x"a4",
           824 => x"33",
           825 => x"70",
           826 => x"51",
           827 => x"38",
           828 => x"08",
           829 => x"70",
           830 => x"81",
           831 => x"06",
           832 => x"53",
           833 => x"99",
           834 => x"a4",
           835 => x"22",
           836 => x"07",
           837 => x"82",
           838 => x"e4",
           839 => x"d0",
           840 => x"a4",
           841 => x"33",
           842 => x"70",
           843 => x"70",
           844 => x"11",
           845 => x"51",
           846 => x"55",
           847 => x"bb",
           848 => x"05",
           849 => x"a4",
           850 => x"33",
           851 => x"a4",
           852 => x"33",
           853 => x"11",
           854 => x"72",
           855 => x"08",
           856 => x"82",
           857 => x"e8",
           858 => x"98",
           859 => x"2c",
           860 => x"72",
           861 => x"38",
           862 => x"82",
           863 => x"e8",
           864 => x"bb",
           865 => x"05",
           866 => x"2a",
           867 => x"51",
           868 => x"fd",
           869 => x"bb",
           870 => x"05",
           871 => x"2b",
           872 => x"70",
           873 => x"88",
           874 => x"51",
           875 => x"82",
           876 => x"ec",
           877 => x"b8",
           878 => x"a4",
           879 => x"22",
           880 => x"70",
           881 => x"51",
           882 => x"2e",
           883 => x"bb",
           884 => x"05",
           885 => x"2b",
           886 => x"51",
           887 => x"8a",
           888 => x"82",
           889 => x"e8",
           890 => x"bb",
           891 => x"05",
           892 => x"82",
           893 => x"c4",
           894 => x"82",
           895 => x"c4",
           896 => x"d8",
           897 => x"38",
           898 => x"08",
           899 => x"70",
           900 => x"9a",
           901 => x"08",
           902 => x"53",
           903 => x"bb",
           904 => x"05",
           905 => x"07",
           906 => x"82",
           907 => x"e4",
           908 => x"bb",
           909 => x"05",
           910 => x"07",
           911 => x"82",
           912 => x"e4",
           913 => x"a8",
           914 => x"a4",
           915 => x"22",
           916 => x"07",
           917 => x"82",
           918 => x"e4",
           919 => x"90",
           920 => x"a4",
           921 => x"22",
           922 => x"07",
           923 => x"82",
           924 => x"e4",
           925 => x"f8",
           926 => x"a4",
           927 => x"22",
           928 => x"51",
           929 => x"bb",
           930 => x"05",
           931 => x"82",
           932 => x"e8",
           933 => x"d8",
           934 => x"a4",
           935 => x"22",
           936 => x"51",
           937 => x"bb",
           938 => x"05",
           939 => x"39",
           940 => x"bb",
           941 => x"05",
           942 => x"a4",
           943 => x"22",
           944 => x"53",
           945 => x"a4",
           946 => x"23",
           947 => x"82",
           948 => x"f8",
           949 => x"a8",
           950 => x"a4",
           951 => x"08",
           952 => x"08",
           953 => x"84",
           954 => x"a4",
           955 => x"0c",
           956 => x"53",
           957 => x"a4",
           958 => x"34",
           959 => x"08",
           960 => x"ff",
           961 => x"72",
           962 => x"08",
           963 => x"8c",
           964 => x"bb",
           965 => x"05",
           966 => x"a4",
           967 => x"08",
           968 => x"bb",
           969 => x"05",
           970 => x"82",
           971 => x"fc",
           972 => x"bb",
           973 => x"05",
           974 => x"2a",
           975 => x"51",
           976 => x"72",
           977 => x"38",
           978 => x"08",
           979 => x"70",
           980 => x"72",
           981 => x"82",
           982 => x"fc",
           983 => x"53",
           984 => x"82",
           985 => x"53",
           986 => x"a4",
           987 => x"23",
           988 => x"bb",
           989 => x"05",
           990 => x"ac",
           991 => x"98",
           992 => x"82",
           993 => x"f4",
           994 => x"bb",
           995 => x"05",
           996 => x"bb",
           997 => x"05",
           998 => x"31",
           999 => x"82",
          1000 => x"ec",
          1001 => x"d8",
          1002 => x"a4",
          1003 => x"08",
          1004 => x"08",
          1005 => x"84",
          1006 => x"a4",
          1007 => x"0c",
          1008 => x"bb",
          1009 => x"05",
          1010 => x"a4",
          1011 => x"22",
          1012 => x"70",
          1013 => x"51",
          1014 => x"80",
          1015 => x"82",
          1016 => x"e8",
          1017 => x"98",
          1018 => x"98",
          1019 => x"bb",
          1020 => x"05",
          1021 => x"ac",
          1022 => x"bb",
          1023 => x"72",
          1024 => x"08",
          1025 => x"99",
          1026 => x"a4",
          1027 => x"08",
          1028 => x"3f",
          1029 => x"08",
          1030 => x"bb",
          1031 => x"05",
          1032 => x"a4",
          1033 => x"22",
          1034 => x"a4",
          1035 => x"22",
          1036 => x"54",
          1037 => x"bb",
          1038 => x"05",
          1039 => x"39",
          1040 => x"08",
          1041 => x"70",
          1042 => x"81",
          1043 => x"53",
          1044 => x"a4",
          1045 => x"a4",
          1046 => x"08",
          1047 => x"08",
          1048 => x"84",
          1049 => x"a4",
          1050 => x"0c",
          1051 => x"bb",
          1052 => x"05",
          1053 => x"39",
          1054 => x"08",
          1055 => x"82",
          1056 => x"90",
          1057 => x"05",
          1058 => x"08",
          1059 => x"70",
          1060 => x"a4",
          1061 => x"0c",
          1062 => x"a4",
          1063 => x"08",
          1064 => x"08",
          1065 => x"82",
          1066 => x"fc",
          1067 => x"25",
          1068 => x"bb",
          1069 => x"05",
          1070 => x"07",
          1071 => x"82",
          1072 => x"e4",
          1073 => x"bb",
          1074 => x"05",
          1075 => x"bb",
          1076 => x"05",
          1077 => x"a4",
          1078 => x"22",
          1079 => x"06",
          1080 => x"82",
          1081 => x"e4",
          1082 => x"af",
          1083 => x"82",
          1084 => x"f4",
          1085 => x"39",
          1086 => x"08",
          1087 => x"70",
          1088 => x"51",
          1089 => x"bb",
          1090 => x"05",
          1091 => x"0b",
          1092 => x"08",
          1093 => x"90",
          1094 => x"a4",
          1095 => x"23",
          1096 => x"08",
          1097 => x"70",
          1098 => x"81",
          1099 => x"53",
          1100 => x"a4",
          1101 => x"a4",
          1102 => x"08",
          1103 => x"08",
          1104 => x"84",
          1105 => x"a4",
          1106 => x"0c",
          1107 => x"bb",
          1108 => x"05",
          1109 => x"39",
          1110 => x"08",
          1111 => x"82",
          1112 => x"90",
          1113 => x"05",
          1114 => x"08",
          1115 => x"70",
          1116 => x"a4",
          1117 => x"0c",
          1118 => x"a4",
          1119 => x"08",
          1120 => x"08",
          1121 => x"82",
          1122 => x"e4",
          1123 => x"cf",
          1124 => x"72",
          1125 => x"08",
          1126 => x"82",
          1127 => x"82",
          1128 => x"f0",
          1129 => x"bb",
          1130 => x"05",
          1131 => x"a4",
          1132 => x"22",
          1133 => x"08",
          1134 => x"71",
          1135 => x"56",
          1136 => x"95",
          1137 => x"98",
          1138 => x"75",
          1139 => x"a4",
          1140 => x"08",
          1141 => x"08",
          1142 => x"82",
          1143 => x"f0",
          1144 => x"33",
          1145 => x"73",
          1146 => x"82",
          1147 => x"f0",
          1148 => x"72",
          1149 => x"bb",
          1150 => x"05",
          1151 => x"df",
          1152 => x"53",
          1153 => x"a4",
          1154 => x"34",
          1155 => x"bb",
          1156 => x"05",
          1157 => x"33",
          1158 => x"53",
          1159 => x"a4",
          1160 => x"34",
          1161 => x"08",
          1162 => x"53",
          1163 => x"08",
          1164 => x"73",
          1165 => x"a4",
          1166 => x"08",
          1167 => x"bb",
          1168 => x"05",
          1169 => x"a4",
          1170 => x"22",
          1171 => x"bb",
          1172 => x"05",
          1173 => x"ad",
          1174 => x"bb",
          1175 => x"82",
          1176 => x"fc",
          1177 => x"82",
          1178 => x"fc",
          1179 => x"2e",
          1180 => x"b2",
          1181 => x"a4",
          1182 => x"08",
          1183 => x"54",
          1184 => x"74",
          1185 => x"51",
          1186 => x"bb",
          1187 => x"05",
          1188 => x"a4",
          1189 => x"22",
          1190 => x"51",
          1191 => x"2e",
          1192 => x"bb",
          1193 => x"05",
          1194 => x"51",
          1195 => x"bb",
          1196 => x"05",
          1197 => x"a4",
          1198 => x"22",
          1199 => x"70",
          1200 => x"51",
          1201 => x"2e",
          1202 => x"82",
          1203 => x"ec",
          1204 => x"90",
          1205 => x"a4",
          1206 => x"0c",
          1207 => x"08",
          1208 => x"90",
          1209 => x"a4",
          1210 => x"0c",
          1211 => x"08",
          1212 => x"51",
          1213 => x"2e",
          1214 => x"95",
          1215 => x"a4",
          1216 => x"08",
          1217 => x"72",
          1218 => x"08",
          1219 => x"93",
          1220 => x"a4",
          1221 => x"08",
          1222 => x"72",
          1223 => x"08",
          1224 => x"82",
          1225 => x"c8",
          1226 => x"bb",
          1227 => x"05",
          1228 => x"a4",
          1229 => x"22",
          1230 => x"70",
          1231 => x"51",
          1232 => x"2e",
          1233 => x"82",
          1234 => x"e8",
          1235 => x"98",
          1236 => x"2c",
          1237 => x"08",
          1238 => x"57",
          1239 => x"72",
          1240 => x"38",
          1241 => x"08",
          1242 => x"70",
          1243 => x"53",
          1244 => x"a4",
          1245 => x"23",
          1246 => x"bb",
          1247 => x"05",
          1248 => x"bb",
          1249 => x"05",
          1250 => x"31",
          1251 => x"82",
          1252 => x"e8",
          1253 => x"bb",
          1254 => x"05",
          1255 => x"2a",
          1256 => x"51",
          1257 => x"80",
          1258 => x"82",
          1259 => x"e8",
          1260 => x"88",
          1261 => x"2b",
          1262 => x"70",
          1263 => x"51",
          1264 => x"72",
          1265 => x"a4",
          1266 => x"22",
          1267 => x"51",
          1268 => x"bb",
          1269 => x"05",
          1270 => x"82",
          1271 => x"fc",
          1272 => x"88",
          1273 => x"2b",
          1274 => x"70",
          1275 => x"51",
          1276 => x"72",
          1277 => x"a4",
          1278 => x"22",
          1279 => x"51",
          1280 => x"bb",
          1281 => x"05",
          1282 => x"a4",
          1283 => x"22",
          1284 => x"06",
          1285 => x"b0",
          1286 => x"a4",
          1287 => x"22",
          1288 => x"54",
          1289 => x"a4",
          1290 => x"23",
          1291 => x"70",
          1292 => x"53",
          1293 => x"90",
          1294 => x"a4",
          1295 => x"08",
          1296 => x"96",
          1297 => x"39",
          1298 => x"08",
          1299 => x"70",
          1300 => x"81",
          1301 => x"53",
          1302 => x"91",
          1303 => x"a4",
          1304 => x"08",
          1305 => x"95",
          1306 => x"c7",
          1307 => x"a4",
          1308 => x"22",
          1309 => x"70",
          1310 => x"51",
          1311 => x"2e",
          1312 => x"bb",
          1313 => x"05",
          1314 => x"51",
          1315 => x"a3",
          1316 => x"a4",
          1317 => x"22",
          1318 => x"70",
          1319 => x"51",
          1320 => x"2e",
          1321 => x"bb",
          1322 => x"05",
          1323 => x"51",
          1324 => x"82",
          1325 => x"e4",
          1326 => x"86",
          1327 => x"06",
          1328 => x"72",
          1329 => x"38",
          1330 => x"08",
          1331 => x"52",
          1332 => x"81",
          1333 => x"a4",
          1334 => x"22",
          1335 => x"2e",
          1336 => x"94",
          1337 => x"a4",
          1338 => x"08",
          1339 => x"a4",
          1340 => x"33",
          1341 => x"3f",
          1342 => x"08",
          1343 => x"70",
          1344 => x"81",
          1345 => x"53",
          1346 => x"b0",
          1347 => x"a4",
          1348 => x"22",
          1349 => x"54",
          1350 => x"a4",
          1351 => x"23",
          1352 => x"70",
          1353 => x"53",
          1354 => x"90",
          1355 => x"a4",
          1356 => x"08",
          1357 => x"94",
          1358 => x"39",
          1359 => x"08",
          1360 => x"70",
          1361 => x"81",
          1362 => x"53",
          1363 => x"b0",
          1364 => x"a4",
          1365 => x"33",
          1366 => x"54",
          1367 => x"a4",
          1368 => x"34",
          1369 => x"70",
          1370 => x"53",
          1371 => x"90",
          1372 => x"a4",
          1373 => x"08",
          1374 => x"93",
          1375 => x"39",
          1376 => x"08",
          1377 => x"70",
          1378 => x"81",
          1379 => x"53",
          1380 => x"82",
          1381 => x"ec",
          1382 => x"11",
          1383 => x"82",
          1384 => x"ec",
          1385 => x"90",
          1386 => x"2c",
          1387 => x"73",
          1388 => x"82",
          1389 => x"88",
          1390 => x"a0",
          1391 => x"3f",
          1392 => x"bb",
          1393 => x"05",
          1394 => x"80",
          1395 => x"81",
          1396 => x"82",
          1397 => x"88",
          1398 => x"82",
          1399 => x"fc",
          1400 => x"92",
          1401 => x"ee",
          1402 => x"a4",
          1403 => x"33",
          1404 => x"f3",
          1405 => x"06",
          1406 => x"82",
          1407 => x"f4",
          1408 => x"11",
          1409 => x"82",
          1410 => x"f4",
          1411 => x"83",
          1412 => x"53",
          1413 => x"ff",
          1414 => x"38",
          1415 => x"08",
          1416 => x"52",
          1417 => x"08",
          1418 => x"70",
          1419 => x"bb",
          1420 => x"05",
          1421 => x"82",
          1422 => x"fc",
          1423 => x"92",
          1424 => x"b7",
          1425 => x"a4",
          1426 => x"33",
          1427 => x"d3",
          1428 => x"06",
          1429 => x"82",
          1430 => x"f4",
          1431 => x"11",
          1432 => x"82",
          1433 => x"f4",
          1434 => x"83",
          1435 => x"53",
          1436 => x"ff",
          1437 => x"38",
          1438 => x"08",
          1439 => x"52",
          1440 => x"08",
          1441 => x"70",
          1442 => x"91",
          1443 => x"bb",
          1444 => x"05",
          1445 => x"82",
          1446 => x"fc",
          1447 => x"b7",
          1448 => x"a4",
          1449 => x"08",
          1450 => x"2e",
          1451 => x"bb",
          1452 => x"05",
          1453 => x"bb",
          1454 => x"05",
          1455 => x"82",
          1456 => x"f0",
          1457 => x"bb",
          1458 => x"05",
          1459 => x"52",
          1460 => x"3f",
          1461 => x"bb",
          1462 => x"05",
          1463 => x"2a",
          1464 => x"51",
          1465 => x"80",
          1466 => x"38",
          1467 => x"08",
          1468 => x"ff",
          1469 => x"72",
          1470 => x"08",
          1471 => x"73",
          1472 => x"90",
          1473 => x"80",
          1474 => x"38",
          1475 => x"08",
          1476 => x"52",
          1477 => x"bd",
          1478 => x"82",
          1479 => x"88",
          1480 => x"82",
          1481 => x"f8",
          1482 => x"90",
          1483 => x"0b",
          1484 => x"08",
          1485 => x"ea",
          1486 => x"bb",
          1487 => x"05",
          1488 => x"a5",
          1489 => x"06",
          1490 => x"0b",
          1491 => x"08",
          1492 => x"80",
          1493 => x"a4",
          1494 => x"23",
          1495 => x"bb",
          1496 => x"05",
          1497 => x"82",
          1498 => x"f4",
          1499 => x"80",
          1500 => x"a4",
          1501 => x"08",
          1502 => x"a4",
          1503 => x"33",
          1504 => x"3f",
          1505 => x"82",
          1506 => x"88",
          1507 => x"11",
          1508 => x"bb",
          1509 => x"05",
          1510 => x"82",
          1511 => x"e0",
          1512 => x"bb",
          1513 => x"3d",
          1514 => x"a4",
          1515 => x"bb",
          1516 => x"82",
          1517 => x"f7",
          1518 => x"0b",
          1519 => x"08",
          1520 => x"82",
          1521 => x"8c",
          1522 => x"80",
          1523 => x"bb",
          1524 => x"05",
          1525 => x"51",
          1526 => x"53",
          1527 => x"a4",
          1528 => x"34",
          1529 => x"06",
          1530 => x"2e",
          1531 => x"91",
          1532 => x"a4",
          1533 => x"08",
          1534 => x"05",
          1535 => x"ce",
          1536 => x"a4",
          1537 => x"33",
          1538 => x"2e",
          1539 => x"a4",
          1540 => x"82",
          1541 => x"f0",
          1542 => x"bb",
          1543 => x"05",
          1544 => x"81",
          1545 => x"70",
          1546 => x"72",
          1547 => x"a4",
          1548 => x"34",
          1549 => x"08",
          1550 => x"53",
          1551 => x"09",
          1552 => x"dc",
          1553 => x"a4",
          1554 => x"08",
          1555 => x"05",
          1556 => x"08",
          1557 => x"33",
          1558 => x"08",
          1559 => x"82",
          1560 => x"f8",
          1561 => x"bb",
          1562 => x"05",
          1563 => x"a4",
          1564 => x"08",
          1565 => x"b6",
          1566 => x"a4",
          1567 => x"08",
          1568 => x"84",
          1569 => x"39",
          1570 => x"bb",
          1571 => x"05",
          1572 => x"a4",
          1573 => x"08",
          1574 => x"05",
          1575 => x"08",
          1576 => x"33",
          1577 => x"08",
          1578 => x"81",
          1579 => x"0b",
          1580 => x"08",
          1581 => x"82",
          1582 => x"88",
          1583 => x"08",
          1584 => x"0c",
          1585 => x"53",
          1586 => x"bb",
          1587 => x"05",
          1588 => x"39",
          1589 => x"08",
          1590 => x"53",
          1591 => x"8d",
          1592 => x"82",
          1593 => x"ec",
          1594 => x"80",
          1595 => x"a4",
          1596 => x"33",
          1597 => x"27",
          1598 => x"bb",
          1599 => x"05",
          1600 => x"b9",
          1601 => x"8d",
          1602 => x"82",
          1603 => x"ec",
          1604 => x"d8",
          1605 => x"82",
          1606 => x"f4",
          1607 => x"39",
          1608 => x"08",
          1609 => x"53",
          1610 => x"90",
          1611 => x"a4",
          1612 => x"33",
          1613 => x"26",
          1614 => x"39",
          1615 => x"bb",
          1616 => x"05",
          1617 => x"39",
          1618 => x"bb",
          1619 => x"05",
          1620 => x"82",
          1621 => x"fc",
          1622 => x"bb",
          1623 => x"05",
          1624 => x"73",
          1625 => x"38",
          1626 => x"08",
          1627 => x"53",
          1628 => x"27",
          1629 => x"bb",
          1630 => x"05",
          1631 => x"51",
          1632 => x"bb",
          1633 => x"05",
          1634 => x"a4",
          1635 => x"33",
          1636 => x"53",
          1637 => x"a4",
          1638 => x"34",
          1639 => x"08",
          1640 => x"53",
          1641 => x"ad",
          1642 => x"a4",
          1643 => x"33",
          1644 => x"53",
          1645 => x"a4",
          1646 => x"34",
          1647 => x"08",
          1648 => x"53",
          1649 => x"8d",
          1650 => x"82",
          1651 => x"ec",
          1652 => x"98",
          1653 => x"a4",
          1654 => x"33",
          1655 => x"08",
          1656 => x"54",
          1657 => x"26",
          1658 => x"0b",
          1659 => x"08",
          1660 => x"80",
          1661 => x"bb",
          1662 => x"05",
          1663 => x"bb",
          1664 => x"05",
          1665 => x"bb",
          1666 => x"05",
          1667 => x"82",
          1668 => x"fc",
          1669 => x"bb",
          1670 => x"05",
          1671 => x"81",
          1672 => x"70",
          1673 => x"52",
          1674 => x"33",
          1675 => x"08",
          1676 => x"fe",
          1677 => x"bb",
          1678 => x"05",
          1679 => x"80",
          1680 => x"82",
          1681 => x"fc",
          1682 => x"82",
          1683 => x"fc",
          1684 => x"bb",
          1685 => x"05",
          1686 => x"a4",
          1687 => x"08",
          1688 => x"81",
          1689 => x"a4",
          1690 => x"0c",
          1691 => x"08",
          1692 => x"82",
          1693 => x"8b",
          1694 => x"bb",
          1695 => x"82",
          1696 => x"02",
          1697 => x"0c",
          1698 => x"82",
          1699 => x"53",
          1700 => x"08",
          1701 => x"52",
          1702 => x"08",
          1703 => x"51",
          1704 => x"82",
          1705 => x"70",
          1706 => x"0c",
          1707 => x"0d",
          1708 => x"0c",
          1709 => x"a4",
          1710 => x"bb",
          1711 => x"3d",
          1712 => x"82",
          1713 => x"f0",
          1714 => x"bb",
          1715 => x"05",
          1716 => x"73",
          1717 => x"a4",
          1718 => x"08",
          1719 => x"53",
          1720 => x"72",
          1721 => x"08",
          1722 => x"72",
          1723 => x"53",
          1724 => x"09",
          1725 => x"38",
          1726 => x"08",
          1727 => x"70",
          1728 => x"71",
          1729 => x"39",
          1730 => x"08",
          1731 => x"53",
          1732 => x"09",
          1733 => x"38",
          1734 => x"bb",
          1735 => x"05",
          1736 => x"a4",
          1737 => x"08",
          1738 => x"05",
          1739 => x"08",
          1740 => x"33",
          1741 => x"08",
          1742 => x"82",
          1743 => x"f8",
          1744 => x"72",
          1745 => x"81",
          1746 => x"38",
          1747 => x"08",
          1748 => x"70",
          1749 => x"71",
          1750 => x"51",
          1751 => x"82",
          1752 => x"f8",
          1753 => x"bb",
          1754 => x"05",
          1755 => x"a4",
          1756 => x"0c",
          1757 => x"08",
          1758 => x"80",
          1759 => x"38",
          1760 => x"08",
          1761 => x"80",
          1762 => x"38",
          1763 => x"90",
          1764 => x"a4",
          1765 => x"34",
          1766 => x"08",
          1767 => x"70",
          1768 => x"71",
          1769 => x"51",
          1770 => x"82",
          1771 => x"f8",
          1772 => x"a4",
          1773 => x"82",
          1774 => x"f4",
          1775 => x"bb",
          1776 => x"05",
          1777 => x"81",
          1778 => x"70",
          1779 => x"72",
          1780 => x"a4",
          1781 => x"34",
          1782 => x"82",
          1783 => x"f8",
          1784 => x"72",
          1785 => x"38",
          1786 => x"bb",
          1787 => x"05",
          1788 => x"39",
          1789 => x"08",
          1790 => x"53",
          1791 => x"90",
          1792 => x"a4",
          1793 => x"33",
          1794 => x"26",
          1795 => x"39",
          1796 => x"bb",
          1797 => x"05",
          1798 => x"39",
          1799 => x"bb",
          1800 => x"05",
          1801 => x"82",
          1802 => x"f8",
          1803 => x"af",
          1804 => x"38",
          1805 => x"08",
          1806 => x"53",
          1807 => x"83",
          1808 => x"80",
          1809 => x"a4",
          1810 => x"0c",
          1811 => x"8a",
          1812 => x"a4",
          1813 => x"34",
          1814 => x"bb",
          1815 => x"05",
          1816 => x"a4",
          1817 => x"33",
          1818 => x"27",
          1819 => x"82",
          1820 => x"f8",
          1821 => x"80",
          1822 => x"94",
          1823 => x"a4",
          1824 => x"33",
          1825 => x"53",
          1826 => x"a4",
          1827 => x"34",
          1828 => x"08",
          1829 => x"d0",
          1830 => x"72",
          1831 => x"08",
          1832 => x"82",
          1833 => x"f8",
          1834 => x"90",
          1835 => x"38",
          1836 => x"08",
          1837 => x"f9",
          1838 => x"72",
          1839 => x"08",
          1840 => x"82",
          1841 => x"f8",
          1842 => x"72",
          1843 => x"38",
          1844 => x"bb",
          1845 => x"05",
          1846 => x"39",
          1847 => x"08",
          1848 => x"82",
          1849 => x"f4",
          1850 => x"54",
          1851 => x"8d",
          1852 => x"82",
          1853 => x"ec",
          1854 => x"f7",
          1855 => x"a4",
          1856 => x"33",
          1857 => x"a4",
          1858 => x"08",
          1859 => x"a4",
          1860 => x"33",
          1861 => x"bb",
          1862 => x"05",
          1863 => x"a4",
          1864 => x"08",
          1865 => x"05",
          1866 => x"08",
          1867 => x"55",
          1868 => x"82",
          1869 => x"f8",
          1870 => x"a5",
          1871 => x"a4",
          1872 => x"33",
          1873 => x"2e",
          1874 => x"bb",
          1875 => x"05",
          1876 => x"bb",
          1877 => x"05",
          1878 => x"a4",
          1879 => x"08",
          1880 => x"08",
          1881 => x"71",
          1882 => x"0b",
          1883 => x"08",
          1884 => x"82",
          1885 => x"ec",
          1886 => x"bb",
          1887 => x"3d",
          1888 => x"a4",
          1889 => x"bb",
          1890 => x"82",
          1891 => x"fb",
          1892 => x"0b",
          1893 => x"08",
          1894 => x"82",
          1895 => x"85",
          1896 => x"81",
          1897 => x"32",
          1898 => x"51",
          1899 => x"53",
          1900 => x"8d",
          1901 => x"82",
          1902 => x"f4",
          1903 => x"92",
          1904 => x"a4",
          1905 => x"08",
          1906 => x"82",
          1907 => x"88",
          1908 => x"05",
          1909 => x"08",
          1910 => x"53",
          1911 => x"a4",
          1912 => x"34",
          1913 => x"06",
          1914 => x"2e",
          1915 => x"d2",
          1916 => x"d2",
          1917 => x"82",
          1918 => x"fc",
          1919 => x"90",
          1920 => x"53",
          1921 => x"bb",
          1922 => x"72",
          1923 => x"b1",
          1924 => x"82",
          1925 => x"f8",
          1926 => x"a5",
          1927 => x"ec",
          1928 => x"ec",
          1929 => x"8a",
          1930 => x"08",
          1931 => x"82",
          1932 => x"53",
          1933 => x"8a",
          1934 => x"82",
          1935 => x"f8",
          1936 => x"bb",
          1937 => x"05",
          1938 => x"bb",
          1939 => x"05",
          1940 => x"bb",
          1941 => x"05",
          1942 => x"98",
          1943 => x"0d",
          1944 => x"0c",
          1945 => x"a4",
          1946 => x"bb",
          1947 => x"3d",
          1948 => x"82",
          1949 => x"f8",
          1950 => x"bb",
          1951 => x"05",
          1952 => x"33",
          1953 => x"70",
          1954 => x"81",
          1955 => x"51",
          1956 => x"80",
          1957 => x"ff",
          1958 => x"a4",
          1959 => x"0c",
          1960 => x"82",
          1961 => x"88",
          1962 => x"72",
          1963 => x"a4",
          1964 => x"08",
          1965 => x"bb",
          1966 => x"05",
          1967 => x"82",
          1968 => x"fc",
          1969 => x"81",
          1970 => x"72",
          1971 => x"38",
          1972 => x"08",
          1973 => x"82",
          1974 => x"8c",
          1975 => x"82",
          1976 => x"fc",
          1977 => x"90",
          1978 => x"53",
          1979 => x"bb",
          1980 => x"72",
          1981 => x"ab",
          1982 => x"82",
          1983 => x"f8",
          1984 => x"9f",
          1985 => x"a4",
          1986 => x"08",
          1987 => x"a4",
          1988 => x"0c",
          1989 => x"a4",
          1990 => x"08",
          1991 => x"0c",
          1992 => x"82",
          1993 => x"04",
          1994 => x"08",
          1995 => x"a4",
          1996 => x"0d",
          1997 => x"08",
          1998 => x"a4",
          1999 => x"08",
          2000 => x"82",
          2001 => x"70",
          2002 => x"0c",
          2003 => x"0d",
          2004 => x"0c",
          2005 => x"a4",
          2006 => x"bb",
          2007 => x"3d",
          2008 => x"a4",
          2009 => x"08",
          2010 => x"70",
          2011 => x"81",
          2012 => x"06",
          2013 => x"51",
          2014 => x"2e",
          2015 => x"0b",
          2016 => x"08",
          2017 => x"81",
          2018 => x"bb",
          2019 => x"05",
          2020 => x"33",
          2021 => x"70",
          2022 => x"51",
          2023 => x"80",
          2024 => x"38",
          2025 => x"08",
          2026 => x"82",
          2027 => x"8c",
          2028 => x"54",
          2029 => x"88",
          2030 => x"9f",
          2031 => x"a4",
          2032 => x"08",
          2033 => x"82",
          2034 => x"88",
          2035 => x"57",
          2036 => x"75",
          2037 => x"81",
          2038 => x"82",
          2039 => x"8c",
          2040 => x"11",
          2041 => x"8c",
          2042 => x"bb",
          2043 => x"05",
          2044 => x"bb",
          2045 => x"05",
          2046 => x"80",
          2047 => x"bb",
          2048 => x"05",
          2049 => x"a4",
          2050 => x"08",
          2051 => x"a4",
          2052 => x"08",
          2053 => x"06",
          2054 => x"08",
          2055 => x"72",
          2056 => x"98",
          2057 => x"a3",
          2058 => x"a4",
          2059 => x"08",
          2060 => x"81",
          2061 => x"0c",
          2062 => x"08",
          2063 => x"70",
          2064 => x"08",
          2065 => x"51",
          2066 => x"ff",
          2067 => x"a4",
          2068 => x"0c",
          2069 => x"08",
          2070 => x"82",
          2071 => x"87",
          2072 => x"bb",
          2073 => x"82",
          2074 => x"02",
          2075 => x"0c",
          2076 => x"82",
          2077 => x"88",
          2078 => x"11",
          2079 => x"32",
          2080 => x"51",
          2081 => x"71",
          2082 => x"38",
          2083 => x"bb",
          2084 => x"05",
          2085 => x"39",
          2086 => x"08",
          2087 => x"85",
          2088 => x"86",
          2089 => x"06",
          2090 => x"52",
          2091 => x"80",
          2092 => x"bb",
          2093 => x"05",
          2094 => x"a4",
          2095 => x"08",
          2096 => x"12",
          2097 => x"bf",
          2098 => x"71",
          2099 => x"82",
          2100 => x"88",
          2101 => x"11",
          2102 => x"8c",
          2103 => x"bb",
          2104 => x"05",
          2105 => x"33",
          2106 => x"a4",
          2107 => x"0c",
          2108 => x"82",
          2109 => x"bb",
          2110 => x"05",
          2111 => x"33",
          2112 => x"70",
          2113 => x"51",
          2114 => x"80",
          2115 => x"38",
          2116 => x"08",
          2117 => x"70",
          2118 => x"82",
          2119 => x"fc",
          2120 => x"52",
          2121 => x"08",
          2122 => x"a9",
          2123 => x"a4",
          2124 => x"08",
          2125 => x"08",
          2126 => x"53",
          2127 => x"33",
          2128 => x"51",
          2129 => x"14",
          2130 => x"82",
          2131 => x"f8",
          2132 => x"d7",
          2133 => x"a4",
          2134 => x"08",
          2135 => x"05",
          2136 => x"81",
          2137 => x"bb",
          2138 => x"05",
          2139 => x"a4",
          2140 => x"08",
          2141 => x"08",
          2142 => x"2d",
          2143 => x"08",
          2144 => x"a4",
          2145 => x"0c",
          2146 => x"a4",
          2147 => x"08",
          2148 => x"f2",
          2149 => x"a4",
          2150 => x"08",
          2151 => x"08",
          2152 => x"82",
          2153 => x"88",
          2154 => x"11",
          2155 => x"a4",
          2156 => x"0c",
          2157 => x"a4",
          2158 => x"08",
          2159 => x"81",
          2160 => x"82",
          2161 => x"f0",
          2162 => x"07",
          2163 => x"bb",
          2164 => x"05",
          2165 => x"82",
          2166 => x"f0",
          2167 => x"07",
          2168 => x"bb",
          2169 => x"05",
          2170 => x"a4",
          2171 => x"08",
          2172 => x"a4",
          2173 => x"33",
          2174 => x"ff",
          2175 => x"a4",
          2176 => x"0c",
          2177 => x"bb",
          2178 => x"05",
          2179 => x"08",
          2180 => x"12",
          2181 => x"a4",
          2182 => x"08",
          2183 => x"06",
          2184 => x"a4",
          2185 => x"0c",
          2186 => x"82",
          2187 => x"f8",
          2188 => x"bb",
          2189 => x"3d",
          2190 => x"a4",
          2191 => x"bb",
          2192 => x"82",
          2193 => x"fd",
          2194 => x"bb",
          2195 => x"05",
          2196 => x"a4",
          2197 => x"0c",
          2198 => x"08",
          2199 => x"82",
          2200 => x"f8",
          2201 => x"bb",
          2202 => x"05",
          2203 => x"82",
          2204 => x"bb",
          2205 => x"05",
          2206 => x"a4",
          2207 => x"08",
          2208 => x"38",
          2209 => x"08",
          2210 => x"82",
          2211 => x"90",
          2212 => x"51",
          2213 => x"08",
          2214 => x"71",
          2215 => x"38",
          2216 => x"08",
          2217 => x"82",
          2218 => x"90",
          2219 => x"82",
          2220 => x"fc",
          2221 => x"bb",
          2222 => x"05",
          2223 => x"a4",
          2224 => x"08",
          2225 => x"a4",
          2226 => x"0c",
          2227 => x"08",
          2228 => x"81",
          2229 => x"a4",
          2230 => x"0c",
          2231 => x"08",
          2232 => x"ff",
          2233 => x"a4",
          2234 => x"0c",
          2235 => x"08",
          2236 => x"80",
          2237 => x"38",
          2238 => x"08",
          2239 => x"ff",
          2240 => x"a4",
          2241 => x"0c",
          2242 => x"08",
          2243 => x"ff",
          2244 => x"a4",
          2245 => x"0c",
          2246 => x"08",
          2247 => x"82",
          2248 => x"f8",
          2249 => x"51",
          2250 => x"34",
          2251 => x"82",
          2252 => x"90",
          2253 => x"05",
          2254 => x"08",
          2255 => x"82",
          2256 => x"90",
          2257 => x"05",
          2258 => x"08",
          2259 => x"82",
          2260 => x"90",
          2261 => x"2e",
          2262 => x"bb",
          2263 => x"05",
          2264 => x"33",
          2265 => x"08",
          2266 => x"81",
          2267 => x"a4",
          2268 => x"0c",
          2269 => x"08",
          2270 => x"52",
          2271 => x"34",
          2272 => x"08",
          2273 => x"81",
          2274 => x"a4",
          2275 => x"0c",
          2276 => x"82",
          2277 => x"88",
          2278 => x"82",
          2279 => x"51",
          2280 => x"82",
          2281 => x"04",
          2282 => x"08",
          2283 => x"a4",
          2284 => x"0d",
          2285 => x"08",
          2286 => x"82",
          2287 => x"fc",
          2288 => x"bb",
          2289 => x"05",
          2290 => x"33",
          2291 => x"08",
          2292 => x"81",
          2293 => x"a4",
          2294 => x"0c",
          2295 => x"06",
          2296 => x"80",
          2297 => x"da",
          2298 => x"a4",
          2299 => x"08",
          2300 => x"bb",
          2301 => x"05",
          2302 => x"a4",
          2303 => x"08",
          2304 => x"08",
          2305 => x"31",
          2306 => x"98",
          2307 => x"3d",
          2308 => x"a4",
          2309 => x"bb",
          2310 => x"82",
          2311 => x"fe",
          2312 => x"bb",
          2313 => x"05",
          2314 => x"a4",
          2315 => x"0c",
          2316 => x"08",
          2317 => x"52",
          2318 => x"bb",
          2319 => x"05",
          2320 => x"82",
          2321 => x"8c",
          2322 => x"bb",
          2323 => x"05",
          2324 => x"70",
          2325 => x"bb",
          2326 => x"05",
          2327 => x"82",
          2328 => x"fc",
          2329 => x"81",
          2330 => x"70",
          2331 => x"38",
          2332 => x"82",
          2333 => x"88",
          2334 => x"82",
          2335 => x"51",
          2336 => x"82",
          2337 => x"04",
          2338 => x"08",
          2339 => x"a4",
          2340 => x"0d",
          2341 => x"08",
          2342 => x"82",
          2343 => x"fc",
          2344 => x"bb",
          2345 => x"05",
          2346 => x"a4",
          2347 => x"0c",
          2348 => x"08",
          2349 => x"80",
          2350 => x"38",
          2351 => x"08",
          2352 => x"81",
          2353 => x"a4",
          2354 => x"0c",
          2355 => x"08",
          2356 => x"ff",
          2357 => x"a4",
          2358 => x"0c",
          2359 => x"08",
          2360 => x"80",
          2361 => x"82",
          2362 => x"f8",
          2363 => x"70",
          2364 => x"a4",
          2365 => x"08",
          2366 => x"bb",
          2367 => x"05",
          2368 => x"a4",
          2369 => x"08",
          2370 => x"71",
          2371 => x"a4",
          2372 => x"08",
          2373 => x"bb",
          2374 => x"05",
          2375 => x"39",
          2376 => x"08",
          2377 => x"70",
          2378 => x"0c",
          2379 => x"0d",
          2380 => x"0c",
          2381 => x"a4",
          2382 => x"bb",
          2383 => x"3d",
          2384 => x"a4",
          2385 => x"08",
          2386 => x"f4",
          2387 => x"a4",
          2388 => x"08",
          2389 => x"82",
          2390 => x"8c",
          2391 => x"05",
          2392 => x"08",
          2393 => x"82",
          2394 => x"88",
          2395 => x"33",
          2396 => x"06",
          2397 => x"51",
          2398 => x"84",
          2399 => x"39",
          2400 => x"08",
          2401 => x"52",
          2402 => x"bb",
          2403 => x"05",
          2404 => x"82",
          2405 => x"88",
          2406 => x"81",
          2407 => x"51",
          2408 => x"80",
          2409 => x"a4",
          2410 => x"0c",
          2411 => x"82",
          2412 => x"90",
          2413 => x"05",
          2414 => x"08",
          2415 => x"82",
          2416 => x"90",
          2417 => x"2e",
          2418 => x"81",
          2419 => x"a4",
          2420 => x"08",
          2421 => x"e8",
          2422 => x"a4",
          2423 => x"08",
          2424 => x"53",
          2425 => x"ff",
          2426 => x"a4",
          2427 => x"0c",
          2428 => x"82",
          2429 => x"8c",
          2430 => x"05",
          2431 => x"08",
          2432 => x"82",
          2433 => x"8c",
          2434 => x"33",
          2435 => x"8c",
          2436 => x"82",
          2437 => x"fc",
          2438 => x"39",
          2439 => x"08",
          2440 => x"70",
          2441 => x"a4",
          2442 => x"08",
          2443 => x"71",
          2444 => x"bb",
          2445 => x"05",
          2446 => x"52",
          2447 => x"39",
          2448 => x"bb",
          2449 => x"05",
          2450 => x"a4",
          2451 => x"08",
          2452 => x"0c",
          2453 => x"82",
          2454 => x"04",
          2455 => x"08",
          2456 => x"a4",
          2457 => x"0d",
          2458 => x"08",
          2459 => x"82",
          2460 => x"f8",
          2461 => x"bb",
          2462 => x"05",
          2463 => x"80",
          2464 => x"a4",
          2465 => x"0c",
          2466 => x"82",
          2467 => x"f8",
          2468 => x"71",
          2469 => x"a4",
          2470 => x"08",
          2471 => x"bb",
          2472 => x"05",
          2473 => x"ff",
          2474 => x"70",
          2475 => x"38",
          2476 => x"08",
          2477 => x"ff",
          2478 => x"a4",
          2479 => x"0c",
          2480 => x"08",
          2481 => x"ff",
          2482 => x"ff",
          2483 => x"bb",
          2484 => x"05",
          2485 => x"82",
          2486 => x"f8",
          2487 => x"bb",
          2488 => x"05",
          2489 => x"a4",
          2490 => x"08",
          2491 => x"bb",
          2492 => x"05",
          2493 => x"bb",
          2494 => x"05",
          2495 => x"98",
          2496 => x"0d",
          2497 => x"0c",
          2498 => x"a4",
          2499 => x"bb",
          2500 => x"3d",
          2501 => x"a4",
          2502 => x"08",
          2503 => x"08",
          2504 => x"82",
          2505 => x"90",
          2506 => x"2e",
          2507 => x"82",
          2508 => x"90",
          2509 => x"05",
          2510 => x"08",
          2511 => x"82",
          2512 => x"90",
          2513 => x"05",
          2514 => x"08",
          2515 => x"82",
          2516 => x"90",
          2517 => x"2e",
          2518 => x"bb",
          2519 => x"05",
          2520 => x"82",
          2521 => x"fc",
          2522 => x"52",
          2523 => x"82",
          2524 => x"fc",
          2525 => x"05",
          2526 => x"08",
          2527 => x"ff",
          2528 => x"bb",
          2529 => x"05",
          2530 => x"bb",
          2531 => x"84",
          2532 => x"bb",
          2533 => x"82",
          2534 => x"02",
          2535 => x"0c",
          2536 => x"80",
          2537 => x"a4",
          2538 => x"0c",
          2539 => x"08",
          2540 => x"80",
          2541 => x"82",
          2542 => x"88",
          2543 => x"82",
          2544 => x"88",
          2545 => x"0b",
          2546 => x"08",
          2547 => x"82",
          2548 => x"fc",
          2549 => x"38",
          2550 => x"bb",
          2551 => x"05",
          2552 => x"a4",
          2553 => x"08",
          2554 => x"08",
          2555 => x"82",
          2556 => x"8c",
          2557 => x"25",
          2558 => x"bb",
          2559 => x"05",
          2560 => x"bb",
          2561 => x"05",
          2562 => x"82",
          2563 => x"f0",
          2564 => x"bb",
          2565 => x"05",
          2566 => x"81",
          2567 => x"a4",
          2568 => x"0c",
          2569 => x"08",
          2570 => x"82",
          2571 => x"fc",
          2572 => x"53",
          2573 => x"08",
          2574 => x"52",
          2575 => x"08",
          2576 => x"51",
          2577 => x"82",
          2578 => x"70",
          2579 => x"08",
          2580 => x"54",
          2581 => x"08",
          2582 => x"80",
          2583 => x"82",
          2584 => x"f8",
          2585 => x"82",
          2586 => x"f8",
          2587 => x"bb",
          2588 => x"05",
          2589 => x"bb",
          2590 => x"89",
          2591 => x"bb",
          2592 => x"82",
          2593 => x"02",
          2594 => x"0c",
          2595 => x"80",
          2596 => x"a4",
          2597 => x"0c",
          2598 => x"08",
          2599 => x"80",
          2600 => x"82",
          2601 => x"88",
          2602 => x"82",
          2603 => x"88",
          2604 => x"0b",
          2605 => x"08",
          2606 => x"82",
          2607 => x"8c",
          2608 => x"25",
          2609 => x"bb",
          2610 => x"05",
          2611 => x"bb",
          2612 => x"05",
          2613 => x"82",
          2614 => x"8c",
          2615 => x"82",
          2616 => x"88",
          2617 => x"81",
          2618 => x"bb",
          2619 => x"82",
          2620 => x"f8",
          2621 => x"82",
          2622 => x"fc",
          2623 => x"2e",
          2624 => x"bb",
          2625 => x"05",
          2626 => x"bb",
          2627 => x"05",
          2628 => x"a4",
          2629 => x"08",
          2630 => x"98",
          2631 => x"3d",
          2632 => x"a4",
          2633 => x"bb",
          2634 => x"82",
          2635 => x"fd",
          2636 => x"53",
          2637 => x"08",
          2638 => x"52",
          2639 => x"08",
          2640 => x"51",
          2641 => x"82",
          2642 => x"70",
          2643 => x"0c",
          2644 => x"0d",
          2645 => x"0c",
          2646 => x"a4",
          2647 => x"bb",
          2648 => x"3d",
          2649 => x"82",
          2650 => x"8c",
          2651 => x"82",
          2652 => x"88",
          2653 => x"93",
          2654 => x"98",
          2655 => x"bb",
          2656 => x"85",
          2657 => x"bb",
          2658 => x"82",
          2659 => x"02",
          2660 => x"0c",
          2661 => x"81",
          2662 => x"a4",
          2663 => x"0c",
          2664 => x"bb",
          2665 => x"05",
          2666 => x"a4",
          2667 => x"08",
          2668 => x"08",
          2669 => x"27",
          2670 => x"bb",
          2671 => x"05",
          2672 => x"ae",
          2673 => x"82",
          2674 => x"8c",
          2675 => x"a2",
          2676 => x"a4",
          2677 => x"08",
          2678 => x"a4",
          2679 => x"0c",
          2680 => x"08",
          2681 => x"10",
          2682 => x"08",
          2683 => x"ff",
          2684 => x"bb",
          2685 => x"05",
          2686 => x"80",
          2687 => x"bb",
          2688 => x"05",
          2689 => x"a4",
          2690 => x"08",
          2691 => x"82",
          2692 => x"88",
          2693 => x"bb",
          2694 => x"05",
          2695 => x"bb",
          2696 => x"05",
          2697 => x"a4",
          2698 => x"08",
          2699 => x"08",
          2700 => x"07",
          2701 => x"08",
          2702 => x"82",
          2703 => x"fc",
          2704 => x"2a",
          2705 => x"08",
          2706 => x"82",
          2707 => x"8c",
          2708 => x"2a",
          2709 => x"08",
          2710 => x"ff",
          2711 => x"bb",
          2712 => x"05",
          2713 => x"93",
          2714 => x"a4",
          2715 => x"08",
          2716 => x"a4",
          2717 => x"0c",
          2718 => x"82",
          2719 => x"f8",
          2720 => x"82",
          2721 => x"f4",
          2722 => x"82",
          2723 => x"f4",
          2724 => x"bb",
          2725 => x"3d",
          2726 => x"a4",
          2727 => x"3d",
          2728 => x"08",
          2729 => x"58",
          2730 => x"80",
          2731 => x"39",
          2732 => x"f1",
          2733 => x"bb",
          2734 => x"78",
          2735 => x"33",
          2736 => x"39",
          2737 => x"73",
          2738 => x"81",
          2739 => x"81",
          2740 => x"39",
          2741 => x"90",
          2742 => x"98",
          2743 => x"52",
          2744 => x"3f",
          2745 => x"08",
          2746 => x"75",
          2747 => x"c5",
          2748 => x"98",
          2749 => x"84",
          2750 => x"73",
          2751 => x"b0",
          2752 => x"70",
          2753 => x"58",
          2754 => x"27",
          2755 => x"54",
          2756 => x"98",
          2757 => x"0d",
          2758 => x"0d",
          2759 => x"93",
          2760 => x"38",
          2761 => x"82",
          2762 => x"52",
          2763 => x"82",
          2764 => x"81",
          2765 => x"9f",
          2766 => x"f9",
          2767 => x"9c",
          2768 => x"39",
          2769 => x"51",
          2770 => x"82",
          2771 => x"80",
          2772 => x"9f",
          2773 => x"dd",
          2774 => x"e4",
          2775 => x"39",
          2776 => x"51",
          2777 => x"82",
          2778 => x"80",
          2779 => x"a0",
          2780 => x"c1",
          2781 => x"bc",
          2782 => x"82",
          2783 => x"b5",
          2784 => x"ec",
          2785 => x"82",
          2786 => x"a9",
          2787 => x"ac",
          2788 => x"82",
          2789 => x"9d",
          2790 => x"e0",
          2791 => x"82",
          2792 => x"91",
          2793 => x"90",
          2794 => x"82",
          2795 => x"85",
          2796 => x"b4",
          2797 => x"3f",
          2798 => x"04",
          2799 => x"77",
          2800 => x"74",
          2801 => x"8a",
          2802 => x"75",
          2803 => x"51",
          2804 => x"e8",
          2805 => x"fa",
          2806 => x"bb",
          2807 => x"75",
          2808 => x"3f",
          2809 => x"08",
          2810 => x"75",
          2811 => x"c4",
          2812 => x"e5",
          2813 => x"0d",
          2814 => x"0d",
          2815 => x"05",
          2816 => x"33",
          2817 => x"68",
          2818 => x"7a",
          2819 => x"51",
          2820 => x"78",
          2821 => x"ff",
          2822 => x"81",
          2823 => x"07",
          2824 => x"06",
          2825 => x"56",
          2826 => x"38",
          2827 => x"52",
          2828 => x"52",
          2829 => x"cf",
          2830 => x"98",
          2831 => x"bb",
          2832 => x"38",
          2833 => x"08",
          2834 => x"88",
          2835 => x"98",
          2836 => x"3d",
          2837 => x"84",
          2838 => x"52",
          2839 => x"88",
          2840 => x"bb",
          2841 => x"82",
          2842 => x"90",
          2843 => x"74",
          2844 => x"38",
          2845 => x"19",
          2846 => x"39",
          2847 => x"05",
          2848 => x"f4",
          2849 => x"70",
          2850 => x"25",
          2851 => x"9f",
          2852 => x"51",
          2853 => x"74",
          2854 => x"38",
          2855 => x"53",
          2856 => x"88",
          2857 => x"51",
          2858 => x"76",
          2859 => x"bb",
          2860 => x"3d",
          2861 => x"3d",
          2862 => x"84",
          2863 => x"33",
          2864 => x"58",
          2865 => x"52",
          2866 => x"ad",
          2867 => x"98",
          2868 => x"76",
          2869 => x"38",
          2870 => x"9a",
          2871 => x"62",
          2872 => x"60",
          2873 => x"98",
          2874 => x"7e",
          2875 => x"82",
          2876 => x"58",
          2877 => x"04",
          2878 => x"98",
          2879 => x"0d",
          2880 => x"0d",
          2881 => x"02",
          2882 => x"cf",
          2883 => x"73",
          2884 => x"5f",
          2885 => x"5e",
          2886 => x"82",
          2887 => x"ff",
          2888 => x"82",
          2889 => x"e0",
          2890 => x"55",
          2891 => x"80",
          2892 => x"90",
          2893 => x"7b",
          2894 => x"38",
          2895 => x"74",
          2896 => x"7a",
          2897 => x"72",
          2898 => x"a2",
          2899 => x"b9",
          2900 => x"39",
          2901 => x"51",
          2902 => x"82",
          2903 => x"c1",
          2904 => x"53",
          2905 => x"8e",
          2906 => x"52",
          2907 => x"51",
          2908 => x"3f",
          2909 => x"a3",
          2910 => x"8a",
          2911 => x"55",
          2912 => x"18",
          2913 => x"27",
          2914 => x"33",
          2915 => x"90",
          2916 => x"c5",
          2917 => x"82",
          2918 => x"df",
          2919 => x"15",
          2920 => x"ec",
          2921 => x"51",
          2922 => x"fe",
          2923 => x"a3",
          2924 => x"d2",
          2925 => x"74",
          2926 => x"c6",
          2927 => x"70",
          2928 => x"80",
          2929 => x"27",
          2930 => x"56",
          2931 => x"74",
          2932 => x"81",
          2933 => x"06",
          2934 => x"06",
          2935 => x"80",
          2936 => x"73",
          2937 => x"8a",
          2938 => x"ec",
          2939 => x"51",
          2940 => x"d2",
          2941 => x"a0",
          2942 => x"3f",
          2943 => x"ff",
          2944 => x"a3",
          2945 => x"fe",
          2946 => x"79",
          2947 => x"a0",
          2948 => x"bb",
          2949 => x"2b",
          2950 => x"51",
          2951 => x"2e",
          2952 => x"aa",
          2953 => x"3f",
          2954 => x"08",
          2955 => x"98",
          2956 => x"32",
          2957 => x"9b",
          2958 => x"70",
          2959 => x"75",
          2960 => x"58",
          2961 => x"51",
          2962 => x"24",
          2963 => x"9b",
          2964 => x"06",
          2965 => x"53",
          2966 => x"1e",
          2967 => x"26",
          2968 => x"ff",
          2969 => x"bb",
          2970 => x"3d",
          2971 => x"3d",
          2972 => x"05",
          2973 => x"a4",
          2974 => x"ac",
          2975 => x"b6",
          2976 => x"b9",
          2977 => x"a9",
          2978 => x"a3",
          2979 => x"a3",
          2980 => x"b9",
          2981 => x"82",
          2982 => x"ff",
          2983 => x"74",
          2984 => x"38",
          2985 => x"86",
          2986 => x"fe",
          2987 => x"c0",
          2988 => x"53",
          2989 => x"81",
          2990 => x"3f",
          2991 => x"51",
          2992 => x"80",
          2993 => x"3f",
          2994 => x"70",
          2995 => x"52",
          2996 => x"92",
          2997 => x"9c",
          2998 => x"a4",
          2999 => x"a9",
          3000 => x"9c",
          3001 => x"82",
          3002 => x"06",
          3003 => x"80",
          3004 => x"81",
          3005 => x"3f",
          3006 => x"51",
          3007 => x"80",
          3008 => x"3f",
          3009 => x"70",
          3010 => x"52",
          3011 => x"92",
          3012 => x"9b",
          3013 => x"a4",
          3014 => x"ed",
          3015 => x"9b",
          3016 => x"84",
          3017 => x"06",
          3018 => x"80",
          3019 => x"81",
          3020 => x"3f",
          3021 => x"51",
          3022 => x"80",
          3023 => x"3f",
          3024 => x"70",
          3025 => x"52",
          3026 => x"92",
          3027 => x"9b",
          3028 => x"a4",
          3029 => x"b1",
          3030 => x"9b",
          3031 => x"86",
          3032 => x"06",
          3033 => x"80",
          3034 => x"81",
          3035 => x"3f",
          3036 => x"51",
          3037 => x"80",
          3038 => x"3f",
          3039 => x"70",
          3040 => x"52",
          3041 => x"92",
          3042 => x"9a",
          3043 => x"a4",
          3044 => x"f5",
          3045 => x"9a",
          3046 => x"88",
          3047 => x"06",
          3048 => x"80",
          3049 => x"81",
          3050 => x"3f",
          3051 => x"51",
          3052 => x"80",
          3053 => x"3f",
          3054 => x"84",
          3055 => x"fb",
          3056 => x"02",
          3057 => x"05",
          3058 => x"56",
          3059 => x"75",
          3060 => x"3f",
          3061 => x"b6",
          3062 => x"73",
          3063 => x"53",
          3064 => x"52",
          3065 => x"51",
          3066 => x"3f",
          3067 => x"08",
          3068 => x"bb",
          3069 => x"80",
          3070 => x"31",
          3071 => x"73",
          3072 => x"b6",
          3073 => x"0b",
          3074 => x"33",
          3075 => x"2e",
          3076 => x"af",
          3077 => x"98",
          3078 => x"75",
          3079 => x"cd",
          3080 => x"98",
          3081 => x"8b",
          3082 => x"98",
          3083 => x"d6",
          3084 => x"82",
          3085 => x"81",
          3086 => x"82",
          3087 => x"82",
          3088 => x"0b",
          3089 => x"94",
          3090 => x"82",
          3091 => x"06",
          3092 => x"a5",
          3093 => x"52",
          3094 => x"95",
          3095 => x"82",
          3096 => x"87",
          3097 => x"cd",
          3098 => x"70",
          3099 => x"94",
          3100 => x"81",
          3101 => x"80",
          3102 => x"82",
          3103 => x"81",
          3104 => x"79",
          3105 => x"81",
          3106 => x"97",
          3107 => x"53",
          3108 => x"52",
          3109 => x"f0",
          3110 => x"79",
          3111 => x"c4",
          3112 => x"82",
          3113 => x"98",
          3114 => x"88",
          3115 => x"ec",
          3116 => x"39",
          3117 => x"5e",
          3118 => x"51",
          3119 => x"97",
          3120 => x"5b",
          3121 => x"7a",
          3122 => x"3f",
          3123 => x"84",
          3124 => x"ca",
          3125 => x"98",
          3126 => x"70",
          3127 => x"5a",
          3128 => x"2e",
          3129 => x"79",
          3130 => x"80",
          3131 => x"ab",
          3132 => x"38",
          3133 => x"a4",
          3134 => x"2e",
          3135 => x"79",
          3136 => x"38",
          3137 => x"ff",
          3138 => x"ed",
          3139 => x"2e",
          3140 => x"79",
          3141 => x"ad",
          3142 => x"39",
          3143 => x"84",
          3144 => x"bd",
          3145 => x"79",
          3146 => x"a6",
          3147 => x"2e",
          3148 => x"8e",
          3149 => x"bf",
          3150 => x"38",
          3151 => x"2e",
          3152 => x"8e",
          3153 => x"80",
          3154 => x"90",
          3155 => x"d5",
          3156 => x"79",
          3157 => x"8c",
          3158 => x"80",
          3159 => x"38",
          3160 => x"2e",
          3161 => x"79",
          3162 => x"8b",
          3163 => x"89",
          3164 => x"d1",
          3165 => x"38",
          3166 => x"2e",
          3167 => x"8d",
          3168 => x"81",
          3169 => x"d1",
          3170 => x"82",
          3171 => x"79",
          3172 => x"8c",
          3173 => x"80",
          3174 => x"80",
          3175 => x"39",
          3176 => x"2e",
          3177 => x"79",
          3178 => x"8d",
          3179 => x"c9",
          3180 => x"ff",
          3181 => x"ff",
          3182 => x"d1",
          3183 => x"bb",
          3184 => x"38",
          3185 => x"51",
          3186 => x"b5",
          3187 => x"11",
          3188 => x"05",
          3189 => x"3f",
          3190 => x"08",
          3191 => x"38",
          3192 => x"83",
          3193 => x"02",
          3194 => x"33",
          3195 => x"d3",
          3196 => x"80",
          3197 => x"82",
          3198 => x"81",
          3199 => x"79",
          3200 => x"a6",
          3201 => x"fe",
          3202 => x"fd",
          3203 => x"a6",
          3204 => x"e7",
          3205 => x"ff",
          3206 => x"ff",
          3207 => x"d1",
          3208 => x"bb",
          3209 => x"2e",
          3210 => x"80",
          3211 => x"02",
          3212 => x"33",
          3213 => x"f7",
          3214 => x"98",
          3215 => x"a6",
          3216 => x"8e",
          3217 => x"ff",
          3218 => x"ff",
          3219 => x"d0",
          3220 => x"bb",
          3221 => x"2e",
          3222 => x"89",
          3223 => x"38",
          3224 => x"fc",
          3225 => x"84",
          3226 => x"c9",
          3227 => x"98",
          3228 => x"82",
          3229 => x"44",
          3230 => x"a6",
          3231 => x"51",
          3232 => x"3f",
          3233 => x"05",
          3234 => x"52",
          3235 => x"29",
          3236 => x"05",
          3237 => x"8e",
          3238 => x"98",
          3239 => x"38",
          3240 => x"51",
          3241 => x"81",
          3242 => x"39",
          3243 => x"84",
          3244 => x"b1",
          3245 => x"98",
          3246 => x"ff",
          3247 => x"5c",
          3248 => x"81",
          3249 => x"98",
          3250 => x"51",
          3251 => x"80",
          3252 => x"3d",
          3253 => x"51",
          3254 => x"82",
          3255 => x"b6",
          3256 => x"05",
          3257 => x"a1",
          3258 => x"98",
          3259 => x"ff",
          3260 => x"5b",
          3261 => x"82",
          3262 => x"b6",
          3263 => x"05",
          3264 => x"85",
          3265 => x"e8",
          3266 => x"bc",
          3267 => x"c8",
          3268 => x"80",
          3269 => x"98",
          3270 => x"06",
          3271 => x"7a",
          3272 => x"f3",
          3273 => x"bb",
          3274 => x"2e",
          3275 => x"82",
          3276 => x"51",
          3277 => x"fa",
          3278 => x"3d",
          3279 => x"53",
          3280 => x"51",
          3281 => x"82",
          3282 => x"80",
          3283 => x"38",
          3284 => x"fc",
          3285 => x"84",
          3286 => x"d9",
          3287 => x"98",
          3288 => x"fa",
          3289 => x"3d",
          3290 => x"53",
          3291 => x"51",
          3292 => x"82",
          3293 => x"86",
          3294 => x"98",
          3295 => x"a6",
          3296 => x"82",
          3297 => x"5d",
          3298 => x"27",
          3299 => x"62",
          3300 => x"70",
          3301 => x"0c",
          3302 => x"f5",
          3303 => x"39",
          3304 => x"80",
          3305 => x"84",
          3306 => x"89",
          3307 => x"98",
          3308 => x"fa",
          3309 => x"3d",
          3310 => x"53",
          3311 => x"51",
          3312 => x"82",
          3313 => x"80",
          3314 => x"38",
          3315 => x"f8",
          3316 => x"84",
          3317 => x"dd",
          3318 => x"98",
          3319 => x"f9",
          3320 => x"a6",
          3321 => x"9e",
          3322 => x"7a",
          3323 => x"88",
          3324 => x"7a",
          3325 => x"5c",
          3326 => x"62",
          3327 => x"eb",
          3328 => x"ff",
          3329 => x"ff",
          3330 => x"cd",
          3331 => x"bb",
          3332 => x"2e",
          3333 => x"b5",
          3334 => x"11",
          3335 => x"05",
          3336 => x"3f",
          3337 => x"08",
          3338 => x"8c",
          3339 => x"fe",
          3340 => x"ff",
          3341 => x"cc",
          3342 => x"bb",
          3343 => x"2e",
          3344 => x"82",
          3345 => x"d2",
          3346 => x"5b",
          3347 => x"a8",
          3348 => x"33",
          3349 => x"5b",
          3350 => x"2e",
          3351 => x"55",
          3352 => x"33",
          3353 => x"82",
          3354 => x"ff",
          3355 => x"81",
          3356 => x"05",
          3357 => x"39",
          3358 => x"51",
          3359 => x"b5",
          3360 => x"11",
          3361 => x"05",
          3362 => x"3f",
          3363 => x"08",
          3364 => x"82",
          3365 => x"5a",
          3366 => x"89",
          3367 => x"bc",
          3368 => x"cd",
          3369 => x"85",
          3370 => x"80",
          3371 => x"82",
          3372 => x"45",
          3373 => x"ba",
          3374 => x"79",
          3375 => x"38",
          3376 => x"08",
          3377 => x"82",
          3378 => x"5a",
          3379 => x"88",
          3380 => x"d4",
          3381 => x"39",
          3382 => x"33",
          3383 => x"2e",
          3384 => x"b9",
          3385 => x"89",
          3386 => x"ec",
          3387 => x"05",
          3388 => x"fe",
          3389 => x"ff",
          3390 => x"cb",
          3391 => x"bb",
          3392 => x"de",
          3393 => x"84",
          3394 => x"80",
          3395 => x"82",
          3396 => x"44",
          3397 => x"82",
          3398 => x"5a",
          3399 => x"88",
          3400 => x"c8",
          3401 => x"39",
          3402 => x"33",
          3403 => x"2e",
          3404 => x"b9",
          3405 => x"aa",
          3406 => x"87",
          3407 => x"80",
          3408 => x"82",
          3409 => x"44",
          3410 => x"ba",
          3411 => x"79",
          3412 => x"38",
          3413 => x"08",
          3414 => x"82",
          3415 => x"88",
          3416 => x"3d",
          3417 => x"53",
          3418 => x"51",
          3419 => x"82",
          3420 => x"80",
          3421 => x"80",
          3422 => x"7b",
          3423 => x"38",
          3424 => x"90",
          3425 => x"70",
          3426 => x"2a",
          3427 => x"51",
          3428 => x"79",
          3429 => x"38",
          3430 => x"83",
          3431 => x"82",
          3432 => x"cf",
          3433 => x"55",
          3434 => x"53",
          3435 => x"51",
          3436 => x"82",
          3437 => x"87",
          3438 => x"3d",
          3439 => x"53",
          3440 => x"51",
          3441 => x"82",
          3442 => x"80",
          3443 => x"38",
          3444 => x"fc",
          3445 => x"84",
          3446 => x"d9",
          3447 => x"98",
          3448 => x"a4",
          3449 => x"02",
          3450 => x"33",
          3451 => x"81",
          3452 => x"3d",
          3453 => x"53",
          3454 => x"51",
          3455 => x"82",
          3456 => x"e1",
          3457 => x"39",
          3458 => x"54",
          3459 => x"d0",
          3460 => x"c5",
          3461 => x"52",
          3462 => x"e3",
          3463 => x"7a",
          3464 => x"ae",
          3465 => x"38",
          3466 => x"9f",
          3467 => x"fe",
          3468 => x"ff",
          3469 => x"c8",
          3470 => x"bb",
          3471 => x"2e",
          3472 => x"5a",
          3473 => x"05",
          3474 => x"64",
          3475 => x"ff",
          3476 => x"a7",
          3477 => x"ae",
          3478 => x"39",
          3479 => x"f4",
          3480 => x"84",
          3481 => x"c6",
          3482 => x"98",
          3483 => x"f4",
          3484 => x"3d",
          3485 => x"53",
          3486 => x"51",
          3487 => x"82",
          3488 => x"80",
          3489 => x"61",
          3490 => x"c2",
          3491 => x"70",
          3492 => x"23",
          3493 => x"3d",
          3494 => x"53",
          3495 => x"51",
          3496 => x"82",
          3497 => x"df",
          3498 => x"39",
          3499 => x"54",
          3500 => x"e4",
          3501 => x"a1",
          3502 => x"52",
          3503 => x"bf",
          3504 => x"7a",
          3505 => x"ae",
          3506 => x"38",
          3507 => x"87",
          3508 => x"05",
          3509 => x"b5",
          3510 => x"11",
          3511 => x"05",
          3512 => x"3f",
          3513 => x"08",
          3514 => x"38",
          3515 => x"80",
          3516 => x"7a",
          3517 => x"5c",
          3518 => x"ff",
          3519 => x"a7",
          3520 => x"82",
          3521 => x"39",
          3522 => x"f4",
          3523 => x"84",
          3524 => x"9a",
          3525 => x"98",
          3526 => x"f3",
          3527 => x"3d",
          3528 => x"53",
          3529 => x"51",
          3530 => x"82",
          3531 => x"80",
          3532 => x"61",
          3533 => x"5a",
          3534 => x"42",
          3535 => x"f0",
          3536 => x"84",
          3537 => x"e6",
          3538 => x"98",
          3539 => x"f2",
          3540 => x"70",
          3541 => x"82",
          3542 => x"ff",
          3543 => x"80",
          3544 => x"51",
          3545 => x"7a",
          3546 => x"5a",
          3547 => x"f2",
          3548 => x"7a",
          3549 => x"b5",
          3550 => x"11",
          3551 => x"05",
          3552 => x"3f",
          3553 => x"08",
          3554 => x"38",
          3555 => x"0c",
          3556 => x"05",
          3557 => x"39",
          3558 => x"51",
          3559 => x"ff",
          3560 => x"a7",
          3561 => x"de",
          3562 => x"98",
          3563 => x"88",
          3564 => x"94",
          3565 => x"3f",
          3566 => x"e0",
          3567 => x"39",
          3568 => x"51",
          3569 => x"84",
          3570 => x"87",
          3571 => x"0c",
          3572 => x"0b",
          3573 => x"94",
          3574 => x"39",
          3575 => x"51",
          3576 => x"8c",
          3577 => x"87",
          3578 => x"0c",
          3579 => x"0b",
          3580 => x"94",
          3581 => x"39",
          3582 => x"80",
          3583 => x"84",
          3584 => x"b1",
          3585 => x"98",
          3586 => x"f1",
          3587 => x"52",
          3588 => x"51",
          3589 => x"3f",
          3590 => x"04",
          3591 => x"80",
          3592 => x"84",
          3593 => x"8d",
          3594 => x"98",
          3595 => x"f1",
          3596 => x"52",
          3597 => x"51",
          3598 => x"3f",
          3599 => x"2d",
          3600 => x"08",
          3601 => x"f0",
          3602 => x"98",
          3603 => x"a9",
          3604 => x"a3",
          3605 => x"e0",
          3606 => x"a8",
          3607 => x"3f",
          3608 => x"3f",
          3609 => x"82",
          3610 => x"ca",
          3611 => x"5a",
          3612 => x"91",
          3613 => x"c0",
          3614 => x"7a",
          3615 => x"80",
          3616 => x"38",
          3617 => x"5a",
          3618 => x"81",
          3619 => x"3d",
          3620 => x"51",
          3621 => x"82",
          3622 => x"5c",
          3623 => x"82",
          3624 => x"7c",
          3625 => x"38",
          3626 => x"8c",
          3627 => x"39",
          3628 => x"b0",
          3629 => x"39",
          3630 => x"56",
          3631 => x"a9",
          3632 => x"53",
          3633 => x"52",
          3634 => x"b0",
          3635 => x"a4",
          3636 => x"39",
          3637 => x"52",
          3638 => x"b0",
          3639 => x"a4",
          3640 => x"39",
          3641 => x"a9",
          3642 => x"53",
          3643 => x"52",
          3644 => x"b0",
          3645 => x"a4",
          3646 => x"39",
          3647 => x"53",
          3648 => x"52",
          3649 => x"b0",
          3650 => x"a4",
          3651 => x"d2",
          3652 => x"b9",
          3653 => x"bb",
          3654 => x"56",
          3655 => x"54",
          3656 => x"53",
          3657 => x"52",
          3658 => x"b0",
          3659 => x"86",
          3660 => x"98",
          3661 => x"98",
          3662 => x"30",
          3663 => x"80",
          3664 => x"5c",
          3665 => x"7c",
          3666 => x"38",
          3667 => x"7b",
          3668 => x"80",
          3669 => x"81",
          3670 => x"ff",
          3671 => x"7c",
          3672 => x"7e",
          3673 => x"81",
          3674 => x"79",
          3675 => x"ff",
          3676 => x"06",
          3677 => x"82",
          3678 => x"c8",
          3679 => x"b8",
          3680 => x"0d",
          3681 => x"bb",
          3682 => x"c0",
          3683 => x"08",
          3684 => x"84",
          3685 => x"51",
          3686 => x"82",
          3687 => x"90",
          3688 => x"55",
          3689 => x"80",
          3690 => x"de",
          3691 => x"82",
          3692 => x"07",
          3693 => x"c0",
          3694 => x"08",
          3695 => x"84",
          3696 => x"51",
          3697 => x"82",
          3698 => x"90",
          3699 => x"55",
          3700 => x"80",
          3701 => x"de",
          3702 => x"82",
          3703 => x"07",
          3704 => x"80",
          3705 => x"c0",
          3706 => x"8c",
          3707 => x"87",
          3708 => x"0c",
          3709 => x"5a",
          3710 => x"5b",
          3711 => x"05",
          3712 => x"80",
          3713 => x"e8",
          3714 => x"70",
          3715 => x"70",
          3716 => x"d2",
          3717 => x"89",
          3718 => x"c1",
          3719 => x"94",
          3720 => x"3f",
          3721 => x"51",
          3722 => x"80",
          3723 => x"92",
          3724 => x"51",
          3725 => x"ec",
          3726 => x"04",
          3727 => x"80",
          3728 => x"71",
          3729 => x"87",
          3730 => x"bb",
          3731 => x"ff",
          3732 => x"ff",
          3733 => x"72",
          3734 => x"38",
          3735 => x"98",
          3736 => x"0d",
          3737 => x"0d",
          3738 => x"54",
          3739 => x"52",
          3740 => x"2e",
          3741 => x"72",
          3742 => x"a0",
          3743 => x"06",
          3744 => x"13",
          3745 => x"72",
          3746 => x"a2",
          3747 => x"06",
          3748 => x"13",
          3749 => x"72",
          3750 => x"2e",
          3751 => x"9f",
          3752 => x"81",
          3753 => x"72",
          3754 => x"70",
          3755 => x"38",
          3756 => x"80",
          3757 => x"73",
          3758 => x"39",
          3759 => x"80",
          3760 => x"54",
          3761 => x"83",
          3762 => x"70",
          3763 => x"38",
          3764 => x"80",
          3765 => x"54",
          3766 => x"09",
          3767 => x"38",
          3768 => x"a2",
          3769 => x"70",
          3770 => x"07",
          3771 => x"70",
          3772 => x"38",
          3773 => x"81",
          3774 => x"71",
          3775 => x"51",
          3776 => x"98",
          3777 => x"0d",
          3778 => x"0d",
          3779 => x"08",
          3780 => x"38",
          3781 => x"05",
          3782 => x"ff",
          3783 => x"82",
          3784 => x"85",
          3785 => x"83",
          3786 => x"72",
          3787 => x"0c",
          3788 => x"04",
          3789 => x"76",
          3790 => x"ff",
          3791 => x"81",
          3792 => x"26",
          3793 => x"83",
          3794 => x"05",
          3795 => x"70",
          3796 => x"8a",
          3797 => x"33",
          3798 => x"70",
          3799 => x"fe",
          3800 => x"33",
          3801 => x"70",
          3802 => x"f2",
          3803 => x"33",
          3804 => x"70",
          3805 => x"e6",
          3806 => x"22",
          3807 => x"74",
          3808 => x"80",
          3809 => x"13",
          3810 => x"52",
          3811 => x"26",
          3812 => x"81",
          3813 => x"98",
          3814 => x"22",
          3815 => x"bc",
          3816 => x"33",
          3817 => x"b8",
          3818 => x"33",
          3819 => x"b4",
          3820 => x"33",
          3821 => x"b0",
          3822 => x"33",
          3823 => x"ac",
          3824 => x"33",
          3825 => x"a8",
          3826 => x"c0",
          3827 => x"73",
          3828 => x"a0",
          3829 => x"87",
          3830 => x"0c",
          3831 => x"82",
          3832 => x"86",
          3833 => x"f3",
          3834 => x"5b",
          3835 => x"9c",
          3836 => x"0c",
          3837 => x"bc",
          3838 => x"7b",
          3839 => x"98",
          3840 => x"79",
          3841 => x"87",
          3842 => x"08",
          3843 => x"1c",
          3844 => x"98",
          3845 => x"79",
          3846 => x"87",
          3847 => x"08",
          3848 => x"1c",
          3849 => x"98",
          3850 => x"79",
          3851 => x"87",
          3852 => x"08",
          3853 => x"1c",
          3854 => x"98",
          3855 => x"79",
          3856 => x"80",
          3857 => x"83",
          3858 => x"59",
          3859 => x"ff",
          3860 => x"1b",
          3861 => x"1b",
          3862 => x"1b",
          3863 => x"1b",
          3864 => x"1b",
          3865 => x"83",
          3866 => x"52",
          3867 => x"51",
          3868 => x"3f",
          3869 => x"04",
          3870 => x"02",
          3871 => x"82",
          3872 => x"70",
          3873 => x"58",
          3874 => x"c0",
          3875 => x"75",
          3876 => x"38",
          3877 => x"94",
          3878 => x"70",
          3879 => x"81",
          3880 => x"52",
          3881 => x"8c",
          3882 => x"2a",
          3883 => x"51",
          3884 => x"38",
          3885 => x"70",
          3886 => x"51",
          3887 => x"8d",
          3888 => x"2a",
          3889 => x"51",
          3890 => x"be",
          3891 => x"ff",
          3892 => x"c0",
          3893 => x"70",
          3894 => x"38",
          3895 => x"90",
          3896 => x"0c",
          3897 => x"98",
          3898 => x"0d",
          3899 => x"0d",
          3900 => x"33",
          3901 => x"9f",
          3902 => x"52",
          3903 => x"b8",
          3904 => x"0d",
          3905 => x"0d",
          3906 => x"33",
          3907 => x"2e",
          3908 => x"87",
          3909 => x"8d",
          3910 => x"82",
          3911 => x"70",
          3912 => x"58",
          3913 => x"94",
          3914 => x"80",
          3915 => x"87",
          3916 => x"53",
          3917 => x"96",
          3918 => x"06",
          3919 => x"72",
          3920 => x"38",
          3921 => x"70",
          3922 => x"53",
          3923 => x"74",
          3924 => x"81",
          3925 => x"72",
          3926 => x"38",
          3927 => x"70",
          3928 => x"53",
          3929 => x"38",
          3930 => x"06",
          3931 => x"94",
          3932 => x"80",
          3933 => x"87",
          3934 => x"54",
          3935 => x"80",
          3936 => x"98",
          3937 => x"0d",
          3938 => x"0d",
          3939 => x"74",
          3940 => x"ff",
          3941 => x"57",
          3942 => x"80",
          3943 => x"81",
          3944 => x"15",
          3945 => x"33",
          3946 => x"06",
          3947 => x"58",
          3948 => x"84",
          3949 => x"2e",
          3950 => x"c0",
          3951 => x"70",
          3952 => x"2a",
          3953 => x"53",
          3954 => x"80",
          3955 => x"71",
          3956 => x"81",
          3957 => x"70",
          3958 => x"81",
          3959 => x"06",
          3960 => x"80",
          3961 => x"71",
          3962 => x"81",
          3963 => x"70",
          3964 => x"74",
          3965 => x"51",
          3966 => x"80",
          3967 => x"2e",
          3968 => x"c0",
          3969 => x"77",
          3970 => x"17",
          3971 => x"81",
          3972 => x"53",
          3973 => x"86",
          3974 => x"bb",
          3975 => x"3d",
          3976 => x"3d",
          3977 => x"b8",
          3978 => x"ff",
          3979 => x"87",
          3980 => x"51",
          3981 => x"86",
          3982 => x"94",
          3983 => x"08",
          3984 => x"70",
          3985 => x"51",
          3986 => x"2e",
          3987 => x"81",
          3988 => x"87",
          3989 => x"52",
          3990 => x"86",
          3991 => x"94",
          3992 => x"08",
          3993 => x"06",
          3994 => x"0c",
          3995 => x"0d",
          3996 => x"3f",
          3997 => x"08",
          3998 => x"82",
          3999 => x"04",
          4000 => x"82",
          4001 => x"70",
          4002 => x"52",
          4003 => x"94",
          4004 => x"80",
          4005 => x"87",
          4006 => x"52",
          4007 => x"82",
          4008 => x"06",
          4009 => x"ff",
          4010 => x"2e",
          4011 => x"81",
          4012 => x"87",
          4013 => x"52",
          4014 => x"86",
          4015 => x"94",
          4016 => x"08",
          4017 => x"70",
          4018 => x"53",
          4019 => x"bb",
          4020 => x"3d",
          4021 => x"3d",
          4022 => x"9e",
          4023 => x"9c",
          4024 => x"51",
          4025 => x"2e",
          4026 => x"87",
          4027 => x"08",
          4028 => x"0c",
          4029 => x"a8",
          4030 => x"c0",
          4031 => x"9e",
          4032 => x"b9",
          4033 => x"c0",
          4034 => x"82",
          4035 => x"87",
          4036 => x"08",
          4037 => x"0c",
          4038 => x"a0",
          4039 => x"d0",
          4040 => x"9e",
          4041 => x"b9",
          4042 => x"c0",
          4043 => x"82",
          4044 => x"87",
          4045 => x"08",
          4046 => x"0c",
          4047 => x"b8",
          4048 => x"e0",
          4049 => x"9e",
          4050 => x"b9",
          4051 => x"c0",
          4052 => x"82",
          4053 => x"87",
          4054 => x"08",
          4055 => x"0c",
          4056 => x"80",
          4057 => x"82",
          4058 => x"87",
          4059 => x"08",
          4060 => x"0c",
          4061 => x"88",
          4062 => x"f8",
          4063 => x"9e",
          4064 => x"b9",
          4065 => x"0b",
          4066 => x"34",
          4067 => x"c0",
          4068 => x"70",
          4069 => x"06",
          4070 => x"70",
          4071 => x"38",
          4072 => x"82",
          4073 => x"80",
          4074 => x"9e",
          4075 => x"88",
          4076 => x"51",
          4077 => x"80",
          4078 => x"81",
          4079 => x"ba",
          4080 => x"0b",
          4081 => x"90",
          4082 => x"80",
          4083 => x"52",
          4084 => x"2e",
          4085 => x"52",
          4086 => x"83",
          4087 => x"87",
          4088 => x"08",
          4089 => x"80",
          4090 => x"52",
          4091 => x"83",
          4092 => x"71",
          4093 => x"34",
          4094 => x"c0",
          4095 => x"70",
          4096 => x"06",
          4097 => x"70",
          4098 => x"38",
          4099 => x"82",
          4100 => x"80",
          4101 => x"9e",
          4102 => x"90",
          4103 => x"51",
          4104 => x"80",
          4105 => x"81",
          4106 => x"ba",
          4107 => x"0b",
          4108 => x"90",
          4109 => x"80",
          4110 => x"52",
          4111 => x"2e",
          4112 => x"52",
          4113 => x"87",
          4114 => x"87",
          4115 => x"08",
          4116 => x"80",
          4117 => x"52",
          4118 => x"83",
          4119 => x"71",
          4120 => x"34",
          4121 => x"c0",
          4122 => x"70",
          4123 => x"06",
          4124 => x"70",
          4125 => x"38",
          4126 => x"82",
          4127 => x"80",
          4128 => x"9e",
          4129 => x"80",
          4130 => x"51",
          4131 => x"80",
          4132 => x"81",
          4133 => x"ba",
          4134 => x"0b",
          4135 => x"90",
          4136 => x"80",
          4137 => x"52",
          4138 => x"83",
          4139 => x"71",
          4140 => x"34",
          4141 => x"90",
          4142 => x"80",
          4143 => x"2a",
          4144 => x"70",
          4145 => x"34",
          4146 => x"c0",
          4147 => x"70",
          4148 => x"51",
          4149 => x"80",
          4150 => x"81",
          4151 => x"ba",
          4152 => x"c0",
          4153 => x"70",
          4154 => x"70",
          4155 => x"51",
          4156 => x"ba",
          4157 => x"0b",
          4158 => x"90",
          4159 => x"06",
          4160 => x"70",
          4161 => x"38",
          4162 => x"82",
          4163 => x"87",
          4164 => x"08",
          4165 => x"51",
          4166 => x"ba",
          4167 => x"3d",
          4168 => x"3d",
          4169 => x"d0",
          4170 => x"da",
          4171 => x"80",
          4172 => x"80",
          4173 => x"82",
          4174 => x"ff",
          4175 => x"82",
          4176 => x"ff",
          4177 => x"82",
          4178 => x"54",
          4179 => x"94",
          4180 => x"dc",
          4181 => x"e0",
          4182 => x"52",
          4183 => x"51",
          4184 => x"3f",
          4185 => x"33",
          4186 => x"2e",
          4187 => x"b9",
          4188 => x"b9",
          4189 => x"54",
          4190 => x"ac",
          4191 => x"d9",
          4192 => x"84",
          4193 => x"80",
          4194 => x"82",
          4195 => x"82",
          4196 => x"11",
          4197 => x"ab",
          4198 => x"90",
          4199 => x"ba",
          4200 => x"73",
          4201 => x"38",
          4202 => x"08",
          4203 => x"08",
          4204 => x"82",
          4205 => x"ff",
          4206 => x"82",
          4207 => x"54",
          4208 => x"94",
          4209 => x"cc",
          4210 => x"d0",
          4211 => x"52",
          4212 => x"51",
          4213 => x"3f",
          4214 => x"33",
          4215 => x"2e",
          4216 => x"ba",
          4217 => x"82",
          4218 => x"ff",
          4219 => x"82",
          4220 => x"54",
          4221 => x"8e",
          4222 => x"90",
          4223 => x"ac",
          4224 => x"8f",
          4225 => x"ba",
          4226 => x"73",
          4227 => x"38",
          4228 => x"33",
          4229 => x"dc",
          4230 => x"bd",
          4231 => x"81",
          4232 => x"80",
          4233 => x"82",
          4234 => x"ff",
          4235 => x"82",
          4236 => x"54",
          4237 => x"89",
          4238 => x"90",
          4239 => x"c6",
          4240 => x"88",
          4241 => x"80",
          4242 => x"82",
          4243 => x"ff",
          4244 => x"82",
          4245 => x"54",
          4246 => x"89",
          4247 => x"a8",
          4248 => x"a2",
          4249 => x"8a",
          4250 => x"80",
          4251 => x"82",
          4252 => x"ff",
          4253 => x"82",
          4254 => x"ff",
          4255 => x"82",
          4256 => x"52",
          4257 => x"51",
          4258 => x"3f",
          4259 => x"08",
          4260 => x"f4",
          4261 => x"c1",
          4262 => x"ec",
          4263 => x"ae",
          4264 => x"8e",
          4265 => x"ae",
          4266 => x"b5",
          4267 => x"b9",
          4268 => x"82",
          4269 => x"ff",
          4270 => x"82",
          4271 => x"56",
          4272 => x"52",
          4273 => x"de",
          4274 => x"98",
          4275 => x"c0",
          4276 => x"31",
          4277 => x"bb",
          4278 => x"82",
          4279 => x"ff",
          4280 => x"82",
          4281 => x"54",
          4282 => x"a9",
          4283 => x"f8",
          4284 => x"84",
          4285 => x"51",
          4286 => x"82",
          4287 => x"bd",
          4288 => x"76",
          4289 => x"54",
          4290 => x"08",
          4291 => x"a0",
          4292 => x"c5",
          4293 => x"82",
          4294 => x"80",
          4295 => x"82",
          4296 => x"56",
          4297 => x"52",
          4298 => x"fa",
          4299 => x"98",
          4300 => x"c0",
          4301 => x"31",
          4302 => x"bb",
          4303 => x"82",
          4304 => x"ff",
          4305 => x"82",
          4306 => x"ff",
          4307 => x"87",
          4308 => x"fe",
          4309 => x"92",
          4310 => x"05",
          4311 => x"26",
          4312 => x"84",
          4313 => x"80",
          4314 => x"08",
          4315 => x"f8",
          4316 => x"82",
          4317 => x"97",
          4318 => x"88",
          4319 => x"82",
          4320 => x"8b",
          4321 => x"94",
          4322 => x"82",
          4323 => x"ff",
          4324 => x"84",
          4325 => x"71",
          4326 => x"04",
          4327 => x"87",
          4328 => x"70",
          4329 => x"80",
          4330 => x"74",
          4331 => x"ba",
          4332 => x"0c",
          4333 => x"04",
          4334 => x"87",
          4335 => x"70",
          4336 => x"94",
          4337 => x"72",
          4338 => x"70",
          4339 => x"08",
          4340 => x"ba",
          4341 => x"0c",
          4342 => x"0d",
          4343 => x"87",
          4344 => x"0c",
          4345 => x"94",
          4346 => x"96",
          4347 => x"fd",
          4348 => x"98",
          4349 => x"2c",
          4350 => x"70",
          4351 => x"10",
          4352 => x"2b",
          4353 => x"54",
          4354 => x"0b",
          4355 => x"12",
          4356 => x"71",
          4357 => x"38",
          4358 => x"11",
          4359 => x"84",
          4360 => x"33",
          4361 => x"52",
          4362 => x"2e",
          4363 => x"83",
          4364 => x"72",
          4365 => x"0c",
          4366 => x"04",
          4367 => x"78",
          4368 => x"9f",
          4369 => x"33",
          4370 => x"71",
          4371 => x"38",
          4372 => x"b5",
          4373 => x"51",
          4374 => x"3f",
          4375 => x"b5",
          4376 => x"33",
          4377 => x"71",
          4378 => x"81",
          4379 => x"db",
          4380 => x"ff",
          4381 => x"73",
          4382 => x"3d",
          4383 => x"3d",
          4384 => x"84",
          4385 => x"33",
          4386 => x"bb",
          4387 => x"ba",
          4388 => x"84",
          4389 => x"98",
          4390 => x"51",
          4391 => x"58",
          4392 => x"2e",
          4393 => x"51",
          4394 => x"82",
          4395 => x"70",
          4396 => x"ba",
          4397 => x"19",
          4398 => x"56",
          4399 => x"3f",
          4400 => x"08",
          4401 => x"ba",
          4402 => x"84",
          4403 => x"98",
          4404 => x"51",
          4405 => x"80",
          4406 => x"75",
          4407 => x"74",
          4408 => x"a4",
          4409 => x"f0",
          4410 => x"55",
          4411 => x"f0",
          4412 => x"ff",
          4413 => x"75",
          4414 => x"80",
          4415 => x"f0",
          4416 => x"2e",
          4417 => x"ba",
          4418 => x"75",
          4419 => x"38",
          4420 => x"33",
          4421 => x"38",
          4422 => x"05",
          4423 => x"78",
          4424 => x"80",
          4425 => x"82",
          4426 => x"52",
          4427 => x"8e",
          4428 => x"ba",
          4429 => x"80",
          4430 => x"8c",
          4431 => x"fd",
          4432 => x"ba",
          4433 => x"54",
          4434 => x"71",
          4435 => x"38",
          4436 => x"8b",
          4437 => x"0c",
          4438 => x"14",
          4439 => x"80",
          4440 => x"80",
          4441 => x"f0",
          4442 => x"ec",
          4443 => x"80",
          4444 => x"71",
          4445 => x"80",
          4446 => x"ec",
          4447 => x"df",
          4448 => x"82",
          4449 => x"85",
          4450 => x"dc",
          4451 => x"57",
          4452 => x"ba",
          4453 => x"80",
          4454 => x"82",
          4455 => x"80",
          4456 => x"ba",
          4457 => x"80",
          4458 => x"3d",
          4459 => x"81",
          4460 => x"82",
          4461 => x"80",
          4462 => x"75",
          4463 => x"e8",
          4464 => x"98",
          4465 => x"0b",
          4466 => x"08",
          4467 => x"82",
          4468 => x"ff",
          4469 => x"55",
          4470 => x"34",
          4471 => x"52",
          4472 => x"b3",
          4473 => x"ff",
          4474 => x"74",
          4475 => x"81",
          4476 => x"38",
          4477 => x"04",
          4478 => x"aa",
          4479 => x"3d",
          4480 => x"81",
          4481 => x"80",
          4482 => x"ec",
          4483 => x"e1",
          4484 => x"bb",
          4485 => x"95",
          4486 => x"82",
          4487 => x"54",
          4488 => x"52",
          4489 => x"52",
          4490 => x"c1",
          4491 => x"98",
          4492 => x"a5",
          4493 => x"ff",
          4494 => x"82",
          4495 => x"81",
          4496 => x"80",
          4497 => x"98",
          4498 => x"38",
          4499 => x"08",
          4500 => x"17",
          4501 => x"74",
          4502 => x"70",
          4503 => x"07",
          4504 => x"55",
          4505 => x"2e",
          4506 => x"ff",
          4507 => x"ba",
          4508 => x"11",
          4509 => x"80",
          4510 => x"82",
          4511 => x"80",
          4512 => x"82",
          4513 => x"ff",
          4514 => x"78",
          4515 => x"81",
          4516 => x"75",
          4517 => x"ff",
          4518 => x"79",
          4519 => x"88",
          4520 => x"08",
          4521 => x"98",
          4522 => x"80",
          4523 => x"bb",
          4524 => x"3d",
          4525 => x"3d",
          4526 => x"71",
          4527 => x"33",
          4528 => x"58",
          4529 => x"09",
          4530 => x"38",
          4531 => x"05",
          4532 => x"27",
          4533 => x"17",
          4534 => x"71",
          4535 => x"55",
          4536 => x"09",
          4537 => x"38",
          4538 => x"ea",
          4539 => x"73",
          4540 => x"ba",
          4541 => x"08",
          4542 => x"b9",
          4543 => x"bb",
          4544 => x"79",
          4545 => x"51",
          4546 => x"3f",
          4547 => x"08",
          4548 => x"84",
          4549 => x"74",
          4550 => x"38",
          4551 => x"88",
          4552 => x"fc",
          4553 => x"39",
          4554 => x"8c",
          4555 => x"53",
          4556 => x"ff",
          4557 => x"82",
          4558 => x"80",
          4559 => x"ff",
          4560 => x"52",
          4561 => x"b0",
          4562 => x"98",
          4563 => x"06",
          4564 => x"38",
          4565 => x"39",
          4566 => x"81",
          4567 => x"54",
          4568 => x"ff",
          4569 => x"54",
          4570 => x"98",
          4571 => x"0d",
          4572 => x"0d",
          4573 => x"b2",
          4574 => x"3d",
          4575 => x"5a",
          4576 => x"3d",
          4577 => x"f0",
          4578 => x"ec",
          4579 => x"73",
          4580 => x"73",
          4581 => x"33",
          4582 => x"83",
          4583 => x"76",
          4584 => x"bc",
          4585 => x"76",
          4586 => x"73",
          4587 => x"ad",
          4588 => x"97",
          4589 => x"bb",
          4590 => x"ba",
          4591 => x"bb",
          4592 => x"2e",
          4593 => x"93",
          4594 => x"82",
          4595 => x"51",
          4596 => x"3f",
          4597 => x"08",
          4598 => x"38",
          4599 => x"51",
          4600 => x"3f",
          4601 => x"82",
          4602 => x"5b",
          4603 => x"08",
          4604 => x"52",
          4605 => x"52",
          4606 => x"f1",
          4607 => x"98",
          4608 => x"bb",
          4609 => x"2e",
          4610 => x"80",
          4611 => x"bb",
          4612 => x"ff",
          4613 => x"82",
          4614 => x"55",
          4615 => x"bb",
          4616 => x"a9",
          4617 => x"98",
          4618 => x"70",
          4619 => x"80",
          4620 => x"53",
          4621 => x"06",
          4622 => x"f8",
          4623 => x"1b",
          4624 => x"06",
          4625 => x"7b",
          4626 => x"80",
          4627 => x"2e",
          4628 => x"ff",
          4629 => x"39",
          4630 => x"e8",
          4631 => x"38",
          4632 => x"08",
          4633 => x"38",
          4634 => x"8f",
          4635 => x"90",
          4636 => x"98",
          4637 => x"70",
          4638 => x"59",
          4639 => x"ee",
          4640 => x"ff",
          4641 => x"c4",
          4642 => x"2b",
          4643 => x"82",
          4644 => x"70",
          4645 => x"97",
          4646 => x"2c",
          4647 => x"29",
          4648 => x"05",
          4649 => x"70",
          4650 => x"51",
          4651 => x"51",
          4652 => x"81",
          4653 => x"2e",
          4654 => x"77",
          4655 => x"38",
          4656 => x"0a",
          4657 => x"0a",
          4658 => x"2c",
          4659 => x"75",
          4660 => x"38",
          4661 => x"52",
          4662 => x"93",
          4663 => x"98",
          4664 => x"06",
          4665 => x"2e",
          4666 => x"82",
          4667 => x"81",
          4668 => x"74",
          4669 => x"29",
          4670 => x"05",
          4671 => x"70",
          4672 => x"56",
          4673 => x"95",
          4674 => x"76",
          4675 => x"77",
          4676 => x"3f",
          4677 => x"08",
          4678 => x"54",
          4679 => x"d3",
          4680 => x"75",
          4681 => x"ca",
          4682 => x"55",
          4683 => x"c4",
          4684 => x"2b",
          4685 => x"82",
          4686 => x"70",
          4687 => x"98",
          4688 => x"11",
          4689 => x"82",
          4690 => x"33",
          4691 => x"51",
          4692 => x"55",
          4693 => x"09",
          4694 => x"92",
          4695 => x"ac",
          4696 => x"0c",
          4697 => x"d2",
          4698 => x"0b",
          4699 => x"34",
          4700 => x"82",
          4701 => x"75",
          4702 => x"34",
          4703 => x"34",
          4704 => x"7e",
          4705 => x"26",
          4706 => x"73",
          4707 => x"9a",
          4708 => x"73",
          4709 => x"d2",
          4710 => x"73",
          4711 => x"cb",
          4712 => x"c8",
          4713 => x"75",
          4714 => x"74",
          4715 => x"98",
          4716 => x"73",
          4717 => x"38",
          4718 => x"73",
          4719 => x"34",
          4720 => x"0a",
          4721 => x"0a",
          4722 => x"2c",
          4723 => x"33",
          4724 => x"df",
          4725 => x"cc",
          4726 => x"56",
          4727 => x"d2",
          4728 => x"1a",
          4729 => x"33",
          4730 => x"d2",
          4731 => x"73",
          4732 => x"38",
          4733 => x"73",
          4734 => x"34",
          4735 => x"33",
          4736 => x"0a",
          4737 => x"0a",
          4738 => x"2c",
          4739 => x"33",
          4740 => x"56",
          4741 => x"a3",
          4742 => x"70",
          4743 => x"ff",
          4744 => x"74",
          4745 => x"29",
          4746 => x"05",
          4747 => x"82",
          4748 => x"56",
          4749 => x"75",
          4750 => x"82",
          4751 => x"70",
          4752 => x"98",
          4753 => x"c8",
          4754 => x"56",
          4755 => x"25",
          4756 => x"88",
          4757 => x"d0",
          4758 => x"80",
          4759 => x"80",
          4760 => x"98",
          4761 => x"c8",
          4762 => x"55",
          4763 => x"e3",
          4764 => x"39",
          4765 => x"80",
          4766 => x"34",
          4767 => x"53",
          4768 => x"a9",
          4769 => x"b4",
          4770 => x"39",
          4771 => x"33",
          4772 => x"06",
          4773 => x"80",
          4774 => x"38",
          4775 => x"33",
          4776 => x"73",
          4777 => x"34",
          4778 => x"73",
          4779 => x"34",
          4780 => x"a8",
          4781 => x"d2",
          4782 => x"98",
          4783 => x"2c",
          4784 => x"33",
          4785 => x"57",
          4786 => x"a8",
          4787 => x"54",
          4788 => x"74",
          4789 => x"51",
          4790 => x"3f",
          4791 => x"0a",
          4792 => x"0a",
          4793 => x"2c",
          4794 => x"33",
          4795 => x"75",
          4796 => x"38",
          4797 => x"a8",
          4798 => x"d2",
          4799 => x"98",
          4800 => x"2c",
          4801 => x"33",
          4802 => x"57",
          4803 => x"fa",
          4804 => x"51",
          4805 => x"3f",
          4806 => x"0a",
          4807 => x"0a",
          4808 => x"2c",
          4809 => x"33",
          4810 => x"75",
          4811 => x"38",
          4812 => x"82",
          4813 => x"7a",
          4814 => x"74",
          4815 => x"ff",
          4816 => x"82",
          4817 => x"79",
          4818 => x"3f",
          4819 => x"08",
          4820 => x"54",
          4821 => x"82",
          4822 => x"54",
          4823 => x"8f",
          4824 => x"73",
          4825 => x"f2",
          4826 => x"39",
          4827 => x"80",
          4828 => x"cc",
          4829 => x"82",
          4830 => x"79",
          4831 => x"0c",
          4832 => x"04",
          4833 => x"33",
          4834 => x"2e",
          4835 => x"88",
          4836 => x"94",
          4837 => x"cc",
          4838 => x"54",
          4839 => x"cc",
          4840 => x"ff",
          4841 => x"39",
          4842 => x"33",
          4843 => x"33",
          4844 => x"75",
          4845 => x"38",
          4846 => x"73",
          4847 => x"34",
          4848 => x"70",
          4849 => x"81",
          4850 => x"51",
          4851 => x"25",
          4852 => x"1a",
          4853 => x"33",
          4854 => x"33",
          4855 => x"c8",
          4856 => x"80",
          4857 => x"80",
          4858 => x"98",
          4859 => x"c8",
          4860 => x"55",
          4861 => x"da",
          4862 => x"ff",
          4863 => x"82",
          4864 => x"70",
          4865 => x"98",
          4866 => x"c8",
          4867 => x"56",
          4868 => x"24",
          4869 => x"88",
          4870 => x"8c",
          4871 => x"80",
          4872 => x"80",
          4873 => x"98",
          4874 => x"c8",
          4875 => x"55",
          4876 => x"e3",
          4877 => x"39",
          4878 => x"33",
          4879 => x"06",
          4880 => x"33",
          4881 => x"74",
          4882 => x"9f",
          4883 => x"54",
          4884 => x"cc",
          4885 => x"70",
          4886 => x"ff",
          4887 => x"82",
          4888 => x"70",
          4889 => x"82",
          4890 => x"58",
          4891 => x"75",
          4892 => x"f7",
          4893 => x"d2",
          4894 => x"52",
          4895 => x"51",
          4896 => x"80",
          4897 => x"cc",
          4898 => x"82",
          4899 => x"f7",
          4900 => x"b0",
          4901 => x"e4",
          4902 => x"80",
          4903 => x"74",
          4904 => x"84",
          4905 => x"98",
          4906 => x"c8",
          4907 => x"98",
          4908 => x"06",
          4909 => x"74",
          4910 => x"ff",
          4911 => x"93",
          4912 => x"39",
          4913 => x"82",
          4914 => x"fc",
          4915 => x"54",
          4916 => x"a7",
          4917 => x"ff",
          4918 => x"82",
          4919 => x"82",
          4920 => x"82",
          4921 => x"81",
          4922 => x"05",
          4923 => x"79",
          4924 => x"94",
          4925 => x"54",
          4926 => x"73",
          4927 => x"80",
          4928 => x"38",
          4929 => x"ad",
          4930 => x"39",
          4931 => x"09",
          4932 => x"38",
          4933 => x"08",
          4934 => x"2e",
          4935 => x"51",
          4936 => x"3f",
          4937 => x"08",
          4938 => x"34",
          4939 => x"08",
          4940 => x"81",
          4941 => x"52",
          4942 => x"ae",
          4943 => x"c3",
          4944 => x"29",
          4945 => x"05",
          4946 => x"54",
          4947 => x"ab",
          4948 => x"ff",
          4949 => x"82",
          4950 => x"82",
          4951 => x"82",
          4952 => x"81",
          4953 => x"05",
          4954 => x"79",
          4955 => x"98",
          4956 => x"54",
          4957 => x"06",
          4958 => x"74",
          4959 => x"34",
          4960 => x"82",
          4961 => x"82",
          4962 => x"52",
          4963 => x"ac",
          4964 => x"39",
          4965 => x"33",
          4966 => x"06",
          4967 => x"33",
          4968 => x"74",
          4969 => x"c3",
          4970 => x"54",
          4971 => x"cc",
          4972 => x"70",
          4973 => x"ff",
          4974 => x"f5",
          4975 => x"d2",
          4976 => x"73",
          4977 => x"a3",
          4978 => x"ff",
          4979 => x"82",
          4980 => x"ff",
          4981 => x"82",
          4982 => x"f5",
          4983 => x"3d",
          4984 => x"80",
          4985 => x"90",
          4986 => x"0b",
          4987 => x"23",
          4988 => x"80",
          4989 => x"80",
          4990 => x"8d",
          4991 => x"90",
          4992 => x"58",
          4993 => x"81",
          4994 => x"15",
          4995 => x"90",
          4996 => x"84",
          4997 => x"85",
          4998 => x"bb",
          4999 => x"77",
          5000 => x"76",
          5001 => x"82",
          5002 => x"82",
          5003 => x"ff",
          5004 => x"80",
          5005 => x"ff",
          5006 => x"88",
          5007 => x"55",
          5008 => x"17",
          5009 => x"17",
          5010 => x"8c",
          5011 => x"29",
          5012 => x"08",
          5013 => x"51",
          5014 => x"82",
          5015 => x"83",
          5016 => x"3d",
          5017 => x"3d",
          5018 => x"81",
          5019 => x"27",
          5020 => x"12",
          5021 => x"11",
          5022 => x"ff",
          5023 => x"51",
          5024 => x"98",
          5025 => x"0d",
          5026 => x"0d",
          5027 => x"22",
          5028 => x"aa",
          5029 => x"05",
          5030 => x"08",
          5031 => x"71",
          5032 => x"2b",
          5033 => x"33",
          5034 => x"71",
          5035 => x"02",
          5036 => x"05",
          5037 => x"ff",
          5038 => x"70",
          5039 => x"51",
          5040 => x"5b",
          5041 => x"54",
          5042 => x"34",
          5043 => x"34",
          5044 => x"08",
          5045 => x"2a",
          5046 => x"82",
          5047 => x"83",
          5048 => x"bb",
          5049 => x"17",
          5050 => x"12",
          5051 => x"2b",
          5052 => x"2b",
          5053 => x"06",
          5054 => x"52",
          5055 => x"83",
          5056 => x"70",
          5057 => x"54",
          5058 => x"12",
          5059 => x"ff",
          5060 => x"83",
          5061 => x"bb",
          5062 => x"56",
          5063 => x"72",
          5064 => x"89",
          5065 => x"fb",
          5066 => x"bb",
          5067 => x"84",
          5068 => x"22",
          5069 => x"72",
          5070 => x"33",
          5071 => x"71",
          5072 => x"83",
          5073 => x"5b",
          5074 => x"52",
          5075 => x"12",
          5076 => x"33",
          5077 => x"07",
          5078 => x"54",
          5079 => x"70",
          5080 => x"73",
          5081 => x"82",
          5082 => x"70",
          5083 => x"33",
          5084 => x"71",
          5085 => x"83",
          5086 => x"59",
          5087 => x"05",
          5088 => x"87",
          5089 => x"88",
          5090 => x"88",
          5091 => x"56",
          5092 => x"13",
          5093 => x"13",
          5094 => x"90",
          5095 => x"33",
          5096 => x"71",
          5097 => x"70",
          5098 => x"06",
          5099 => x"53",
          5100 => x"53",
          5101 => x"70",
          5102 => x"87",
          5103 => x"fa",
          5104 => x"a2",
          5105 => x"bb",
          5106 => x"83",
          5107 => x"70",
          5108 => x"33",
          5109 => x"07",
          5110 => x"15",
          5111 => x"12",
          5112 => x"2b",
          5113 => x"07",
          5114 => x"55",
          5115 => x"57",
          5116 => x"80",
          5117 => x"38",
          5118 => x"ab",
          5119 => x"90",
          5120 => x"70",
          5121 => x"33",
          5122 => x"71",
          5123 => x"74",
          5124 => x"81",
          5125 => x"88",
          5126 => x"83",
          5127 => x"f8",
          5128 => x"54",
          5129 => x"58",
          5130 => x"74",
          5131 => x"52",
          5132 => x"34",
          5133 => x"34",
          5134 => x"08",
          5135 => x"33",
          5136 => x"71",
          5137 => x"83",
          5138 => x"59",
          5139 => x"05",
          5140 => x"12",
          5141 => x"2b",
          5142 => x"ff",
          5143 => x"88",
          5144 => x"52",
          5145 => x"74",
          5146 => x"15",
          5147 => x"0d",
          5148 => x"0d",
          5149 => x"08",
          5150 => x"9e",
          5151 => x"83",
          5152 => x"82",
          5153 => x"12",
          5154 => x"2b",
          5155 => x"07",
          5156 => x"52",
          5157 => x"05",
          5158 => x"13",
          5159 => x"2b",
          5160 => x"05",
          5161 => x"71",
          5162 => x"2a",
          5163 => x"53",
          5164 => x"34",
          5165 => x"34",
          5166 => x"08",
          5167 => x"33",
          5168 => x"71",
          5169 => x"83",
          5170 => x"59",
          5171 => x"05",
          5172 => x"83",
          5173 => x"88",
          5174 => x"88",
          5175 => x"56",
          5176 => x"13",
          5177 => x"13",
          5178 => x"90",
          5179 => x"11",
          5180 => x"33",
          5181 => x"07",
          5182 => x"0c",
          5183 => x"3d",
          5184 => x"3d",
          5185 => x"bb",
          5186 => x"83",
          5187 => x"ff",
          5188 => x"53",
          5189 => x"a7",
          5190 => x"90",
          5191 => x"2b",
          5192 => x"11",
          5193 => x"33",
          5194 => x"71",
          5195 => x"75",
          5196 => x"81",
          5197 => x"98",
          5198 => x"2b",
          5199 => x"40",
          5200 => x"58",
          5201 => x"72",
          5202 => x"38",
          5203 => x"52",
          5204 => x"9d",
          5205 => x"39",
          5206 => x"85",
          5207 => x"8b",
          5208 => x"2b",
          5209 => x"79",
          5210 => x"51",
          5211 => x"76",
          5212 => x"75",
          5213 => x"56",
          5214 => x"34",
          5215 => x"08",
          5216 => x"12",
          5217 => x"33",
          5218 => x"07",
          5219 => x"54",
          5220 => x"53",
          5221 => x"34",
          5222 => x"34",
          5223 => x"08",
          5224 => x"0b",
          5225 => x"80",
          5226 => x"34",
          5227 => x"08",
          5228 => x"14",
          5229 => x"14",
          5230 => x"90",
          5231 => x"33",
          5232 => x"71",
          5233 => x"70",
          5234 => x"07",
          5235 => x"53",
          5236 => x"54",
          5237 => x"72",
          5238 => x"8b",
          5239 => x"ff",
          5240 => x"52",
          5241 => x"08",
          5242 => x"f2",
          5243 => x"2e",
          5244 => x"51",
          5245 => x"83",
          5246 => x"f5",
          5247 => x"7e",
          5248 => x"e2",
          5249 => x"98",
          5250 => x"ff",
          5251 => x"90",
          5252 => x"33",
          5253 => x"71",
          5254 => x"70",
          5255 => x"58",
          5256 => x"ff",
          5257 => x"2e",
          5258 => x"75",
          5259 => x"70",
          5260 => x"33",
          5261 => x"07",
          5262 => x"ff",
          5263 => x"70",
          5264 => x"06",
          5265 => x"52",
          5266 => x"59",
          5267 => x"27",
          5268 => x"80",
          5269 => x"75",
          5270 => x"84",
          5271 => x"16",
          5272 => x"2b",
          5273 => x"75",
          5274 => x"81",
          5275 => x"85",
          5276 => x"59",
          5277 => x"83",
          5278 => x"90",
          5279 => x"33",
          5280 => x"71",
          5281 => x"70",
          5282 => x"06",
          5283 => x"56",
          5284 => x"75",
          5285 => x"81",
          5286 => x"79",
          5287 => x"cc",
          5288 => x"74",
          5289 => x"c4",
          5290 => x"2e",
          5291 => x"89",
          5292 => x"f8",
          5293 => x"ac",
          5294 => x"80",
          5295 => x"75",
          5296 => x"3f",
          5297 => x"08",
          5298 => x"11",
          5299 => x"33",
          5300 => x"71",
          5301 => x"53",
          5302 => x"74",
          5303 => x"70",
          5304 => x"06",
          5305 => x"5c",
          5306 => x"78",
          5307 => x"76",
          5308 => x"57",
          5309 => x"34",
          5310 => x"08",
          5311 => x"71",
          5312 => x"86",
          5313 => x"12",
          5314 => x"2b",
          5315 => x"2a",
          5316 => x"53",
          5317 => x"73",
          5318 => x"75",
          5319 => x"82",
          5320 => x"70",
          5321 => x"33",
          5322 => x"71",
          5323 => x"83",
          5324 => x"5d",
          5325 => x"05",
          5326 => x"15",
          5327 => x"15",
          5328 => x"90",
          5329 => x"71",
          5330 => x"33",
          5331 => x"71",
          5332 => x"70",
          5333 => x"5a",
          5334 => x"54",
          5335 => x"34",
          5336 => x"34",
          5337 => x"08",
          5338 => x"54",
          5339 => x"98",
          5340 => x"0d",
          5341 => x"0d",
          5342 => x"bb",
          5343 => x"38",
          5344 => x"71",
          5345 => x"2e",
          5346 => x"51",
          5347 => x"82",
          5348 => x"53",
          5349 => x"98",
          5350 => x"0d",
          5351 => x"0d",
          5352 => x"5c",
          5353 => x"40",
          5354 => x"08",
          5355 => x"81",
          5356 => x"f4",
          5357 => x"8e",
          5358 => x"ff",
          5359 => x"bb",
          5360 => x"83",
          5361 => x"8b",
          5362 => x"fc",
          5363 => x"54",
          5364 => x"7e",
          5365 => x"3f",
          5366 => x"08",
          5367 => x"06",
          5368 => x"08",
          5369 => x"83",
          5370 => x"ff",
          5371 => x"83",
          5372 => x"70",
          5373 => x"33",
          5374 => x"07",
          5375 => x"70",
          5376 => x"06",
          5377 => x"fc",
          5378 => x"29",
          5379 => x"81",
          5380 => x"88",
          5381 => x"90",
          5382 => x"4e",
          5383 => x"52",
          5384 => x"41",
          5385 => x"5b",
          5386 => x"8f",
          5387 => x"ff",
          5388 => x"31",
          5389 => x"ff",
          5390 => x"82",
          5391 => x"17",
          5392 => x"2b",
          5393 => x"29",
          5394 => x"81",
          5395 => x"98",
          5396 => x"2b",
          5397 => x"45",
          5398 => x"73",
          5399 => x"38",
          5400 => x"70",
          5401 => x"06",
          5402 => x"7b",
          5403 => x"38",
          5404 => x"73",
          5405 => x"81",
          5406 => x"78",
          5407 => x"3f",
          5408 => x"ff",
          5409 => x"e5",
          5410 => x"38",
          5411 => x"89",
          5412 => x"f6",
          5413 => x"a5",
          5414 => x"55",
          5415 => x"80",
          5416 => x"1d",
          5417 => x"83",
          5418 => x"88",
          5419 => x"57",
          5420 => x"3f",
          5421 => x"51",
          5422 => x"82",
          5423 => x"83",
          5424 => x"7e",
          5425 => x"70",
          5426 => x"bb",
          5427 => x"84",
          5428 => x"59",
          5429 => x"3f",
          5430 => x"08",
          5431 => x"75",
          5432 => x"06",
          5433 => x"85",
          5434 => x"54",
          5435 => x"80",
          5436 => x"51",
          5437 => x"82",
          5438 => x"1d",
          5439 => x"83",
          5440 => x"88",
          5441 => x"43",
          5442 => x"3f",
          5443 => x"51",
          5444 => x"82",
          5445 => x"83",
          5446 => x"7e",
          5447 => x"70",
          5448 => x"bb",
          5449 => x"84",
          5450 => x"59",
          5451 => x"3f",
          5452 => x"08",
          5453 => x"60",
          5454 => x"55",
          5455 => x"ff",
          5456 => x"a9",
          5457 => x"52",
          5458 => x"3f",
          5459 => x"08",
          5460 => x"98",
          5461 => x"93",
          5462 => x"73",
          5463 => x"98",
          5464 => x"9e",
          5465 => x"51",
          5466 => x"7a",
          5467 => x"27",
          5468 => x"53",
          5469 => x"51",
          5470 => x"7a",
          5471 => x"82",
          5472 => x"05",
          5473 => x"f6",
          5474 => x"54",
          5475 => x"98",
          5476 => x"0d",
          5477 => x"0d",
          5478 => x"70",
          5479 => x"d5",
          5480 => x"98",
          5481 => x"bb",
          5482 => x"2e",
          5483 => x"53",
          5484 => x"bb",
          5485 => x"ff",
          5486 => x"74",
          5487 => x"0c",
          5488 => x"04",
          5489 => x"02",
          5490 => x"51",
          5491 => x"72",
          5492 => x"82",
          5493 => x"33",
          5494 => x"bb",
          5495 => x"3d",
          5496 => x"3d",
          5497 => x"05",
          5498 => x"05",
          5499 => x"56",
          5500 => x"72",
          5501 => x"e0",
          5502 => x"2b",
          5503 => x"8c",
          5504 => x"88",
          5505 => x"2e",
          5506 => x"88",
          5507 => x"0c",
          5508 => x"8c",
          5509 => x"71",
          5510 => x"87",
          5511 => x"0c",
          5512 => x"08",
          5513 => x"51",
          5514 => x"2e",
          5515 => x"c0",
          5516 => x"51",
          5517 => x"71",
          5518 => x"80",
          5519 => x"92",
          5520 => x"98",
          5521 => x"70",
          5522 => x"38",
          5523 => x"94",
          5524 => x"bb",
          5525 => x"51",
          5526 => x"98",
          5527 => x"0d",
          5528 => x"0d",
          5529 => x"02",
          5530 => x"05",
          5531 => x"58",
          5532 => x"52",
          5533 => x"3f",
          5534 => x"08",
          5535 => x"54",
          5536 => x"be",
          5537 => x"75",
          5538 => x"c0",
          5539 => x"87",
          5540 => x"12",
          5541 => x"84",
          5542 => x"40",
          5543 => x"85",
          5544 => x"98",
          5545 => x"7d",
          5546 => x"0c",
          5547 => x"85",
          5548 => x"06",
          5549 => x"71",
          5550 => x"38",
          5551 => x"71",
          5552 => x"05",
          5553 => x"19",
          5554 => x"a2",
          5555 => x"71",
          5556 => x"38",
          5557 => x"83",
          5558 => x"38",
          5559 => x"8a",
          5560 => x"98",
          5561 => x"71",
          5562 => x"c0",
          5563 => x"52",
          5564 => x"87",
          5565 => x"80",
          5566 => x"81",
          5567 => x"c0",
          5568 => x"53",
          5569 => x"82",
          5570 => x"71",
          5571 => x"1a",
          5572 => x"84",
          5573 => x"19",
          5574 => x"06",
          5575 => x"79",
          5576 => x"38",
          5577 => x"80",
          5578 => x"87",
          5579 => x"26",
          5580 => x"73",
          5581 => x"06",
          5582 => x"2e",
          5583 => x"52",
          5584 => x"82",
          5585 => x"8f",
          5586 => x"f3",
          5587 => x"62",
          5588 => x"05",
          5589 => x"57",
          5590 => x"83",
          5591 => x"52",
          5592 => x"3f",
          5593 => x"08",
          5594 => x"54",
          5595 => x"2e",
          5596 => x"81",
          5597 => x"74",
          5598 => x"c0",
          5599 => x"87",
          5600 => x"12",
          5601 => x"84",
          5602 => x"5f",
          5603 => x"0b",
          5604 => x"8c",
          5605 => x"0c",
          5606 => x"80",
          5607 => x"70",
          5608 => x"81",
          5609 => x"54",
          5610 => x"8c",
          5611 => x"81",
          5612 => x"7c",
          5613 => x"58",
          5614 => x"70",
          5615 => x"52",
          5616 => x"8a",
          5617 => x"98",
          5618 => x"71",
          5619 => x"c0",
          5620 => x"52",
          5621 => x"87",
          5622 => x"80",
          5623 => x"81",
          5624 => x"c0",
          5625 => x"53",
          5626 => x"82",
          5627 => x"71",
          5628 => x"19",
          5629 => x"81",
          5630 => x"ff",
          5631 => x"19",
          5632 => x"78",
          5633 => x"38",
          5634 => x"80",
          5635 => x"87",
          5636 => x"26",
          5637 => x"73",
          5638 => x"06",
          5639 => x"2e",
          5640 => x"52",
          5641 => x"82",
          5642 => x"8f",
          5643 => x"fa",
          5644 => x"02",
          5645 => x"05",
          5646 => x"05",
          5647 => x"71",
          5648 => x"57",
          5649 => x"82",
          5650 => x"81",
          5651 => x"54",
          5652 => x"38",
          5653 => x"c0",
          5654 => x"81",
          5655 => x"2e",
          5656 => x"71",
          5657 => x"38",
          5658 => x"87",
          5659 => x"11",
          5660 => x"80",
          5661 => x"80",
          5662 => x"83",
          5663 => x"38",
          5664 => x"72",
          5665 => x"2a",
          5666 => x"51",
          5667 => x"80",
          5668 => x"87",
          5669 => x"08",
          5670 => x"38",
          5671 => x"8c",
          5672 => x"96",
          5673 => x"0c",
          5674 => x"8c",
          5675 => x"08",
          5676 => x"51",
          5677 => x"38",
          5678 => x"56",
          5679 => x"80",
          5680 => x"85",
          5681 => x"77",
          5682 => x"83",
          5683 => x"75",
          5684 => x"bb",
          5685 => x"3d",
          5686 => x"3d",
          5687 => x"11",
          5688 => x"71",
          5689 => x"82",
          5690 => x"53",
          5691 => x"0d",
          5692 => x"0d",
          5693 => x"33",
          5694 => x"71",
          5695 => x"88",
          5696 => x"14",
          5697 => x"07",
          5698 => x"33",
          5699 => x"bb",
          5700 => x"53",
          5701 => x"52",
          5702 => x"04",
          5703 => x"73",
          5704 => x"92",
          5705 => x"52",
          5706 => x"81",
          5707 => x"70",
          5708 => x"70",
          5709 => x"3d",
          5710 => x"3d",
          5711 => x"52",
          5712 => x"70",
          5713 => x"34",
          5714 => x"51",
          5715 => x"81",
          5716 => x"70",
          5717 => x"70",
          5718 => x"05",
          5719 => x"88",
          5720 => x"72",
          5721 => x"0d",
          5722 => x"0d",
          5723 => x"54",
          5724 => x"80",
          5725 => x"71",
          5726 => x"53",
          5727 => x"81",
          5728 => x"ff",
          5729 => x"39",
          5730 => x"04",
          5731 => x"75",
          5732 => x"52",
          5733 => x"70",
          5734 => x"34",
          5735 => x"70",
          5736 => x"3d",
          5737 => x"3d",
          5738 => x"79",
          5739 => x"74",
          5740 => x"56",
          5741 => x"81",
          5742 => x"71",
          5743 => x"16",
          5744 => x"52",
          5745 => x"86",
          5746 => x"2e",
          5747 => x"82",
          5748 => x"86",
          5749 => x"fe",
          5750 => x"76",
          5751 => x"39",
          5752 => x"8a",
          5753 => x"51",
          5754 => x"71",
          5755 => x"33",
          5756 => x"0c",
          5757 => x"04",
          5758 => x"bb",
          5759 => x"80",
          5760 => x"98",
          5761 => x"3d",
          5762 => x"80",
          5763 => x"33",
          5764 => x"7a",
          5765 => x"38",
          5766 => x"16",
          5767 => x"16",
          5768 => x"17",
          5769 => x"fa",
          5770 => x"bb",
          5771 => x"2e",
          5772 => x"b7",
          5773 => x"98",
          5774 => x"34",
          5775 => x"70",
          5776 => x"31",
          5777 => x"59",
          5778 => x"77",
          5779 => x"82",
          5780 => x"74",
          5781 => x"81",
          5782 => x"81",
          5783 => x"53",
          5784 => x"16",
          5785 => x"e3",
          5786 => x"81",
          5787 => x"bb",
          5788 => x"3d",
          5789 => x"3d",
          5790 => x"56",
          5791 => x"74",
          5792 => x"2e",
          5793 => x"51",
          5794 => x"82",
          5795 => x"57",
          5796 => x"08",
          5797 => x"54",
          5798 => x"16",
          5799 => x"33",
          5800 => x"3f",
          5801 => x"08",
          5802 => x"38",
          5803 => x"57",
          5804 => x"0c",
          5805 => x"98",
          5806 => x"0d",
          5807 => x"0d",
          5808 => x"57",
          5809 => x"82",
          5810 => x"58",
          5811 => x"08",
          5812 => x"76",
          5813 => x"83",
          5814 => x"06",
          5815 => x"84",
          5816 => x"78",
          5817 => x"81",
          5818 => x"38",
          5819 => x"82",
          5820 => x"52",
          5821 => x"52",
          5822 => x"3f",
          5823 => x"52",
          5824 => x"51",
          5825 => x"84",
          5826 => x"d2",
          5827 => x"fc",
          5828 => x"8a",
          5829 => x"52",
          5830 => x"51",
          5831 => x"90",
          5832 => x"84",
          5833 => x"fc",
          5834 => x"17",
          5835 => x"a0",
          5836 => x"86",
          5837 => x"08",
          5838 => x"b0",
          5839 => x"55",
          5840 => x"81",
          5841 => x"f8",
          5842 => x"84",
          5843 => x"53",
          5844 => x"17",
          5845 => x"d7",
          5846 => x"98",
          5847 => x"83",
          5848 => x"77",
          5849 => x"0c",
          5850 => x"04",
          5851 => x"77",
          5852 => x"12",
          5853 => x"55",
          5854 => x"56",
          5855 => x"8d",
          5856 => x"22",
          5857 => x"ac",
          5858 => x"57",
          5859 => x"bb",
          5860 => x"3d",
          5861 => x"3d",
          5862 => x"70",
          5863 => x"57",
          5864 => x"81",
          5865 => x"98",
          5866 => x"81",
          5867 => x"74",
          5868 => x"72",
          5869 => x"f5",
          5870 => x"24",
          5871 => x"81",
          5872 => x"81",
          5873 => x"83",
          5874 => x"38",
          5875 => x"76",
          5876 => x"70",
          5877 => x"16",
          5878 => x"74",
          5879 => x"96",
          5880 => x"98",
          5881 => x"38",
          5882 => x"06",
          5883 => x"33",
          5884 => x"89",
          5885 => x"08",
          5886 => x"54",
          5887 => x"fc",
          5888 => x"bb",
          5889 => x"fe",
          5890 => x"ff",
          5891 => x"11",
          5892 => x"2b",
          5893 => x"81",
          5894 => x"2a",
          5895 => x"51",
          5896 => x"e2",
          5897 => x"ff",
          5898 => x"da",
          5899 => x"2a",
          5900 => x"05",
          5901 => x"fc",
          5902 => x"bb",
          5903 => x"c6",
          5904 => x"83",
          5905 => x"05",
          5906 => x"f9",
          5907 => x"bb",
          5908 => x"ff",
          5909 => x"ae",
          5910 => x"2a",
          5911 => x"05",
          5912 => x"fc",
          5913 => x"bb",
          5914 => x"38",
          5915 => x"83",
          5916 => x"05",
          5917 => x"f8",
          5918 => x"bb",
          5919 => x"0a",
          5920 => x"39",
          5921 => x"82",
          5922 => x"89",
          5923 => x"f8",
          5924 => x"7c",
          5925 => x"56",
          5926 => x"77",
          5927 => x"38",
          5928 => x"08",
          5929 => x"38",
          5930 => x"72",
          5931 => x"9d",
          5932 => x"24",
          5933 => x"81",
          5934 => x"82",
          5935 => x"83",
          5936 => x"38",
          5937 => x"76",
          5938 => x"70",
          5939 => x"18",
          5940 => x"76",
          5941 => x"9e",
          5942 => x"98",
          5943 => x"bb",
          5944 => x"d9",
          5945 => x"ff",
          5946 => x"05",
          5947 => x"81",
          5948 => x"54",
          5949 => x"80",
          5950 => x"77",
          5951 => x"f0",
          5952 => x"8f",
          5953 => x"51",
          5954 => x"34",
          5955 => x"17",
          5956 => x"2a",
          5957 => x"05",
          5958 => x"fa",
          5959 => x"bb",
          5960 => x"82",
          5961 => x"81",
          5962 => x"83",
          5963 => x"b4",
          5964 => x"2a",
          5965 => x"8f",
          5966 => x"2a",
          5967 => x"f0",
          5968 => x"06",
          5969 => x"72",
          5970 => x"ec",
          5971 => x"2a",
          5972 => x"05",
          5973 => x"fa",
          5974 => x"bb",
          5975 => x"82",
          5976 => x"80",
          5977 => x"83",
          5978 => x"52",
          5979 => x"fe",
          5980 => x"b4",
          5981 => x"a4",
          5982 => x"76",
          5983 => x"17",
          5984 => x"75",
          5985 => x"3f",
          5986 => x"08",
          5987 => x"98",
          5988 => x"77",
          5989 => x"77",
          5990 => x"fc",
          5991 => x"b4",
          5992 => x"51",
          5993 => x"c9",
          5994 => x"98",
          5995 => x"06",
          5996 => x"72",
          5997 => x"3f",
          5998 => x"17",
          5999 => x"bb",
          6000 => x"3d",
          6001 => x"3d",
          6002 => x"7e",
          6003 => x"56",
          6004 => x"75",
          6005 => x"74",
          6006 => x"27",
          6007 => x"80",
          6008 => x"ff",
          6009 => x"75",
          6010 => x"3f",
          6011 => x"08",
          6012 => x"98",
          6013 => x"38",
          6014 => x"54",
          6015 => x"81",
          6016 => x"39",
          6017 => x"08",
          6018 => x"39",
          6019 => x"51",
          6020 => x"82",
          6021 => x"58",
          6022 => x"08",
          6023 => x"c7",
          6024 => x"98",
          6025 => x"d2",
          6026 => x"98",
          6027 => x"cf",
          6028 => x"74",
          6029 => x"fc",
          6030 => x"bb",
          6031 => x"38",
          6032 => x"fe",
          6033 => x"08",
          6034 => x"74",
          6035 => x"38",
          6036 => x"17",
          6037 => x"33",
          6038 => x"73",
          6039 => x"77",
          6040 => x"26",
          6041 => x"80",
          6042 => x"bb",
          6043 => x"3d",
          6044 => x"3d",
          6045 => x"71",
          6046 => x"5b",
          6047 => x"8c",
          6048 => x"77",
          6049 => x"38",
          6050 => x"78",
          6051 => x"81",
          6052 => x"79",
          6053 => x"f9",
          6054 => x"55",
          6055 => x"98",
          6056 => x"e0",
          6057 => x"98",
          6058 => x"bb",
          6059 => x"2e",
          6060 => x"98",
          6061 => x"bb",
          6062 => x"82",
          6063 => x"58",
          6064 => x"70",
          6065 => x"80",
          6066 => x"38",
          6067 => x"09",
          6068 => x"e2",
          6069 => x"56",
          6070 => x"76",
          6071 => x"82",
          6072 => x"7a",
          6073 => x"3f",
          6074 => x"bb",
          6075 => x"2e",
          6076 => x"86",
          6077 => x"98",
          6078 => x"bb",
          6079 => x"70",
          6080 => x"07",
          6081 => x"7c",
          6082 => x"98",
          6083 => x"51",
          6084 => x"81",
          6085 => x"bb",
          6086 => x"2e",
          6087 => x"17",
          6088 => x"74",
          6089 => x"73",
          6090 => x"27",
          6091 => x"58",
          6092 => x"80",
          6093 => x"56",
          6094 => x"98",
          6095 => x"26",
          6096 => x"56",
          6097 => x"81",
          6098 => x"52",
          6099 => x"c6",
          6100 => x"98",
          6101 => x"b8",
          6102 => x"82",
          6103 => x"81",
          6104 => x"06",
          6105 => x"bb",
          6106 => x"82",
          6107 => x"09",
          6108 => x"72",
          6109 => x"70",
          6110 => x"51",
          6111 => x"80",
          6112 => x"78",
          6113 => x"06",
          6114 => x"73",
          6115 => x"39",
          6116 => x"52",
          6117 => x"f7",
          6118 => x"98",
          6119 => x"98",
          6120 => x"82",
          6121 => x"07",
          6122 => x"55",
          6123 => x"2e",
          6124 => x"80",
          6125 => x"75",
          6126 => x"76",
          6127 => x"3f",
          6128 => x"08",
          6129 => x"38",
          6130 => x"0c",
          6131 => x"fe",
          6132 => x"08",
          6133 => x"74",
          6134 => x"ff",
          6135 => x"0c",
          6136 => x"81",
          6137 => x"84",
          6138 => x"39",
          6139 => x"81",
          6140 => x"8c",
          6141 => x"8c",
          6142 => x"98",
          6143 => x"39",
          6144 => x"55",
          6145 => x"98",
          6146 => x"0d",
          6147 => x"0d",
          6148 => x"55",
          6149 => x"82",
          6150 => x"58",
          6151 => x"bb",
          6152 => x"d8",
          6153 => x"74",
          6154 => x"3f",
          6155 => x"08",
          6156 => x"08",
          6157 => x"59",
          6158 => x"77",
          6159 => x"70",
          6160 => x"c8",
          6161 => x"84",
          6162 => x"56",
          6163 => x"58",
          6164 => x"97",
          6165 => x"75",
          6166 => x"52",
          6167 => x"51",
          6168 => x"82",
          6169 => x"80",
          6170 => x"8a",
          6171 => x"32",
          6172 => x"72",
          6173 => x"2a",
          6174 => x"56",
          6175 => x"98",
          6176 => x"0d",
          6177 => x"0d",
          6178 => x"08",
          6179 => x"74",
          6180 => x"26",
          6181 => x"74",
          6182 => x"72",
          6183 => x"74",
          6184 => x"88",
          6185 => x"73",
          6186 => x"33",
          6187 => x"27",
          6188 => x"16",
          6189 => x"9b",
          6190 => x"2a",
          6191 => x"88",
          6192 => x"58",
          6193 => x"80",
          6194 => x"16",
          6195 => x"0c",
          6196 => x"8a",
          6197 => x"89",
          6198 => x"72",
          6199 => x"38",
          6200 => x"51",
          6201 => x"82",
          6202 => x"54",
          6203 => x"08",
          6204 => x"38",
          6205 => x"bb",
          6206 => x"8b",
          6207 => x"08",
          6208 => x"08",
          6209 => x"82",
          6210 => x"74",
          6211 => x"cb",
          6212 => x"75",
          6213 => x"3f",
          6214 => x"08",
          6215 => x"73",
          6216 => x"98",
          6217 => x"82",
          6218 => x"2e",
          6219 => x"39",
          6220 => x"39",
          6221 => x"13",
          6222 => x"74",
          6223 => x"16",
          6224 => x"18",
          6225 => x"77",
          6226 => x"0c",
          6227 => x"04",
          6228 => x"7a",
          6229 => x"12",
          6230 => x"59",
          6231 => x"80",
          6232 => x"86",
          6233 => x"98",
          6234 => x"14",
          6235 => x"55",
          6236 => x"81",
          6237 => x"83",
          6238 => x"77",
          6239 => x"81",
          6240 => x"0c",
          6241 => x"55",
          6242 => x"76",
          6243 => x"17",
          6244 => x"74",
          6245 => x"9b",
          6246 => x"39",
          6247 => x"ff",
          6248 => x"2a",
          6249 => x"81",
          6250 => x"52",
          6251 => x"e6",
          6252 => x"98",
          6253 => x"55",
          6254 => x"bb",
          6255 => x"80",
          6256 => x"55",
          6257 => x"08",
          6258 => x"f4",
          6259 => x"08",
          6260 => x"08",
          6261 => x"38",
          6262 => x"77",
          6263 => x"84",
          6264 => x"39",
          6265 => x"52",
          6266 => x"86",
          6267 => x"98",
          6268 => x"55",
          6269 => x"08",
          6270 => x"c4",
          6271 => x"82",
          6272 => x"81",
          6273 => x"81",
          6274 => x"98",
          6275 => x"b0",
          6276 => x"98",
          6277 => x"51",
          6278 => x"82",
          6279 => x"a0",
          6280 => x"15",
          6281 => x"75",
          6282 => x"3f",
          6283 => x"08",
          6284 => x"76",
          6285 => x"77",
          6286 => x"9c",
          6287 => x"55",
          6288 => x"98",
          6289 => x"0d",
          6290 => x"0d",
          6291 => x"08",
          6292 => x"80",
          6293 => x"fc",
          6294 => x"bb",
          6295 => x"82",
          6296 => x"80",
          6297 => x"bb",
          6298 => x"98",
          6299 => x"78",
          6300 => x"3f",
          6301 => x"08",
          6302 => x"98",
          6303 => x"38",
          6304 => x"08",
          6305 => x"70",
          6306 => x"58",
          6307 => x"2e",
          6308 => x"83",
          6309 => x"82",
          6310 => x"55",
          6311 => x"81",
          6312 => x"07",
          6313 => x"2e",
          6314 => x"16",
          6315 => x"2e",
          6316 => x"88",
          6317 => x"82",
          6318 => x"56",
          6319 => x"51",
          6320 => x"82",
          6321 => x"54",
          6322 => x"08",
          6323 => x"9b",
          6324 => x"2e",
          6325 => x"83",
          6326 => x"73",
          6327 => x"0c",
          6328 => x"04",
          6329 => x"76",
          6330 => x"54",
          6331 => x"82",
          6332 => x"83",
          6333 => x"76",
          6334 => x"53",
          6335 => x"2e",
          6336 => x"90",
          6337 => x"51",
          6338 => x"82",
          6339 => x"90",
          6340 => x"53",
          6341 => x"98",
          6342 => x"0d",
          6343 => x"0d",
          6344 => x"83",
          6345 => x"54",
          6346 => x"55",
          6347 => x"3f",
          6348 => x"51",
          6349 => x"2e",
          6350 => x"8b",
          6351 => x"2a",
          6352 => x"51",
          6353 => x"86",
          6354 => x"f7",
          6355 => x"7d",
          6356 => x"75",
          6357 => x"98",
          6358 => x"2e",
          6359 => x"98",
          6360 => x"78",
          6361 => x"3f",
          6362 => x"08",
          6363 => x"98",
          6364 => x"38",
          6365 => x"70",
          6366 => x"73",
          6367 => x"58",
          6368 => x"8b",
          6369 => x"bf",
          6370 => x"ff",
          6371 => x"53",
          6372 => x"34",
          6373 => x"08",
          6374 => x"e5",
          6375 => x"81",
          6376 => x"2e",
          6377 => x"70",
          6378 => x"57",
          6379 => x"9e",
          6380 => x"2e",
          6381 => x"bb",
          6382 => x"df",
          6383 => x"72",
          6384 => x"81",
          6385 => x"76",
          6386 => x"2e",
          6387 => x"52",
          6388 => x"fc",
          6389 => x"98",
          6390 => x"bb",
          6391 => x"38",
          6392 => x"fe",
          6393 => x"39",
          6394 => x"16",
          6395 => x"bb",
          6396 => x"3d",
          6397 => x"3d",
          6398 => x"08",
          6399 => x"52",
          6400 => x"c5",
          6401 => x"98",
          6402 => x"bb",
          6403 => x"38",
          6404 => x"52",
          6405 => x"de",
          6406 => x"98",
          6407 => x"bb",
          6408 => x"38",
          6409 => x"bb",
          6410 => x"9c",
          6411 => x"ea",
          6412 => x"53",
          6413 => x"9c",
          6414 => x"ea",
          6415 => x"0b",
          6416 => x"74",
          6417 => x"0c",
          6418 => x"04",
          6419 => x"75",
          6420 => x"12",
          6421 => x"53",
          6422 => x"9a",
          6423 => x"98",
          6424 => x"9c",
          6425 => x"e5",
          6426 => x"0b",
          6427 => x"85",
          6428 => x"fa",
          6429 => x"7a",
          6430 => x"0b",
          6431 => x"98",
          6432 => x"2e",
          6433 => x"80",
          6434 => x"55",
          6435 => x"17",
          6436 => x"33",
          6437 => x"51",
          6438 => x"2e",
          6439 => x"85",
          6440 => x"06",
          6441 => x"e5",
          6442 => x"2e",
          6443 => x"8b",
          6444 => x"70",
          6445 => x"34",
          6446 => x"71",
          6447 => x"05",
          6448 => x"15",
          6449 => x"27",
          6450 => x"15",
          6451 => x"80",
          6452 => x"34",
          6453 => x"52",
          6454 => x"88",
          6455 => x"17",
          6456 => x"52",
          6457 => x"3f",
          6458 => x"08",
          6459 => x"12",
          6460 => x"3f",
          6461 => x"08",
          6462 => x"98",
          6463 => x"da",
          6464 => x"98",
          6465 => x"23",
          6466 => x"04",
          6467 => x"7f",
          6468 => x"5b",
          6469 => x"33",
          6470 => x"73",
          6471 => x"38",
          6472 => x"80",
          6473 => x"38",
          6474 => x"8c",
          6475 => x"08",
          6476 => x"aa",
          6477 => x"41",
          6478 => x"33",
          6479 => x"73",
          6480 => x"81",
          6481 => x"81",
          6482 => x"dc",
          6483 => x"70",
          6484 => x"07",
          6485 => x"73",
          6486 => x"88",
          6487 => x"70",
          6488 => x"73",
          6489 => x"38",
          6490 => x"ab",
          6491 => x"52",
          6492 => x"91",
          6493 => x"98",
          6494 => x"98",
          6495 => x"61",
          6496 => x"5a",
          6497 => x"a0",
          6498 => x"e7",
          6499 => x"70",
          6500 => x"79",
          6501 => x"73",
          6502 => x"81",
          6503 => x"38",
          6504 => x"33",
          6505 => x"ae",
          6506 => x"70",
          6507 => x"82",
          6508 => x"51",
          6509 => x"54",
          6510 => x"79",
          6511 => x"74",
          6512 => x"57",
          6513 => x"af",
          6514 => x"70",
          6515 => x"51",
          6516 => x"dc",
          6517 => x"73",
          6518 => x"38",
          6519 => x"82",
          6520 => x"19",
          6521 => x"54",
          6522 => x"82",
          6523 => x"54",
          6524 => x"78",
          6525 => x"81",
          6526 => x"54",
          6527 => x"81",
          6528 => x"af",
          6529 => x"77",
          6530 => x"70",
          6531 => x"25",
          6532 => x"07",
          6533 => x"51",
          6534 => x"2e",
          6535 => x"39",
          6536 => x"80",
          6537 => x"33",
          6538 => x"73",
          6539 => x"81",
          6540 => x"81",
          6541 => x"dc",
          6542 => x"70",
          6543 => x"07",
          6544 => x"73",
          6545 => x"b5",
          6546 => x"2e",
          6547 => x"83",
          6548 => x"76",
          6549 => x"07",
          6550 => x"2e",
          6551 => x"8b",
          6552 => x"77",
          6553 => x"30",
          6554 => x"71",
          6555 => x"53",
          6556 => x"55",
          6557 => x"38",
          6558 => x"5c",
          6559 => x"75",
          6560 => x"73",
          6561 => x"38",
          6562 => x"06",
          6563 => x"11",
          6564 => x"75",
          6565 => x"3f",
          6566 => x"08",
          6567 => x"38",
          6568 => x"33",
          6569 => x"54",
          6570 => x"e6",
          6571 => x"bb",
          6572 => x"2e",
          6573 => x"ff",
          6574 => x"74",
          6575 => x"38",
          6576 => x"75",
          6577 => x"17",
          6578 => x"57",
          6579 => x"a7",
          6580 => x"82",
          6581 => x"e5",
          6582 => x"bb",
          6583 => x"38",
          6584 => x"54",
          6585 => x"89",
          6586 => x"70",
          6587 => x"57",
          6588 => x"54",
          6589 => x"81",
          6590 => x"f7",
          6591 => x"7e",
          6592 => x"2e",
          6593 => x"33",
          6594 => x"e5",
          6595 => x"06",
          6596 => x"7a",
          6597 => x"a0",
          6598 => x"38",
          6599 => x"55",
          6600 => x"84",
          6601 => x"39",
          6602 => x"8b",
          6603 => x"7b",
          6604 => x"7a",
          6605 => x"3f",
          6606 => x"08",
          6607 => x"98",
          6608 => x"38",
          6609 => x"52",
          6610 => x"aa",
          6611 => x"98",
          6612 => x"bb",
          6613 => x"c2",
          6614 => x"08",
          6615 => x"55",
          6616 => x"ff",
          6617 => x"15",
          6618 => x"54",
          6619 => x"34",
          6620 => x"70",
          6621 => x"81",
          6622 => x"58",
          6623 => x"8b",
          6624 => x"74",
          6625 => x"3f",
          6626 => x"08",
          6627 => x"38",
          6628 => x"51",
          6629 => x"ff",
          6630 => x"ab",
          6631 => x"55",
          6632 => x"bb",
          6633 => x"2e",
          6634 => x"80",
          6635 => x"85",
          6636 => x"06",
          6637 => x"58",
          6638 => x"80",
          6639 => x"75",
          6640 => x"73",
          6641 => x"b5",
          6642 => x"0b",
          6643 => x"80",
          6644 => x"39",
          6645 => x"54",
          6646 => x"85",
          6647 => x"75",
          6648 => x"81",
          6649 => x"73",
          6650 => x"1b",
          6651 => x"2a",
          6652 => x"51",
          6653 => x"80",
          6654 => x"90",
          6655 => x"ff",
          6656 => x"05",
          6657 => x"f5",
          6658 => x"bb",
          6659 => x"1c",
          6660 => x"39",
          6661 => x"98",
          6662 => x"0d",
          6663 => x"0d",
          6664 => x"7b",
          6665 => x"73",
          6666 => x"55",
          6667 => x"2e",
          6668 => x"75",
          6669 => x"57",
          6670 => x"26",
          6671 => x"ba",
          6672 => x"70",
          6673 => x"ba",
          6674 => x"06",
          6675 => x"73",
          6676 => x"70",
          6677 => x"51",
          6678 => x"89",
          6679 => x"82",
          6680 => x"ff",
          6681 => x"56",
          6682 => x"2e",
          6683 => x"80",
          6684 => x"d0",
          6685 => x"08",
          6686 => x"76",
          6687 => x"58",
          6688 => x"81",
          6689 => x"ff",
          6690 => x"53",
          6691 => x"26",
          6692 => x"13",
          6693 => x"06",
          6694 => x"9f",
          6695 => x"99",
          6696 => x"e0",
          6697 => x"ff",
          6698 => x"72",
          6699 => x"2a",
          6700 => x"72",
          6701 => x"06",
          6702 => x"ff",
          6703 => x"30",
          6704 => x"70",
          6705 => x"07",
          6706 => x"9f",
          6707 => x"54",
          6708 => x"80",
          6709 => x"81",
          6710 => x"59",
          6711 => x"25",
          6712 => x"8b",
          6713 => x"24",
          6714 => x"76",
          6715 => x"78",
          6716 => x"82",
          6717 => x"51",
          6718 => x"98",
          6719 => x"0d",
          6720 => x"0d",
          6721 => x"0b",
          6722 => x"ff",
          6723 => x"0c",
          6724 => x"51",
          6725 => x"84",
          6726 => x"98",
          6727 => x"38",
          6728 => x"51",
          6729 => x"82",
          6730 => x"83",
          6731 => x"54",
          6732 => x"82",
          6733 => x"09",
          6734 => x"e3",
          6735 => x"b4",
          6736 => x"57",
          6737 => x"2e",
          6738 => x"83",
          6739 => x"74",
          6740 => x"70",
          6741 => x"25",
          6742 => x"51",
          6743 => x"38",
          6744 => x"2e",
          6745 => x"b5",
          6746 => x"82",
          6747 => x"80",
          6748 => x"e0",
          6749 => x"bb",
          6750 => x"82",
          6751 => x"80",
          6752 => x"85",
          6753 => x"94",
          6754 => x"16",
          6755 => x"3f",
          6756 => x"08",
          6757 => x"98",
          6758 => x"83",
          6759 => x"74",
          6760 => x"0c",
          6761 => x"04",
          6762 => x"61",
          6763 => x"80",
          6764 => x"58",
          6765 => x"0c",
          6766 => x"e1",
          6767 => x"98",
          6768 => x"56",
          6769 => x"bb",
          6770 => x"86",
          6771 => x"bb",
          6772 => x"29",
          6773 => x"05",
          6774 => x"53",
          6775 => x"80",
          6776 => x"38",
          6777 => x"76",
          6778 => x"74",
          6779 => x"72",
          6780 => x"38",
          6781 => x"51",
          6782 => x"82",
          6783 => x"81",
          6784 => x"81",
          6785 => x"72",
          6786 => x"80",
          6787 => x"38",
          6788 => x"70",
          6789 => x"53",
          6790 => x"86",
          6791 => x"a7",
          6792 => x"34",
          6793 => x"34",
          6794 => x"14",
          6795 => x"b2",
          6796 => x"98",
          6797 => x"06",
          6798 => x"54",
          6799 => x"72",
          6800 => x"76",
          6801 => x"38",
          6802 => x"70",
          6803 => x"53",
          6804 => x"85",
          6805 => x"70",
          6806 => x"5b",
          6807 => x"82",
          6808 => x"81",
          6809 => x"76",
          6810 => x"81",
          6811 => x"38",
          6812 => x"56",
          6813 => x"83",
          6814 => x"70",
          6815 => x"80",
          6816 => x"83",
          6817 => x"dc",
          6818 => x"bb",
          6819 => x"76",
          6820 => x"05",
          6821 => x"16",
          6822 => x"56",
          6823 => x"d7",
          6824 => x"8d",
          6825 => x"72",
          6826 => x"54",
          6827 => x"57",
          6828 => x"95",
          6829 => x"73",
          6830 => x"3f",
          6831 => x"08",
          6832 => x"57",
          6833 => x"89",
          6834 => x"56",
          6835 => x"d7",
          6836 => x"76",
          6837 => x"f1",
          6838 => x"76",
          6839 => x"e9",
          6840 => x"51",
          6841 => x"82",
          6842 => x"83",
          6843 => x"53",
          6844 => x"2e",
          6845 => x"84",
          6846 => x"ca",
          6847 => x"da",
          6848 => x"98",
          6849 => x"ff",
          6850 => x"8d",
          6851 => x"14",
          6852 => x"3f",
          6853 => x"08",
          6854 => x"15",
          6855 => x"14",
          6856 => x"34",
          6857 => x"33",
          6858 => x"81",
          6859 => x"54",
          6860 => x"72",
          6861 => x"91",
          6862 => x"ff",
          6863 => x"29",
          6864 => x"33",
          6865 => x"72",
          6866 => x"72",
          6867 => x"38",
          6868 => x"06",
          6869 => x"2e",
          6870 => x"56",
          6871 => x"80",
          6872 => x"da",
          6873 => x"bb",
          6874 => x"82",
          6875 => x"88",
          6876 => x"8f",
          6877 => x"56",
          6878 => x"38",
          6879 => x"51",
          6880 => x"82",
          6881 => x"83",
          6882 => x"55",
          6883 => x"80",
          6884 => x"da",
          6885 => x"bb",
          6886 => x"80",
          6887 => x"da",
          6888 => x"bb",
          6889 => x"ff",
          6890 => x"8d",
          6891 => x"2e",
          6892 => x"88",
          6893 => x"14",
          6894 => x"05",
          6895 => x"75",
          6896 => x"38",
          6897 => x"52",
          6898 => x"51",
          6899 => x"3f",
          6900 => x"08",
          6901 => x"98",
          6902 => x"82",
          6903 => x"bb",
          6904 => x"ff",
          6905 => x"26",
          6906 => x"57",
          6907 => x"f5",
          6908 => x"82",
          6909 => x"f5",
          6910 => x"81",
          6911 => x"8d",
          6912 => x"2e",
          6913 => x"82",
          6914 => x"16",
          6915 => x"16",
          6916 => x"70",
          6917 => x"7a",
          6918 => x"0c",
          6919 => x"83",
          6920 => x"06",
          6921 => x"de",
          6922 => x"ae",
          6923 => x"98",
          6924 => x"ff",
          6925 => x"56",
          6926 => x"38",
          6927 => x"38",
          6928 => x"51",
          6929 => x"82",
          6930 => x"a8",
          6931 => x"82",
          6932 => x"39",
          6933 => x"80",
          6934 => x"38",
          6935 => x"15",
          6936 => x"53",
          6937 => x"8d",
          6938 => x"15",
          6939 => x"76",
          6940 => x"51",
          6941 => x"13",
          6942 => x"8d",
          6943 => x"15",
          6944 => x"c5",
          6945 => x"90",
          6946 => x"0b",
          6947 => x"ff",
          6948 => x"15",
          6949 => x"2e",
          6950 => x"81",
          6951 => x"e4",
          6952 => x"b6",
          6953 => x"98",
          6954 => x"ff",
          6955 => x"81",
          6956 => x"06",
          6957 => x"81",
          6958 => x"51",
          6959 => x"82",
          6960 => x"80",
          6961 => x"bb",
          6962 => x"15",
          6963 => x"14",
          6964 => x"3f",
          6965 => x"08",
          6966 => x"06",
          6967 => x"d4",
          6968 => x"81",
          6969 => x"38",
          6970 => x"d8",
          6971 => x"bb",
          6972 => x"8b",
          6973 => x"2e",
          6974 => x"b3",
          6975 => x"14",
          6976 => x"3f",
          6977 => x"08",
          6978 => x"e4",
          6979 => x"81",
          6980 => x"84",
          6981 => x"d7",
          6982 => x"bb",
          6983 => x"15",
          6984 => x"14",
          6985 => x"3f",
          6986 => x"08",
          6987 => x"76",
          6988 => x"d2",
          6989 => x"05",
          6990 => x"d2",
          6991 => x"86",
          6992 => x"0b",
          6993 => x"80",
          6994 => x"bb",
          6995 => x"3d",
          6996 => x"3d",
          6997 => x"89",
          6998 => x"2e",
          6999 => x"08",
          7000 => x"2e",
          7001 => x"33",
          7002 => x"2e",
          7003 => x"13",
          7004 => x"22",
          7005 => x"76",
          7006 => x"06",
          7007 => x"13",
          7008 => x"c0",
          7009 => x"98",
          7010 => x"52",
          7011 => x"71",
          7012 => x"55",
          7013 => x"53",
          7014 => x"0c",
          7015 => x"bb",
          7016 => x"3d",
          7017 => x"3d",
          7018 => x"05",
          7019 => x"89",
          7020 => x"52",
          7021 => x"3f",
          7022 => x"0b",
          7023 => x"08",
          7024 => x"82",
          7025 => x"84",
          7026 => x"d0",
          7027 => x"55",
          7028 => x"2e",
          7029 => x"74",
          7030 => x"73",
          7031 => x"38",
          7032 => x"78",
          7033 => x"54",
          7034 => x"92",
          7035 => x"89",
          7036 => x"84",
          7037 => x"b0",
          7038 => x"98",
          7039 => x"82",
          7040 => x"88",
          7041 => x"eb",
          7042 => x"02",
          7043 => x"e7",
          7044 => x"59",
          7045 => x"80",
          7046 => x"38",
          7047 => x"70",
          7048 => x"d0",
          7049 => x"3d",
          7050 => x"58",
          7051 => x"82",
          7052 => x"55",
          7053 => x"08",
          7054 => x"7a",
          7055 => x"8c",
          7056 => x"56",
          7057 => x"82",
          7058 => x"55",
          7059 => x"08",
          7060 => x"80",
          7061 => x"70",
          7062 => x"57",
          7063 => x"83",
          7064 => x"77",
          7065 => x"73",
          7066 => x"ab",
          7067 => x"2e",
          7068 => x"84",
          7069 => x"06",
          7070 => x"51",
          7071 => x"82",
          7072 => x"55",
          7073 => x"b2",
          7074 => x"06",
          7075 => x"b8",
          7076 => x"2a",
          7077 => x"51",
          7078 => x"2e",
          7079 => x"55",
          7080 => x"77",
          7081 => x"74",
          7082 => x"77",
          7083 => x"81",
          7084 => x"73",
          7085 => x"af",
          7086 => x"7a",
          7087 => x"3f",
          7088 => x"08",
          7089 => x"b2",
          7090 => x"8e",
          7091 => x"ea",
          7092 => x"a0",
          7093 => x"34",
          7094 => x"52",
          7095 => x"bd",
          7096 => x"62",
          7097 => x"d4",
          7098 => x"54",
          7099 => x"15",
          7100 => x"2e",
          7101 => x"7a",
          7102 => x"51",
          7103 => x"75",
          7104 => x"d4",
          7105 => x"be",
          7106 => x"98",
          7107 => x"bb",
          7108 => x"ca",
          7109 => x"74",
          7110 => x"02",
          7111 => x"70",
          7112 => x"81",
          7113 => x"56",
          7114 => x"86",
          7115 => x"82",
          7116 => x"81",
          7117 => x"06",
          7118 => x"80",
          7119 => x"75",
          7120 => x"73",
          7121 => x"38",
          7122 => x"92",
          7123 => x"7a",
          7124 => x"3f",
          7125 => x"08",
          7126 => x"8c",
          7127 => x"55",
          7128 => x"08",
          7129 => x"77",
          7130 => x"81",
          7131 => x"73",
          7132 => x"38",
          7133 => x"07",
          7134 => x"11",
          7135 => x"0c",
          7136 => x"0c",
          7137 => x"52",
          7138 => x"3f",
          7139 => x"08",
          7140 => x"08",
          7141 => x"63",
          7142 => x"5a",
          7143 => x"82",
          7144 => x"82",
          7145 => x"8c",
          7146 => x"7a",
          7147 => x"17",
          7148 => x"23",
          7149 => x"34",
          7150 => x"1a",
          7151 => x"9c",
          7152 => x"0b",
          7153 => x"77",
          7154 => x"81",
          7155 => x"73",
          7156 => x"8d",
          7157 => x"98",
          7158 => x"81",
          7159 => x"bb",
          7160 => x"1a",
          7161 => x"22",
          7162 => x"7b",
          7163 => x"a8",
          7164 => x"78",
          7165 => x"3f",
          7166 => x"08",
          7167 => x"98",
          7168 => x"83",
          7169 => x"82",
          7170 => x"ff",
          7171 => x"06",
          7172 => x"55",
          7173 => x"56",
          7174 => x"76",
          7175 => x"51",
          7176 => x"27",
          7177 => x"70",
          7178 => x"5a",
          7179 => x"76",
          7180 => x"74",
          7181 => x"83",
          7182 => x"73",
          7183 => x"38",
          7184 => x"51",
          7185 => x"82",
          7186 => x"85",
          7187 => x"8e",
          7188 => x"2a",
          7189 => x"08",
          7190 => x"0c",
          7191 => x"79",
          7192 => x"73",
          7193 => x"0c",
          7194 => x"04",
          7195 => x"60",
          7196 => x"40",
          7197 => x"80",
          7198 => x"3d",
          7199 => x"78",
          7200 => x"3f",
          7201 => x"08",
          7202 => x"98",
          7203 => x"91",
          7204 => x"74",
          7205 => x"38",
          7206 => x"c4",
          7207 => x"33",
          7208 => x"87",
          7209 => x"2e",
          7210 => x"95",
          7211 => x"91",
          7212 => x"56",
          7213 => x"81",
          7214 => x"34",
          7215 => x"a0",
          7216 => x"08",
          7217 => x"31",
          7218 => x"27",
          7219 => x"5c",
          7220 => x"82",
          7221 => x"19",
          7222 => x"ff",
          7223 => x"74",
          7224 => x"7e",
          7225 => x"ff",
          7226 => x"2a",
          7227 => x"79",
          7228 => x"87",
          7229 => x"08",
          7230 => x"98",
          7231 => x"78",
          7232 => x"3f",
          7233 => x"08",
          7234 => x"27",
          7235 => x"74",
          7236 => x"a3",
          7237 => x"1a",
          7238 => x"08",
          7239 => x"d4",
          7240 => x"bb",
          7241 => x"2e",
          7242 => x"82",
          7243 => x"1a",
          7244 => x"59",
          7245 => x"2e",
          7246 => x"77",
          7247 => x"11",
          7248 => x"55",
          7249 => x"85",
          7250 => x"31",
          7251 => x"76",
          7252 => x"81",
          7253 => x"ca",
          7254 => x"bb",
          7255 => x"d7",
          7256 => x"11",
          7257 => x"74",
          7258 => x"38",
          7259 => x"77",
          7260 => x"78",
          7261 => x"84",
          7262 => x"16",
          7263 => x"08",
          7264 => x"2b",
          7265 => x"cf",
          7266 => x"89",
          7267 => x"39",
          7268 => x"0c",
          7269 => x"83",
          7270 => x"80",
          7271 => x"55",
          7272 => x"83",
          7273 => x"9c",
          7274 => x"7e",
          7275 => x"3f",
          7276 => x"08",
          7277 => x"75",
          7278 => x"08",
          7279 => x"1f",
          7280 => x"7c",
          7281 => x"3f",
          7282 => x"7e",
          7283 => x"0c",
          7284 => x"1b",
          7285 => x"1c",
          7286 => x"fd",
          7287 => x"56",
          7288 => x"98",
          7289 => x"0d",
          7290 => x"0d",
          7291 => x"64",
          7292 => x"58",
          7293 => x"90",
          7294 => x"52",
          7295 => x"d2",
          7296 => x"98",
          7297 => x"bb",
          7298 => x"38",
          7299 => x"55",
          7300 => x"86",
          7301 => x"83",
          7302 => x"18",
          7303 => x"2a",
          7304 => x"51",
          7305 => x"56",
          7306 => x"83",
          7307 => x"39",
          7308 => x"19",
          7309 => x"83",
          7310 => x"0b",
          7311 => x"81",
          7312 => x"39",
          7313 => x"7c",
          7314 => x"74",
          7315 => x"38",
          7316 => x"7b",
          7317 => x"ec",
          7318 => x"08",
          7319 => x"06",
          7320 => x"81",
          7321 => x"8a",
          7322 => x"05",
          7323 => x"06",
          7324 => x"bf",
          7325 => x"38",
          7326 => x"55",
          7327 => x"7a",
          7328 => x"98",
          7329 => x"77",
          7330 => x"3f",
          7331 => x"08",
          7332 => x"98",
          7333 => x"82",
          7334 => x"81",
          7335 => x"38",
          7336 => x"ff",
          7337 => x"98",
          7338 => x"18",
          7339 => x"74",
          7340 => x"7e",
          7341 => x"08",
          7342 => x"2e",
          7343 => x"8d",
          7344 => x"ce",
          7345 => x"bb",
          7346 => x"ee",
          7347 => x"08",
          7348 => x"d1",
          7349 => x"bb",
          7350 => x"2e",
          7351 => x"82",
          7352 => x"1b",
          7353 => x"5a",
          7354 => x"2e",
          7355 => x"78",
          7356 => x"11",
          7357 => x"55",
          7358 => x"85",
          7359 => x"31",
          7360 => x"76",
          7361 => x"81",
          7362 => x"c8",
          7363 => x"bb",
          7364 => x"a6",
          7365 => x"11",
          7366 => x"56",
          7367 => x"27",
          7368 => x"80",
          7369 => x"08",
          7370 => x"2b",
          7371 => x"b4",
          7372 => x"b5",
          7373 => x"80",
          7374 => x"34",
          7375 => x"56",
          7376 => x"8c",
          7377 => x"19",
          7378 => x"38",
          7379 => x"b6",
          7380 => x"98",
          7381 => x"38",
          7382 => x"12",
          7383 => x"9c",
          7384 => x"18",
          7385 => x"06",
          7386 => x"31",
          7387 => x"76",
          7388 => x"7b",
          7389 => x"08",
          7390 => x"cd",
          7391 => x"bb",
          7392 => x"b6",
          7393 => x"7c",
          7394 => x"08",
          7395 => x"1f",
          7396 => x"cb",
          7397 => x"55",
          7398 => x"16",
          7399 => x"31",
          7400 => x"7f",
          7401 => x"94",
          7402 => x"70",
          7403 => x"8c",
          7404 => x"58",
          7405 => x"76",
          7406 => x"75",
          7407 => x"19",
          7408 => x"39",
          7409 => x"80",
          7410 => x"74",
          7411 => x"80",
          7412 => x"bb",
          7413 => x"3d",
          7414 => x"3d",
          7415 => x"3d",
          7416 => x"70",
          7417 => x"ea",
          7418 => x"98",
          7419 => x"bb",
          7420 => x"fb",
          7421 => x"33",
          7422 => x"70",
          7423 => x"55",
          7424 => x"2e",
          7425 => x"a0",
          7426 => x"78",
          7427 => x"3f",
          7428 => x"08",
          7429 => x"98",
          7430 => x"38",
          7431 => x"8b",
          7432 => x"07",
          7433 => x"8b",
          7434 => x"16",
          7435 => x"52",
          7436 => x"dd",
          7437 => x"16",
          7438 => x"15",
          7439 => x"3f",
          7440 => x"0a",
          7441 => x"51",
          7442 => x"76",
          7443 => x"51",
          7444 => x"78",
          7445 => x"83",
          7446 => x"51",
          7447 => x"82",
          7448 => x"90",
          7449 => x"bf",
          7450 => x"73",
          7451 => x"76",
          7452 => x"0c",
          7453 => x"04",
          7454 => x"76",
          7455 => x"fe",
          7456 => x"bb",
          7457 => x"82",
          7458 => x"9c",
          7459 => x"fc",
          7460 => x"51",
          7461 => x"82",
          7462 => x"53",
          7463 => x"08",
          7464 => x"bb",
          7465 => x"0c",
          7466 => x"98",
          7467 => x"0d",
          7468 => x"0d",
          7469 => x"e6",
          7470 => x"52",
          7471 => x"bb",
          7472 => x"8b",
          7473 => x"98",
          7474 => x"e4",
          7475 => x"71",
          7476 => x"0c",
          7477 => x"04",
          7478 => x"80",
          7479 => x"d0",
          7480 => x"3d",
          7481 => x"3f",
          7482 => x"08",
          7483 => x"98",
          7484 => x"38",
          7485 => x"52",
          7486 => x"05",
          7487 => x"3f",
          7488 => x"08",
          7489 => x"98",
          7490 => x"02",
          7491 => x"33",
          7492 => x"55",
          7493 => x"25",
          7494 => x"7a",
          7495 => x"54",
          7496 => x"a2",
          7497 => x"84",
          7498 => x"06",
          7499 => x"73",
          7500 => x"38",
          7501 => x"70",
          7502 => x"a8",
          7503 => x"98",
          7504 => x"0c",
          7505 => x"bb",
          7506 => x"2e",
          7507 => x"83",
          7508 => x"74",
          7509 => x"0c",
          7510 => x"04",
          7511 => x"6f",
          7512 => x"80",
          7513 => x"53",
          7514 => x"b8",
          7515 => x"3d",
          7516 => x"3f",
          7517 => x"08",
          7518 => x"98",
          7519 => x"38",
          7520 => x"7c",
          7521 => x"47",
          7522 => x"54",
          7523 => x"81",
          7524 => x"52",
          7525 => x"52",
          7526 => x"3f",
          7527 => x"08",
          7528 => x"98",
          7529 => x"38",
          7530 => x"51",
          7531 => x"82",
          7532 => x"57",
          7533 => x"08",
          7534 => x"69",
          7535 => x"da",
          7536 => x"bb",
          7537 => x"76",
          7538 => x"d5",
          7539 => x"bb",
          7540 => x"82",
          7541 => x"82",
          7542 => x"52",
          7543 => x"eb",
          7544 => x"98",
          7545 => x"bb",
          7546 => x"38",
          7547 => x"51",
          7548 => x"73",
          7549 => x"08",
          7550 => x"76",
          7551 => x"d6",
          7552 => x"bb",
          7553 => x"82",
          7554 => x"80",
          7555 => x"76",
          7556 => x"81",
          7557 => x"82",
          7558 => x"39",
          7559 => x"38",
          7560 => x"bc",
          7561 => x"51",
          7562 => x"76",
          7563 => x"11",
          7564 => x"51",
          7565 => x"73",
          7566 => x"38",
          7567 => x"55",
          7568 => x"16",
          7569 => x"56",
          7570 => x"38",
          7571 => x"73",
          7572 => x"90",
          7573 => x"2e",
          7574 => x"16",
          7575 => x"ff",
          7576 => x"ff",
          7577 => x"58",
          7578 => x"74",
          7579 => x"75",
          7580 => x"18",
          7581 => x"58",
          7582 => x"fe",
          7583 => x"7b",
          7584 => x"06",
          7585 => x"18",
          7586 => x"58",
          7587 => x"80",
          7588 => x"e4",
          7589 => x"29",
          7590 => x"05",
          7591 => x"33",
          7592 => x"56",
          7593 => x"2e",
          7594 => x"16",
          7595 => x"33",
          7596 => x"73",
          7597 => x"16",
          7598 => x"26",
          7599 => x"55",
          7600 => x"91",
          7601 => x"54",
          7602 => x"70",
          7603 => x"34",
          7604 => x"ec",
          7605 => x"70",
          7606 => x"34",
          7607 => x"09",
          7608 => x"38",
          7609 => x"39",
          7610 => x"19",
          7611 => x"33",
          7612 => x"05",
          7613 => x"78",
          7614 => x"80",
          7615 => x"82",
          7616 => x"9e",
          7617 => x"f7",
          7618 => x"7d",
          7619 => x"05",
          7620 => x"57",
          7621 => x"3f",
          7622 => x"08",
          7623 => x"98",
          7624 => x"38",
          7625 => x"53",
          7626 => x"38",
          7627 => x"54",
          7628 => x"92",
          7629 => x"33",
          7630 => x"70",
          7631 => x"54",
          7632 => x"38",
          7633 => x"15",
          7634 => x"70",
          7635 => x"58",
          7636 => x"82",
          7637 => x"8a",
          7638 => x"89",
          7639 => x"53",
          7640 => x"b7",
          7641 => x"ff",
          7642 => x"e3",
          7643 => x"bb",
          7644 => x"15",
          7645 => x"53",
          7646 => x"e3",
          7647 => x"bb",
          7648 => x"26",
          7649 => x"30",
          7650 => x"70",
          7651 => x"77",
          7652 => x"18",
          7653 => x"51",
          7654 => x"88",
          7655 => x"73",
          7656 => x"52",
          7657 => x"ca",
          7658 => x"98",
          7659 => x"bb",
          7660 => x"2e",
          7661 => x"82",
          7662 => x"ff",
          7663 => x"38",
          7664 => x"08",
          7665 => x"73",
          7666 => x"73",
          7667 => x"9c",
          7668 => x"27",
          7669 => x"75",
          7670 => x"16",
          7671 => x"17",
          7672 => x"33",
          7673 => x"70",
          7674 => x"55",
          7675 => x"80",
          7676 => x"73",
          7677 => x"cc",
          7678 => x"bb",
          7679 => x"82",
          7680 => x"94",
          7681 => x"98",
          7682 => x"39",
          7683 => x"51",
          7684 => x"82",
          7685 => x"54",
          7686 => x"be",
          7687 => x"27",
          7688 => x"53",
          7689 => x"08",
          7690 => x"73",
          7691 => x"ff",
          7692 => x"15",
          7693 => x"16",
          7694 => x"ff",
          7695 => x"80",
          7696 => x"73",
          7697 => x"c6",
          7698 => x"bb",
          7699 => x"38",
          7700 => x"16",
          7701 => x"80",
          7702 => x"0b",
          7703 => x"81",
          7704 => x"75",
          7705 => x"bb",
          7706 => x"58",
          7707 => x"54",
          7708 => x"74",
          7709 => x"73",
          7710 => x"90",
          7711 => x"c0",
          7712 => x"90",
          7713 => x"83",
          7714 => x"72",
          7715 => x"38",
          7716 => x"08",
          7717 => x"77",
          7718 => x"80",
          7719 => x"bb",
          7720 => x"3d",
          7721 => x"3d",
          7722 => x"89",
          7723 => x"2e",
          7724 => x"80",
          7725 => x"fc",
          7726 => x"3d",
          7727 => x"e1",
          7728 => x"bb",
          7729 => x"82",
          7730 => x"80",
          7731 => x"76",
          7732 => x"75",
          7733 => x"3f",
          7734 => x"08",
          7735 => x"98",
          7736 => x"38",
          7737 => x"70",
          7738 => x"57",
          7739 => x"a2",
          7740 => x"33",
          7741 => x"70",
          7742 => x"55",
          7743 => x"2e",
          7744 => x"16",
          7745 => x"51",
          7746 => x"82",
          7747 => x"88",
          7748 => x"54",
          7749 => x"84",
          7750 => x"52",
          7751 => x"e5",
          7752 => x"98",
          7753 => x"84",
          7754 => x"06",
          7755 => x"55",
          7756 => x"80",
          7757 => x"80",
          7758 => x"54",
          7759 => x"98",
          7760 => x"0d",
          7761 => x"0d",
          7762 => x"fc",
          7763 => x"52",
          7764 => x"3f",
          7765 => x"08",
          7766 => x"bb",
          7767 => x"0c",
          7768 => x"04",
          7769 => x"77",
          7770 => x"fc",
          7771 => x"53",
          7772 => x"de",
          7773 => x"98",
          7774 => x"bb",
          7775 => x"df",
          7776 => x"38",
          7777 => x"08",
          7778 => x"cd",
          7779 => x"bb",
          7780 => x"80",
          7781 => x"bb",
          7782 => x"73",
          7783 => x"3f",
          7784 => x"08",
          7785 => x"98",
          7786 => x"09",
          7787 => x"38",
          7788 => x"39",
          7789 => x"08",
          7790 => x"52",
          7791 => x"b3",
          7792 => x"73",
          7793 => x"3f",
          7794 => x"08",
          7795 => x"30",
          7796 => x"9f",
          7797 => x"bb",
          7798 => x"51",
          7799 => x"72",
          7800 => x"0c",
          7801 => x"04",
          7802 => x"65",
          7803 => x"89",
          7804 => x"96",
          7805 => x"df",
          7806 => x"bb",
          7807 => x"82",
          7808 => x"b2",
          7809 => x"75",
          7810 => x"3f",
          7811 => x"08",
          7812 => x"98",
          7813 => x"02",
          7814 => x"33",
          7815 => x"55",
          7816 => x"25",
          7817 => x"55",
          7818 => x"80",
          7819 => x"76",
          7820 => x"d4",
          7821 => x"82",
          7822 => x"94",
          7823 => x"f0",
          7824 => x"65",
          7825 => x"53",
          7826 => x"05",
          7827 => x"51",
          7828 => x"82",
          7829 => x"5b",
          7830 => x"08",
          7831 => x"7c",
          7832 => x"08",
          7833 => x"fe",
          7834 => x"08",
          7835 => x"55",
          7836 => x"91",
          7837 => x"0c",
          7838 => x"81",
          7839 => x"39",
          7840 => x"c7",
          7841 => x"98",
          7842 => x"55",
          7843 => x"2e",
          7844 => x"bf",
          7845 => x"5f",
          7846 => x"92",
          7847 => x"51",
          7848 => x"82",
          7849 => x"ff",
          7850 => x"82",
          7851 => x"81",
          7852 => x"82",
          7853 => x"30",
          7854 => x"98",
          7855 => x"25",
          7856 => x"19",
          7857 => x"5a",
          7858 => x"08",
          7859 => x"38",
          7860 => x"a4",
          7861 => x"bb",
          7862 => x"58",
          7863 => x"77",
          7864 => x"7d",
          7865 => x"bf",
          7866 => x"bb",
          7867 => x"82",
          7868 => x"80",
          7869 => x"70",
          7870 => x"ff",
          7871 => x"56",
          7872 => x"2e",
          7873 => x"9e",
          7874 => x"51",
          7875 => x"3f",
          7876 => x"08",
          7877 => x"06",
          7878 => x"80",
          7879 => x"19",
          7880 => x"54",
          7881 => x"14",
          7882 => x"c5",
          7883 => x"98",
          7884 => x"06",
          7885 => x"80",
          7886 => x"19",
          7887 => x"54",
          7888 => x"06",
          7889 => x"79",
          7890 => x"78",
          7891 => x"79",
          7892 => x"84",
          7893 => x"07",
          7894 => x"84",
          7895 => x"82",
          7896 => x"92",
          7897 => x"f9",
          7898 => x"8a",
          7899 => x"53",
          7900 => x"e3",
          7901 => x"bb",
          7902 => x"82",
          7903 => x"81",
          7904 => x"17",
          7905 => x"81",
          7906 => x"17",
          7907 => x"2a",
          7908 => x"51",
          7909 => x"55",
          7910 => x"81",
          7911 => x"17",
          7912 => x"8c",
          7913 => x"81",
          7914 => x"9b",
          7915 => x"98",
          7916 => x"17",
          7917 => x"51",
          7918 => x"82",
          7919 => x"74",
          7920 => x"56",
          7921 => x"98",
          7922 => x"76",
          7923 => x"c6",
          7924 => x"98",
          7925 => x"09",
          7926 => x"38",
          7927 => x"bb",
          7928 => x"2e",
          7929 => x"85",
          7930 => x"a3",
          7931 => x"38",
          7932 => x"bb",
          7933 => x"15",
          7934 => x"38",
          7935 => x"53",
          7936 => x"08",
          7937 => x"c3",
          7938 => x"bb",
          7939 => x"94",
          7940 => x"18",
          7941 => x"33",
          7942 => x"54",
          7943 => x"34",
          7944 => x"85",
          7945 => x"18",
          7946 => x"74",
          7947 => x"0c",
          7948 => x"04",
          7949 => x"82",
          7950 => x"ff",
          7951 => x"a1",
          7952 => x"e4",
          7953 => x"98",
          7954 => x"bb",
          7955 => x"f5",
          7956 => x"a1",
          7957 => x"95",
          7958 => x"58",
          7959 => x"82",
          7960 => x"55",
          7961 => x"08",
          7962 => x"02",
          7963 => x"33",
          7964 => x"70",
          7965 => x"55",
          7966 => x"73",
          7967 => x"75",
          7968 => x"80",
          7969 => x"bd",
          7970 => x"d6",
          7971 => x"81",
          7972 => x"87",
          7973 => x"ad",
          7974 => x"78",
          7975 => x"3f",
          7976 => x"08",
          7977 => x"70",
          7978 => x"55",
          7979 => x"2e",
          7980 => x"78",
          7981 => x"98",
          7982 => x"08",
          7983 => x"38",
          7984 => x"bb",
          7985 => x"76",
          7986 => x"70",
          7987 => x"b5",
          7988 => x"98",
          7989 => x"bb",
          7990 => x"e9",
          7991 => x"98",
          7992 => x"51",
          7993 => x"82",
          7994 => x"55",
          7995 => x"08",
          7996 => x"55",
          7997 => x"82",
          7998 => x"84",
          7999 => x"82",
          8000 => x"80",
          8001 => x"51",
          8002 => x"82",
          8003 => x"82",
          8004 => x"30",
          8005 => x"98",
          8006 => x"25",
          8007 => x"75",
          8008 => x"38",
          8009 => x"8f",
          8010 => x"75",
          8011 => x"c1",
          8012 => x"bb",
          8013 => x"74",
          8014 => x"51",
          8015 => x"3f",
          8016 => x"08",
          8017 => x"bb",
          8018 => x"3d",
          8019 => x"3d",
          8020 => x"99",
          8021 => x"52",
          8022 => x"d8",
          8023 => x"bb",
          8024 => x"82",
          8025 => x"82",
          8026 => x"5e",
          8027 => x"3d",
          8028 => x"cf",
          8029 => x"bb",
          8030 => x"82",
          8031 => x"86",
          8032 => x"82",
          8033 => x"bb",
          8034 => x"2e",
          8035 => x"82",
          8036 => x"80",
          8037 => x"70",
          8038 => x"06",
          8039 => x"54",
          8040 => x"38",
          8041 => x"52",
          8042 => x"52",
          8043 => x"3f",
          8044 => x"08",
          8045 => x"82",
          8046 => x"83",
          8047 => x"82",
          8048 => x"81",
          8049 => x"06",
          8050 => x"54",
          8051 => x"08",
          8052 => x"81",
          8053 => x"81",
          8054 => x"39",
          8055 => x"38",
          8056 => x"08",
          8057 => x"c4",
          8058 => x"bb",
          8059 => x"82",
          8060 => x"81",
          8061 => x"53",
          8062 => x"19",
          8063 => x"8c",
          8064 => x"ae",
          8065 => x"34",
          8066 => x"0b",
          8067 => x"82",
          8068 => x"52",
          8069 => x"51",
          8070 => x"3f",
          8071 => x"b4",
          8072 => x"c9",
          8073 => x"53",
          8074 => x"53",
          8075 => x"51",
          8076 => x"3f",
          8077 => x"0b",
          8078 => x"34",
          8079 => x"80",
          8080 => x"51",
          8081 => x"78",
          8082 => x"83",
          8083 => x"51",
          8084 => x"82",
          8085 => x"54",
          8086 => x"08",
          8087 => x"88",
          8088 => x"64",
          8089 => x"ff",
          8090 => x"75",
          8091 => x"78",
          8092 => x"3f",
          8093 => x"0b",
          8094 => x"78",
          8095 => x"83",
          8096 => x"51",
          8097 => x"3f",
          8098 => x"08",
          8099 => x"80",
          8100 => x"76",
          8101 => x"ae",
          8102 => x"bb",
          8103 => x"3d",
          8104 => x"3d",
          8105 => x"84",
          8106 => x"f1",
          8107 => x"a8",
          8108 => x"05",
          8109 => x"51",
          8110 => x"82",
          8111 => x"55",
          8112 => x"08",
          8113 => x"78",
          8114 => x"08",
          8115 => x"70",
          8116 => x"b8",
          8117 => x"98",
          8118 => x"bb",
          8119 => x"b9",
          8120 => x"9b",
          8121 => x"a0",
          8122 => x"55",
          8123 => x"38",
          8124 => x"3d",
          8125 => x"3d",
          8126 => x"51",
          8127 => x"3f",
          8128 => x"52",
          8129 => x"52",
          8130 => x"dd",
          8131 => x"08",
          8132 => x"cb",
          8133 => x"bb",
          8134 => x"82",
          8135 => x"95",
          8136 => x"2e",
          8137 => x"88",
          8138 => x"3d",
          8139 => x"38",
          8140 => x"e5",
          8141 => x"98",
          8142 => x"09",
          8143 => x"b8",
          8144 => x"c9",
          8145 => x"bb",
          8146 => x"82",
          8147 => x"81",
          8148 => x"56",
          8149 => x"3d",
          8150 => x"52",
          8151 => x"ff",
          8152 => x"02",
          8153 => x"8b",
          8154 => x"16",
          8155 => x"2a",
          8156 => x"51",
          8157 => x"89",
          8158 => x"07",
          8159 => x"17",
          8160 => x"81",
          8161 => x"34",
          8162 => x"70",
          8163 => x"81",
          8164 => x"55",
          8165 => x"80",
          8166 => x"64",
          8167 => x"38",
          8168 => x"51",
          8169 => x"82",
          8170 => x"52",
          8171 => x"b7",
          8172 => x"55",
          8173 => x"08",
          8174 => x"dd",
          8175 => x"98",
          8176 => x"51",
          8177 => x"3f",
          8178 => x"08",
          8179 => x"11",
          8180 => x"82",
          8181 => x"80",
          8182 => x"16",
          8183 => x"ae",
          8184 => x"06",
          8185 => x"53",
          8186 => x"51",
          8187 => x"78",
          8188 => x"83",
          8189 => x"39",
          8190 => x"08",
          8191 => x"51",
          8192 => x"82",
          8193 => x"55",
          8194 => x"08",
          8195 => x"51",
          8196 => x"3f",
          8197 => x"08",
          8198 => x"bb",
          8199 => x"3d",
          8200 => x"3d",
          8201 => x"db",
          8202 => x"84",
          8203 => x"05",
          8204 => x"82",
          8205 => x"d0",
          8206 => x"3d",
          8207 => x"3f",
          8208 => x"08",
          8209 => x"98",
          8210 => x"38",
          8211 => x"52",
          8212 => x"05",
          8213 => x"3f",
          8214 => x"08",
          8215 => x"98",
          8216 => x"02",
          8217 => x"33",
          8218 => x"54",
          8219 => x"aa",
          8220 => x"06",
          8221 => x"8b",
          8222 => x"06",
          8223 => x"07",
          8224 => x"56",
          8225 => x"34",
          8226 => x"0b",
          8227 => x"78",
          8228 => x"a9",
          8229 => x"98",
          8230 => x"82",
          8231 => x"95",
          8232 => x"ef",
          8233 => x"56",
          8234 => x"3d",
          8235 => x"94",
          8236 => x"f4",
          8237 => x"98",
          8238 => x"bb",
          8239 => x"cb",
          8240 => x"63",
          8241 => x"d4",
          8242 => x"c0",
          8243 => x"98",
          8244 => x"bb",
          8245 => x"38",
          8246 => x"05",
          8247 => x"06",
          8248 => x"73",
          8249 => x"16",
          8250 => x"22",
          8251 => x"07",
          8252 => x"1f",
          8253 => x"c2",
          8254 => x"81",
          8255 => x"34",
          8256 => x"b3",
          8257 => x"bb",
          8258 => x"74",
          8259 => x"0c",
          8260 => x"04",
          8261 => x"69",
          8262 => x"80",
          8263 => x"d0",
          8264 => x"3d",
          8265 => x"3f",
          8266 => x"08",
          8267 => x"08",
          8268 => x"bb",
          8269 => x"80",
          8270 => x"57",
          8271 => x"81",
          8272 => x"70",
          8273 => x"55",
          8274 => x"80",
          8275 => x"5d",
          8276 => x"52",
          8277 => x"52",
          8278 => x"a9",
          8279 => x"98",
          8280 => x"bb",
          8281 => x"d1",
          8282 => x"73",
          8283 => x"3f",
          8284 => x"08",
          8285 => x"98",
          8286 => x"82",
          8287 => x"82",
          8288 => x"65",
          8289 => x"78",
          8290 => x"7b",
          8291 => x"55",
          8292 => x"34",
          8293 => x"8a",
          8294 => x"38",
          8295 => x"1a",
          8296 => x"34",
          8297 => x"9e",
          8298 => x"70",
          8299 => x"51",
          8300 => x"a0",
          8301 => x"8e",
          8302 => x"2e",
          8303 => x"86",
          8304 => x"34",
          8305 => x"30",
          8306 => x"80",
          8307 => x"7a",
          8308 => x"c1",
          8309 => x"2e",
          8310 => x"a0",
          8311 => x"51",
          8312 => x"3f",
          8313 => x"08",
          8314 => x"98",
          8315 => x"7b",
          8316 => x"55",
          8317 => x"73",
          8318 => x"38",
          8319 => x"73",
          8320 => x"38",
          8321 => x"15",
          8322 => x"ff",
          8323 => x"82",
          8324 => x"7b",
          8325 => x"bb",
          8326 => x"3d",
          8327 => x"3d",
          8328 => x"9c",
          8329 => x"05",
          8330 => x"51",
          8331 => x"82",
          8332 => x"82",
          8333 => x"56",
          8334 => x"98",
          8335 => x"38",
          8336 => x"52",
          8337 => x"52",
          8338 => x"c0",
          8339 => x"70",
          8340 => x"ff",
          8341 => x"55",
          8342 => x"27",
          8343 => x"78",
          8344 => x"ff",
          8345 => x"05",
          8346 => x"55",
          8347 => x"3f",
          8348 => x"08",
          8349 => x"38",
          8350 => x"70",
          8351 => x"ff",
          8352 => x"82",
          8353 => x"80",
          8354 => x"74",
          8355 => x"07",
          8356 => x"4e",
          8357 => x"82",
          8358 => x"55",
          8359 => x"70",
          8360 => x"06",
          8361 => x"99",
          8362 => x"e0",
          8363 => x"ff",
          8364 => x"54",
          8365 => x"27",
          8366 => x"b3",
          8367 => x"55",
          8368 => x"a3",
          8369 => x"82",
          8370 => x"ff",
          8371 => x"82",
          8372 => x"93",
          8373 => x"75",
          8374 => x"76",
          8375 => x"38",
          8376 => x"77",
          8377 => x"86",
          8378 => x"39",
          8379 => x"27",
          8380 => x"88",
          8381 => x"78",
          8382 => x"5a",
          8383 => x"57",
          8384 => x"81",
          8385 => x"81",
          8386 => x"33",
          8387 => x"06",
          8388 => x"57",
          8389 => x"fe",
          8390 => x"3d",
          8391 => x"55",
          8392 => x"2e",
          8393 => x"76",
          8394 => x"38",
          8395 => x"55",
          8396 => x"33",
          8397 => x"a0",
          8398 => x"06",
          8399 => x"17",
          8400 => x"38",
          8401 => x"43",
          8402 => x"3d",
          8403 => x"ff",
          8404 => x"82",
          8405 => x"54",
          8406 => x"08",
          8407 => x"81",
          8408 => x"ff",
          8409 => x"82",
          8410 => x"54",
          8411 => x"08",
          8412 => x"80",
          8413 => x"54",
          8414 => x"80",
          8415 => x"bb",
          8416 => x"2e",
          8417 => x"80",
          8418 => x"54",
          8419 => x"80",
          8420 => x"52",
          8421 => x"bd",
          8422 => x"bb",
          8423 => x"82",
          8424 => x"b1",
          8425 => x"82",
          8426 => x"52",
          8427 => x"ab",
          8428 => x"54",
          8429 => x"15",
          8430 => x"78",
          8431 => x"ff",
          8432 => x"79",
          8433 => x"83",
          8434 => x"51",
          8435 => x"3f",
          8436 => x"08",
          8437 => x"74",
          8438 => x"0c",
          8439 => x"04",
          8440 => x"60",
          8441 => x"05",
          8442 => x"33",
          8443 => x"05",
          8444 => x"40",
          8445 => x"da",
          8446 => x"98",
          8447 => x"bb",
          8448 => x"bd",
          8449 => x"33",
          8450 => x"b5",
          8451 => x"2e",
          8452 => x"1a",
          8453 => x"90",
          8454 => x"33",
          8455 => x"70",
          8456 => x"55",
          8457 => x"38",
          8458 => x"97",
          8459 => x"82",
          8460 => x"58",
          8461 => x"7e",
          8462 => x"70",
          8463 => x"55",
          8464 => x"56",
          8465 => x"de",
          8466 => x"7d",
          8467 => x"70",
          8468 => x"2a",
          8469 => x"08",
          8470 => x"08",
          8471 => x"5d",
          8472 => x"77",
          8473 => x"98",
          8474 => x"26",
          8475 => x"57",
          8476 => x"59",
          8477 => x"52",
          8478 => x"ae",
          8479 => x"15",
          8480 => x"98",
          8481 => x"26",
          8482 => x"55",
          8483 => x"08",
          8484 => x"99",
          8485 => x"98",
          8486 => x"ff",
          8487 => x"bb",
          8488 => x"38",
          8489 => x"75",
          8490 => x"81",
          8491 => x"93",
          8492 => x"80",
          8493 => x"2e",
          8494 => x"ff",
          8495 => x"58",
          8496 => x"7d",
          8497 => x"38",
          8498 => x"55",
          8499 => x"b4",
          8500 => x"56",
          8501 => x"09",
          8502 => x"38",
          8503 => x"53",
          8504 => x"51",
          8505 => x"3f",
          8506 => x"08",
          8507 => x"98",
          8508 => x"38",
          8509 => x"ff",
          8510 => x"5c",
          8511 => x"84",
          8512 => x"5c",
          8513 => x"12",
          8514 => x"80",
          8515 => x"78",
          8516 => x"7c",
          8517 => x"90",
          8518 => x"c0",
          8519 => x"90",
          8520 => x"15",
          8521 => x"90",
          8522 => x"54",
          8523 => x"91",
          8524 => x"31",
          8525 => x"84",
          8526 => x"07",
          8527 => x"16",
          8528 => x"73",
          8529 => x"0c",
          8530 => x"04",
          8531 => x"6b",
          8532 => x"05",
          8533 => x"33",
          8534 => x"5a",
          8535 => x"bd",
          8536 => x"80",
          8537 => x"98",
          8538 => x"f8",
          8539 => x"98",
          8540 => x"82",
          8541 => x"70",
          8542 => x"74",
          8543 => x"38",
          8544 => x"82",
          8545 => x"81",
          8546 => x"81",
          8547 => x"ff",
          8548 => x"82",
          8549 => x"81",
          8550 => x"81",
          8551 => x"83",
          8552 => x"c0",
          8553 => x"2a",
          8554 => x"51",
          8555 => x"74",
          8556 => x"99",
          8557 => x"53",
          8558 => x"51",
          8559 => x"3f",
          8560 => x"08",
          8561 => x"55",
          8562 => x"92",
          8563 => x"80",
          8564 => x"38",
          8565 => x"06",
          8566 => x"2e",
          8567 => x"48",
          8568 => x"87",
          8569 => x"79",
          8570 => x"78",
          8571 => x"26",
          8572 => x"19",
          8573 => x"74",
          8574 => x"38",
          8575 => x"e4",
          8576 => x"2a",
          8577 => x"70",
          8578 => x"59",
          8579 => x"7a",
          8580 => x"56",
          8581 => x"80",
          8582 => x"51",
          8583 => x"74",
          8584 => x"99",
          8585 => x"53",
          8586 => x"51",
          8587 => x"3f",
          8588 => x"bb",
          8589 => x"ac",
          8590 => x"2a",
          8591 => x"82",
          8592 => x"43",
          8593 => x"83",
          8594 => x"66",
          8595 => x"60",
          8596 => x"90",
          8597 => x"31",
          8598 => x"80",
          8599 => x"8a",
          8600 => x"56",
          8601 => x"26",
          8602 => x"77",
          8603 => x"81",
          8604 => x"74",
          8605 => x"38",
          8606 => x"55",
          8607 => x"83",
          8608 => x"81",
          8609 => x"80",
          8610 => x"38",
          8611 => x"55",
          8612 => x"5e",
          8613 => x"89",
          8614 => x"5a",
          8615 => x"09",
          8616 => x"e1",
          8617 => x"38",
          8618 => x"57",
          8619 => x"b6",
          8620 => x"5a",
          8621 => x"9d",
          8622 => x"26",
          8623 => x"b6",
          8624 => x"10",
          8625 => x"22",
          8626 => x"74",
          8627 => x"38",
          8628 => x"ee",
          8629 => x"66",
          8630 => x"ca",
          8631 => x"98",
          8632 => x"84",
          8633 => x"89",
          8634 => x"a0",
          8635 => x"82",
          8636 => x"fc",
          8637 => x"56",
          8638 => x"f0",
          8639 => x"80",
          8640 => x"d3",
          8641 => x"38",
          8642 => x"57",
          8643 => x"b5",
          8644 => x"5a",
          8645 => x"9d",
          8646 => x"26",
          8647 => x"b5",
          8648 => x"10",
          8649 => x"22",
          8650 => x"74",
          8651 => x"38",
          8652 => x"ee",
          8653 => x"66",
          8654 => x"ea",
          8655 => x"98",
          8656 => x"05",
          8657 => x"98",
          8658 => x"26",
          8659 => x"0b",
          8660 => x"08",
          8661 => x"98",
          8662 => x"11",
          8663 => x"05",
          8664 => x"83",
          8665 => x"2a",
          8666 => x"a0",
          8667 => x"7d",
          8668 => x"69",
          8669 => x"05",
          8670 => x"72",
          8671 => x"5c",
          8672 => x"59",
          8673 => x"2e",
          8674 => x"89",
          8675 => x"60",
          8676 => x"84",
          8677 => x"5d",
          8678 => x"18",
          8679 => x"68",
          8680 => x"74",
          8681 => x"af",
          8682 => x"31",
          8683 => x"53",
          8684 => x"52",
          8685 => x"ee",
          8686 => x"98",
          8687 => x"83",
          8688 => x"06",
          8689 => x"bb",
          8690 => x"ff",
          8691 => x"dd",
          8692 => x"83",
          8693 => x"2a",
          8694 => x"be",
          8695 => x"39",
          8696 => x"09",
          8697 => x"c5",
          8698 => x"f5",
          8699 => x"98",
          8700 => x"38",
          8701 => x"79",
          8702 => x"80",
          8703 => x"38",
          8704 => x"96",
          8705 => x"06",
          8706 => x"2e",
          8707 => x"5e",
          8708 => x"82",
          8709 => x"9f",
          8710 => x"38",
          8711 => x"38",
          8712 => x"81",
          8713 => x"fc",
          8714 => x"ab",
          8715 => x"7d",
          8716 => x"81",
          8717 => x"7d",
          8718 => x"78",
          8719 => x"74",
          8720 => x"8e",
          8721 => x"9c",
          8722 => x"53",
          8723 => x"51",
          8724 => x"3f",
          8725 => x"b4",
          8726 => x"51",
          8727 => x"3f",
          8728 => x"8b",
          8729 => x"a1",
          8730 => x"8d",
          8731 => x"83",
          8732 => x"52",
          8733 => x"ff",
          8734 => x"81",
          8735 => x"34",
          8736 => x"70",
          8737 => x"2a",
          8738 => x"54",
          8739 => x"1b",
          8740 => x"88",
          8741 => x"74",
          8742 => x"26",
          8743 => x"83",
          8744 => x"52",
          8745 => x"ff",
          8746 => x"8a",
          8747 => x"a0",
          8748 => x"a1",
          8749 => x"0b",
          8750 => x"bf",
          8751 => x"51",
          8752 => x"3f",
          8753 => x"9a",
          8754 => x"a0",
          8755 => x"52",
          8756 => x"ff",
          8757 => x"7d",
          8758 => x"81",
          8759 => x"38",
          8760 => x"0a",
          8761 => x"1b",
          8762 => x"ce",
          8763 => x"a4",
          8764 => x"a0",
          8765 => x"52",
          8766 => x"ff",
          8767 => x"81",
          8768 => x"51",
          8769 => x"3f",
          8770 => x"1b",
          8771 => x"8c",
          8772 => x"0b",
          8773 => x"34",
          8774 => x"c2",
          8775 => x"53",
          8776 => x"52",
          8777 => x"51",
          8778 => x"88",
          8779 => x"a7",
          8780 => x"a0",
          8781 => x"83",
          8782 => x"52",
          8783 => x"ff",
          8784 => x"ff",
          8785 => x"1c",
          8786 => x"a6",
          8787 => x"53",
          8788 => x"52",
          8789 => x"ff",
          8790 => x"82",
          8791 => x"83",
          8792 => x"52",
          8793 => x"b4",
          8794 => x"60",
          8795 => x"7e",
          8796 => x"d7",
          8797 => x"82",
          8798 => x"83",
          8799 => x"83",
          8800 => x"06",
          8801 => x"75",
          8802 => x"05",
          8803 => x"7e",
          8804 => x"b7",
          8805 => x"53",
          8806 => x"51",
          8807 => x"3f",
          8808 => x"a4",
          8809 => x"51",
          8810 => x"3f",
          8811 => x"e4",
          8812 => x"e4",
          8813 => x"9f",
          8814 => x"18",
          8815 => x"1b",
          8816 => x"f6",
          8817 => x"83",
          8818 => x"ff",
          8819 => x"82",
          8820 => x"78",
          8821 => x"c4",
          8822 => x"60",
          8823 => x"7a",
          8824 => x"ff",
          8825 => x"75",
          8826 => x"53",
          8827 => x"51",
          8828 => x"3f",
          8829 => x"52",
          8830 => x"9f",
          8831 => x"56",
          8832 => x"83",
          8833 => x"06",
          8834 => x"52",
          8835 => x"9e",
          8836 => x"52",
          8837 => x"ff",
          8838 => x"f0",
          8839 => x"1b",
          8840 => x"87",
          8841 => x"55",
          8842 => x"83",
          8843 => x"74",
          8844 => x"ff",
          8845 => x"7c",
          8846 => x"74",
          8847 => x"38",
          8848 => x"54",
          8849 => x"52",
          8850 => x"99",
          8851 => x"bb",
          8852 => x"87",
          8853 => x"53",
          8854 => x"08",
          8855 => x"ff",
          8856 => x"76",
          8857 => x"31",
          8858 => x"cd",
          8859 => x"58",
          8860 => x"ff",
          8861 => x"55",
          8862 => x"83",
          8863 => x"61",
          8864 => x"26",
          8865 => x"57",
          8866 => x"53",
          8867 => x"51",
          8868 => x"3f",
          8869 => x"08",
          8870 => x"76",
          8871 => x"31",
          8872 => x"db",
          8873 => x"7d",
          8874 => x"38",
          8875 => x"83",
          8876 => x"8a",
          8877 => x"7d",
          8878 => x"38",
          8879 => x"81",
          8880 => x"80",
          8881 => x"80",
          8882 => x"7a",
          8883 => x"bc",
          8884 => x"d5",
          8885 => x"ff",
          8886 => x"83",
          8887 => x"77",
          8888 => x"0b",
          8889 => x"81",
          8890 => x"34",
          8891 => x"34",
          8892 => x"34",
          8893 => x"56",
          8894 => x"52",
          8895 => x"bc",
          8896 => x"0b",
          8897 => x"82",
          8898 => x"82",
          8899 => x"56",
          8900 => x"34",
          8901 => x"08",
          8902 => x"60",
          8903 => x"1b",
          8904 => x"96",
          8905 => x"83",
          8906 => x"ff",
          8907 => x"81",
          8908 => x"7a",
          8909 => x"ff",
          8910 => x"81",
          8911 => x"98",
          8912 => x"80",
          8913 => x"7e",
          8914 => x"e3",
          8915 => x"82",
          8916 => x"90",
          8917 => x"8e",
          8918 => x"81",
          8919 => x"82",
          8920 => x"56",
          8921 => x"98",
          8922 => x"0d",
          8923 => x"0d",
          8924 => x"59",
          8925 => x"ff",
          8926 => x"57",
          8927 => x"b4",
          8928 => x"f8",
          8929 => x"81",
          8930 => x"52",
          8931 => x"dc",
          8932 => x"2e",
          8933 => x"9c",
          8934 => x"33",
          8935 => x"2e",
          8936 => x"76",
          8937 => x"58",
          8938 => x"57",
          8939 => x"09",
          8940 => x"38",
          8941 => x"78",
          8942 => x"38",
          8943 => x"82",
          8944 => x"8d",
          8945 => x"f7",
          8946 => x"02",
          8947 => x"05",
          8948 => x"77",
          8949 => x"81",
          8950 => x"8d",
          8951 => x"e7",
          8952 => x"08",
          8953 => x"24",
          8954 => x"17",
          8955 => x"8c",
          8956 => x"77",
          8957 => x"16",
          8958 => x"25",
          8959 => x"3d",
          8960 => x"75",
          8961 => x"52",
          8962 => x"cb",
          8963 => x"76",
          8964 => x"70",
          8965 => x"2a",
          8966 => x"51",
          8967 => x"84",
          8968 => x"19",
          8969 => x"8b",
          8970 => x"f9",
          8971 => x"84",
          8972 => x"56",
          8973 => x"a7",
          8974 => x"fc",
          8975 => x"53",
          8976 => x"75",
          8977 => x"a1",
          8978 => x"98",
          8979 => x"84",
          8980 => x"2e",
          8981 => x"87",
          8982 => x"08",
          8983 => x"ff",
          8984 => x"bb",
          8985 => x"3d",
          8986 => x"3d",
          8987 => x"80",
          8988 => x"52",
          8989 => x"9a",
          8990 => x"74",
          8991 => x"0d",
          8992 => x"0d",
          8993 => x"05",
          8994 => x"86",
          8995 => x"54",
          8996 => x"73",
          8997 => x"fe",
          8998 => x"51",
          8999 => x"98",
          9000 => x"00",
          9001 => x"ff",
          9002 => x"ff",
          9003 => x"ff",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"00",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"00",
          9136 => x"00",
          9137 => x"00",
          9138 => x"00",
          9139 => x"00",
          9140 => x"64",
          9141 => x"74",
          9142 => x"64",
          9143 => x"74",
          9144 => x"66",
          9145 => x"74",
          9146 => x"66",
          9147 => x"64",
          9148 => x"66",
          9149 => x"63",
          9150 => x"6d",
          9151 => x"61",
          9152 => x"6d",
          9153 => x"79",
          9154 => x"6d",
          9155 => x"66",
          9156 => x"6d",
          9157 => x"70",
          9158 => x"6d",
          9159 => x"6d",
          9160 => x"6d",
          9161 => x"68",
          9162 => x"68",
          9163 => x"68",
          9164 => x"68",
          9165 => x"63",
          9166 => x"00",
          9167 => x"6a",
          9168 => x"72",
          9169 => x"61",
          9170 => x"72",
          9171 => x"74",
          9172 => x"69",
          9173 => x"00",
          9174 => x"74",
          9175 => x"00",
          9176 => x"74",
          9177 => x"69",
          9178 => x"6d",
          9179 => x"69",
          9180 => x"6b",
          9181 => x"00",
          9182 => x"65",
          9183 => x"44",
          9184 => x"20",
          9185 => x"6f",
          9186 => x"49",
          9187 => x"72",
          9188 => x"20",
          9189 => x"6f",
          9190 => x"00",
          9191 => x"44",
          9192 => x"20",
          9193 => x"20",
          9194 => x"64",
          9195 => x"00",
          9196 => x"4e",
          9197 => x"69",
          9198 => x"66",
          9199 => x"64",
          9200 => x"4e",
          9201 => x"61",
          9202 => x"66",
          9203 => x"64",
          9204 => x"49",
          9205 => x"6c",
          9206 => x"66",
          9207 => x"6e",
          9208 => x"2e",
          9209 => x"41",
          9210 => x"73",
          9211 => x"65",
          9212 => x"64",
          9213 => x"46",
          9214 => x"20",
          9215 => x"65",
          9216 => x"20",
          9217 => x"73",
          9218 => x"0a",
          9219 => x"46",
          9220 => x"20",
          9221 => x"64",
          9222 => x"69",
          9223 => x"6c",
          9224 => x"0a",
          9225 => x"53",
          9226 => x"73",
          9227 => x"69",
          9228 => x"70",
          9229 => x"65",
          9230 => x"64",
          9231 => x"44",
          9232 => x"65",
          9233 => x"6d",
          9234 => x"20",
          9235 => x"69",
          9236 => x"6c",
          9237 => x"0a",
          9238 => x"44",
          9239 => x"20",
          9240 => x"20",
          9241 => x"62",
          9242 => x"2e",
          9243 => x"4e",
          9244 => x"6f",
          9245 => x"74",
          9246 => x"65",
          9247 => x"6c",
          9248 => x"73",
          9249 => x"20",
          9250 => x"6e",
          9251 => x"6e",
          9252 => x"73",
          9253 => x"00",
          9254 => x"46",
          9255 => x"61",
          9256 => x"62",
          9257 => x"65",
          9258 => x"00",
          9259 => x"54",
          9260 => x"6f",
          9261 => x"20",
          9262 => x"72",
          9263 => x"6f",
          9264 => x"61",
          9265 => x"6c",
          9266 => x"2e",
          9267 => x"46",
          9268 => x"20",
          9269 => x"6c",
          9270 => x"65",
          9271 => x"00",
          9272 => x"49",
          9273 => x"66",
          9274 => x"69",
          9275 => x"20",
          9276 => x"6f",
          9277 => x"0a",
          9278 => x"54",
          9279 => x"6d",
          9280 => x"20",
          9281 => x"6e",
          9282 => x"6c",
          9283 => x"0a",
          9284 => x"50",
          9285 => x"6d",
          9286 => x"72",
          9287 => x"6e",
          9288 => x"72",
          9289 => x"2e",
          9290 => x"53",
          9291 => x"65",
          9292 => x"0a",
          9293 => x"55",
          9294 => x"6f",
          9295 => x"65",
          9296 => x"72",
          9297 => x"0a",
          9298 => x"20",
          9299 => x"65",
          9300 => x"73",
          9301 => x"20",
          9302 => x"20",
          9303 => x"65",
          9304 => x"65",
          9305 => x"00",
          9306 => x"72",
          9307 => x"00",
          9308 => x"25",
          9309 => x"00",
          9310 => x"3a",
          9311 => x"25",
          9312 => x"00",
          9313 => x"20",
          9314 => x"20",
          9315 => x"00",
          9316 => x"25",
          9317 => x"00",
          9318 => x"20",
          9319 => x"20",
          9320 => x"7c",
          9321 => x"5a",
          9322 => x"41",
          9323 => x"0a",
          9324 => x"25",
          9325 => x"00",
          9326 => x"30",
          9327 => x"35",
          9328 => x"32",
          9329 => x"76",
          9330 => x"32",
          9331 => x"20",
          9332 => x"2c",
          9333 => x"76",
          9334 => x"32",
          9335 => x"25",
          9336 => x"73",
          9337 => x"0a",
          9338 => x"5a",
          9339 => x"41",
          9340 => x"74",
          9341 => x"75",
          9342 => x"48",
          9343 => x"6c",
          9344 => x"00",
          9345 => x"54",
          9346 => x"72",
          9347 => x"74",
          9348 => x"75",
          9349 => x"00",
          9350 => x"50",
          9351 => x"69",
          9352 => x"72",
          9353 => x"74",
          9354 => x"49",
          9355 => x"4c",
          9356 => x"20",
          9357 => x"65",
          9358 => x"70",
          9359 => x"49",
          9360 => x"4c",
          9361 => x"20",
          9362 => x"65",
          9363 => x"70",
          9364 => x"55",
          9365 => x"30",
          9366 => x"20",
          9367 => x"65",
          9368 => x"70",
          9369 => x"55",
          9370 => x"30",
          9371 => x"20",
          9372 => x"65",
          9373 => x"70",
          9374 => x"55",
          9375 => x"31",
          9376 => x"20",
          9377 => x"65",
          9378 => x"70",
          9379 => x"55",
          9380 => x"31",
          9381 => x"20",
          9382 => x"65",
          9383 => x"70",
          9384 => x"53",
          9385 => x"69",
          9386 => x"75",
          9387 => x"69",
          9388 => x"2e",
          9389 => x"00",
          9390 => x"45",
          9391 => x"6c",
          9392 => x"20",
          9393 => x"65",
          9394 => x"2e",
          9395 => x"61",
          9396 => x"65",
          9397 => x"2e",
          9398 => x"00",
          9399 => x"7a",
          9400 => x"61",
          9401 => x"74",
          9402 => x"30",
          9403 => x"46",
          9404 => x"65",
          9405 => x"6f",
          9406 => x"69",
          9407 => x"6c",
          9408 => x"20",
          9409 => x"63",
          9410 => x"20",
          9411 => x"70",
          9412 => x"73",
          9413 => x"6e",
          9414 => x"6d",
          9415 => x"61",
          9416 => x"2e",
          9417 => x"2a",
          9418 => x"42",
          9419 => x"64",
          9420 => x"20",
          9421 => x"00",
          9422 => x"49",
          9423 => x"69",
          9424 => x"73",
          9425 => x"0a",
          9426 => x"46",
          9427 => x"65",
          9428 => x"6f",
          9429 => x"69",
          9430 => x"6c",
          9431 => x"2e",
          9432 => x"72",
          9433 => x"64",
          9434 => x"25",
          9435 => x"43",
          9436 => x"72",
          9437 => x"2e",
          9438 => x"00",
          9439 => x"43",
          9440 => x"69",
          9441 => x"2e",
          9442 => x"43",
          9443 => x"61",
          9444 => x"67",
          9445 => x"00",
          9446 => x"25",
          9447 => x"78",
          9448 => x"38",
          9449 => x"3e",
          9450 => x"6c",
          9451 => x"30",
          9452 => x"0a",
          9453 => x"44",
          9454 => x"20",
          9455 => x"6f",
          9456 => x"00",
          9457 => x"0a",
          9458 => x"70",
          9459 => x"65",
          9460 => x"25",
          9461 => x"20",
          9462 => x"58",
          9463 => x"3f",
          9464 => x"00",
          9465 => x"25",
          9466 => x"20",
          9467 => x"58",
          9468 => x"25",
          9469 => x"20",
          9470 => x"58",
          9471 => x"44",
          9472 => x"62",
          9473 => x"67",
          9474 => x"74",
          9475 => x"75",
          9476 => x"0a",
          9477 => x"45",
          9478 => x"6c",
          9479 => x"20",
          9480 => x"65",
          9481 => x"70",
          9482 => x"00",
          9483 => x"44",
          9484 => x"62",
          9485 => x"20",
          9486 => x"74",
          9487 => x"66",
          9488 => x"45",
          9489 => x"6c",
          9490 => x"20",
          9491 => x"74",
          9492 => x"66",
          9493 => x"45",
          9494 => x"75",
          9495 => x"67",
          9496 => x"64",
          9497 => x"20",
          9498 => x"78",
          9499 => x"2e",
          9500 => x"43",
          9501 => x"69",
          9502 => x"63",
          9503 => x"20",
          9504 => x"30",
          9505 => x"2e",
          9506 => x"00",
          9507 => x"43",
          9508 => x"20",
          9509 => x"75",
          9510 => x"64",
          9511 => x"64",
          9512 => x"25",
          9513 => x"0a",
          9514 => x"52",
          9515 => x"61",
          9516 => x"6e",
          9517 => x"70",
          9518 => x"63",
          9519 => x"6f",
          9520 => x"2e",
          9521 => x"43",
          9522 => x"20",
          9523 => x"6f",
          9524 => x"6e",
          9525 => x"2e",
          9526 => x"5a",
          9527 => x"62",
          9528 => x"25",
          9529 => x"25",
          9530 => x"73",
          9531 => x"00",
          9532 => x"25",
          9533 => x"25",
          9534 => x"73",
          9535 => x"25",
          9536 => x"25",
          9537 => x"42",
          9538 => x"63",
          9539 => x"61",
          9540 => x"00",
          9541 => x"52",
          9542 => x"69",
          9543 => x"2e",
          9544 => x"45",
          9545 => x"6c",
          9546 => x"20",
          9547 => x"65",
          9548 => x"70",
          9549 => x"2e",
          9550 => x"25",
          9551 => x"64",
          9552 => x"20",
          9553 => x"25",
          9554 => x"64",
          9555 => x"25",
          9556 => x"53",
          9557 => x"43",
          9558 => x"69",
          9559 => x"61",
          9560 => x"6e",
          9561 => x"20",
          9562 => x"6f",
          9563 => x"6f",
          9564 => x"6f",
          9565 => x"67",
          9566 => x"3a",
          9567 => x"76",
          9568 => x"73",
          9569 => x"70",
          9570 => x"65",
          9571 => x"64",
          9572 => x"20",
          9573 => x"57",
          9574 => x"44",
          9575 => x"20",
          9576 => x"30",
          9577 => x"25",
          9578 => x"29",
          9579 => x"20",
          9580 => x"53",
          9581 => x"4d",
          9582 => x"20",
          9583 => x"30",
          9584 => x"25",
          9585 => x"29",
          9586 => x"20",
          9587 => x"49",
          9588 => x"20",
          9589 => x"4d",
          9590 => x"30",
          9591 => x"25",
          9592 => x"29",
          9593 => x"20",
          9594 => x"42",
          9595 => x"20",
          9596 => x"20",
          9597 => x"30",
          9598 => x"25",
          9599 => x"29",
          9600 => x"20",
          9601 => x"52",
          9602 => x"20",
          9603 => x"20",
          9604 => x"30",
          9605 => x"25",
          9606 => x"29",
          9607 => x"20",
          9608 => x"53",
          9609 => x"41",
          9610 => x"20",
          9611 => x"65",
          9612 => x"65",
          9613 => x"25",
          9614 => x"29",
          9615 => x"20",
          9616 => x"54",
          9617 => x"52",
          9618 => x"20",
          9619 => x"69",
          9620 => x"73",
          9621 => x"25",
          9622 => x"29",
          9623 => x"20",
          9624 => x"49",
          9625 => x"20",
          9626 => x"4c",
          9627 => x"68",
          9628 => x"65",
          9629 => x"25",
          9630 => x"29",
          9631 => x"20",
          9632 => x"57",
          9633 => x"42",
          9634 => x"20",
          9635 => x"0a",
          9636 => x"20",
          9637 => x"57",
          9638 => x"32",
          9639 => x"20",
          9640 => x"49",
          9641 => x"4c",
          9642 => x"20",
          9643 => x"50",
          9644 => x"00",
          9645 => x"20",
          9646 => x"53",
          9647 => x"00",
          9648 => x"41",
          9649 => x"65",
          9650 => x"73",
          9651 => x"20",
          9652 => x"43",
          9653 => x"52",
          9654 => x"74",
          9655 => x"63",
          9656 => x"20",
          9657 => x"72",
          9658 => x"20",
          9659 => x"30",
          9660 => x"00",
          9661 => x"20",
          9662 => x"43",
          9663 => x"4d",
          9664 => x"72",
          9665 => x"74",
          9666 => x"20",
          9667 => x"72",
          9668 => x"20",
          9669 => x"30",
          9670 => x"00",
          9671 => x"20",
          9672 => x"53",
          9673 => x"6b",
          9674 => x"61",
          9675 => x"41",
          9676 => x"65",
          9677 => x"20",
          9678 => x"20",
          9679 => x"30",
          9680 => x"00",
          9681 => x"4d",
          9682 => x"3a",
          9683 => x"20",
          9684 => x"5a",
          9685 => x"49",
          9686 => x"20",
          9687 => x"20",
          9688 => x"20",
          9689 => x"20",
          9690 => x"20",
          9691 => x"30",
          9692 => x"00",
          9693 => x"20",
          9694 => x"53",
          9695 => x"65",
          9696 => x"6c",
          9697 => x"20",
          9698 => x"71",
          9699 => x"20",
          9700 => x"20",
          9701 => x"64",
          9702 => x"34",
          9703 => x"7a",
          9704 => x"20",
          9705 => x"53",
          9706 => x"4d",
          9707 => x"6f",
          9708 => x"46",
          9709 => x"20",
          9710 => x"20",
          9711 => x"20",
          9712 => x"64",
          9713 => x"34",
          9714 => x"7a",
          9715 => x"20",
          9716 => x"57",
          9717 => x"62",
          9718 => x"20",
          9719 => x"41",
          9720 => x"6c",
          9721 => x"20",
          9722 => x"71",
          9723 => x"64",
          9724 => x"34",
          9725 => x"7a",
          9726 => x"53",
          9727 => x"6c",
          9728 => x"4d",
          9729 => x"75",
          9730 => x"46",
          9731 => x"00",
          9732 => x"45",
          9733 => x"45",
          9734 => x"69",
          9735 => x"55",
          9736 => x"6f",
          9737 => x"00",
          9738 => x"01",
          9739 => x"00",
          9740 => x"00",
          9741 => x"01",
          9742 => x"00",
          9743 => x"00",
          9744 => x"01",
          9745 => x"00",
          9746 => x"00",
          9747 => x"01",
          9748 => x"00",
          9749 => x"00",
          9750 => x"01",
          9751 => x"00",
          9752 => x"00",
          9753 => x"01",
          9754 => x"00",
          9755 => x"00",
          9756 => x"01",
          9757 => x"00",
          9758 => x"00",
          9759 => x"01",
          9760 => x"00",
          9761 => x"00",
          9762 => x"01",
          9763 => x"00",
          9764 => x"00",
          9765 => x"01",
          9766 => x"00",
          9767 => x"00",
          9768 => x"01",
          9769 => x"00",
          9770 => x"00",
          9771 => x"04",
          9772 => x"00",
          9773 => x"00",
          9774 => x"04",
          9775 => x"00",
          9776 => x"00",
          9777 => x"04",
          9778 => x"00",
          9779 => x"00",
          9780 => x"03",
          9781 => x"00",
          9782 => x"00",
          9783 => x"04",
          9784 => x"00",
          9785 => x"00",
          9786 => x"04",
          9787 => x"00",
          9788 => x"00",
          9789 => x"04",
          9790 => x"00",
          9791 => x"00",
          9792 => x"03",
          9793 => x"00",
          9794 => x"00",
          9795 => x"03",
          9796 => x"00",
          9797 => x"00",
          9798 => x"03",
          9799 => x"00",
          9800 => x"00",
          9801 => x"03",
          9802 => x"00",
          9803 => x"1b",
          9804 => x"1b",
          9805 => x"1b",
          9806 => x"1b",
          9807 => x"1b",
          9808 => x"1b",
          9809 => x"1b",
          9810 => x"1b",
          9811 => x"1b",
          9812 => x"1b",
          9813 => x"1b",
          9814 => x"10",
          9815 => x"0e",
          9816 => x"0d",
          9817 => x"0b",
          9818 => x"08",
          9819 => x"06",
          9820 => x"05",
          9821 => x"04",
          9822 => x"03",
          9823 => x"02",
          9824 => x"01",
          9825 => x"68",
          9826 => x"6f",
          9827 => x"68",
          9828 => x"00",
          9829 => x"21",
          9830 => x"25",
          9831 => x"20",
          9832 => x"0a",
          9833 => x"46",
          9834 => x"65",
          9835 => x"6f",
          9836 => x"73",
          9837 => x"74",
          9838 => x"68",
          9839 => x"6f",
          9840 => x"66",
          9841 => x"20",
          9842 => x"45",
          9843 => x"0a",
          9844 => x"43",
          9845 => x"6f",
          9846 => x"70",
          9847 => x"63",
          9848 => x"74",
          9849 => x"69",
          9850 => x"72",
          9851 => x"69",
          9852 => x"20",
          9853 => x"61",
          9854 => x"6e",
          9855 => x"53",
          9856 => x"22",
          9857 => x"3a",
          9858 => x"3e",
          9859 => x"7c",
          9860 => x"46",
          9861 => x"46",
          9862 => x"32",
          9863 => x"eb",
          9864 => x"53",
          9865 => x"35",
          9866 => x"4e",
          9867 => x"41",
          9868 => x"20",
          9869 => x"41",
          9870 => x"20",
          9871 => x"4e",
          9872 => x"41",
          9873 => x"20",
          9874 => x"41",
          9875 => x"20",
          9876 => x"00",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"80",
          9881 => x"8e",
          9882 => x"45",
          9883 => x"49",
          9884 => x"90",
          9885 => x"99",
          9886 => x"59",
          9887 => x"9c",
          9888 => x"41",
          9889 => x"a5",
          9890 => x"a8",
          9891 => x"ac",
          9892 => x"b0",
          9893 => x"b4",
          9894 => x"b8",
          9895 => x"bc",
          9896 => x"c0",
          9897 => x"c4",
          9898 => x"c8",
          9899 => x"cc",
          9900 => x"d0",
          9901 => x"d4",
          9902 => x"d8",
          9903 => x"dc",
          9904 => x"e0",
          9905 => x"e4",
          9906 => x"e8",
          9907 => x"ec",
          9908 => x"f0",
          9909 => x"f4",
          9910 => x"f8",
          9911 => x"fc",
          9912 => x"2b",
          9913 => x"3d",
          9914 => x"5c",
          9915 => x"3c",
          9916 => x"7f",
          9917 => x"00",
          9918 => x"00",
          9919 => x"01",
          9920 => x"00",
          9921 => x"00",
          9922 => x"00",
          9923 => x"00",
          9924 => x"00",
          9925 => x"00",
          9926 => x"00",
          9927 => x"01",
          9928 => x"00",
          9929 => x"00",
          9930 => x"00",
          9931 => x"01",
          9932 => x"00",
          9933 => x"00",
          9934 => x"00",
          9935 => x"01",
          9936 => x"00",
          9937 => x"00",
          9938 => x"00",
          9939 => x"01",
          9940 => x"00",
          9941 => x"00",
          9942 => x"00",
          9943 => x"01",
          9944 => x"00",
          9945 => x"00",
          9946 => x"00",
          9947 => x"01",
          9948 => x"00",
          9949 => x"00",
          9950 => x"00",
          9951 => x"01",
          9952 => x"00",
          9953 => x"00",
          9954 => x"00",
          9955 => x"01",
          9956 => x"00",
          9957 => x"00",
          9958 => x"00",
          9959 => x"01",
          9960 => x"00",
          9961 => x"00",
          9962 => x"00",
          9963 => x"01",
          9964 => x"00",
          9965 => x"00",
          9966 => x"00",
          9967 => x"01",
          9968 => x"00",
          9969 => x"00",
          9970 => x"00",
          9971 => x"01",
          9972 => x"00",
          9973 => x"00",
          9974 => x"00",
          9975 => x"01",
          9976 => x"00",
          9977 => x"00",
          9978 => x"00",
          9979 => x"01",
          9980 => x"00",
          9981 => x"00",
          9982 => x"00",
          9983 => x"01",
          9984 => x"00",
          9985 => x"00",
          9986 => x"00",
          9987 => x"01",
          9988 => x"00",
          9989 => x"00",
          9990 => x"00",
          9991 => x"01",
          9992 => x"00",
          9993 => x"00",
          9994 => x"00",
          9995 => x"01",
          9996 => x"00",
          9997 => x"00",
          9998 => x"00",
          9999 => x"01",
         10000 => x"00",
         10001 => x"00",
         10002 => x"00",
         10003 => x"01",
         10004 => x"00",
         10005 => x"00",
         10006 => x"00",
         10007 => x"01",
         10008 => x"00",
         10009 => x"00",
         10010 => x"00",
         10011 => x"01",
         10012 => x"00",
         10013 => x"00",
         10014 => x"00",
         10015 => x"01",
         10016 => x"00",
         10017 => x"00",
         10018 => x"00",
         10019 => x"01",
         10020 => x"00",
         10021 => x"00",
         10022 => x"00",
         10023 => x"01",
         10024 => x"00",
         10025 => x"00",
         10026 => x"00",
         10027 => x"01",
         10028 => x"00",
         10029 => x"00",
         10030 => x"00",
         10031 => x"00",
         10032 => x"00",
         10033 => x"00",
         10034 => x"00",
         10035 => x"00",
         10036 => x"00",
         10037 => x"00",
         10038 => x"00",
         10039 => x"01",
         10040 => x"01",
         10041 => x"00",
         10042 => x"00",
         10043 => x"00",
         10044 => x"00",
         10045 => x"05",
         10046 => x"05",
         10047 => x"05",
         10048 => x"00",
         10049 => x"01",
         10050 => x"01",
         10051 => x"01",
         10052 => x"01",
         10053 => x"00",
         10054 => x"00",
         10055 => x"00",
         10056 => x"00",
         10057 => x"00",
         10058 => x"00",
         10059 => x"00",
         10060 => x"00",
         10061 => x"00",
         10062 => x"00",
         10063 => x"00",
         10064 => x"00",
         10065 => x"00",
         10066 => x"00",
         10067 => x"00",
         10068 => x"00",
         10069 => x"00",
         10070 => x"00",
         10071 => x"00",
         10072 => x"00",
         10073 => x"00",
         10074 => x"00",
         10075 => x"00",
         10076 => x"00",
         10077 => x"00",
         10078 => x"01",
         10079 => x"00",
         10080 => x"01",
         10081 => x"00",
         10082 => x"02",
         10083 => x"00",
         10084 => x"00",
         10085 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
