-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b87fa",
             1 => x"f80d0b0b",
             2 => x"0b93e904",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"cd040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b93b0",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b83bd",
           162 => x"f4738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93b50400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0bac",
           171 => x"cc2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0bab",
           179 => x"ab2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"96040b0b",
           269 => x"0b8ca604",
           270 => x"0b0b0b8c",
           271 => x"b6040b0b",
           272 => x"0b8cc604",
           273 => x"0b0b0b8c",
           274 => x"d6040b0b",
           275 => x"0b8ce604",
           276 => x"0b0b0b8c",
           277 => x"f6040b0b",
           278 => x"0b8d8604",
           279 => x"0b0b0b8d",
           280 => x"96040b0b",
           281 => x"0b8da604",
           282 => x"0b0b0b8d",
           283 => x"b6040b0b",
           284 => x"0b8dc604",
           285 => x"0b0b0b8d",
           286 => x"d7040b0b",
           287 => x"0b8de804",
           288 => x"0b0b0b8d",
           289 => x"f9040b0b",
           290 => x"0b8e8a04",
           291 => x"0b0b0b8e",
           292 => x"9b040b0b",
           293 => x"0b8eac04",
           294 => x"0b0b0b8e",
           295 => x"bd040b0b",
           296 => x"0b8ece04",
           297 => x"0b0b0b8e",
           298 => x"df040b0b",
           299 => x"0b8ef004",
           300 => x"0b0b0b8f",
           301 => x"81040b0b",
           302 => x"0b8f9204",
           303 => x"0b0b0b8f",
           304 => x"a3040b0b",
           305 => x"0b8fb404",
           306 => x"0b0b0b8f",
           307 => x"c5040b0b",
           308 => x"0b8fd604",
           309 => x"0b0b0b8f",
           310 => x"e7040b0b",
           311 => x"0b8ff804",
           312 => x"0b0b0b90",
           313 => x"89040b0b",
           314 => x"0b909a04",
           315 => x"0b0b0b90",
           316 => x"ab040b0b",
           317 => x"0b90bc04",
           318 => x"0b0b0b90",
           319 => x"cd040b0b",
           320 => x"0b90de04",
           321 => x"0b0b0b90",
           322 => x"ef040b0b",
           323 => x"0b918004",
           324 => x"0b0b0b91",
           325 => x"91040b0b",
           326 => x"0b91a204",
           327 => x"0b0b0b91",
           328 => x"b3040b0b",
           329 => x"0b91c404",
           330 => x"0b0b0b91",
           331 => x"d5040b0b",
           332 => x"0b91e604",
           333 => x"0b0b0b91",
           334 => x"f7040b0b",
           335 => x"0b928804",
           336 => x"0b0b0b92",
           337 => x"99040b0b",
           338 => x"0b92aa04",
           339 => x"0b0b0b92",
           340 => x"bb040b0b",
           341 => x"0b92cb04",
           342 => x"0b0b0b92",
           343 => x"dc040b0b",
           344 => x"0b92ed04",
           345 => x"0b0b0b92",
           346 => x"fe04ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0484b9d4",
           386 => x"0c80d687",
           387 => x"2d84b9d4",
           388 => x"0880c080",
           389 => x"900484b9",
           390 => x"d40ca2ee",
           391 => x"2d84b9d4",
           392 => x"0880c080",
           393 => x"900484b9",
           394 => x"d40ca0f3",
           395 => x"2d84b9d4",
           396 => x"0880c080",
           397 => x"900484b9",
           398 => x"d40ca0e0",
           399 => x"2d84b9d4",
           400 => x"0880c080",
           401 => x"900484b9",
           402 => x"d40c94a3",
           403 => x"2d84b9d4",
           404 => x"0880c080",
           405 => x"900484b9",
           406 => x"d40ca1f6",
           407 => x"2d84b9d4",
           408 => x"0880c080",
           409 => x"900484b9",
           410 => x"d40caf86",
           411 => x"2d84b9d4",
           412 => x"0880c080",
           413 => x"900484b9",
           414 => x"d40cad82",
           415 => x"2d84b9d4",
           416 => x"0880c080",
           417 => x"900484b9",
           418 => x"d40c9488",
           419 => x"2d84b9d4",
           420 => x"0880c080",
           421 => x"900484b9",
           422 => x"d40c95a8",
           423 => x"2d84b9d4",
           424 => x"0880c080",
           425 => x"900484b9",
           426 => x"d40c95d1",
           427 => x"2d84b9d4",
           428 => x"0880c080",
           429 => x"900484b9",
           430 => x"d40cb18a",
           431 => x"2d84b9d4",
           432 => x"0880c080",
           433 => x"900484b9",
           434 => x"d40c80d4",
           435 => x"ec2d84b9",
           436 => x"d40880c0",
           437 => x"80900484",
           438 => x"b9d40c80",
           439 => x"d5d12d84",
           440 => x"b9d40880",
           441 => x"c0809004",
           442 => x"84b9d40c",
           443 => x"80d2a82d",
           444 => x"84b9d408",
           445 => x"80c08090",
           446 => x"0484b9d4",
           447 => x"0c80d3db",
           448 => x"2d84b9d4",
           449 => x"0880c080",
           450 => x"900484b9",
           451 => x"d40c82c9",
           452 => x"ae2d84b9",
           453 => x"d40880c0",
           454 => x"80900484",
           455 => x"b9d40c82",
           456 => x"e3802d84",
           457 => x"b9d40880",
           458 => x"c0809004",
           459 => x"84b9d40c",
           460 => x"82d29e2d",
           461 => x"84b9d408",
           462 => x"80c08090",
           463 => x"0484b9d4",
           464 => x"0c82d7c0",
           465 => x"2d84b9d4",
           466 => x"0880c080",
           467 => x"900484b9",
           468 => x"d40c82ed",
           469 => x"9d2d84b9",
           470 => x"d40880c0",
           471 => x"80900484",
           472 => x"b9d40c82",
           473 => x"faa52d84",
           474 => x"b9d40880",
           475 => x"c0809004",
           476 => x"84b9d40c",
           477 => x"82df872d",
           478 => x"84b9d408",
           479 => x"80c08090",
           480 => x"0484b9d4",
           481 => x"0c82f1be",
           482 => x"2d84b9d4",
           483 => x"0880c080",
           484 => x"900484b9",
           485 => x"d40c82f3",
           486 => x"8b2d84b9",
           487 => x"d40880c0",
           488 => x"80900484",
           489 => x"b9d40c82",
           490 => x"f3e02d84",
           491 => x"b9d40880",
           492 => x"c0809004",
           493 => x"84b9d40c",
           494 => x"8384a22d",
           495 => x"84b9d408",
           496 => x"80c08090",
           497 => x"0484b9d4",
           498 => x"0c82fee7",
           499 => x"2d84b9d4",
           500 => x"0880c080",
           501 => x"900484b9",
           502 => x"d40c838b",
           503 => x"862d84b9",
           504 => x"d40880c0",
           505 => x"80900484",
           506 => x"b9d40c82",
           507 => x"f5bd2d84",
           508 => x"b9d40880",
           509 => x"c0809004",
           510 => x"84b9d40c",
           511 => x"8393fd2d",
           512 => x"84b9d408",
           513 => x"80c08090",
           514 => x"0484b9d4",
           515 => x"0c839588",
           516 => x"2d84b9d4",
           517 => x"0880c080",
           518 => x"900484b9",
           519 => x"d40c82e5",
           520 => x"d02d84b9",
           521 => x"d40880c0",
           522 => x"80900484",
           523 => x"b9d40c82",
           524 => x"e3e72d84",
           525 => x"b9d40880",
           526 => x"c0809004",
           527 => x"84b9d40c",
           528 => x"82e78e2d",
           529 => x"84b9d408",
           530 => x"80c08090",
           531 => x"0484b9d4",
           532 => x"0c82f6a7",
           533 => x"2d84b9d4",
           534 => x"0880c080",
           535 => x"900484b9",
           536 => x"d40c8396",
           537 => x"9a2d84b9",
           538 => x"d40880c0",
           539 => x"80900484",
           540 => x"b9d40c83",
           541 => x"99f72d84",
           542 => x"b9d40880",
           543 => x"c0809004",
           544 => x"84b9d40c",
           545 => x"83a0e92d",
           546 => x"84b9d408",
           547 => x"80c08090",
           548 => x"0484b9d4",
           549 => x"0c82c6ff",
           550 => x"2d84b9d4",
           551 => x"0880c080",
           552 => x"900484b9",
           553 => x"d40c83a4",
           554 => x"922d84b9",
           555 => x"d40880c0",
           556 => x"80900484",
           557 => x"b9d40c83",
           558 => x"b9932d84",
           559 => x"b9d40880",
           560 => x"c0809004",
           561 => x"84b9d40c",
           562 => x"83b7c52d",
           563 => x"84b9d408",
           564 => x"80c08090",
           565 => x"0484b9d4",
           566 => x"0c81f3e3",
           567 => x"2d84b9d4",
           568 => x"0880c080",
           569 => x"900484b9",
           570 => x"d40c81f4",
           571 => x"e22d84b9",
           572 => x"d40880c0",
           573 => x"80900484",
           574 => x"b9d40c81",
           575 => x"f5e12d84",
           576 => x"b9d40880",
           577 => x"c0809004",
           578 => x"84b9d40c",
           579 => x"80d0aa2d",
           580 => x"84b9d408",
           581 => x"80c08090",
           582 => x"0484b9d4",
           583 => x"0c80d1fa",
           584 => x"2d84b9d4",
           585 => x"0880c080",
           586 => x"900484b9",
           587 => x"d40c80d7",
           588 => x"a52d84b9",
           589 => x"d40880c0",
           590 => x"80900484",
           591 => x"b9d40cb1",
           592 => x"9a2d84b9",
           593 => x"d40880c0",
           594 => x"80900484",
           595 => x"b9d40c81",
           596 => x"db812d84",
           597 => x"b9d40880",
           598 => x"c0809004",
           599 => x"84b9d40c",
           600 => x"81dcbc2d",
           601 => x"84b9d408",
           602 => x"80c08090",
           603 => x"0484b9d4",
           604 => x"0c81f1bd",
           605 => x"2d84b9d4",
           606 => x"0880c080",
           607 => x"900484b9",
           608 => x"d40c81d5",
           609 => x"912d84b9",
           610 => x"d40880c0",
           611 => x"8090043c",
           612 => x"04101010",
           613 => x"10101010",
           614 => x"10101010",
           615 => x"10101010",
           616 => x"10101010",
           617 => x"10101010",
           618 => x"10101010",
           619 => x"10101010",
           620 => x"53510400",
           621 => x"007381ff",
           622 => x"06738306",
           623 => x"09810583",
           624 => x"05101010",
           625 => x"2b0772fc",
           626 => x"060c5151",
           627 => x"04727280",
           628 => x"728106ff",
           629 => x"05097206",
           630 => x"05711052",
           631 => x"720a100a",
           632 => x"5372ed38",
           633 => x"51515351",
           634 => x"0484b9c8",
           635 => x"7084d5b4",
           636 => x"278e3880",
           637 => x"71708405",
           638 => x"530c0b0b",
           639 => x"0b93ec04",
           640 => x"8c815180",
           641 => x"ceba0400",
           642 => x"fc3d0d87",
           643 => x"3d707084",
           644 => x"05520856",
           645 => x"53745284",
           646 => x"d5ac0851",
           647 => x"81c53f86",
           648 => x"3d0d04fa",
           649 => x"3d0d787a",
           650 => x"7c851133",
           651 => x"81328106",
           652 => x"80732507",
           653 => x"56585557",
           654 => x"80527272",
           655 => x"2e098106",
           656 => x"80d338ff",
           657 => x"1477748a",
           658 => x"32703070",
           659 => x"72079f2a",
           660 => x"51555556",
           661 => x"54807425",
           662 => x"b7387180",
           663 => x"2eb23875",
           664 => x"518efa3f",
           665 => x"84b9c808",
           666 => x"5384b9c8",
           667 => x"08ff2eae",
           668 => x"3884b9c8",
           669 => x"08757081",
           670 => x"055734ff",
           671 => x"14738a32",
           672 => x"70307072",
           673 => x"079f2a51",
           674 => x"54545473",
           675 => x"8024cb38",
           676 => x"80753476",
           677 => x"527184b9",
           678 => x"c80c883d",
           679 => x"0d04800b",
           680 => x"84b9c80c",
           681 => x"883d0d04",
           682 => x"f53d0d7d",
           683 => x"54860284",
           684 => x"05990534",
           685 => x"7356fe0a",
           686 => x"588e3d88",
           687 => x"05537e52",
           688 => x"8d3de405",
           689 => x"519d3f73",
           690 => x"19548074",
           691 => x"348d3d0d",
           692 => x"04fd3d0d",
           693 => x"863d8805",
           694 => x"53765275",
           695 => x"51853f85",
           696 => x"3d0d04f1",
           697 => x"3d0d6163",
           698 => x"65425d5d",
           699 => x"80708c1f",
           700 => x"0c851e33",
           701 => x"70812a81",
           702 => x"32810655",
           703 => x"555bff54",
           704 => x"727b2e09",
           705 => x"810680d2",
           706 => x"387b3357",
           707 => x"767b2e80",
           708 => x"c538811c",
           709 => x"7b810654",
           710 => x"5c72802e",
           711 => x"818138d0",
           712 => x"175f7e89",
           713 => x"2681a338",
           714 => x"76b03270",
           715 => x"30708025",
           716 => x"51545578",
           717 => x"ae387280",
           718 => x"2ea9387a",
           719 => x"832a7081",
           720 => x"32810640",
           721 => x"547e802e",
           722 => x"9e387a82",
           723 => x"80075b7b",
           724 => x"335776ff",
           725 => x"bd388c1d",
           726 => x"08547384",
           727 => x"b9c80c91",
           728 => x"3d0d047a",
           729 => x"832a5478",
           730 => x"10101079",
           731 => x"10057098",
           732 => x"2b70982c",
           733 => x"19708180",
           734 => x"0a298b0a",
           735 => x"0570982c",
           736 => x"525a5b56",
           737 => x"5f807924",
           738 => x"81863873",
           739 => x"81065372",
           740 => x"ffbd3878",
           741 => x"7c335858",
           742 => x"76fef738",
           743 => x"ffb83976",
           744 => x"a52e0981",
           745 => x"06933881",
           746 => x"73745a5a",
           747 => x"5b8a7c33",
           748 => x"585a76fe",
           749 => x"dd38ff9e",
           750 => x"397c5276",
           751 => x"518baf3f",
           752 => x"7b335776",
           753 => x"fecc38ff",
           754 => x"8d397a83",
           755 => x"2a708106",
           756 => x"5455788a",
           757 => x"38817074",
           758 => x"0640547e",
           759 => x"9538e017",
           760 => x"537280d8",
           761 => x"26973872",
           762 => x"101083ca",
           763 => x"84055473",
           764 => x"080473e0",
           765 => x"18545980",
           766 => x"d87327eb",
           767 => x"387c5276",
           768 => x"518aeb3f",
           769 => x"807c3358",
           770 => x"5b76fe86",
           771 => x"38fec739",
           772 => x"80ff59fe",
           773 => x"f639885a",
           774 => x"7f608405",
           775 => x"71087d83",
           776 => x"ffcf065e",
           777 => x"58415484",
           778 => x"b9d85e79",
           779 => x"52755193",
           780 => x"9a3f84b9",
           781 => x"c80881ff",
           782 => x"0684b9c8",
           783 => x"0818df05",
           784 => x"56537289",
           785 => x"26883884",
           786 => x"b9c808b0",
           787 => x"0555747e",
           788 => x"70810540",
           789 => x"34795275",
           790 => x"5190ca3f",
           791 => x"84b9c808",
           792 => x"5684b9c8",
           793 => x"08c5387d",
           794 => x"84b9d831",
           795 => x"982b7bb2",
           796 => x"0640567e",
           797 => x"802e8f38",
           798 => x"77848080",
           799 => x"29fc8080",
           800 => x"0570902c",
           801 => x"59557a86",
           802 => x"2a708106",
           803 => x"555f7380",
           804 => x"2e9e3877",
           805 => x"84808029",
           806 => x"f8808005",
           807 => x"5379902e",
           808 => x"8b387784",
           809 => x"808029fc",
           810 => x"80800553",
           811 => x"72902c58",
           812 => x"7a832a70",
           813 => x"81065455",
           814 => x"72802e9e",
           815 => x"3875982c",
           816 => x"7081ff06",
           817 => x"54547873",
           818 => x"2486cc38",
           819 => x"7a83fff7",
           820 => x"0670832a",
           821 => x"71862a41",
           822 => x"565b7481",
           823 => x"06547380",
           824 => x"2e85f038",
           825 => x"77793190",
           826 => x"2b70902c",
           827 => x"7c838006",
           828 => x"56595373",
           829 => x"802e8596",
           830 => x"387a812a",
           831 => x"81065473",
           832 => x"85eb387a",
           833 => x"842a8106",
           834 => x"54738698",
           835 => x"387a852a",
           836 => x"81065473",
           837 => x"8697387e",
           838 => x"81065473",
           839 => x"858f387a",
           840 => x"882a8106",
           841 => x"5f7e802e",
           842 => x"b2387778",
           843 => x"84808029",
           844 => x"fc808005",
           845 => x"70902c5a",
           846 => x"40548074",
           847 => x"259d387c",
           848 => x"52b05188",
           849 => x"a93f7778",
           850 => x"84808029",
           851 => x"fc808005",
           852 => x"70902c5a",
           853 => x"40547380",
           854 => x"24e53874",
           855 => x"81065372",
           856 => x"802eb238",
           857 => x"78798180",
           858 => x"0a2981ff",
           859 => x"0a057098",
           860 => x"2c5b5555",
           861 => x"8075259d",
           862 => x"387c52b0",
           863 => x"5187ef3f",
           864 => x"78798180",
           865 => x"0a2981ff",
           866 => x"0a057098",
           867 => x"2c5b5555",
           868 => x"748024e5",
           869 => x"387a872a",
           870 => x"7081065c",
           871 => x"557a802e",
           872 => x"81b93876",
           873 => x"80e32e84",
           874 => x"d8387680",
           875 => x"f32e81ca",
           876 => x"387680d3",
           877 => x"2e81e238",
           878 => x"7d84b9d8",
           879 => x"2e96387c",
           880 => x"52ff1e70",
           881 => x"33525e87",
           882 => x"a53f7d84",
           883 => x"b9d82e09",
           884 => x"8106ec38",
           885 => x"7481065b",
           886 => x"7a802efc",
           887 => x"a7387778",
           888 => x"84808029",
           889 => x"fc808005",
           890 => x"70902c5a",
           891 => x"40558075",
           892 => x"25fc9138",
           893 => x"7c52a051",
           894 => x"86f43fe2",
           895 => x"397a9007",
           896 => x"5b7aa007",
           897 => x"7c33585b",
           898 => x"76fa8738",
           899 => x"fac8397a",
           900 => x"80c0075b",
           901 => x"80f85790",
           902 => x"60618405",
           903 => x"71087e83",
           904 => x"ffcf065f",
           905 => x"5942555a",
           906 => x"fbfd397f",
           907 => x"60840577",
           908 => x"fe800a06",
           909 => x"83133370",
           910 => x"982b7207",
           911 => x"7c848080",
           912 => x"29fc8080",
           913 => x"0570902c",
           914 => x"5e525a56",
           915 => x"57415f7a",
           916 => x"872a7081",
           917 => x"065c557a",
           918 => x"fec93877",
           919 => x"78848080",
           920 => x"29fc8080",
           921 => x"0570902c",
           922 => x"5a545f80",
           923 => x"7f25feb3",
           924 => x"387c52a0",
           925 => x"5185f73f",
           926 => x"e239ff1a",
           927 => x"7083ffff",
           928 => x"065b5779",
           929 => x"83ffff2e",
           930 => x"feca387c",
           931 => x"52757081",
           932 => x"05573351",
           933 => x"85d83fe2",
           934 => x"39ff1a70",
           935 => x"83ffff06",
           936 => x"5b547983",
           937 => x"ffff2efe",
           938 => x"ab387c52",
           939 => x"75708105",
           940 => x"57335185",
           941 => x"b93fe239",
           942 => x"75fc0a06",
           943 => x"81fc0a07",
           944 => x"78848080",
           945 => x"29fc8080",
           946 => x"0570902c",
           947 => x"5a585680",
           948 => x"e37b872a",
           949 => x"7081065d",
           950 => x"56577afd",
           951 => x"c638fefb",
           952 => x"397f6084",
           953 => x"05710870",
           954 => x"53404156",
           955 => x"807e2482",
           956 => x"df387a83",
           957 => x"ffbf065b",
           958 => x"84b9d85e",
           959 => x"faad397a",
           960 => x"84077c33",
           961 => x"585b76f8",
           962 => x"8938f8ca",
           963 => x"397a8807",
           964 => x"5b807c33",
           965 => x"585976f7",
           966 => x"f938f8ba",
           967 => x"397f6084",
           968 => x"05710877",
           969 => x"81065658",
           970 => x"415f7282",
           971 => x"8a387551",
           972 => x"87f63f84",
           973 => x"b9c80883",
           974 => x"ffff0678",
           975 => x"7131902b",
           976 => x"545a7290",
           977 => x"2c58fe87",
           978 => x"397a80c0",
           979 => x"077c3358",
           980 => x"5b76f7be",
           981 => x"38f7ff39",
           982 => x"7f608405",
           983 => x"71087781",
           984 => x"065d5841",
           985 => x"547981cf",
           986 => x"38755187",
           987 => x"bb3f84b9",
           988 => x"c80883ff",
           989 => x"ff067871",
           990 => x"31902b54",
           991 => x"5ac4397a",
           992 => x"8180077c",
           993 => x"33585b76",
           994 => x"f78838f7",
           995 => x"c9397778",
           996 => x"84808029",
           997 => x"fc808005",
           998 => x"70902c5a",
           999 => x"54548074",
          1000 => x"25fad638",
          1001 => x"7c52a051",
          1002 => x"83c43fe2",
          1003 => x"397c52b0",
          1004 => x"5183bb3f",
          1005 => x"79902e09",
          1006 => x"8106fae3",
          1007 => x"387c5276",
          1008 => x"5183ab3f",
          1009 => x"7a882a81",
          1010 => x"065f7e80",
          1011 => x"2efb8c38",
          1012 => x"fad83975",
          1013 => x"982c7871",
          1014 => x"31902b70",
          1015 => x"902c7d83",
          1016 => x"8006575a",
          1017 => x"515373fa",
          1018 => x"9038ffa2",
          1019 => x"397c52ad",
          1020 => x"5182fb3f",
          1021 => x"7e810654",
          1022 => x"73802efa",
          1023 => x"a238ffad",
          1024 => x"397c5275",
          1025 => x"982a5182",
          1026 => x"e53f7481",
          1027 => x"065b7a80",
          1028 => x"2ef7f138",
          1029 => x"fbc83978",
          1030 => x"7431982b",
          1031 => x"70982c5a",
          1032 => x"53f9b739",
          1033 => x"7c52ab51",
          1034 => x"82c43fc8",
          1035 => x"397c52a0",
          1036 => x"5182bb3f",
          1037 => x"ffbe3978",
          1038 => x"52755188",
          1039 => x"8b3f84b9",
          1040 => x"c80883ff",
          1041 => x"ff067871",
          1042 => x"31902b54",
          1043 => x"5afdf339",
          1044 => x"7a82077e",
          1045 => x"307183ff",
          1046 => x"bf065257",
          1047 => x"5bfd9939",
          1048 => x"fe3d0d84",
          1049 => x"d5a80853",
          1050 => x"75527451",
          1051 => x"f3b53f84",
          1052 => x"3d0d04fa",
          1053 => x"3d0d7855",
          1054 => x"800b84d5",
          1055 => x"ac088511",
          1056 => x"3370812a",
          1057 => x"81327081",
          1058 => x"06515658",
          1059 => x"5557ff56",
          1060 => x"72772e09",
          1061 => x"810680d5",
          1062 => x"38747081",
          1063 => x"05563353",
          1064 => x"72772eb0",
          1065 => x"3884d5ac",
          1066 => x"08527251",
          1067 => x"90140853",
          1068 => x"722d84b9",
          1069 => x"c808802e",
          1070 => x"8338ff57",
          1071 => x"74708105",
          1072 => x"56335372",
          1073 => x"802e8838",
          1074 => x"84d5ac08",
          1075 => x"54d73984",
          1076 => x"d5ac0854",
          1077 => x"84d5ac08",
          1078 => x"528a5190",
          1079 => x"14085574",
          1080 => x"2d84b9c8",
          1081 => x"08802e83",
          1082 => x"38ff5776",
          1083 => x"567584b9",
          1084 => x"c80c883d",
          1085 => x"0d04fa3d",
          1086 => x"0d787a56",
          1087 => x"54800b85",
          1088 => x"16337081",
          1089 => x"2a813270",
          1090 => x"81065155",
          1091 => x"5757ff56",
          1092 => x"72772e09",
          1093 => x"81069238",
          1094 => x"73708105",
          1095 => x"55335372",
          1096 => x"772e0981",
          1097 => x"06983876",
          1098 => x"567584b9",
          1099 => x"c80c883d",
          1100 => x"0d047370",
          1101 => x"81055533",
          1102 => x"5372802e",
          1103 => x"ea387452",
          1104 => x"72519015",
          1105 => x"0853722d",
          1106 => x"84b9c808",
          1107 => x"802ee338",
          1108 => x"ff747081",
          1109 => x"05563354",
          1110 => x"5772e338",
          1111 => x"ca39ff3d",
          1112 => x"0d84d5ac",
          1113 => x"08527351",
          1114 => x"853f833d",
          1115 => x"0d04fa3d",
          1116 => x"0d787a85",
          1117 => x"11337081",
          1118 => x"2a813281",
          1119 => x"06565656",
          1120 => x"57ff5672",
          1121 => x"ae387382",
          1122 => x"2a810654",
          1123 => x"73802eac",
          1124 => x"388c1508",
          1125 => x"53728816",
          1126 => x"08259138",
          1127 => x"74085676",
          1128 => x"76347408",
          1129 => x"8105750c",
          1130 => x"8c150853",
          1131 => x"81138c16",
          1132 => x"0c765675",
          1133 => x"84b9c80c",
          1134 => x"883d0d04",
          1135 => x"74527681",
          1136 => x"ff065190",
          1137 => x"15085473",
          1138 => x"2dff5684",
          1139 => x"b9c808e3",
          1140 => x"388c1508",
          1141 => x"81058c16",
          1142 => x"0c7656d7",
          1143 => x"39fb3d0d",
          1144 => x"77851133",
          1145 => x"7081ff06",
          1146 => x"70813281",
          1147 => x"06555556",
          1148 => x"56ff5471",
          1149 => x"b3387286",
          1150 => x"2a810652",
          1151 => x"71b33872",
          1152 => x"822a8106",
          1153 => x"5271802e",
          1154 => x"80c33875",
          1155 => x"08703353",
          1156 => x"5371802e",
          1157 => x"80f03881",
          1158 => x"13760c8c",
          1159 => x"16088105",
          1160 => x"8c170c71",
          1161 => x"81ff0654",
          1162 => x"7384b9c8",
          1163 => x"0c873d0d",
          1164 => x"0474ffbf",
          1165 => x"06537285",
          1166 => x"17348c16",
          1167 => x"0881058c",
          1168 => x"170c8416",
          1169 => x"3384b9c8",
          1170 => x"0c873d0d",
          1171 => x"04755194",
          1172 => x"16085574",
          1173 => x"2d84b9c8",
          1174 => x"085284b9",
          1175 => x"c8088025",
          1176 => x"ffb93885",
          1177 => x"16337090",
          1178 => x"07545284",
          1179 => x"b9c808ff",
          1180 => x"2e853871",
          1181 => x"a0075372",
          1182 => x"851734ff",
          1183 => x"547384b9",
          1184 => x"c80c873d",
          1185 => x"0d0474a0",
          1186 => x"07537285",
          1187 => x"1734ff54",
          1188 => x"ec39fd3d",
          1189 => x"0d757771",
          1190 => x"54545471",
          1191 => x"70810553",
          1192 => x"335170f7",
          1193 => x"38ff1252",
          1194 => x"72708105",
          1195 => x"54335170",
          1196 => x"72708105",
          1197 => x"543470f0",
          1198 => x"387384b9",
          1199 => x"c80c853d",
          1200 => x"0d04fc3d",
          1201 => x"0d767971",
          1202 => x"7a555552",
          1203 => x"5470802e",
          1204 => x"9d387372",
          1205 => x"27a13870",
          1206 => x"802e9338",
          1207 => x"71708105",
          1208 => x"53337370",
          1209 => x"81055534",
          1210 => x"ff115170",
          1211 => x"ef387384",
          1212 => x"b9c80c86",
          1213 => x"3d0d0470",
          1214 => x"12557375",
          1215 => x"27d93870",
          1216 => x"14755353",
          1217 => x"ff13ff13",
          1218 => x"53537133",
          1219 => x"7334ff11",
          1220 => x"5170802e",
          1221 => x"d938ff13",
          1222 => x"ff135353",
          1223 => x"71337334",
          1224 => x"ff115170",
          1225 => x"df38c739",
          1226 => x"fe3d0d74",
          1227 => x"70535371",
          1228 => x"70810553",
          1229 => x"335170f7",
          1230 => x"38ff1270",
          1231 => x"743184b9",
          1232 => x"c80c5184",
          1233 => x"3d0d04fd",
          1234 => x"3d0d7577",
          1235 => x"71545454",
          1236 => x"72708105",
          1237 => x"54335170",
          1238 => x"72708105",
          1239 => x"543470f0",
          1240 => x"387384b9",
          1241 => x"c80c853d",
          1242 => x"0d04fd3d",
          1243 => x"0d757871",
          1244 => x"79555552",
          1245 => x"5470802e",
          1246 => x"93387170",
          1247 => x"81055333",
          1248 => x"73708105",
          1249 => x"5534ff11",
          1250 => x"5170ef38",
          1251 => x"7384b9c8",
          1252 => x"0c853d0d",
          1253 => x"04fc3d0d",
          1254 => x"76787a55",
          1255 => x"56547280",
          1256 => x"2ea13873",
          1257 => x"33757081",
          1258 => x"05573352",
          1259 => x"5271712e",
          1260 => x"0981069a",
          1261 => x"38811454",
          1262 => x"71802eb7",
          1263 => x"38ff1353",
          1264 => x"72e13880",
          1265 => x"517084b9",
          1266 => x"c80c863d",
          1267 => x"0d047280",
          1268 => x"2ef13873",
          1269 => x"3353ff51",
          1270 => x"72802ee9",
          1271 => x"38ff1533",
          1272 => x"52815171",
          1273 => x"802ede38",
          1274 => x"72723184",
          1275 => x"b9c80c86",
          1276 => x"3d0d0471",
          1277 => x"84b9c80c",
          1278 => x"863d0d04",
          1279 => x"fb3d0d77",
          1280 => x"79537052",
          1281 => x"5680c13f",
          1282 => x"84b9c808",
          1283 => x"84b9c808",
          1284 => x"81055255",
          1285 => x"81b2ea3f",
          1286 => x"84b9c808",
          1287 => x"5484b9c8",
          1288 => x"08802e9b",
          1289 => x"3884b9c8",
          1290 => x"08155480",
          1291 => x"74347453",
          1292 => x"755284b9",
          1293 => x"c80851fe",
          1294 => x"b13f84b9",
          1295 => x"c8085473",
          1296 => x"84b9c80c",
          1297 => x"873d0d04",
          1298 => x"fd3d0d75",
          1299 => x"77717154",
          1300 => x"55535471",
          1301 => x"802e9f38",
          1302 => x"72708105",
          1303 => x"54335170",
          1304 => x"802e8c38",
          1305 => x"ff125271",
          1306 => x"ff2e0981",
          1307 => x"06ea38ff",
          1308 => x"13707531",
          1309 => x"52527084",
          1310 => x"b9c80c85",
          1311 => x"3d0d04fd",
          1312 => x"3d0d7577",
          1313 => x"79725553",
          1314 => x"54547080",
          1315 => x"2e8e3872",
          1316 => x"72708105",
          1317 => x"5434ff11",
          1318 => x"5170f438",
          1319 => x"7384b9c8",
          1320 => x"0c853d0d",
          1321 => x"04fa3d0d",
          1322 => x"787a5854",
          1323 => x"a0527680",
          1324 => x"2e8b3876",
          1325 => x"5180f53f",
          1326 => x"84b9c808",
          1327 => x"52e01253",
          1328 => x"73802e8d",
          1329 => x"38735180",
          1330 => x"e33f7184",
          1331 => x"b9c80831",
          1332 => x"53805272",
          1333 => x"9f2680cb",
          1334 => x"38735272",
          1335 => x"9f2e80c3",
          1336 => x"38811374",
          1337 => x"712aa072",
          1338 => x"3176712b",
          1339 => x"57545455",
          1340 => x"80567476",
          1341 => x"2ea83872",
          1342 => x"10749f2a",
          1343 => x"07741077",
          1344 => x"07787231",
          1345 => x"ff119f2c",
          1346 => x"7081067b",
          1347 => x"72067571",
          1348 => x"31ff1c5c",
          1349 => x"56525255",
          1350 => x"58555374",
          1351 => x"da387310",
          1352 => x"76075271",
          1353 => x"84b9c80c",
          1354 => x"883d0d04",
          1355 => x"fc3d0d76",
          1356 => x"70fc8080",
          1357 => x"06703070",
          1358 => x"72078025",
          1359 => x"70842b90",
          1360 => x"71317571",
          1361 => x"2a7083fe",
          1362 => x"80067030",
          1363 => x"70802583",
          1364 => x"2b887131",
          1365 => x"74712a70",
          1366 => x"81f00670",
          1367 => x"30708025",
          1368 => x"822b8471",
          1369 => x"3174712a",
          1370 => x"5553751b",
          1371 => x"05738c06",
          1372 => x"70307080",
          1373 => x"25108271",
          1374 => x"3177712a",
          1375 => x"70812a81",
          1376 => x"32708106",
          1377 => x"70308274",
          1378 => x"31067519",
          1379 => x"0584b9c8",
          1380 => x"0c515254",
          1381 => x"55515456",
          1382 => x"5a535555",
          1383 => x"55515656",
          1384 => x"56565158",
          1385 => x"56545286",
          1386 => x"3d0d04fd",
          1387 => x"3d0d7577",
          1388 => x"70547153",
          1389 => x"54548194",
          1390 => x"3f84b9c8",
          1391 => x"08732974",
          1392 => x"713184b9",
          1393 => x"c80c5385",
          1394 => x"3d0d04fa",
          1395 => x"3d0d787a",
          1396 => x"5854a053",
          1397 => x"76802e8b",
          1398 => x"387651fe",
          1399 => x"cf3f84b9",
          1400 => x"c80853e0",
          1401 => x"13527380",
          1402 => x"2e8d3873",
          1403 => x"51febd3f",
          1404 => x"7284b9c8",
          1405 => x"08315273",
          1406 => x"53719f26",
          1407 => x"80c53880",
          1408 => x"53719f2e",
          1409 => x"be388112",
          1410 => x"74712aa0",
          1411 => x"72317671",
          1412 => x"2b575454",
          1413 => x"55805674",
          1414 => x"762ea838",
          1415 => x"7210749f",
          1416 => x"2a077410",
          1417 => x"77077872",
          1418 => x"31ff119f",
          1419 => x"2c708106",
          1420 => x"7b720675",
          1421 => x"7131ff1c",
          1422 => x"5c565252",
          1423 => x"55585553",
          1424 => x"74da3872",
          1425 => x"84b9c80c",
          1426 => x"883d0d04",
          1427 => x"fa3d0d78",
          1428 => x"9f2c7a9f",
          1429 => x"2c7a9f2c",
          1430 => x"7b327c9f",
          1431 => x"2c7d3273",
          1432 => x"73327174",
          1433 => x"31577275",
          1434 => x"31565956",
          1435 => x"595556fc",
          1436 => x"b43f84b9",
          1437 => x"c8087532",
          1438 => x"753184b9",
          1439 => x"c80c883d",
          1440 => x"0d04f73d",
          1441 => x"0d7b7d5b",
          1442 => x"5780707b",
          1443 => x"0c770870",
          1444 => x"33565659",
          1445 => x"73a02e09",
          1446 => x"81068f38",
          1447 => x"81157078",
          1448 => x"0c703355",
          1449 => x"5573a02e",
          1450 => x"f33873ad",
          1451 => x"2e80f538",
          1452 => x"73b02e81",
          1453 => x"8338d014",
          1454 => x"58805677",
          1455 => x"892680db",
          1456 => x"388a5880",
          1457 => x"56a07427",
          1458 => x"80c43880",
          1459 => x"e0742789",
          1460 => x"38e01470",
          1461 => x"81ff0655",
          1462 => x"53d01470",
          1463 => x"81ff0651",
          1464 => x"53907327",
          1465 => x"8f38f913",
          1466 => x"7081ff06",
          1467 => x"54548973",
          1468 => x"27818938",
          1469 => x"72782781",
          1470 => x"83387776",
          1471 => x"29138116",
          1472 => x"70790c70",
          1473 => x"33565656",
          1474 => x"73a026ff",
          1475 => x"be387880",
          1476 => x"2e843875",
          1477 => x"3056757a",
          1478 => x"0c815675",
          1479 => x"84b9c80c",
          1480 => x"8b3d0d04",
          1481 => x"81701670",
          1482 => x"790c7033",
          1483 => x"56565973",
          1484 => x"b02e0981",
          1485 => x"06feff38",
          1486 => x"81157078",
          1487 => x"0c703355",
          1488 => x"557380e2",
          1489 => x"2ea63890",
          1490 => x"587380f8",
          1491 => x"2ea03881",
          1492 => x"56a07427",
          1493 => x"c638d014",
          1494 => x"53805688",
          1495 => x"58897327",
          1496 => x"fee13875",
          1497 => x"84b9c80c",
          1498 => x"8b3d0d04",
          1499 => x"82588115",
          1500 => x"70780c70",
          1501 => x"33555580",
          1502 => x"56feca39",
          1503 => x"800b84b9",
          1504 => x"c80c8b3d",
          1505 => x"0d04f73d",
          1506 => x"0d7b7d5b",
          1507 => x"5780707b",
          1508 => x"0c770870",
          1509 => x"33565659",
          1510 => x"73a02e09",
          1511 => x"81068f38",
          1512 => x"81157078",
          1513 => x"0c703355",
          1514 => x"5573a02e",
          1515 => x"f33873ad",
          1516 => x"2e80f538",
          1517 => x"73b02e81",
          1518 => x"8338d014",
          1519 => x"58805677",
          1520 => x"892680db",
          1521 => x"388a5880",
          1522 => x"56a07427",
          1523 => x"80c43880",
          1524 => x"e0742789",
          1525 => x"38e01470",
          1526 => x"81ff0655",
          1527 => x"53d01470",
          1528 => x"81ff0651",
          1529 => x"53907327",
          1530 => x"8f38f913",
          1531 => x"7081ff06",
          1532 => x"54548973",
          1533 => x"27818938",
          1534 => x"72782781",
          1535 => x"83387776",
          1536 => x"29138116",
          1537 => x"70790c70",
          1538 => x"33565656",
          1539 => x"73a026ff",
          1540 => x"be387880",
          1541 => x"2e843875",
          1542 => x"3056757a",
          1543 => x"0c815675",
          1544 => x"84b9c80c",
          1545 => x"8b3d0d04",
          1546 => x"81701670",
          1547 => x"790c7033",
          1548 => x"56565973",
          1549 => x"b02e0981",
          1550 => x"06feff38",
          1551 => x"81157078",
          1552 => x"0c703355",
          1553 => x"557380e2",
          1554 => x"2ea63890",
          1555 => x"587380f8",
          1556 => x"2ea03881",
          1557 => x"56a07427",
          1558 => x"c638d014",
          1559 => x"53805688",
          1560 => x"58897327",
          1561 => x"fee13875",
          1562 => x"84b9c80c",
          1563 => x"8b3d0d04",
          1564 => x"82588115",
          1565 => x"70780c70",
          1566 => x"33555580",
          1567 => x"56feca39",
          1568 => x"800b84b9",
          1569 => x"c80c8b3d",
          1570 => x"0d0480d6",
          1571 => x"e23f84b9",
          1572 => x"c80881ff",
          1573 => x"0684b9c8",
          1574 => x"0c04ff3d",
          1575 => x"0d735271",
          1576 => x"93268c38",
          1577 => x"71101083",
          1578 => x"be840552",
          1579 => x"71080483",
          1580 => x"ce9c51ef",
          1581 => x"be3f833d",
          1582 => x"0d0483ce",
          1583 => x"ac51efb3",
          1584 => x"3f833d0d",
          1585 => x"0483cec4",
          1586 => x"51efa83f",
          1587 => x"833d0d04",
          1588 => x"83cedc51",
          1589 => x"ef9d3f83",
          1590 => x"3d0d0483",
          1591 => x"cef451ef",
          1592 => x"923f833d",
          1593 => x"0d0483cf",
          1594 => x"8451ef87",
          1595 => x"3f833d0d",
          1596 => x"0483cfa4",
          1597 => x"51eefc3f",
          1598 => x"833d0d04",
          1599 => x"83cfb451",
          1600 => x"eef13f83",
          1601 => x"3d0d0483",
          1602 => x"cfdc51ee",
          1603 => x"e63f833d",
          1604 => x"0d0483cf",
          1605 => x"f051eedb",
          1606 => x"3f833d0d",
          1607 => x"0483d08c",
          1608 => x"51eed03f",
          1609 => x"833d0d04",
          1610 => x"83d0a451",
          1611 => x"eec53f83",
          1612 => x"3d0d0483",
          1613 => x"d0bc51ee",
          1614 => x"ba3f833d",
          1615 => x"0d0483d0",
          1616 => x"d451eeaf",
          1617 => x"3f833d0d",
          1618 => x"0483d0e4",
          1619 => x"51eea43f",
          1620 => x"833d0d04",
          1621 => x"83d0f851",
          1622 => x"ee993f83",
          1623 => x"3d0d0483",
          1624 => x"d18851ee",
          1625 => x"8e3f833d",
          1626 => x"0d0483d1",
          1627 => x"9851ee83",
          1628 => x"3f833d0d",
          1629 => x"0483d1a8",
          1630 => x"51edf83f",
          1631 => x"833d0d04",
          1632 => x"83d1b851",
          1633 => x"eded3f83",
          1634 => x"3d0d0483",
          1635 => x"d1c451ed",
          1636 => x"e23f833d",
          1637 => x"0d04ec3d",
          1638 => x"0d660284",
          1639 => x"0580e305",
          1640 => x"335b5880",
          1641 => x"68793070",
          1642 => x"7b077325",
          1643 => x"51575759",
          1644 => x"78577587",
          1645 => x"ff268338",
          1646 => x"81577477",
          1647 => x"077081ff",
          1648 => x"06515593",
          1649 => x"577480e2",
          1650 => x"38815377",
          1651 => x"528c3d70",
          1652 => x"52588295",
          1653 => x"d93f84b9",
          1654 => x"c8085784",
          1655 => x"b9c80880",
          1656 => x"2e80d038",
          1657 => x"775182af",
          1658 => x"973f7630",
          1659 => x"70780780",
          1660 => x"257b3070",
          1661 => x"9f2a7206",
          1662 => x"53575758",
          1663 => x"77802eaa",
          1664 => x"3887c098",
          1665 => x"88085574",
          1666 => x"87e72680",
          1667 => x"e0387452",
          1668 => x"7887e829",
          1669 => x"51f58e3f",
          1670 => x"84b9c808",
          1671 => x"5483d1f4",
          1672 => x"53785283",
          1673 => x"d1d051df",
          1674 => x"df3f7684",
          1675 => x"b9c80c96",
          1676 => x"3d0d0484",
          1677 => x"b9c80887",
          1678 => x"c098880c",
          1679 => x"84b9c808",
          1680 => x"59963dd4",
          1681 => x"05548480",
          1682 => x"53755277",
          1683 => x"51829dce",
          1684 => x"3f84b9c8",
          1685 => x"085784b9",
          1686 => x"c808ff88",
          1687 => x"387a5574",
          1688 => x"802eff80",
          1689 => x"38741975",
          1690 => x"175759d5",
          1691 => x"3987e852",
          1692 => x"7451f4b1",
          1693 => x"3f84b9c8",
          1694 => x"08527851",
          1695 => x"f4a73f84",
          1696 => x"b9c80854",
          1697 => x"83d1f453",
          1698 => x"785283d1",
          1699 => x"d051def8",
          1700 => x"3fff9739",
          1701 => x"f83d0d7c",
          1702 => x"028405b7",
          1703 => x"05335859",
          1704 => x"ff588053",
          1705 => x"7b527a51",
          1706 => x"fdec3f84",
          1707 => x"b9c8088b",
          1708 => x"3876802e",
          1709 => x"91387681",
          1710 => x"2e8a3877",
          1711 => x"84b9c80c",
          1712 => x"8a3d0d04",
          1713 => x"780484d5",
          1714 => x"a8566155",
          1715 => x"605484b9",
          1716 => x"c8537f52",
          1717 => x"7e51782d",
          1718 => x"84b9c808",
          1719 => x"84b9c80c",
          1720 => x"8a3d0d04",
          1721 => x"f33d0d7f",
          1722 => x"6163028c",
          1723 => x"0580cf05",
          1724 => x"33737315",
          1725 => x"68415f5c",
          1726 => x"5c5f5d5e",
          1727 => x"78802e83",
          1728 => x"82387a52",
          1729 => x"83d1fc51",
          1730 => x"ddfe3f83",
          1731 => x"d28451dd",
          1732 => x"f73f8054",
          1733 => x"737927b2",
          1734 => x"387c902e",
          1735 => x"81ed387c",
          1736 => x"a02e82a8",
          1737 => x"38731853",
          1738 => x"727a2781",
          1739 => x"a7387233",
          1740 => x"5283d288",
          1741 => x"51ddd13f",
          1742 => x"811484d5",
          1743 => x"ac085354",
          1744 => x"a051ecaa",
          1745 => x"3f787426",
          1746 => x"dc3883d2",
          1747 => x"9051ddb8",
          1748 => x"3f805675",
          1749 => x"792780c0",
          1750 => x"38751870",
          1751 => x"33555380",
          1752 => x"55727a27",
          1753 => x"83388155",
          1754 => x"80539f74",
          1755 => x"27833881",
          1756 => x"53747306",
          1757 => x"7081ff06",
          1758 => x"56577480",
          1759 => x"2e883880",
          1760 => x"fe742781",
          1761 => x"ee3884d5",
          1762 => x"ac0852a0",
          1763 => x"51ebdf3f",
          1764 => x"81165678",
          1765 => x"7626c238",
          1766 => x"83d29451",
          1767 => x"e9d53f78",
          1768 => x"18791c5c",
          1769 => x"5880519d",
          1770 => x"c33f84b9",
          1771 => x"c808982b",
          1772 => x"70982c58",
          1773 => x"5476a02e",
          1774 => x"81ee3876",
          1775 => x"9b2e82c3",
          1776 => x"387b1e57",
          1777 => x"767826fe",
          1778 => x"b938ff0b",
          1779 => x"84b9c80c",
          1780 => x"8f3d0d04",
          1781 => x"83d29851",
          1782 => x"dcae3f81",
          1783 => x"1484d5ac",
          1784 => x"085354a0",
          1785 => x"51eb873f",
          1786 => x"787426fe",
          1787 => x"b838feda",
          1788 => x"3983d2a8",
          1789 => x"51dc913f",
          1790 => x"821484d5",
          1791 => x"ac085354",
          1792 => x"a051eaea",
          1793 => x"3f737927",
          1794 => x"fec03873",
          1795 => x"1853727a",
          1796 => x"27df3872",
          1797 => x"225283d2",
          1798 => x"9c51dbec",
          1799 => x"3f821484",
          1800 => x"d5ac0853",
          1801 => x"54a051ea",
          1802 => x"c53f7874",
          1803 => x"26dd38fe",
          1804 => x"993983d2",
          1805 => x"a451dbd0",
          1806 => x"3f841484",
          1807 => x"d5ac0853",
          1808 => x"54a051ea",
          1809 => x"a93f7379",
          1810 => x"27fdff38",
          1811 => x"73185372",
          1812 => x"7a27df38",
          1813 => x"72085283",
          1814 => x"d1fc51db",
          1815 => x"ab3f8414",
          1816 => x"84d5ac08",
          1817 => x"5354a051",
          1818 => x"ea843f78",
          1819 => x"7426dd38",
          1820 => x"fdd83984",
          1821 => x"d5ac0852",
          1822 => x"7351e9f2",
          1823 => x"3f811656",
          1824 => x"fe913980",
          1825 => x"cee93f84",
          1826 => x"b9c80881",
          1827 => x"ff065388",
          1828 => x"5972a82e",
          1829 => x"fcec38a0",
          1830 => x"597280d0",
          1831 => x"2e098106",
          1832 => x"fce03890",
          1833 => x"59fcdb39",
          1834 => x"80519bc0",
          1835 => x"3f84b9c8",
          1836 => x"08982b70",
          1837 => x"982c70a0",
          1838 => x"32703072",
          1839 => x"9b327030",
          1840 => x"70720773",
          1841 => x"75070651",
          1842 => x"55585957",
          1843 => x"58537280",
          1844 => x"25fde838",
          1845 => x"80519b94",
          1846 => x"3f84b9c8",
          1847 => x"08982b70",
          1848 => x"982c70a0",
          1849 => x"32703072",
          1850 => x"9b327030",
          1851 => x"70720773",
          1852 => x"75070651",
          1853 => x"55585957",
          1854 => x"58538073",
          1855 => x"24ffa938",
          1856 => x"fdb93980",
          1857 => x"0b84b9c8",
          1858 => x"0c8f3d0d",
          1859 => x"04fe3d0d",
          1860 => x"87c09680",
          1861 => x"0853aad7",
          1862 => x"3f81519d",
          1863 => x"883f83d3",
          1864 => x"c0519d99",
          1865 => x"3f80519c",
          1866 => x"fc3f7281",
          1867 => x"2a708106",
          1868 => x"51527182",
          1869 => x"b7387282",
          1870 => x"2a708106",
          1871 => x"51527182",
          1872 => x"89387283",
          1873 => x"2a708106",
          1874 => x"51527181",
          1875 => x"db387284",
          1876 => x"2a708106",
          1877 => x"51527181",
          1878 => x"ad387285",
          1879 => x"2a708106",
          1880 => x"51527180",
          1881 => x"ff387286",
          1882 => x"2a708106",
          1883 => x"51527180",
          1884 => x"d2387287",
          1885 => x"2a708106",
          1886 => x"515271a9",
          1887 => x"3872882a",
          1888 => x"81065372",
          1889 => x"8838a9ef",
          1890 => x"3f843d0d",
          1891 => x"0481519c",
          1892 => x"943f83d3",
          1893 => x"d8519ca5",
          1894 => x"3f80519c",
          1895 => x"883fa9d7",
          1896 => x"3f843d0d",
          1897 => x"0481519b",
          1898 => x"fc3f83d3",
          1899 => x"ec519c8d",
          1900 => x"3f80519b",
          1901 => x"f03f7288",
          1902 => x"2a810653",
          1903 => x"72802ec6",
          1904 => x"38cb3981",
          1905 => x"519bde3f",
          1906 => x"83d48051",
          1907 => x"9bef3f80",
          1908 => x"519bd23f",
          1909 => x"72872a70",
          1910 => x"81065152",
          1911 => x"71802eff",
          1912 => x"9c38c239",
          1913 => x"81519bbd",
          1914 => x"3f83d494",
          1915 => x"519bce3f",
          1916 => x"80519bb1",
          1917 => x"3f72862a",
          1918 => x"70810651",
          1919 => x"5271802e",
          1920 => x"fef038ff",
          1921 => x"be398151",
          1922 => x"9b9b3f83",
          1923 => x"d4a8519b",
          1924 => x"ac3f8051",
          1925 => x"9b8f3f72",
          1926 => x"852a7081",
          1927 => x"06515271",
          1928 => x"802efec2",
          1929 => x"38ffbd39",
          1930 => x"81519af9",
          1931 => x"3f83d4bc",
          1932 => x"519b8a3f",
          1933 => x"80519aed",
          1934 => x"3f72842a",
          1935 => x"70810651",
          1936 => x"5271802e",
          1937 => x"fe9438ff",
          1938 => x"bd398151",
          1939 => x"9ad73f83",
          1940 => x"d4d0519a",
          1941 => x"e83f8051",
          1942 => x"9acb3f72",
          1943 => x"832a7081",
          1944 => x"06515271",
          1945 => x"802efde6",
          1946 => x"38ffbd39",
          1947 => x"81519ab5",
          1948 => x"3f83d4e0",
          1949 => x"519ac63f",
          1950 => x"80519aa9",
          1951 => x"3f72822a",
          1952 => x"70810651",
          1953 => x"5271802e",
          1954 => x"fdb838ff",
          1955 => x"bd39ca3d",
          1956 => x"0d807041",
          1957 => x"41ff6184",
          1958 => x"d0d40c42",
          1959 => x"81526051",
          1960 => x"81b68c3f",
          1961 => x"84b9c808",
          1962 => x"81ff069b",
          1963 => x"3d405978",
          1964 => x"612e84b1",
          1965 => x"3883d5b4",
          1966 => x"51e3b83f",
          1967 => x"983d4383",
          1968 => x"d5ec51d6",
          1969 => x"c33f7e48",
          1970 => x"80f85380",
          1971 => x"527e51eb",
          1972 => x"ae3f0b0b",
          1973 => x"83eebc33",
          1974 => x"7081ff06",
          1975 => x"5b597980",
          1976 => x"2e82f138",
          1977 => x"79812e83",
          1978 => x"88387881",
          1979 => x"ff065e7d",
          1980 => x"822e83c1",
          1981 => x"3867705a",
          1982 => x"5a79802e",
          1983 => x"83dc3879",
          1984 => x"335c7ba0",
          1985 => x"2e098106",
          1986 => x"8c38811a",
          1987 => x"70335d5a",
          1988 => x"7ba02ef6",
          1989 => x"38805c7b",
          1990 => x"9b26be38",
          1991 => x"7b902983",
          1992 => x"eec00570",
          1993 => x"08525be7",
          1994 => x"ff3f84b9",
          1995 => x"c80884b9",
          1996 => x"c808547a",
          1997 => x"537b0852",
          1998 => x"5de8da3f",
          1999 => x"84b9c808",
          2000 => x"8b38841b",
          2001 => x"335e7d81",
          2002 => x"2e838038",
          2003 => x"811c7081",
          2004 => x"ff065d5b",
          2005 => x"9b7c27c4",
          2006 => x"389a3d33",
          2007 => x"5c7b802e",
          2008 => x"fedd3880",
          2009 => x"f8527e51",
          2010 => x"e9923f84",
          2011 => x"b9c8085e",
          2012 => x"84b9c808",
          2013 => x"802e8dc9",
          2014 => x"3884b9c8",
          2015 => x"0848b83d",
          2016 => x"ff800551",
          2017 => x"91a43f84",
          2018 => x"b9c80860",
          2019 => x"62065c5c",
          2020 => x"7a802e81",
          2021 => x"843884b9",
          2022 => x"c80851e7",
          2023 => x"8b3f84b9",
          2024 => x"c8088f26",
          2025 => x"80f33881",
          2026 => x"0ba53d5e",
          2027 => x"5b7a822e",
          2028 => x"8d85387a",
          2029 => x"82248ce2",
          2030 => x"387a812e",
          2031 => x"82e4387b",
          2032 => x"54805383",
          2033 => x"d5f0527c",
          2034 => x"51d5dd3f",
          2035 => x"83f28458",
          2036 => x"84b9f857",
          2037 => x"7d566755",
          2038 => x"80549080",
          2039 => x"0a539080",
          2040 => x"0a527c51",
          2041 => x"f5ae3f84",
          2042 => x"b9c80884",
          2043 => x"b9c80809",
          2044 => x"70307072",
          2045 => x"07802551",
          2046 => x"5b5b4280",
          2047 => x"5a7a8326",
          2048 => x"8338815a",
          2049 => x"787a0659",
          2050 => x"78802e8d",
          2051 => x"38811b70",
          2052 => x"81ff065c",
          2053 => x"5a7aff95",
          2054 => x"387f8132",
          2055 => x"61813207",
          2056 => x"5d7c81ee",
          2057 => x"3861ff2e",
          2058 => x"81e8387d",
          2059 => x"518194e1",
          2060 => x"3f83d5ec",
          2061 => x"51d3d13f",
          2062 => x"7e4880f8",
          2063 => x"5380527e",
          2064 => x"51e8bc3f",
          2065 => x"0b0b83ee",
          2066 => x"bc337081",
          2067 => x"ff065b59",
          2068 => x"79fd9138",
          2069 => x"815383d5",
          2070 => x"985284d0",
          2071 => x"d8518288",
          2072 => x"cd3f84b9",
          2073 => x"c80880c5",
          2074 => x"38810b0b",
          2075 => x"0b83eebc",
          2076 => x"3484d0d8",
          2077 => x"5380f852",
          2078 => x"7e5182f6",
          2079 => x"c83f84b9",
          2080 => x"c808802e",
          2081 => x"a03884b9",
          2082 => x"c80851df",
          2083 => x"e63f0b0b",
          2084 => x"83eebc33",
          2085 => x"7081ff06",
          2086 => x"5f597d82",
          2087 => x"2e098106",
          2088 => x"fcd33891",
          2089 => x"3984d0d8",
          2090 => x"5182a1d4",
          2091 => x"3f820b0b",
          2092 => x"0b83eebc",
          2093 => x"3483d5a8",
          2094 => x"5380f852",
          2095 => x"7e51a7d4",
          2096 => x"3f67705a",
          2097 => x"5a79fcb7",
          2098 => x"3890397c",
          2099 => x"1a630c85",
          2100 => x"1b335978",
          2101 => x"818926fd",
          2102 => x"80387810",
          2103 => x"1083bed4",
          2104 => x"055a7908",
          2105 => x"04835383",
          2106 => x"d5f8527e",
          2107 => x"51e4fb3f",
          2108 => x"60537e52",
          2109 => x"84baf451",
          2110 => x"8285843f",
          2111 => x"84b9c808",
          2112 => x"612e0981",
          2113 => x"06fbae38",
          2114 => x"81709a3d",
          2115 => x"454141fb",
          2116 => x"ae3983d5",
          2117 => x"fc51dedb",
          2118 => x"3f7d5181",
          2119 => x"92f33ffe",
          2120 => x"903983d6",
          2121 => x"8c567b55",
          2122 => x"83d69054",
          2123 => x"805383d6",
          2124 => x"94527c51",
          2125 => x"d2f23ffd",
          2126 => x"9339818c",
          2127 => x"ab3ffaff",
          2128 => x"399af83f",
          2129 => x"faf93981",
          2130 => x"528351bf",
          2131 => x"a43ffaef",
          2132 => x"39818dd6",
          2133 => x"3ffae839",
          2134 => x"83d6a451",
          2135 => x"de953f80",
          2136 => x"59780483",
          2137 => x"d6b851de",
          2138 => x"8a3fd0fd",
          2139 => x"3ffad039",
          2140 => x"b83dff84",
          2141 => x"1153ff80",
          2142 => x"0551ec8a",
          2143 => x"3f84b9c8",
          2144 => x"08802efa",
          2145 => x"ba386852",
          2146 => x"83d6d451",
          2147 => x"d0fa3f68",
          2148 => x"5a792d84",
          2149 => x"b9c80880",
          2150 => x"2efaa438",
          2151 => x"84b9c808",
          2152 => x"5283d6f0",
          2153 => x"51d0e13f",
          2154 => x"fa9539b8",
          2155 => x"3dff8411",
          2156 => x"53ff8005",
          2157 => x"51ebcf3f",
          2158 => x"84b9c808",
          2159 => x"802ef9ff",
          2160 => x"38685283",
          2161 => x"d78c51d0",
          2162 => x"bf3f6859",
          2163 => x"7804b83d",
          2164 => x"fef41153",
          2165 => x"ff800551",
          2166 => x"e9a83f84",
          2167 => x"b9c80880",
          2168 => x"2ef9dc38",
          2169 => x"b83dfef0",
          2170 => x"1153ff80",
          2171 => x"0551e992",
          2172 => x"3f84b9c8",
          2173 => x"0886d038",
          2174 => x"64597808",
          2175 => x"53785283",
          2176 => x"d7a851d0",
          2177 => x"833f84d5",
          2178 => x"a8085380",
          2179 => x"f8527e51",
          2180 => x"d0913f7e",
          2181 => x"487e3359",
          2182 => x"78ae2ef9",
          2183 => x"a238789f",
          2184 => x"2687d338",
          2185 => x"64840570",
          2186 => x"4659cf39",
          2187 => x"b83dfef4",
          2188 => x"1153ff80",
          2189 => x"0551e8ca",
          2190 => x"3f84b9c8",
          2191 => x"08802ef8",
          2192 => x"fe38b83d",
          2193 => x"fef01153",
          2194 => x"ff800551",
          2195 => x"e8b43f84",
          2196 => x"b9c80886",
          2197 => x"b0386459",
          2198 => x"78225378",
          2199 => x"5283d7b8",
          2200 => x"51cfa53f",
          2201 => x"84d5a808",
          2202 => x"5380f852",
          2203 => x"7e51cfb3",
          2204 => x"3f7e487e",
          2205 => x"335978ae",
          2206 => x"2ef8c438",
          2207 => x"789f2687",
          2208 => x"ca386482",
          2209 => x"05704659",
          2210 => x"cf39b83d",
          2211 => x"ff841153",
          2212 => x"ff800551",
          2213 => x"e9f03f84",
          2214 => x"b9c80880",
          2215 => x"2ef8a038",
          2216 => x"b83dfefc",
          2217 => x"1153ff80",
          2218 => x"0551e9da",
          2219 => x"3f84b9c8",
          2220 => x"08802ef8",
          2221 => x"8a38b83d",
          2222 => x"fef81153",
          2223 => x"ff800551",
          2224 => x"e9c43f84",
          2225 => x"b9c80880",
          2226 => x"2ef7f438",
          2227 => x"83d7c451",
          2228 => x"ceb63f68",
          2229 => x"675d5978",
          2230 => x"7c27838d",
          2231 => x"38657033",
          2232 => x"7a335f5c",
          2233 => x"5a7a7d2e",
          2234 => x"95387a55",
          2235 => x"79547833",
          2236 => x"53785283",
          2237 => x"d7d451ce",
          2238 => x"8f3f6666",
          2239 => x"5b5c8119",
          2240 => x"811b4759",
          2241 => x"d239b83d",
          2242 => x"ff841153",
          2243 => x"ff800551",
          2244 => x"e8f43f84",
          2245 => x"b9c80880",
          2246 => x"2ef7a438",
          2247 => x"b83dfefc",
          2248 => x"1153ff80",
          2249 => x"0551e8de",
          2250 => x"3f84b9c8",
          2251 => x"08802ef7",
          2252 => x"8e38b83d",
          2253 => x"fef81153",
          2254 => x"ff800551",
          2255 => x"e8c83f84",
          2256 => x"b9c80880",
          2257 => x"2ef6f838",
          2258 => x"83d7f051",
          2259 => x"cdba3f68",
          2260 => x"5a796727",
          2261 => x"82933865",
          2262 => x"5c797081",
          2263 => x"055b337c",
          2264 => x"34658105",
          2265 => x"46eb39b8",
          2266 => x"3dff8411",
          2267 => x"53ff8005",
          2268 => x"51e8933f",
          2269 => x"84b9c808",
          2270 => x"802ef6c3",
          2271 => x"38b83dfe",
          2272 => x"fc1153ff",
          2273 => x"800551e7",
          2274 => x"fd3f84b9",
          2275 => x"c808b138",
          2276 => x"68703354",
          2277 => x"5283d7fc",
          2278 => x"51cced3f",
          2279 => x"84d5a808",
          2280 => x"5380f852",
          2281 => x"7e51ccfb",
          2282 => x"3f7e487e",
          2283 => x"335978ae",
          2284 => x"2ef68c38",
          2285 => x"789f2684",
          2286 => x"97386881",
          2287 => x"0549d139",
          2288 => x"68590280",
          2289 => x"db053379",
          2290 => x"34688105",
          2291 => x"49b83dfe",
          2292 => x"fc1153ff",
          2293 => x"800551e7",
          2294 => x"ad3f84b9",
          2295 => x"c808802e",
          2296 => x"f5dd3868",
          2297 => x"590280db",
          2298 => x"05337934",
          2299 => x"68810549",
          2300 => x"b83dfefc",
          2301 => x"1153ff80",
          2302 => x"0551e78a",
          2303 => x"3f84b9c8",
          2304 => x"08ffbd38",
          2305 => x"f5b939b8",
          2306 => x"3dff8411",
          2307 => x"53ff8005",
          2308 => x"51e6f33f",
          2309 => x"84b9c808",
          2310 => x"802ef5a3",
          2311 => x"38b83dfe",
          2312 => x"fc1153ff",
          2313 => x"800551e6",
          2314 => x"dd3f84b9",
          2315 => x"c808802e",
          2316 => x"f58d38b8",
          2317 => x"3dfef811",
          2318 => x"53ff8005",
          2319 => x"51e6c73f",
          2320 => x"84b9c808",
          2321 => x"863884b9",
          2322 => x"c8084683",
          2323 => x"d88851cb",
          2324 => x"b73f6867",
          2325 => x"5b59787a",
          2326 => x"278f3865",
          2327 => x"5b7a7970",
          2328 => x"84055b0c",
          2329 => x"797926f5",
          2330 => x"388a51d9",
          2331 => x"f13ff4cf",
          2332 => x"39b83dff",
          2333 => x"80055187",
          2334 => x"b13f84b9",
          2335 => x"c808b93d",
          2336 => x"ff800552",
          2337 => x"5988f33f",
          2338 => x"815384b9",
          2339 => x"c8085278",
          2340 => x"51ea833f",
          2341 => x"84b9c808",
          2342 => x"802ef4a3",
          2343 => x"3884b9c8",
          2344 => x"0851e7f6",
          2345 => x"3ff49839",
          2346 => x"b83dff84",
          2347 => x"1153ff80",
          2348 => x"0551e5d2",
          2349 => x"3f84b9c8",
          2350 => x"08913883",
          2351 => x"f2cc335a",
          2352 => x"79802e83",
          2353 => x"c03883f2",
          2354 => x"840849b8",
          2355 => x"3dfefc11",
          2356 => x"53ff8005",
          2357 => x"51e5af3f",
          2358 => x"84b9c808",
          2359 => x"913883f2",
          2360 => x"cc335a79",
          2361 => x"802e838a",
          2362 => x"3883f288",
          2363 => x"0847b83d",
          2364 => x"fef81153",
          2365 => x"ff800551",
          2366 => x"e58c3f84",
          2367 => x"b9c80880",
          2368 => x"2ea53880",
          2369 => x"665c5c7a",
          2370 => x"882e8338",
          2371 => x"815c7a90",
          2372 => x"32703070",
          2373 => x"72079f2a",
          2374 => x"7e065c5f",
          2375 => x"5d79802e",
          2376 => x"88387aa0",
          2377 => x"2e833888",
          2378 => x"4683d898",
          2379 => x"51d6c43f",
          2380 => x"80556854",
          2381 => x"65536652",
          2382 => x"6851eba8",
          2383 => x"3f83d8a4",
          2384 => x"51d6b03f",
          2385 => x"f2f93964",
          2386 => x"64710c59",
          2387 => x"64840545",
          2388 => x"b83dfef0",
          2389 => x"1153ff80",
          2390 => x"0551e2a6",
          2391 => x"3f84b9c8",
          2392 => x"08802ef2",
          2393 => x"da386464",
          2394 => x"710c5964",
          2395 => x"840545b8",
          2396 => x"3dfef011",
          2397 => x"53ff8005",
          2398 => x"51e2873f",
          2399 => x"84b9c808",
          2400 => x"c638f2bb",
          2401 => x"39645e02",
          2402 => x"80ce0522",
          2403 => x"7e708205",
          2404 => x"40237d45",
          2405 => x"b83dfef0",
          2406 => x"1153ff80",
          2407 => x"0551e1e2",
          2408 => x"3f84b9c8",
          2409 => x"08802ef2",
          2410 => x"9638645e",
          2411 => x"0280ce05",
          2412 => x"227e7082",
          2413 => x"0540237d",
          2414 => x"45b83dfe",
          2415 => x"f01153ff",
          2416 => x"800551e1",
          2417 => x"bd3f84b9",
          2418 => x"c808ffb9",
          2419 => x"38f1f039",
          2420 => x"b83dfefc",
          2421 => x"1153ff80",
          2422 => x"0551e3aa",
          2423 => x"3f84b9c8",
          2424 => x"08802e81",
          2425 => x"dc38685c",
          2426 => x"0280db05",
          2427 => x"337c3468",
          2428 => x"810549fb",
          2429 => x"9b39b83d",
          2430 => x"fef01153",
          2431 => x"ff800551",
          2432 => x"e1803f84",
          2433 => x"b9c80880",
          2434 => x"2e819838",
          2435 => x"6464710c",
          2436 => x"5d648405",
          2437 => x"704659f7",
          2438 => x"e1397a83",
          2439 => x"2e098106",
          2440 => x"f39d387b",
          2441 => x"5583d690",
          2442 => x"54805383",
          2443 => x"d8b0527c",
          2444 => x"51c8f53f",
          2445 => x"f396397b",
          2446 => x"527c51da",
          2447 => x"8a3ff38c",
          2448 => x"3983d8bc",
          2449 => x"51d4ac3f",
          2450 => x"f0f539b8",
          2451 => x"3dfef011",
          2452 => x"53ff8005",
          2453 => x"51e0ab3f",
          2454 => x"84b9c808",
          2455 => x"802eb838",
          2456 => x"64590280",
          2457 => x"ce052279",
          2458 => x"7082055b",
          2459 => x"237845f7",
          2460 => x"e73983f2",
          2461 => x"cd335c7b",
          2462 => x"802e80cf",
          2463 => x"3883f290",
          2464 => x"0847fcea",
          2465 => x"3983f2cd",
          2466 => x"335c7b80",
          2467 => x"2ea13883",
          2468 => x"f28c0849",
          2469 => x"fcb53983",
          2470 => x"d8e851d3",
          2471 => x"d63f6459",
          2472 => x"f7b63983",
          2473 => x"d8e851d3",
          2474 => x"ca3f6459",
          2475 => x"f6cc3983",
          2476 => x"f2ce3359",
          2477 => x"78802ea5",
          2478 => x"3883f294",
          2479 => x"0849fc8b",
          2480 => x"3983d8e8",
          2481 => x"51d3ac3f",
          2482 => x"f9c63983",
          2483 => x"f2ce3359",
          2484 => x"78802e9b",
          2485 => x"3883f298",
          2486 => x"0847fc92",
          2487 => x"3983f2cf",
          2488 => x"335e7d80",
          2489 => x"2e9b3883",
          2490 => x"f29c0849",
          2491 => x"fbdd3983",
          2492 => x"f2cf335e",
          2493 => x"7d802e9b",
          2494 => x"3883f2a0",
          2495 => x"0847fbee",
          2496 => x"3983f2ca",
          2497 => x"335d7c80",
          2498 => x"2e9b3883",
          2499 => x"f2a40849",
          2500 => x"fbb93983",
          2501 => x"f2ca335d",
          2502 => x"7c802e94",
          2503 => x"3883f2a8",
          2504 => x"0847fbca",
          2505 => x"3983f2b4",
          2506 => x"08fc8005",
          2507 => x"49fb9c39",
          2508 => x"83f2b408",
          2509 => x"880547fb",
          2510 => x"b539f33d",
          2511 => x"0d800b84",
          2512 => x"b9f83487",
          2513 => x"c0948c70",
          2514 => x"08565787",
          2515 => x"84805274",
          2516 => x"51dad23f",
          2517 => x"84b9c808",
          2518 => x"902b7708",
          2519 => x"57558784",
          2520 => x"80527551",
          2521 => x"dabf3f74",
          2522 => x"84b9c808",
          2523 => x"07770c87",
          2524 => x"c0949c70",
          2525 => x"08565787",
          2526 => x"84805274",
          2527 => x"51daa63f",
          2528 => x"84b9c808",
          2529 => x"902b7708",
          2530 => x"57558784",
          2531 => x"80527551",
          2532 => x"da933f74",
          2533 => x"84b9c808",
          2534 => x"07770c8c",
          2535 => x"80830b87",
          2536 => x"c094840c",
          2537 => x"8c80830b",
          2538 => x"87c09494",
          2539 => x"0c81bcf2",
          2540 => x"5c81c7f1",
          2541 => x"5d830284",
          2542 => x"05a10534",
          2543 => x"805e84d5",
          2544 => x"a80b893d",
          2545 => x"7088130c",
          2546 => x"70720c84",
          2547 => x"d5ac0c56",
          2548 => x"b7853f89",
          2549 => x"9e3f9597",
          2550 => x"3fba8d51",
          2551 => x"958c3f83",
          2552 => x"d2b05283",
          2553 => x"d2b451c4",
          2554 => x"9f3f83f2",
          2555 => x"b8702252",
          2556 => x"5594973f",
          2557 => x"83d2bc54",
          2558 => x"83d2c853",
          2559 => x"81153352",
          2560 => x"83d2d051",
          2561 => x"c4823f8d",
          2562 => x"b23f83d2",
          2563 => x"ec51d0e3",
          2564 => x"3f805283",
          2565 => x"d2f051c3",
          2566 => x"ef3f9080",
          2567 => x"0a5283d3",
          2568 => x"9851c3e4",
          2569 => x"3fece73f",
          2570 => x"8004fb3d",
          2571 => x"0d777008",
          2572 => x"56568075",
          2573 => x"52537473",
          2574 => x"2e818338",
          2575 => x"74337081",
          2576 => x"ff065252",
          2577 => x"70a02e09",
          2578 => x"81069138",
          2579 => x"81157033",
          2580 => x"7081ff06",
          2581 => x"53535570",
          2582 => x"a02ef138",
          2583 => x"7181ff06",
          2584 => x"5473a22e",
          2585 => x"81823874",
          2586 => x"5272812e",
          2587 => x"80e73880",
          2588 => x"72337081",
          2589 => x"ff065354",
          2590 => x"5470a02e",
          2591 => x"83388154",
          2592 => x"70802e8b",
          2593 => x"3873802e",
          2594 => x"86388112",
          2595 => x"52e13980",
          2596 => x"7381ff06",
          2597 => x"525470a0",
          2598 => x"2e098106",
          2599 => x"83388154",
          2600 => x"70a23270",
          2601 => x"30708025",
          2602 => x"76075252",
          2603 => x"5372802e",
          2604 => x"88388072",
          2605 => x"70810554",
          2606 => x"3471760c",
          2607 => x"74517084",
          2608 => x"b9c80c87",
          2609 => x"3d0d0470",
          2610 => x"802ec438",
          2611 => x"73802eff",
          2612 => x"be388112",
          2613 => x"52807233",
          2614 => x"7081ff06",
          2615 => x"53545470",
          2616 => x"a22ee438",
          2617 => x"8154e039",
          2618 => x"81155581",
          2619 => x"75535372",
          2620 => x"812e0981",
          2621 => x"06fef838",
          2622 => x"dc39fc3d",
          2623 => x"0d765372",
          2624 => x"088b3880",
          2625 => x"0b84b9c8",
          2626 => x"0c863d0d",
          2627 => x"04863dfc",
          2628 => x"05527251",
          2629 => x"daec3f84",
          2630 => x"b9c80880",
          2631 => x"2ee53874",
          2632 => x"84b9c80c",
          2633 => x"863d0d04",
          2634 => x"fc3d0d76",
          2635 => x"821133ff",
          2636 => x"05525381",
          2637 => x"52708b26",
          2638 => x"81983883",
          2639 => x"1333ff05",
          2640 => x"54825273",
          2641 => x"9e26818a",
          2642 => x"38841333",
          2643 => x"51835270",
          2644 => x"972680fe",
          2645 => x"38851333",
          2646 => x"54845273",
          2647 => x"bb2680f2",
          2648 => x"38861333",
          2649 => x"55855274",
          2650 => x"bb2680e6",
          2651 => x"38881322",
          2652 => x"55865274",
          2653 => x"87e72680",
          2654 => x"d9388a13",
          2655 => x"22548752",
          2656 => x"7387e726",
          2657 => x"80cc3881",
          2658 => x"0b87c098",
          2659 => x"9c0c7222",
          2660 => x"87c098bc",
          2661 => x"0c821333",
          2662 => x"87c098b8",
          2663 => x"0c831333",
          2664 => x"87c098b4",
          2665 => x"0c841333",
          2666 => x"87c098b0",
          2667 => x"0c851333",
          2668 => x"87c098ac",
          2669 => x"0c861333",
          2670 => x"87c098a8",
          2671 => x"0c7487c0",
          2672 => x"98a40c73",
          2673 => x"87c098a0",
          2674 => x"0c800b87",
          2675 => x"c0989c0c",
          2676 => x"80527184",
          2677 => x"b9c80c86",
          2678 => x"3d0d04f3",
          2679 => x"3d0d7f5b",
          2680 => x"87c0989c",
          2681 => x"5d817d0c",
          2682 => x"87c098bc",
          2683 => x"085e7d7b",
          2684 => x"2387c098",
          2685 => x"b8085c7b",
          2686 => x"821c3487",
          2687 => x"c098b408",
          2688 => x"5a79831c",
          2689 => x"3487c098",
          2690 => x"b0085c7b",
          2691 => x"841c3487",
          2692 => x"c098ac08",
          2693 => x"5a79851c",
          2694 => x"3487c098",
          2695 => x"a8085c7b",
          2696 => x"861c3487",
          2697 => x"c098a408",
          2698 => x"5c7b881c",
          2699 => x"2387c098",
          2700 => x"a0085a79",
          2701 => x"8a1c2380",
          2702 => x"7d0c7983",
          2703 => x"ffff0659",
          2704 => x"7b83ffff",
          2705 => x"0658861b",
          2706 => x"3357851b",
          2707 => x"3356841b",
          2708 => x"3355831b",
          2709 => x"3354821b",
          2710 => x"33537d83",
          2711 => x"ffff0652",
          2712 => x"83d8ec51",
          2713 => x"ffbfa13f",
          2714 => x"8f3d0d04",
          2715 => x"fe3d0d02",
          2716 => x"93053353",
          2717 => x"72812ea8",
          2718 => x"38725180",
          2719 => x"e8a63f84",
          2720 => x"b9c80898",
          2721 => x"2b70982c",
          2722 => x"515271ff",
          2723 => x"2e098106",
          2724 => x"86387283",
          2725 => x"2ee33871",
          2726 => x"84b9c80c",
          2727 => x"843d0d04",
          2728 => x"725180e7",
          2729 => x"ff3f84b9",
          2730 => x"c808982b",
          2731 => x"70982c51",
          2732 => x"5271ff2e",
          2733 => x"098106df",
          2734 => x"38725180",
          2735 => x"e7e63f84",
          2736 => x"b9c80898",
          2737 => x"2b70982c",
          2738 => x"515271ff",
          2739 => x"2ed238c7",
          2740 => x"39fd3d0d",
          2741 => x"80705452",
          2742 => x"71882b54",
          2743 => x"815180e7",
          2744 => x"c33f84b9",
          2745 => x"c808982b",
          2746 => x"70982c51",
          2747 => x"5271ff2e",
          2748 => x"eb387372",
          2749 => x"07811454",
          2750 => x"52837325",
          2751 => x"db387184",
          2752 => x"b9c80c85",
          2753 => x"3d0d04fc",
          2754 => x"3d0d029b",
          2755 => x"053383f2",
          2756 => x"80337081",
          2757 => x"ff065355",
          2758 => x"5570802e",
          2759 => x"80f43887",
          2760 => x"c0949408",
          2761 => x"70962a70",
          2762 => x"81065354",
          2763 => x"5270802e",
          2764 => x"8c387191",
          2765 => x"2a708106",
          2766 => x"515170e3",
          2767 => x"38728132",
          2768 => x"81065372",
          2769 => x"802e8a38",
          2770 => x"71932a81",
          2771 => x"065271cf",
          2772 => x"387381ff",
          2773 => x"065187c0",
          2774 => x"94805270",
          2775 => x"802e8638",
          2776 => x"87c09490",
          2777 => x"5274720c",
          2778 => x"7484b9c8",
          2779 => x"0c863d0d",
          2780 => x"0471912a",
          2781 => x"70810651",
          2782 => x"51709738",
          2783 => x"72813281",
          2784 => x"06537280",
          2785 => x"2ecb3871",
          2786 => x"932a8106",
          2787 => x"5271802e",
          2788 => x"c03887c0",
          2789 => x"94840870",
          2790 => x"962a7081",
          2791 => x"06535452",
          2792 => x"70cf38d8",
          2793 => x"39ff3d0d",
          2794 => x"028f0533",
          2795 => x"7030709f",
          2796 => x"2a515252",
          2797 => x"7083f280",
          2798 => x"34833d0d",
          2799 => x"04fa3d0d",
          2800 => x"78558075",
          2801 => x"33705652",
          2802 => x"5770772e",
          2803 => x"80e73881",
          2804 => x"1583f280",
          2805 => x"337081ff",
          2806 => x"06545755",
          2807 => x"71802e80",
          2808 => x"ff3887c0",
          2809 => x"94940870",
          2810 => x"962a7081",
          2811 => x"06535452",
          2812 => x"70802e8c",
          2813 => x"3871912a",
          2814 => x"70810651",
          2815 => x"5170e338",
          2816 => x"72813281",
          2817 => x"06537280",
          2818 => x"2e8a3871",
          2819 => x"932a8106",
          2820 => x"5271cf38",
          2821 => x"7581ff06",
          2822 => x"5187c094",
          2823 => x"80527080",
          2824 => x"2e863887",
          2825 => x"c0949052",
          2826 => x"73720c81",
          2827 => x"17753355",
          2828 => x"5773ff9b",
          2829 => x"387684b9",
          2830 => x"c80c883d",
          2831 => x"0d047191",
          2832 => x"2a708106",
          2833 => x"51517098",
          2834 => x"38728132",
          2835 => x"81065372",
          2836 => x"802ec138",
          2837 => x"71932a81",
          2838 => x"06527180",
          2839 => x"2effb538",
          2840 => x"87c09484",
          2841 => x"0870962a",
          2842 => x"70810653",
          2843 => x"545270ce",
          2844 => x"38d739ff",
          2845 => x"3d0d87c0",
          2846 => x"9e800870",
          2847 => x"9c2a8a06",
          2848 => x"52527080",
          2849 => x"2e84ab38",
          2850 => x"87c09ea4",
          2851 => x"0883f284",
          2852 => x"0c87c09e",
          2853 => x"a80883f2",
          2854 => x"880c87c0",
          2855 => x"9e940883",
          2856 => x"f28c0c87",
          2857 => x"c09e9808",
          2858 => x"83f2900c",
          2859 => x"87c09e9c",
          2860 => x"0883f294",
          2861 => x"0c87c09e",
          2862 => x"a00883f2",
          2863 => x"980c87c0",
          2864 => x"9eac0883",
          2865 => x"f29c0c87",
          2866 => x"c09eb008",
          2867 => x"83f2a00c",
          2868 => x"87c09eb4",
          2869 => x"0883f2a4",
          2870 => x"0c87c09e",
          2871 => x"b80883f2",
          2872 => x"a80c87c0",
          2873 => x"9ebc0883",
          2874 => x"f2ac0c87",
          2875 => x"c09ec008",
          2876 => x"83f2b00c",
          2877 => x"87c09ec4",
          2878 => x"0883f2b4",
          2879 => x"0c87c09e",
          2880 => x"80085271",
          2881 => x"83f2b823",
          2882 => x"87c09e84",
          2883 => x"0883f2bc",
          2884 => x"0c87c09e",
          2885 => x"880883f2",
          2886 => x"c00c87c0",
          2887 => x"9e8c0883",
          2888 => x"f2c40c81",
          2889 => x"0b83f2c8",
          2890 => x"34800b87",
          2891 => x"c09e9008",
          2892 => x"7084800a",
          2893 => x"06515252",
          2894 => x"7082fb38",
          2895 => x"7183f2c9",
          2896 => x"34800b87",
          2897 => x"c09e9008",
          2898 => x"7088800a",
          2899 => x"06515252",
          2900 => x"70802e83",
          2901 => x"38815271",
          2902 => x"83f2ca34",
          2903 => x"800b87c0",
          2904 => x"9e900870",
          2905 => x"90800a06",
          2906 => x"51525270",
          2907 => x"802e8338",
          2908 => x"81527183",
          2909 => x"f2cb3480",
          2910 => x"0b87c09e",
          2911 => x"90087088",
          2912 => x"80800651",
          2913 => x"52527080",
          2914 => x"2e833881",
          2915 => x"527183f2",
          2916 => x"cc34800b",
          2917 => x"87c09e90",
          2918 => x"0870a080",
          2919 => x"80065152",
          2920 => x"5270802e",
          2921 => x"83388152",
          2922 => x"7183f2cd",
          2923 => x"34800b87",
          2924 => x"c09e9008",
          2925 => x"70908080",
          2926 => x"06515252",
          2927 => x"70802e83",
          2928 => x"38815271",
          2929 => x"83f2ce34",
          2930 => x"800b87c0",
          2931 => x"9e900870",
          2932 => x"84808006",
          2933 => x"51525270",
          2934 => x"802e8338",
          2935 => x"81527183",
          2936 => x"f2cf3480",
          2937 => x"0b87c09e",
          2938 => x"90087082",
          2939 => x"80800651",
          2940 => x"52527080",
          2941 => x"2e833881",
          2942 => x"527183f2",
          2943 => x"d034800b",
          2944 => x"87c09e90",
          2945 => x"08708180",
          2946 => x"80065152",
          2947 => x"5270802e",
          2948 => x"83388152",
          2949 => x"7183f2d1",
          2950 => x"34800b87",
          2951 => x"c09e9008",
          2952 => x"7080c080",
          2953 => x"06515252",
          2954 => x"70802e83",
          2955 => x"38815271",
          2956 => x"83f2d234",
          2957 => x"800b87c0",
          2958 => x"9e900870",
          2959 => x"a0800651",
          2960 => x"52527080",
          2961 => x"2e833881",
          2962 => x"527183f2",
          2963 => x"d33487c0",
          2964 => x"9e900898",
          2965 => x"8006708a",
          2966 => x"2a535171",
          2967 => x"83f2d434",
          2968 => x"800b87c0",
          2969 => x"9e900870",
          2970 => x"84800651",
          2971 => x"52527080",
          2972 => x"2e833881",
          2973 => x"527183f2",
          2974 => x"d53487c0",
          2975 => x"9e900883",
          2976 => x"f0067084",
          2977 => x"2a535171",
          2978 => x"83f2d634",
          2979 => x"800b87c0",
          2980 => x"9e900870",
          2981 => x"88065152",
          2982 => x"5270802e",
          2983 => x"83388152",
          2984 => x"7183f2d7",
          2985 => x"3487c09e",
          2986 => x"90088706",
          2987 => x"517083f2",
          2988 => x"d834833d",
          2989 => x"0d048152",
          2990 => x"fd8239fb",
          2991 => x"3d0d83d9",
          2992 => x"8451ffb6",
          2993 => x"c33f83f2",
          2994 => x"c8335473",
          2995 => x"869f3883",
          2996 => x"d99851c3",
          2997 => x"9e3f83f2",
          2998 => x"ca335574",
          2999 => x"85ef3883",
          3000 => x"f2cf3354",
          3001 => x"7385c638",
          3002 => x"83f2cc33",
          3003 => x"5675859d",
          3004 => x"3883f2cd",
          3005 => x"33557484",
          3006 => x"f43883f2",
          3007 => x"ce335473",
          3008 => x"84cb3883",
          3009 => x"f2d33356",
          3010 => x"7584a838",
          3011 => x"83f2d733",
          3012 => x"54738485",
          3013 => x"3883f2d5",
          3014 => x"33557483",
          3015 => x"e23883f2",
          3016 => x"c9335675",
          3017 => x"83c43883",
          3018 => x"f2cb3354",
          3019 => x"7383a638",
          3020 => x"83f2d033",
          3021 => x"55748388",
          3022 => x"3883f2d1",
          3023 => x"33567582",
          3024 => x"e93883f2",
          3025 => x"d2335473",
          3026 => x"81e13883",
          3027 => x"d9b051c2",
          3028 => x"a23f83f2",
          3029 => x"ac085283",
          3030 => x"d9bc51ff",
          3031 => x"b5aa3f83",
          3032 => x"f2b00852",
          3033 => x"83d9e451",
          3034 => x"ffb59d3f",
          3035 => x"83f2b408",
          3036 => x"5283da8c",
          3037 => x"51ffb590",
          3038 => x"3f83dab4",
          3039 => x"51c1f43f",
          3040 => x"83f2b822",
          3041 => x"5283dabc",
          3042 => x"51ffb4fc",
          3043 => x"3f83f2bc",
          3044 => x"0856bd84",
          3045 => x"c0527551",
          3046 => x"ca8b3f84",
          3047 => x"b9c808bd",
          3048 => x"84c02976",
          3049 => x"71315454",
          3050 => x"84b9c808",
          3051 => x"5283dae4",
          3052 => x"51ffb4d4",
          3053 => x"3f83f2cf",
          3054 => x"335574b9",
          3055 => x"3883f2ca",
          3056 => x"33557485",
          3057 => x"38873d0d",
          3058 => x"0483f2c4",
          3059 => x"0856bd84",
          3060 => x"c0527551",
          3061 => x"c9cf3f84",
          3062 => x"b9c808bd",
          3063 => x"84c02976",
          3064 => x"71315454",
          3065 => x"84b9c808",
          3066 => x"5283db90",
          3067 => x"51ffb498",
          3068 => x"3f873d0d",
          3069 => x"0483f2c0",
          3070 => x"0856bd84",
          3071 => x"c0527551",
          3072 => x"c9a33f84",
          3073 => x"b9c808bd",
          3074 => x"84c02976",
          3075 => x"71315454",
          3076 => x"84b9c808",
          3077 => x"5283dbbc",
          3078 => x"51ffb3ec",
          3079 => x"3f83f2ca",
          3080 => x"33557480",
          3081 => x"2eff9e38",
          3082 => x"ff9f3983",
          3083 => x"dbe851c0",
          3084 => x"c23f83d9",
          3085 => x"b051c0bb",
          3086 => x"3f83f2ac",
          3087 => x"085283d9",
          3088 => x"bc51ffb3",
          3089 => x"c33f83f2",
          3090 => x"b0085283",
          3091 => x"d9e451ff",
          3092 => x"b3b63f83",
          3093 => x"f2b40852",
          3094 => x"83da8c51",
          3095 => x"ffb3a93f",
          3096 => x"83dab451",
          3097 => x"c08d3f83",
          3098 => x"f2b82252",
          3099 => x"83dabc51",
          3100 => x"ffb3953f",
          3101 => x"83f2bc08",
          3102 => x"56bd84c0",
          3103 => x"527551c8",
          3104 => x"a43f84b9",
          3105 => x"c808bd84",
          3106 => x"c0297671",
          3107 => x"31545484",
          3108 => x"b9c80852",
          3109 => x"83dae451",
          3110 => x"ffb2ed3f",
          3111 => x"83f2cf33",
          3112 => x"5574802e",
          3113 => x"fe9738fe",
          3114 => x"cc3983db",
          3115 => x"f051ffbf",
          3116 => x"c23f83f2",
          3117 => x"d2335473",
          3118 => x"802efd8f",
          3119 => x"38feec39",
          3120 => x"83dbf851",
          3121 => x"ffbfac3f",
          3122 => x"83f2d133",
          3123 => x"5675802e",
          3124 => x"fcf038d6",
          3125 => x"3983dc84",
          3126 => x"51ffbf97",
          3127 => x"3f83f2d0",
          3128 => x"33557480",
          3129 => x"2efcd238",
          3130 => x"d73983dc",
          3131 => x"9051ffbf",
          3132 => x"823f83f2",
          3133 => x"cb335473",
          3134 => x"802efcb4",
          3135 => x"38d73983",
          3136 => x"f2d63352",
          3137 => x"83dca451",
          3138 => x"ffb1fd3f",
          3139 => x"83f2c933",
          3140 => x"5675802e",
          3141 => x"fc9138d2",
          3142 => x"3983f2d8",
          3143 => x"335283dc",
          3144 => x"c451ffb1",
          3145 => x"e33f83f2",
          3146 => x"d5335574",
          3147 => x"802efbee",
          3148 => x"38cd3983",
          3149 => x"f2d43352",
          3150 => x"83dce451",
          3151 => x"ffb1c93f",
          3152 => x"83f2d733",
          3153 => x"5473802e",
          3154 => x"fbcb38cd",
          3155 => x"3983f294",
          3156 => x"0883f298",
          3157 => x"08115452",
          3158 => x"83dd8451",
          3159 => x"ffb1a93f",
          3160 => x"83f2d333",
          3161 => x"5675802e",
          3162 => x"fba238c7",
          3163 => x"3983f28c",
          3164 => x"0883f290",
          3165 => x"08115452",
          3166 => x"83dda051",
          3167 => x"ffb1893f",
          3168 => x"83f2ce33",
          3169 => x"5473802e",
          3170 => x"faf938c1",
          3171 => x"3983f284",
          3172 => x"0883f288",
          3173 => x"08115452",
          3174 => x"83ddbc51",
          3175 => x"ffb0e93f",
          3176 => x"83f2cd33",
          3177 => x"5574802e",
          3178 => x"fad038c1",
          3179 => x"3983f29c",
          3180 => x"0883f2a0",
          3181 => x"08115452",
          3182 => x"83ddd851",
          3183 => x"ffb0c93f",
          3184 => x"83f2cc33",
          3185 => x"5675802e",
          3186 => x"faa738c1",
          3187 => x"3983f2a4",
          3188 => x"0883f2a8",
          3189 => x"08115452",
          3190 => x"83ddf451",
          3191 => x"ffb0a93f",
          3192 => x"83f2cf33",
          3193 => x"5473802e",
          3194 => x"f9fe38c1",
          3195 => x"3983de90",
          3196 => x"51ffb094",
          3197 => x"3f83d998",
          3198 => x"51ffbcf7",
          3199 => x"3f83f2ca",
          3200 => x"33557480",
          3201 => x"2ef9d838",
          3202 => x"c439ff3d",
          3203 => x"0d028e05",
          3204 => x"33527185",
          3205 => x"268c3871",
          3206 => x"101083c2",
          3207 => x"fc055271",
          3208 => x"080483de",
          3209 => x"a451ffaf",
          3210 => x"df3f833d",
          3211 => x"0d0483de",
          3212 => x"ac51ffaf",
          3213 => x"d33f833d",
          3214 => x"0d0483de",
          3215 => x"b451ffaf",
          3216 => x"c73f833d",
          3217 => x"0d0483de",
          3218 => x"bc51ffaf",
          3219 => x"bb3f833d",
          3220 => x"0d0483de",
          3221 => x"c451ffaf",
          3222 => x"af3f833d",
          3223 => x"0d0483de",
          3224 => x"cc51ffaf",
          3225 => x"a33f833d",
          3226 => x"0d047188",
          3227 => x"800c0480",
          3228 => x"0b87c096",
          3229 => x"840c0483",
          3230 => x"f2dc0887",
          3231 => x"c096840c",
          3232 => x"04d93d0d",
          3233 => x"aa3d08ad",
          3234 => x"3d085a5a",
          3235 => x"81705758",
          3236 => x"805283f3",
          3237 => x"b4085182",
          3238 => x"88833f84",
          3239 => x"b9c80880",
          3240 => x"ed388b3d",
          3241 => x"57ff0b83",
          3242 => x"f3b40854",
          3243 => x"5580f852",
          3244 => x"765182d2",
          3245 => x"903f84b9",
          3246 => x"c808802e",
          3247 => x"a4387651",
          3248 => x"c0e63f84",
          3249 => x"b9c80881",
          3250 => x"17575580",
          3251 => x"0b84b9c8",
          3252 => x"08258e38",
          3253 => x"84b9c808",
          3254 => x"ff057018",
          3255 => x"55558074",
          3256 => x"34740970",
          3257 => x"30707207",
          3258 => x"9f2a5155",
          3259 => x"5578762e",
          3260 => x"853873ff",
          3261 => x"b03883f3",
          3262 => x"b4088c11",
          3263 => x"08535182",
          3264 => x"879b3f84",
          3265 => x"b9c8088f",
          3266 => x"3878762e",
          3267 => x"9a387784",
          3268 => x"b9c80ca9",
          3269 => x"3d0d0483",
          3270 => x"e1fc51ff",
          3271 => x"adea3f78",
          3272 => x"762e0981",
          3273 => x"06e83876",
          3274 => x"527951c0",
          3275 => x"9a3f7951",
          3276 => x"ffbff53f",
          3277 => x"ab3d0856",
          3278 => x"84b9c808",
          3279 => x"76347652",
          3280 => x"83e2a851",
          3281 => x"ffadc13f",
          3282 => x"800b84b9",
          3283 => x"c80ca93d",
          3284 => x"0d04d83d",
          3285 => x"0dab3d08",
          3286 => x"ad3d0871",
          3287 => x"725d7233",
          3288 => x"57575a57",
          3289 => x"73a02e81",
          3290 => x"9138800b",
          3291 => x"8d3d5956",
          3292 => x"75101010",
          3293 => x"83f3bc05",
          3294 => x"70085254",
          3295 => x"ffbfa93f",
          3296 => x"84b9c808",
          3297 => x"53795273",
          3298 => x"0851c089",
          3299 => x"3f84b9c8",
          3300 => x"08903884",
          3301 => x"14335473",
          3302 => x"812e8188",
          3303 => x"3873822e",
          3304 => x"99388116",
          3305 => x"7081ff06",
          3306 => x"57548276",
          3307 => x"27c23880",
          3308 => x"547384b9",
          3309 => x"c80caa3d",
          3310 => x"0d04811a",
          3311 => x"5aaa3dff",
          3312 => x"841153ff",
          3313 => x"800551c7",
          3314 => x"bd3f84b9",
          3315 => x"c808802e",
          3316 => x"d138ff1b",
          3317 => x"53785276",
          3318 => x"51fda63f",
          3319 => x"84b9c808",
          3320 => x"81ff0654",
          3321 => x"73802ec9",
          3322 => x"38811670",
          3323 => x"81ff0657",
          3324 => x"54827627",
          3325 => x"fefa38ff",
          3326 => x"b6397833",
          3327 => x"77055676",
          3328 => x"7627fee6",
          3329 => x"38811570",
          3330 => x"5b703355",
          3331 => x"5573a02e",
          3332 => x"098106fe",
          3333 => x"d5387575",
          3334 => x"26eb3880",
          3335 => x"0b8d3d59",
          3336 => x"56fecd39",
          3337 => x"7384b9c8",
          3338 => x"085383f3",
          3339 => x"b4085256",
          3340 => x"8284ea3f",
          3341 => x"84b9c808",
          3342 => x"80d03883",
          3343 => x"f3b40853",
          3344 => x"80f85277",
          3345 => x"5182cefd",
          3346 => x"3f84b9c8",
          3347 => x"08802eba",
          3348 => x"387751ff",
          3349 => x"bdd23f84",
          3350 => x"b9c80855",
          3351 => x"800b84b9",
          3352 => x"c808259d",
          3353 => x"3884b9c8",
          3354 => x"08ff0570",
          3355 => x"19585580",
          3356 => x"77347753",
          3357 => x"75528116",
          3358 => x"83e1f052",
          3359 => x"56ffab88",
          3360 => x"3f74ff2e",
          3361 => x"098106ff",
          3362 => x"b238810b",
          3363 => x"84b9c80c",
          3364 => x"aa3d0d04",
          3365 => x"ce3d0db5",
          3366 => x"3d08b73d",
          3367 => x"08b93d08",
          3368 => x"5a415c80",
          3369 => x"0bb43d34",
          3370 => x"83f3b833",
          3371 => x"83f3b408",
          3372 => x"565d749e",
          3373 => x"387483f3",
          3374 => x"b0335656",
          3375 => x"74802e82",
          3376 => x"cb387780",
          3377 => x"2e918d38",
          3378 => x"81707706",
          3379 => x"5a577890",
          3380 => x"a0387780",
          3381 => x"2e90fd38",
          3382 => x"933db43d",
          3383 => x"5f5f8051",
          3384 => x"eb8a3f84",
          3385 => x"b9c80898",
          3386 => x"2b70982c",
          3387 => x"5b5679ff",
          3388 => x"2eec3879",
          3389 => x"81ff0684",
          3390 => x"d1843370",
          3391 => x"982b7098",
          3392 => x"2c84d180",
          3393 => x"3370982b",
          3394 => x"70972c71",
          3395 => x"982c0570",
          3396 => x"101083de",
          3397 => x"d0057008",
          3398 => x"15703352",
          3399 => x"535c5d46",
          3400 => x"525b585c",
          3401 => x"59815774",
          3402 => x"792e80cd",
          3403 => x"38787527",
          3404 => x"81873875",
          3405 => x"81800a29",
          3406 => x"81ff0a05",
          3407 => x"70982c57",
          3408 => x"55807624",
          3409 => x"81cb3875",
          3410 => x"10167082",
          3411 => x"2b565780",
          3412 => x"0b83ded4",
          3413 => x"16334257",
          3414 => x"77612591",
          3415 => x"3883ded0",
          3416 => x"15081870",
          3417 => x"33564178",
          3418 => x"752e8195",
          3419 => x"3876802e",
          3420 => x"c2387584",
          3421 => x"d1803481",
          3422 => x"5776802e",
          3423 => x"81993881",
          3424 => x"1b70982b",
          3425 => x"70982c84",
          3426 => x"d1803370",
          3427 => x"982b7097",
          3428 => x"2c71982c",
          3429 => x"0570822b",
          3430 => x"83ded411",
          3431 => x"335f535f",
          3432 => x"5d585d57",
          3433 => x"577a782e",
          3434 => x"81903876",
          3435 => x"84d18434",
          3436 => x"feac3981",
          3437 => x"5776ffba",
          3438 => x"38758180",
          3439 => x"0a298180",
          3440 => x"0a057098",
          3441 => x"2c7081ff",
          3442 => x"06595741",
          3443 => x"76952680",
          3444 => x"c0387510",
          3445 => x"1670822b",
          3446 => x"5155800b",
          3447 => x"83ded416",
          3448 => x"33425777",
          3449 => x"6125ce38",
          3450 => x"83ded015",
          3451 => x"08187033",
          3452 => x"42557861",
          3453 => x"2effbc38",
          3454 => x"76802eff",
          3455 => x"bc38fef2",
          3456 => x"39815776",
          3457 => x"802efeab",
          3458 => x"38fee739",
          3459 => x"8156fdb2",
          3460 => x"39805776",
          3461 => x"fee93876",
          3462 => x"84d18434",
          3463 => x"7684d180",
          3464 => x"34797e34",
          3465 => x"767f0c62",
          3466 => x"55749526",
          3467 => x"fdb03874",
          3468 => x"101083c3",
          3469 => x"94055776",
          3470 => x"080483de",
          3471 => x"d815087f",
          3472 => x"0c800b84",
          3473 => x"d1843480",
          3474 => x"0b84d180",
          3475 => x"34d93984",
          3476 => x"d18c3356",
          3477 => x"75802efd",
          3478 => x"853884d5",
          3479 => x"ac085288",
          3480 => x"51ffb68a",
          3481 => x"3f84d18c",
          3482 => x"33ff0557",
          3483 => x"7684d18c",
          3484 => x"34fceb39",
          3485 => x"84d18c33",
          3486 => x"7081ff06",
          3487 => x"84d18833",
          3488 => x"5b575575",
          3489 => x"7927fcd6",
          3490 => x"3884d5ac",
          3491 => x"08528115",
          3492 => x"587784d1",
          3493 => x"8c347b16",
          3494 => x"70335255",
          3495 => x"ffb5cf3f",
          3496 => x"fcbc397c",
          3497 => x"932e8bda",
          3498 => x"387c1010",
          3499 => x"83f2e405",
          3500 => x"70085759",
          3501 => x"758f8338",
          3502 => x"7584d188",
          3503 => x"34757c34",
          3504 => x"84d18833",
          3505 => x"84d18c33",
          3506 => x"56567480",
          3507 => x"2eb63884",
          3508 => x"d5ac0852",
          3509 => x"8851ffb5",
          3510 => x"953f84d5",
          3511 => x"ac0852a0",
          3512 => x"51ffb58a",
          3513 => x"3f84d5ac",
          3514 => x"08528851",
          3515 => x"ffb4ff3f",
          3516 => x"84d18c33",
          3517 => x"ff055b7a",
          3518 => x"84d18c34",
          3519 => x"7a81ff06",
          3520 => x"5574cc38",
          3521 => x"7b51ffa5",
          3522 => x"ff3f7584",
          3523 => x"d18c34fb",
          3524 => x"cd397c8a",
          3525 => x"3883f3ac",
          3526 => x"0856758d",
          3527 => x"9e387c10",
          3528 => x"1083f2e0",
          3529 => x"05fc1108",
          3530 => x"5755758e",
          3531 => x"f9387408",
          3532 => x"5675802e",
          3533 => x"fba83875",
          3534 => x"51ffb7ec",
          3535 => x"3f84b9c8",
          3536 => x"0884d188",
          3537 => x"3484b9c8",
          3538 => x"0881ff06",
          3539 => x"81055375",
          3540 => x"527b51ff",
          3541 => x"b8943f84",
          3542 => x"d1883384",
          3543 => x"d18c3356",
          3544 => x"5674802e",
          3545 => x"ff9e3884",
          3546 => x"d5ac0852",
          3547 => x"8851ffb3",
          3548 => x"fd3f84d5",
          3549 => x"ac0852a0",
          3550 => x"51ffb3f2",
          3551 => x"3f84d5ac",
          3552 => x"08528851",
          3553 => x"ffb3e73f",
          3554 => x"84d18c33",
          3555 => x"ff055574",
          3556 => x"84d18c34",
          3557 => x"7481ff06",
          3558 => x"55c73984",
          3559 => x"d18c3370",
          3560 => x"81ff0684",
          3561 => x"d188335b",
          3562 => x"57557579",
          3563 => x"27faaf38",
          3564 => x"84d5ac08",
          3565 => x"52811557",
          3566 => x"7684d18c",
          3567 => x"347b1670",
          3568 => x"335255ff",
          3569 => x"b3a83f84",
          3570 => x"d18c3370",
          3571 => x"81ff0684",
          3572 => x"d188335a",
          3573 => x"57557578",
          3574 => x"27fa8338",
          3575 => x"84d5ac08",
          3576 => x"52811557",
          3577 => x"7684d18c",
          3578 => x"347b1670",
          3579 => x"335255ff",
          3580 => x"b2fc3f84",
          3581 => x"d18c3370",
          3582 => x"81ff0684",
          3583 => x"d188335a",
          3584 => x"57557776",
          3585 => x"26ffa938",
          3586 => x"f9d43984",
          3587 => x"d18c3384",
          3588 => x"d1883356",
          3589 => x"5674762e",
          3590 => x"f9c438ff",
          3591 => x"155b7a84",
          3592 => x"d1883475",
          3593 => x"982b7098",
          3594 => x"2c7c81ff",
          3595 => x"0643575a",
          3596 => x"60762480",
          3597 => x"ef3884d5",
          3598 => x"ac0852a0",
          3599 => x"51ffb2ae",
          3600 => x"3f84d18c",
          3601 => x"3370982b",
          3602 => x"70982c84",
          3603 => x"d188335a",
          3604 => x"57574174",
          3605 => x"7724f986",
          3606 => x"3884d5ac",
          3607 => x"08528851",
          3608 => x"ffb28b3f",
          3609 => x"7481800a",
          3610 => x"2981800a",
          3611 => x"0570982c",
          3612 => x"84d18833",
          3613 => x"5d565a74",
          3614 => x"7b24f8e2",
          3615 => x"3884d5ac",
          3616 => x"08528851",
          3617 => x"ffb1e73f",
          3618 => x"7481800a",
          3619 => x"2981800a",
          3620 => x"0570982c",
          3621 => x"84d18833",
          3622 => x"5d565a7a",
          3623 => x"7525ffb9",
          3624 => x"38f8bb39",
          3625 => x"7b165881",
          3626 => x"18337834",
          3627 => x"84d5ac08",
          3628 => x"52773351",
          3629 => x"ffb1b73f",
          3630 => x"7581800a",
          3631 => x"2981800a",
          3632 => x"0570982c",
          3633 => x"84d18833",
          3634 => x"5b575575",
          3635 => x"7925fee6",
          3636 => x"387b1658",
          3637 => x"81183378",
          3638 => x"3484d5ac",
          3639 => x"08527733",
          3640 => x"51ffb18a",
          3641 => x"3f758180",
          3642 => x"0a298180",
          3643 => x"0a057098",
          3644 => x"2c84d188",
          3645 => x"335b5755",
          3646 => x"787624ff",
          3647 => x"a738feb6",
          3648 => x"3984d18c",
          3649 => x"33557480",
          3650 => x"2ef7d338",
          3651 => x"84d5ac08",
          3652 => x"528851ff",
          3653 => x"b0d83f84",
          3654 => x"d18c33ff",
          3655 => x"05577684",
          3656 => x"d18c3476",
          3657 => x"81ff0655",
          3658 => x"dd3984d1",
          3659 => x"88337c05",
          3660 => x"5f807f34",
          3661 => x"84d5ac08",
          3662 => x"528a51ff",
          3663 => x"b0b03f84",
          3664 => x"d188527b",
          3665 => x"51f48b3f",
          3666 => x"84b9c808",
          3667 => x"81ff0658",
          3668 => x"7789cf38",
          3669 => x"84d18833",
          3670 => x"5776802e",
          3671 => x"80d83883",
          3672 => x"f3b83370",
          3673 => x"101083f2",
          3674 => x"e0057008",
          3675 => x"575e5674",
          3676 => x"8ba03875",
          3677 => x"822b87fc",
          3678 => x"0683f2e0",
          3679 => x"05811870",
          3680 => x"53575b80",
          3681 => x"e7fb3f84",
          3682 => x"b9c8087b",
          3683 => x"0c83f3b8",
          3684 => x"33701010",
          3685 => x"83f2e005",
          3686 => x"70085741",
          3687 => x"41748bad",
          3688 => x"3883f3b4",
          3689 => x"08567580",
          3690 => x"2e8c3883",
          3691 => x"f3b03358",
          3692 => x"77802e8b",
          3693 => x"bc38800b",
          3694 => x"84d18c34",
          3695 => x"800b84d1",
          3696 => x"88347b84",
          3697 => x"b9c80cb4",
          3698 => x"3d0d0484",
          3699 => x"d18c3355",
          3700 => x"74802eb6",
          3701 => x"3884d5ac",
          3702 => x"08528851",
          3703 => x"ffaf8f3f",
          3704 => x"84d5ac08",
          3705 => x"52a051ff",
          3706 => x"af843f84",
          3707 => x"d5ac0852",
          3708 => x"8851ffae",
          3709 => x"f93f84d1",
          3710 => x"8c33ff05",
          3711 => x"567584d1",
          3712 => x"8c347581",
          3713 => x"ff065574",
          3714 => x"cc3883d1",
          3715 => x"f051ff9f",
          3716 => x"f73f800b",
          3717 => x"84d18c34",
          3718 => x"800b84d1",
          3719 => x"8834f5be",
          3720 => x"39837c34",
          3721 => x"800b811d",
          3722 => x"3484d18c",
          3723 => x"33557480",
          3724 => x"2eb63884",
          3725 => x"d5ac0852",
          3726 => x"8851ffae",
          3727 => x"b13f84d5",
          3728 => x"ac0852a0",
          3729 => x"51ffaea6",
          3730 => x"3f84d5ac",
          3731 => x"08528851",
          3732 => x"ffae9b3f",
          3733 => x"84d18c33",
          3734 => x"ff055d7c",
          3735 => x"84d18c34",
          3736 => x"7c81ff06",
          3737 => x"5574cc38",
          3738 => x"83d1f051",
          3739 => x"ff9f993f",
          3740 => x"800b84d1",
          3741 => x"8c34800b",
          3742 => x"84d18834",
          3743 => x"7b84b9c8",
          3744 => x"0cb43d0d",
          3745 => x"0484d18c",
          3746 => x"337081ff",
          3747 => x"065c567a",
          3748 => x"802ef4ca",
          3749 => x"3884d188",
          3750 => x"33ff0559",
          3751 => x"7884d188",
          3752 => x"34ff1658",
          3753 => x"7784d18c",
          3754 => x"3484d5ac",
          3755 => x"08528851",
          3756 => x"ffadbb3f",
          3757 => x"84d18c33",
          3758 => x"70982b70",
          3759 => x"982c84d1",
          3760 => x"88335a52",
          3761 => x"5b567676",
          3762 => x"2480ef38",
          3763 => x"84d5ac08",
          3764 => x"52a051ff",
          3765 => x"ad983f84",
          3766 => x"d18c3370",
          3767 => x"982b7098",
          3768 => x"2c84d188",
          3769 => x"335d5759",
          3770 => x"56747a24",
          3771 => x"f3f03884",
          3772 => x"d5ac0852",
          3773 => x"8851ffac",
          3774 => x"f53f7481",
          3775 => x"800a2981",
          3776 => x"800a0570",
          3777 => x"982c84d1",
          3778 => x"88335b51",
          3779 => x"55747924",
          3780 => x"f3cc3884",
          3781 => x"d5ac0852",
          3782 => x"8851ffac",
          3783 => x"d13f7481",
          3784 => x"800a2981",
          3785 => x"800a0570",
          3786 => x"982c84d1",
          3787 => x"88335b51",
          3788 => x"55787525",
          3789 => x"ffb938f3",
          3790 => x"a5397b16",
          3791 => x"57811733",
          3792 => x"773484d5",
          3793 => x"ac085276",
          3794 => x"3351ffac",
          3795 => x"a13f7581",
          3796 => x"800a2981",
          3797 => x"800a0570",
          3798 => x"982c84d1",
          3799 => x"88334357",
          3800 => x"5b756125",
          3801 => x"fee6387b",
          3802 => x"16578117",
          3803 => x"33773484",
          3804 => x"d5ac0852",
          3805 => x"763351ff",
          3806 => x"abf43f75",
          3807 => x"81800a29",
          3808 => x"81800a05",
          3809 => x"70982c84",
          3810 => x"d1883343",
          3811 => x"575b6076",
          3812 => x"24ffa738",
          3813 => x"feb63984",
          3814 => x"d18c3370",
          3815 => x"81ff0658",
          3816 => x"5876602e",
          3817 => x"f2b83884",
          3818 => x"d1883355",
          3819 => x"767527ae",
          3820 => x"3874982b",
          3821 => x"70982c57",
          3822 => x"41767624",
          3823 => x"a1387b16",
          3824 => x"5b7a3381",
          3825 => x"1c347581",
          3826 => x"800a2981",
          3827 => x"ff0a0570",
          3828 => x"982c84d1",
          3829 => x"8c335257",
          3830 => x"58757825",
          3831 => x"e1388118",
          3832 => x"557484d1",
          3833 => x"8c347781",
          3834 => x"ff067c05",
          3835 => x"5ab33d33",
          3836 => x"7a3484d1",
          3837 => x"88335776",
          3838 => x"60258b38",
          3839 => x"81175675",
          3840 => x"84d18834",
          3841 => x"755784d1",
          3842 => x"8c337081",
          3843 => x"800a2981",
          3844 => x"ff0a0570",
          3845 => x"982c7981",
          3846 => x"ff064458",
          3847 => x"5c586076",
          3848 => x"2481ef38",
          3849 => x"77982b70",
          3850 => x"982c7881",
          3851 => x"ff065c57",
          3852 => x"59757a25",
          3853 => x"f1a83884",
          3854 => x"d5ac0852",
          3855 => x"8851ffaa",
          3856 => x"ad3f7581",
          3857 => x"800a2981",
          3858 => x"800a0570",
          3859 => x"982c84d1",
          3860 => x"88335757",
          3861 => x"41757525",
          3862 => x"f1843884",
          3863 => x"d5ac0852",
          3864 => x"8851ffaa",
          3865 => x"893f7581",
          3866 => x"800a2981",
          3867 => x"800a0570",
          3868 => x"982c84d1",
          3869 => x"88335757",
          3870 => x"41747624",
          3871 => x"ffb938f0",
          3872 => x"dd3983f2",
          3873 => x"e0085675",
          3874 => x"802ef49d",
          3875 => x"387551ff",
          3876 => x"ad963f84",
          3877 => x"b9c80884",
          3878 => x"d1883484",
          3879 => x"b9c80881",
          3880 => x"ff068105",
          3881 => x"5375527b",
          3882 => x"51ffadbe",
          3883 => x"3f84d188",
          3884 => x"3384d18c",
          3885 => x"33565674",
          3886 => x"802ef4c8",
          3887 => x"3884d5ac",
          3888 => x"08528851",
          3889 => x"ffa9a73f",
          3890 => x"84d5ac08",
          3891 => x"52a051ff",
          3892 => x"a99c3f84",
          3893 => x"d5ac0852",
          3894 => x"8851ffa9",
          3895 => x"913f84d1",
          3896 => x"8c33ff05",
          3897 => x"5b7a84d1",
          3898 => x"8c347a81",
          3899 => x"ff0655c7",
          3900 => x"39a85180",
          3901 => x"e18b3f84",
          3902 => x"b9c80883",
          3903 => x"f3b40c84",
          3904 => x"b9c80885",
          3905 => x"a5387683",
          3906 => x"f3b03477",
          3907 => x"efca3880",
          3908 => x"c33984d5",
          3909 => x"ac08527b",
          3910 => x"16703352",
          3911 => x"58ffa8ce",
          3912 => x"3f758180",
          3913 => x"0a298180",
          3914 => x"0a057098",
          3915 => x"2c84d188",
          3916 => x"33525757",
          3917 => x"767624da",
          3918 => x"3884d18c",
          3919 => x"3370982b",
          3920 => x"70982c79",
          3921 => x"81ff065d",
          3922 => x"585a5875",
          3923 => x"7a25ef8e",
          3924 => x"38fde439",
          3925 => x"83f3b408",
          3926 => x"802eeefc",
          3927 => x"3883f2e0",
          3928 => x"57935676",
          3929 => x"085574bb",
          3930 => x"38ff1684",
          3931 => x"18585675",
          3932 => x"8025f038",
          3933 => x"800b83f3",
          3934 => x"b83483f3",
          3935 => x"b4085574",
          3936 => x"802eeed4",
          3937 => x"38745181",
          3938 => x"e7f63f83",
          3939 => x"f3b40851",
          3940 => x"80d9fe3f",
          3941 => x"800b83f3",
          3942 => x"b40c933d",
          3943 => x"b43d5f5f",
          3944 => x"eebc3974",
          3945 => x"5180d9e9",
          3946 => x"3f80770c",
          3947 => x"ff168418",
          3948 => x"58567580",
          3949 => x"25ffac38",
          3950 => x"ffba3975",
          3951 => x"51ffaae8",
          3952 => x"3f84b9c8",
          3953 => x"0884d188",
          3954 => x"3484b9c8",
          3955 => x"0881ff06",
          3956 => x"81055375",
          3957 => x"527b51ff",
          3958 => x"ab903f93",
          3959 => x"0b84d188",
          3960 => x"3384d18c",
          3961 => x"3357575d",
          3962 => x"74802ef2",
          3963 => x"973884d5",
          3964 => x"ac085288",
          3965 => x"51ffa6f6",
          3966 => x"3f84d5ac",
          3967 => x"0852a051",
          3968 => x"ffa6eb3f",
          3969 => x"84d5ac08",
          3970 => x"528851ff",
          3971 => x"a6e03f84",
          3972 => x"d18c33ff",
          3973 => x"055a7984",
          3974 => x"d18c3479",
          3975 => x"81ff0655",
          3976 => x"c739807c",
          3977 => x"34800b84",
          3978 => x"d18c3480",
          3979 => x"0b84d188",
          3980 => x"347b84b9",
          3981 => x"c80cb43d",
          3982 => x"0d047551",
          3983 => x"ffa9e93f",
          3984 => x"84b9c808",
          3985 => x"84d18834",
          3986 => x"84b9c808",
          3987 => x"81ff0681",
          3988 => x"05537552",
          3989 => x"7b51ffaa",
          3990 => x"913f811d",
          3991 => x"7081ff06",
          3992 => x"84d18833",
          3993 => x"84d18c33",
          3994 => x"58525e56",
          3995 => x"74802ef1",
          3996 => x"933884d5",
          3997 => x"ac085288",
          3998 => x"51ffa5f2",
          3999 => x"3f84d5ac",
          4000 => x"0852a051",
          4001 => x"ffa5e73f",
          4002 => x"84d5ac08",
          4003 => x"528851ff",
          4004 => x"a5dc3f84",
          4005 => x"d18c33ff",
          4006 => x"05577684",
          4007 => x"d18c3476",
          4008 => x"81ff0655",
          4009 => x"c7397551",
          4010 => x"ffa8fd3f",
          4011 => x"84b9c808",
          4012 => x"84d18834",
          4013 => x"84b9c808",
          4014 => x"81ff0681",
          4015 => x"05537552",
          4016 => x"7b51ffa9",
          4017 => x"a53fff1d",
          4018 => x"7081ff06",
          4019 => x"84d18833",
          4020 => x"84d18c33",
          4021 => x"58585e58",
          4022 => x"74802ef0",
          4023 => x"a73884d5",
          4024 => x"ac085288",
          4025 => x"51ffa586",
          4026 => x"3f84d5ac",
          4027 => x"0852a051",
          4028 => x"ffa4fb3f",
          4029 => x"84d5ac08",
          4030 => x"528851ff",
          4031 => x"a4f03f84",
          4032 => x"d18c33ff",
          4033 => x"05416084",
          4034 => x"d18c3460",
          4035 => x"81ff0655",
          4036 => x"c7397451",
          4037 => x"80d6fa3f",
          4038 => x"83f3b833",
          4039 => x"70822b87",
          4040 => x"fc0683f2",
          4041 => x"e0058119",
          4042 => x"7054525c",
          4043 => x"5680dcd1",
          4044 => x"3f84b9c8",
          4045 => x"087b0c83",
          4046 => x"f3b83370",
          4047 => x"101083f2",
          4048 => x"e0057008",
          4049 => x"57414174",
          4050 => x"802ef4d5",
          4051 => x"3875537b",
          4052 => x"527451ff",
          4053 => x"a8943f83",
          4054 => x"f3b83381",
          4055 => x"057081ff",
          4056 => x"065a5693",
          4057 => x"792782f2",
          4058 => x"387783f3",
          4059 => x"b834f4b1",
          4060 => x"39b43dfe",
          4061 => x"f8055476",
          4062 => x"537b5275",
          4063 => x"5181d8c0",
          4064 => x"3f83f3b4",
          4065 => x"08528a51",
          4066 => x"82ba883f",
          4067 => x"83f3b408",
          4068 => x"5181dff3",
          4069 => x"3f800b84",
          4070 => x"d18c3480",
          4071 => x"0b84d188",
          4072 => x"347b84b9",
          4073 => x"c80cb43d",
          4074 => x"0d049353",
          4075 => x"775284b9",
          4076 => x"c8085181",
          4077 => x"c9f83f84",
          4078 => x"b9c80882",
          4079 => x"a53884b9",
          4080 => x"c808963d",
          4081 => x"5c5d83f3",
          4082 => x"b4085380",
          4083 => x"f8527a51",
          4084 => x"82b7f23f",
          4085 => x"84b9c808",
          4086 => x"5a84b9c8",
          4087 => x"087b2e09",
          4088 => x"8106e9ee",
          4089 => x"3884b9c8",
          4090 => x"0851ffa6",
          4091 => x"bb3f84b9",
          4092 => x"c8085680",
          4093 => x"0b84b9c8",
          4094 => x"082580e3",
          4095 => x"3884b9c8",
          4096 => x"08ff0570",
          4097 => x"1b585680",
          4098 => x"77347581",
          4099 => x"ff0683f3",
          4100 => x"b8337010",
          4101 => x"1083f2e0",
          4102 => x"05700858",
          4103 => x"40585974",
          4104 => x"80f23876",
          4105 => x"822b87fc",
          4106 => x"0683f2e0",
          4107 => x"05811a70",
          4108 => x"53585580",
          4109 => x"dacb3f84",
          4110 => x"b9c80875",
          4111 => x"0c83f3b8",
          4112 => x"33701010",
          4113 => x"83f2e005",
          4114 => x"70085740",
          4115 => x"4174a038",
          4116 => x"811d7081",
          4117 => x"ff065e57",
          4118 => x"937d2783",
          4119 => x"38805d75",
          4120 => x"ff2e0981",
          4121 => x"06fedf38",
          4122 => x"77e8ed38",
          4123 => x"f9e63976",
          4124 => x"53795274",
          4125 => x"51ffa5f2",
          4126 => x"3f83f3b8",
          4127 => x"33810570",
          4128 => x"81ff065b",
          4129 => x"57937a27",
          4130 => x"80c83880",
          4131 => x"0b83f3b8",
          4132 => x"34ffbd39",
          4133 => x"745180d3",
          4134 => x"f83f83f3",
          4135 => x"b8337082",
          4136 => x"2b87fc06",
          4137 => x"83f2e005",
          4138 => x"811b7054",
          4139 => x"52565780",
          4140 => x"d9cf3f84",
          4141 => x"b9c80875",
          4142 => x"0c83f3b8",
          4143 => x"33701010",
          4144 => x"83f2e005",
          4145 => x"70085740",
          4146 => x"4174802e",
          4147 => x"ff8238ff",
          4148 => x"9e397683",
          4149 => x"f3b834fe",
          4150 => x"f7397583",
          4151 => x"f3b834f1",
          4152 => x"c03983e1",
          4153 => x"b051ff9f",
          4154 => x"8a3f77e7",
          4155 => x"eb38f8e4",
          4156 => x"39f23d0d",
          4157 => x"0280c305",
          4158 => x"33028405",
          4159 => x"80c70533",
          4160 => x"5b537283",
          4161 => x"26818d38",
          4162 => x"72812e81",
          4163 => x"8b388173",
          4164 => x"25839e38",
          4165 => x"72822e82",
          4166 => x"a83886a7",
          4167 => x"a0805986",
          4168 => x"a7b08070",
          4169 => x"5e578056",
          4170 => x"9fa05879",
          4171 => x"762e9038",
          4172 => x"7583f8f8",
          4173 => x"347583f8",
          4174 => x"f9347583",
          4175 => x"f8f62383",
          4176 => x"f8f43370",
          4177 => x"982b7190",
          4178 => x"2b077188",
          4179 => x"2b077107",
          4180 => x"7a7f5656",
          4181 => x"565b7877",
          4182 => x"27943880",
          4183 => x"74708405",
          4184 => x"560c7473",
          4185 => x"70840555",
          4186 => x"0c767426",
          4187 => x"ee387578",
          4188 => x"27a23883",
          4189 => x"f8f43384",
          4190 => x"989a1779",
          4191 => x"78315555",
          4192 => x"55a00be0",
          4193 => x"e0153474",
          4194 => x"74708105",
          4195 => x"5634ff13",
          4196 => x"5372ee38",
          4197 => x"903d0d04",
          4198 => x"86a7a080",
          4199 => x"0b83f8f8",
          4200 => x"33701010",
          4201 => x"1183f8f9",
          4202 => x"33719029",
          4203 => x"1174055b",
          4204 => x"41584059",
          4205 => x"86a7b080",
          4206 => x"0b84b7bc",
          4207 => x"337081ff",
          4208 => x"0684b7bb",
          4209 => x"337081ff",
          4210 => x"0683f8f6",
          4211 => x"227083ff",
          4212 => x"ff067075",
          4213 => x"295d595d",
          4214 => x"585e575b",
          4215 => x"5d737326",
          4216 => x"87387274",
          4217 => x"31752956",
          4218 => x"7981ff06",
          4219 => x"7e81ff06",
          4220 => x"7c81ff06",
          4221 => x"7a83ffff",
          4222 => x"066281ff",
          4223 => x"06707529",
          4224 => x"145d4257",
          4225 => x"575b5c74",
          4226 => x"74268f38",
          4227 => x"83f8f833",
          4228 => x"74763105",
          4229 => x"707d291b",
          4230 => x"595f7683",
          4231 => x"065c7b80",
          4232 => x"2efe9c38",
          4233 => x"787d5553",
          4234 => x"727726fe",
          4235 => x"c1388073",
          4236 => x"70810555",
          4237 => x"3483f8f4",
          4238 => x"33747081",
          4239 => x"055634e8",
          4240 => x"3986a7a0",
          4241 => x"805986a7",
          4242 => x"b0807084",
          4243 => x"b7bc3370",
          4244 => x"81ff0684",
          4245 => x"b7bb3370",
          4246 => x"81ff0683",
          4247 => x"f8f62270",
          4248 => x"74295d5b",
          4249 => x"5d575e56",
          4250 => x"5e577478",
          4251 => x"2781df38",
          4252 => x"7381ff06",
          4253 => x"7381ff06",
          4254 => x"71712918",
          4255 => x"5a545479",
          4256 => x"802efdbb",
          4257 => x"38800b83",
          4258 => x"f8f83480",
          4259 => x"0b83f8f9",
          4260 => x"3483f8f4",
          4261 => x"3370982b",
          4262 => x"71902b07",
          4263 => x"71882b07",
          4264 => x"71077a7f",
          4265 => x"5656565b",
          4266 => x"767926fd",
          4267 => x"ae38fdbe",
          4268 => x"3972fce6",
          4269 => x"3883f8f8",
          4270 => x"337081ff",
          4271 => x"06701010",
          4272 => x"1183f8f9",
          4273 => x"33719029",
          4274 => x"1186a7a0",
          4275 => x"80115e57",
          4276 => x"5b56565f",
          4277 => x"86a7b080",
          4278 => x"701484b7",
          4279 => x"bc337081",
          4280 => x"ff0684b7",
          4281 => x"bb337081",
          4282 => x"ff0683f8",
          4283 => x"f6227083",
          4284 => x"ffff067c",
          4285 => x"75296005",
          4286 => x"5e5a415f",
          4287 => x"585f405e",
          4288 => x"57797326",
          4289 => x"8b38727a",
          4290 => x"3115707d",
          4291 => x"29195753",
          4292 => x"7d81ff06",
          4293 => x"7481ff06",
          4294 => x"7171297d",
          4295 => x"83ffff06",
          4296 => x"6281ff06",
          4297 => x"70752958",
          4298 => x"5f5b5c5d",
          4299 => x"557b7826",
          4300 => x"85387775",
          4301 => x"29537973",
          4302 => x"31167983",
          4303 => x"065b5879",
          4304 => x"fde23876",
          4305 => x"83065c7b",
          4306 => x"fdda38fb",
          4307 => x"f2397478",
          4308 => x"317b2956",
          4309 => x"fe9a39fb",
          4310 => x"3d0d878e",
          4311 => x"808c53ff",
          4312 => x"8a733487",
          4313 => x"73348573",
          4314 => x"34817334",
          4315 => x"878e809c",
          4316 => x"5580f475",
          4317 => x"34ffb075",
          4318 => x"34878e80",
          4319 => x"98568076",
          4320 => x"34807634",
          4321 => x"878e8094",
          4322 => x"548a7434",
          4323 => x"807434ff",
          4324 => x"80753481",
          4325 => x"528351fa",
          4326 => x"d83f86a0",
          4327 => x"87e07008",
          4328 => x"545481f8",
          4329 => x"5686a081",
          4330 => x"f8737706",
          4331 => x"84075455",
          4332 => x"72753473",
          4333 => x"087080ff",
          4334 => x"0680c007",
          4335 => x"51537275",
          4336 => x"3486a087",
          4337 => x"cc087077",
          4338 => x"06810751",
          4339 => x"537286a0",
          4340 => x"81f33473",
          4341 => x"0881f706",
          4342 => x"88075372",
          4343 => x"753480d0",
          4344 => x"0b84b7bc",
          4345 => x"34800b84",
          4346 => x"b9c80c87",
          4347 => x"3d0d0484",
          4348 => x"b7bc3384",
          4349 => x"b9c80c04",
          4350 => x"f73d0d02",
          4351 => x"af053302",
          4352 => x"8405b305",
          4353 => x"3384b7bb",
          4354 => x"335b5956",
          4355 => x"81537579",
          4356 => x"2682da38",
          4357 => x"84b7bc33",
          4358 => x"83f8f933",
          4359 => x"83f8f833",
          4360 => x"72712912",
          4361 => x"86a7a080",
          4362 => x"1183f8f6",
          4363 => x"225f5157",
          4364 => x"59717c29",
          4365 => x"057083ff",
          4366 => x"ff0683f7",
          4367 => x"ce335357",
          4368 => x"58537281",
          4369 => x"2e83c438",
          4370 => x"83f8f622",
          4371 => x"76055574",
          4372 => x"83f8f623",
          4373 => x"83f8f833",
          4374 => x"76057081",
          4375 => x"ff067a81",
          4376 => x"ff06555b",
          4377 => x"55727a26",
          4378 => x"828c38ff",
          4379 => x"19537283",
          4380 => x"f8f83483",
          4381 => x"f8f62270",
          4382 => x"83ffff06",
          4383 => x"84b7ba33",
          4384 => x"5c555779",
          4385 => x"74268289",
          4386 => x"3884b7bc",
          4387 => x"33767129",
          4388 => x"54588054",
          4389 => x"729f9f26",
          4390 => x"ac388498",
          4391 => x"9a701454",
          4392 => x"55e0e013",
          4393 => x"33e0e016",
          4394 => x"34727081",
          4395 => x"05543375",
          4396 => x"70810557",
          4397 => x"34811454",
          4398 => x"84b7b973",
          4399 => x"27e33873",
          4400 => x"9f9f26a1",
          4401 => x"3883f8f4",
          4402 => x"3384989a",
          4403 => x"155455a0",
          4404 => x"0be0e014",
          4405 => x"34747370",
          4406 => x"81055534",
          4407 => x"8114549f",
          4408 => x"9f7427eb",
          4409 => x"3884b7ba",
          4410 => x"33ff0556",
          4411 => x"7583f8f6",
          4412 => x"23755778",
          4413 => x"81ff0677",
          4414 => x"83ffff06",
          4415 => x"54547373",
          4416 => x"2681fd38",
          4417 => x"72743181",
          4418 => x"0584b7bc",
          4419 => x"33717129",
          4420 => x"58555775",
          4421 => x"5586a7a0",
          4422 => x"805886a7",
          4423 => x"b0807981",
          4424 => x"ff067581",
          4425 => x"ff067171",
          4426 => x"29195c5c",
          4427 => x"54577579",
          4428 => x"27b93884",
          4429 => x"989a1654",
          4430 => x"e0e01433",
          4431 => x"5384b7c4",
          4432 => x"13337870",
          4433 => x"81055a34",
          4434 => x"73708105",
          4435 => x"55337770",
          4436 => x"81055934",
          4437 => x"811584b7",
          4438 => x"bc3384b7",
          4439 => x"bb337171",
          4440 => x"2919565c",
          4441 => x"5a557275",
          4442 => x"26ce3880",
          4443 => x"537284b9",
          4444 => x"c80c8b3d",
          4445 => x"0d047483",
          4446 => x"f8f83483",
          4447 => x"f8f62270",
          4448 => x"83ffff06",
          4449 => x"84b7ba33",
          4450 => x"5c555773",
          4451 => x"7a27fdf9",
          4452 => x"3877802e",
          4453 => x"fedd3878",
          4454 => x"81ff06ff",
          4455 => x"0583f8f8",
          4456 => x"33565372",
          4457 => x"752e0981",
          4458 => x"06fec838",
          4459 => x"73763181",
          4460 => x"0584b7bc",
          4461 => x"33717129",
          4462 => x"78722911",
          4463 => x"56525954",
          4464 => x"737327fe",
          4465 => x"ae3883f8",
          4466 => x"f4338498",
          4467 => x"9a157476",
          4468 => x"31555656",
          4469 => x"a00be0e0",
          4470 => x"16347575",
          4471 => x"70810557",
          4472 => x"34ff1353",
          4473 => x"72802efe",
          4474 => x"8a38a00b",
          4475 => x"e0e01634",
          4476 => x"75757081",
          4477 => x"055734ff",
          4478 => x"135372d8",
          4479 => x"38fdf439",
          4480 => x"800b84b7",
          4481 => x"bc335556",
          4482 => x"fe893983",
          4483 => x"f8fa1533",
          4484 => x"5984b7c4",
          4485 => x"19337434",
          4486 => x"84b7bb33",
          4487 => x"59fca939",
          4488 => x"fc3d0d76",
          4489 => x"0284059f",
          4490 => x"05335351",
          4491 => x"7086269b",
          4492 => x"38701010",
          4493 => x"83c3ec05",
          4494 => x"51700804",
          4495 => x"84b7bc33",
          4496 => x"51717127",
          4497 => x"86387183",
          4498 => x"f8f93480",
          4499 => x"0b84b9c8",
          4500 => x"0c863d0d",
          4501 => x"04800b83",
          4502 => x"f8f93483",
          4503 => x"f8f83370",
          4504 => x"81ff0654",
          4505 => x"5272802e",
          4506 => x"e238ff12",
          4507 => x"517083f8",
          4508 => x"f834800b",
          4509 => x"84b9c80c",
          4510 => x"863d0d04",
          4511 => x"83f8f833",
          4512 => x"70733170",
          4513 => x"09709f2c",
          4514 => x"72065455",
          4515 => x"53547083",
          4516 => x"f8f834de",
          4517 => x"3983f8f8",
          4518 => x"33720584",
          4519 => x"b7bb33ff",
          4520 => x"11555651",
          4521 => x"70752583",
          4522 => x"38705372",
          4523 => x"83f8f834",
          4524 => x"800b84b9",
          4525 => x"c80c863d",
          4526 => x"0d0483f8",
          4527 => x"f9337073",
          4528 => x"31700970",
          4529 => x"9f2c7206",
          4530 => x"54565355",
          4531 => x"7083f8f9",
          4532 => x"34800b84",
          4533 => x"b9c80c86",
          4534 => x"3d0d0483",
          4535 => x"f8f93372",
          4536 => x"0584b7bc",
          4537 => x"33ff1155",
          4538 => x"55517074",
          4539 => x"25833870",
          4540 => x"537283f8",
          4541 => x"f934800b",
          4542 => x"84b9c80c",
          4543 => x"863d0d04",
          4544 => x"800b83f8",
          4545 => x"f93483f8",
          4546 => x"f83384b7",
          4547 => x"bb33ff05",
          4548 => x"56527175",
          4549 => x"25feb438",
          4550 => x"81125170",
          4551 => x"83f8f834",
          4552 => x"fed039ff",
          4553 => x"3d0d028f",
          4554 => x"05335170",
          4555 => x"b126b338",
          4556 => x"70101083",
          4557 => x"c4880551",
          4558 => x"70080483",
          4559 => x"f8f43370",
          4560 => x"80f00671",
          4561 => x"842b80f0",
          4562 => x"06707284",
          4563 => x"2a075152",
          4564 => x"53517180",
          4565 => x"f02e0981",
          4566 => x"069c3880",
          4567 => x"f20b83f8",
          4568 => x"f434800b",
          4569 => x"84b9c80c",
          4570 => x"833d0d04",
          4571 => x"83f8f433",
          4572 => x"819f0690",
          4573 => x"07517083",
          4574 => x"f8f43480",
          4575 => x"0b84b9c8",
          4576 => x"0c833d0d",
          4577 => x"0483f8f4",
          4578 => x"3380f007",
          4579 => x"517083f8",
          4580 => x"f434e839",
          4581 => x"83f8f433",
          4582 => x"81fe0686",
          4583 => x"07517083",
          4584 => x"f8f434d7",
          4585 => x"3980f10b",
          4586 => x"83f8f434",
          4587 => x"800b84b9",
          4588 => x"c80c833d",
          4589 => x"0d0483f8",
          4590 => x"f43381fc",
          4591 => x"06840751",
          4592 => x"7083f8f4",
          4593 => x"34ffb439",
          4594 => x"83f8f433",
          4595 => x"87075170",
          4596 => x"83f8f434",
          4597 => x"ffa53983",
          4598 => x"f8f43381",
          4599 => x"fd068507",
          4600 => x"517083f8",
          4601 => x"f434ff93",
          4602 => x"3983f8f4",
          4603 => x"3381fb06",
          4604 => x"83075170",
          4605 => x"83f8f434",
          4606 => x"ff813983",
          4607 => x"f8f43381",
          4608 => x"f9068107",
          4609 => x"517083f8",
          4610 => x"f434feef",
          4611 => x"3983f8f4",
          4612 => x"3381f806",
          4613 => x"517083f8",
          4614 => x"f434fedf",
          4615 => x"3983f8f4",
          4616 => x"3381df06",
          4617 => x"80d00751",
          4618 => x"7083f8f4",
          4619 => x"34fecc39",
          4620 => x"83f8f433",
          4621 => x"81bf06b0",
          4622 => x"07517083",
          4623 => x"f8f434fe",
          4624 => x"ba3983f8",
          4625 => x"f43381ef",
          4626 => x"0680e007",
          4627 => x"517083f8",
          4628 => x"f434fea7",
          4629 => x"3983f8f4",
          4630 => x"3381cf06",
          4631 => x"80c00751",
          4632 => x"7083f8f4",
          4633 => x"34fe9439",
          4634 => x"83f8f433",
          4635 => x"81af06a0",
          4636 => x"07517083",
          4637 => x"f8f434fe",
          4638 => x"823983f8",
          4639 => x"f433818f",
          4640 => x"06517083",
          4641 => x"f8f434fd",
          4642 => x"f23983f8",
          4643 => x"f43381fa",
          4644 => x"06820751",
          4645 => x"7083f8f4",
          4646 => x"34fde039",
          4647 => x"f33d0d02",
          4648 => x"bf053302",
          4649 => x"840580c3",
          4650 => x"053383f8",
          4651 => x"f83383f8",
          4652 => x"f73383f8",
          4653 => x"f93384b7",
          4654 => x"be334341",
          4655 => x"5f5d5b59",
          4656 => x"78822e82",
          4657 => x"a1387882",
          4658 => x"24a53878",
          4659 => x"812e8182",
          4660 => x"387d84b7",
          4661 => x"be34800b",
          4662 => x"84b7c034",
          4663 => x"7a83f8f8",
          4664 => x"347b83f8",
          4665 => x"f6237c83",
          4666 => x"f8f9348f",
          4667 => x"3d0d0478",
          4668 => x"832e0981",
          4669 => x"06db3880",
          4670 => x"0b84b7be",
          4671 => x"34810b84",
          4672 => x"b7c03482",
          4673 => x"0b83f8f8",
          4674 => x"34a80b83",
          4675 => x"f8f93482",
          4676 => x"0b83f8f6",
          4677 => x"23795884",
          4678 => x"b7bc3357",
          4679 => x"84b7bb33",
          4680 => x"5684b7ba",
          4681 => x"33557b54",
          4682 => x"7c537a52",
          4683 => x"83e3bc51",
          4684 => x"ff81d53f",
          4685 => x"7d84b7be",
          4686 => x"34800b84",
          4687 => x"b7c0347a",
          4688 => x"83f8f834",
          4689 => x"7b83f8f6",
          4690 => x"237c83f8",
          4691 => x"f9348f3d",
          4692 => x"0d04800b",
          4693 => x"84b7be34",
          4694 => x"810b84b7",
          4695 => x"c034800b",
          4696 => x"83f8f834",
          4697 => x"a80b83f8",
          4698 => x"f934800b",
          4699 => x"83f8f623",
          4700 => x"84b8cb33",
          4701 => x"5884b8ca",
          4702 => x"335784b8",
          4703 => x"c9335679",
          4704 => x"557b547c",
          4705 => x"537a5283",
          4706 => x"e3d851ff",
          4707 => x"80fa3f80",
          4708 => x"0b84b8c9",
          4709 => x"335a5a79",
          4710 => x"7927a538",
          4711 => x"791084b9",
          4712 => x"9c057022",
          4713 => x"535983e3",
          4714 => x"f051ff80",
          4715 => x"db3f811a",
          4716 => x"7081ff06",
          4717 => x"84b8c933",
          4718 => x"525b5978",
          4719 => x"7a26dd38",
          4720 => x"83d2a451",
          4721 => x"ff80c13f",
          4722 => x"7d84b7be",
          4723 => x"34800b84",
          4724 => x"b7c0347a",
          4725 => x"83f8f834",
          4726 => x"7b83f8f6",
          4727 => x"237c83f8",
          4728 => x"f9348f3d",
          4729 => x"0d04800b",
          4730 => x"84b7be34",
          4731 => x"810b84b7",
          4732 => x"c034810b",
          4733 => x"83f8f834",
          4734 => x"a80b83f8",
          4735 => x"f934810b",
          4736 => x"83f8f623",
          4737 => x"83f7ac51",
          4738 => x"ff929d3f",
          4739 => x"84b9c808",
          4740 => x"5283e3f4",
          4741 => x"51fefff0",
          4742 => x"3f805983",
          4743 => x"f7ac51ff",
          4744 => x"92863f78",
          4745 => x"84b9c808",
          4746 => x"27fda638",
          4747 => x"83f7ac19",
          4748 => x"335283e3",
          4749 => x"fc51feff",
          4750 => x"cf3f8119",
          4751 => x"7081ff06",
          4752 => x"5a5ad839",
          4753 => x"f93d0d7a",
          4754 => x"028405a7",
          4755 => x"053384b7",
          4756 => x"bc3383f8",
          4757 => x"f93383f8",
          4758 => x"f8337271",
          4759 => x"291286a7",
          4760 => x"a0801183",
          4761 => x"f8f62253",
          4762 => x"51595c71",
          4763 => x"7c290570",
          4764 => x"83ffff06",
          4765 => x"83f7ce33",
          4766 => x"52595155",
          4767 => x"57577281",
          4768 => x"2e81e938",
          4769 => x"75892e81",
          4770 => x"f9387589",
          4771 => x"2481b938",
          4772 => x"75812e83",
          4773 => x"85387588",
          4774 => x"2e82d538",
          4775 => x"84b7bc33",
          4776 => x"83f8f833",
          4777 => x"83f8f933",
          4778 => x"72722905",
          4779 => x"55565484",
          4780 => x"b7c41633",
          4781 => x"86a7a080",
          4782 => x"143484b7",
          4783 => x"bc3383f8",
          4784 => x"f93383f8",
          4785 => x"f6227271",
          4786 => x"29125a5a",
          4787 => x"56537583",
          4788 => x"f8fa1834",
          4789 => x"83f8f833",
          4790 => x"73712916",
          4791 => x"585483f8",
          4792 => x"f43386a7",
          4793 => x"b0801834",
          4794 => x"84b7bc33",
          4795 => x"7081ff06",
          4796 => x"83f8f622",
          4797 => x"83f8f933",
          4798 => x"72722911",
          4799 => x"575b5755",
          4800 => x"5783f8f4",
          4801 => x"3384989a",
          4802 => x"14348118",
          4803 => x"7081ff06",
          4804 => x"59557378",
          4805 => x"26819938",
          4806 => x"84b7bd33",
          4807 => x"587781ea",
          4808 => x"38ff1753",
          4809 => x"7283f8f9",
          4810 => x"3484b7bf",
          4811 => x"33537280",
          4812 => x"2e8c3884",
          4813 => x"b7c03357",
          4814 => x"76802e80",
          4815 => x"fb38800b",
          4816 => x"84b9c80c",
          4817 => x"893d0d04",
          4818 => x"758d2e97",
          4819 => x"38758d24",
          4820 => x"80f73875",
          4821 => x"8a2e0981",
          4822 => x"06fec138",
          4823 => x"81528151",
          4824 => x"f1963f80",
          4825 => x"0b83f8f9",
          4826 => x"34ffbe39",
          4827 => x"83f8fa15",
          4828 => x"335384b7",
          4829 => x"c4133374",
          4830 => x"3475892e",
          4831 => x"098106fe",
          4832 => x"89388053",
          4833 => x"7652a051",
          4834 => x"fdba3f81",
          4835 => x"137081ff",
          4836 => x"06545472",
          4837 => x"8326ff91",
          4838 => x"387652a0",
          4839 => x"51fda53f",
          4840 => x"81137081",
          4841 => x"ff065454",
          4842 => x"837327d8",
          4843 => x"38fefa39",
          4844 => x"7483f8f9",
          4845 => x"34fef239",
          4846 => x"75528351",
          4847 => x"f9de3f80",
          4848 => x"0b84b9c8",
          4849 => x"0c893d0d",
          4850 => x"047580ff",
          4851 => x"2e098106",
          4852 => x"fdca3883",
          4853 => x"f8f93370",
          4854 => x"81ff0655",
          4855 => x"ff055373",
          4856 => x"83387353",
          4857 => x"7283f8f9",
          4858 => x"347652a0",
          4859 => x"51fcd53f",
          4860 => x"83f8f933",
          4861 => x"7081ff06",
          4862 => x"55ff0553",
          4863 => x"73fea538",
          4864 => x"73537283",
          4865 => x"f8f934fe",
          4866 => x"a039800b",
          4867 => x"83f8f934",
          4868 => x"81528151",
          4869 => x"efe23ffe",
          4870 => x"90398052",
          4871 => x"7551efd8",
          4872 => x"3ffe8639",
          4873 => x"e63d0d02",
          4874 => x"80f30533",
          4875 => x"84b8c408",
          4876 => x"57597581",
          4877 => x"2e81b838",
          4878 => x"75822e83",
          4879 => x"8238788a",
          4880 => x"2e84b538",
          4881 => x"788a2482",
          4882 => x"d1387888",
          4883 => x"2e84b938",
          4884 => x"78892e88",
          4885 => x"8f3884b7",
          4886 => x"bc3383f8",
          4887 => x"f83383f8",
          4888 => x"f9337272",
          4889 => x"2905585e",
          4890 => x"5c84b7c4",
          4891 => x"193386a7",
          4892 => x"a0801734",
          4893 => x"84b7bc33",
          4894 => x"83f8f933",
          4895 => x"83f8f622",
          4896 => x"72712912",
          4897 => x"5a5a4240",
          4898 => x"7883f8fa",
          4899 => x"183483f8",
          4900 => x"f8336071",
          4901 => x"29620540",
          4902 => x"5a83f8f4",
          4903 => x"337f86a7",
          4904 => x"b0800534",
          4905 => x"84b7bc33",
          4906 => x"7081ff06",
          4907 => x"83f8f622",
          4908 => x"83f8f933",
          4909 => x"72722911",
          4910 => x"42405d58",
          4911 => x"5983f8f4",
          4912 => x"3384989a",
          4913 => x"1f34811d",
          4914 => x"7081ff06",
          4915 => x"42587661",
          4916 => x"2681b838",
          4917 => x"84b7bd33",
          4918 => x"5a7986f1",
          4919 => x"38ff1956",
          4920 => x"7583f8f9",
          4921 => x"34800b84",
          4922 => x"b9c80c9c",
          4923 => x"3d0d0478",
          4924 => x"b72e848a",
          4925 => x"38b77925",
          4926 => x"81fd3878",
          4927 => x"b82e9bb3",
          4928 => x"387880db",
          4929 => x"2e89cc38",
          4930 => x"800b84b8",
          4931 => x"c40c84b7",
          4932 => x"bc3383f8",
          4933 => x"f83383f8",
          4934 => x"f9337272",
          4935 => x"29055e40",
          4936 => x"4084b7c4",
          4937 => x"193386a7",
          4938 => x"a0801d34",
          4939 => x"84b7bc33",
          4940 => x"83f8f933",
          4941 => x"83f8f622",
          4942 => x"72712912",
          4943 => x"415f5956",
          4944 => x"7883f8fa",
          4945 => x"1f3483f8",
          4946 => x"f8337671",
          4947 => x"29195b57",
          4948 => x"83f8f433",
          4949 => x"86a7b080",
          4950 => x"1b3484b7",
          4951 => x"bc337081",
          4952 => x"ff0683f8",
          4953 => x"f62283f8",
          4954 => x"f9337272",
          4955 => x"29114442",
          4956 => x"43585983",
          4957 => x"f8f43360",
          4958 => x"84989a05",
          4959 => x"34811f58",
          4960 => x"7781ff06",
          4961 => x"41607727",
          4962 => x"feca3877",
          4963 => x"83f8f934",
          4964 => x"800b84b9",
          4965 => x"c80c9c3d",
          4966 => x"0d04789b",
          4967 => x"2e82b738",
          4968 => x"789b2483",
          4969 => x"8138788d",
          4970 => x"2e098106",
          4971 => x"fda83880",
          4972 => x"0b83f8f9",
          4973 => x"34800b84",
          4974 => x"b9c80c9c",
          4975 => x"3d0d0478",
          4976 => x"9b2e82aa",
          4977 => x"38d01956",
          4978 => x"75892684",
          4979 => x"d03884b8",
          4980 => x"c8338111",
          4981 => x"59577784",
          4982 => x"b8c83478",
          4983 => x"84b8cc18",
          4984 => x"347781ff",
          4985 => x"0659800b",
          4986 => x"84b8cc1a",
          4987 => x"34800b84",
          4988 => x"b9c80c9c",
          4989 => x"3d0d0478",
          4990 => x"9b2efde9",
          4991 => x"38800b84",
          4992 => x"b8c40c84",
          4993 => x"b7bc3383",
          4994 => x"f8f83383",
          4995 => x"f8f93372",
          4996 => x"7229055e",
          4997 => x"404084b7",
          4998 => x"c4193386",
          4999 => x"a7a0801d",
          5000 => x"3484b7bc",
          5001 => x"3383f8f9",
          5002 => x"3383f8f6",
          5003 => x"22727129",
          5004 => x"12415f59",
          5005 => x"567883f8",
          5006 => x"fa1f3483",
          5007 => x"f8f83376",
          5008 => x"7129195b",
          5009 => x"5783f8f4",
          5010 => x"3386a7b0",
          5011 => x"801b3484",
          5012 => x"b7bc3370",
          5013 => x"81ff0683",
          5014 => x"f8f62283",
          5015 => x"f8f93372",
          5016 => x"72291144",
          5017 => x"42435859",
          5018 => x"83f8f433",
          5019 => x"6084989a",
          5020 => x"0534811f",
          5021 => x"58fe8939",
          5022 => x"81528151",
          5023 => x"eafa3f80",
          5024 => x"0b83f8f9",
          5025 => x"34feae39",
          5026 => x"84b7bc33",
          5027 => x"83f8f933",
          5028 => x"7081ff06",
          5029 => x"83f8f833",
          5030 => x"73712912",
          5031 => x"86a7a080",
          5032 => x"0583f8f6",
          5033 => x"2240515d",
          5034 => x"727e2905",
          5035 => x"7083ffff",
          5036 => x"0683f7ce",
          5037 => x"335a5159",
          5038 => x"5a5c7581",
          5039 => x"2e86a438",
          5040 => x"7881ff06",
          5041 => x"ff1a5757",
          5042 => x"76fc9538",
          5043 => x"76567583",
          5044 => x"f8f934fc",
          5045 => x"9039800b",
          5046 => x"84b8c834",
          5047 => x"800b84b8",
          5048 => x"c934800b",
          5049 => x"84b8ca34",
          5050 => x"800b84b8",
          5051 => x"cb34810b",
          5052 => x"84b8c40c",
          5053 => x"800b84b9",
          5054 => x"c80c9c3d",
          5055 => x"0d0483f8",
          5056 => x"f83384b9",
          5057 => x"b03483f8",
          5058 => x"f93384b9",
          5059 => x"b13483f8",
          5060 => x"f73384b9",
          5061 => x"b234800b",
          5062 => x"84b8c40c",
          5063 => x"800b84b9",
          5064 => x"c80c9c3d",
          5065 => x"0d047880",
          5066 => x"ff2e0981",
          5067 => x"06faa738",
          5068 => x"83f8f833",
          5069 => x"84b7bc33",
          5070 => x"7081ff06",
          5071 => x"83f8f933",
          5072 => x"7081ff06",
          5073 => x"72752911",
          5074 => x"86a7a080",
          5075 => x"0583f8f6",
          5076 => x"225c4072",
          5077 => x"7b290570",
          5078 => x"83ffff06",
          5079 => x"83f7ce33",
          5080 => x"445c435c",
          5081 => x"425b5c7d",
          5082 => x"812e85fe",
          5083 => x"387881ff",
          5084 => x"06ff1a58",
          5085 => x"56758338",
          5086 => x"75577683",
          5087 => x"f8f9347b",
          5088 => x"81ff067a",
          5089 => x"81ff0678",
          5090 => x"81ff0672",
          5091 => x"7229055f",
          5092 => x"405b84b7",
          5093 => x"e43386a7",
          5094 => x"a0801e34",
          5095 => x"84b7bc33",
          5096 => x"83f8f933",
          5097 => x"83f8f622",
          5098 => x"72712912",
          5099 => x"5a5e4240",
          5100 => x"a00b83f8",
          5101 => x"fa183483",
          5102 => x"f8f83360",
          5103 => x"71296205",
          5104 => x"5a5683f8",
          5105 => x"f43386a7",
          5106 => x"b0801a34",
          5107 => x"84b7bc33",
          5108 => x"7081ff06",
          5109 => x"83f8f622",
          5110 => x"83f8f933",
          5111 => x"72722911",
          5112 => x"435d5a5e",
          5113 => x"5983f8f4",
          5114 => x"337f8498",
          5115 => x"9a053481",
          5116 => x"1a7081ff",
          5117 => x"065c587c",
          5118 => x"7b2695ea",
          5119 => x"3884b7bd",
          5120 => x"335a7996",
          5121 => x"d038ff19",
          5122 => x"587783f8",
          5123 => x"f93483f8",
          5124 => x"f9337081",
          5125 => x"ff0658ff",
          5126 => x"0556fdac",
          5127 => x"3978bb2e",
          5128 => x"95d83878",
          5129 => x"bd2e83d7",
          5130 => x"3878bf2e",
          5131 => x"95a83884",
          5132 => x"b8c8335f",
          5133 => x"7e83f938",
          5134 => x"ffbf1956",
          5135 => x"75b42684",
          5136 => x"c8387510",
          5137 => x"1083c5d0",
          5138 => x"05587708",
          5139 => x"04800b83",
          5140 => x"f8f93480",
          5141 => x"528151e7",
          5142 => x"9f3f800b",
          5143 => x"84b9c80c",
          5144 => x"9c3d0d04",
          5145 => x"83f8f833",
          5146 => x"84b7bc33",
          5147 => x"7081ff06",
          5148 => x"83f8f933",
          5149 => x"7081ff06",
          5150 => x"72752911",
          5151 => x"86a7a080",
          5152 => x"0583f8f6",
          5153 => x"225c4172",
          5154 => x"7b290570",
          5155 => x"83ffff06",
          5156 => x"83f7ce33",
          5157 => x"4653455c",
          5158 => x"595b5b7f",
          5159 => x"812e82ef",
          5160 => x"38805c7a",
          5161 => x"81ff067a",
          5162 => x"81ff067a",
          5163 => x"81ff0672",
          5164 => x"7229055c",
          5165 => x"584084b7",
          5166 => x"e43386a7",
          5167 => x"a0801b34",
          5168 => x"84b7bc33",
          5169 => x"83f8f933",
          5170 => x"83f8f622",
          5171 => x"72712912",
          5172 => x"5e415e56",
          5173 => x"a00b83f8",
          5174 => x"fa1c3483",
          5175 => x"f8f83376",
          5176 => x"71291e5a",
          5177 => x"5e83f8f4",
          5178 => x"3386a7b0",
          5179 => x"801a3484",
          5180 => x"b7bc3370",
          5181 => x"81ff0683",
          5182 => x"f8f62283",
          5183 => x"f8f93372",
          5184 => x"7229115b",
          5185 => x"445a4059",
          5186 => x"83f8f433",
          5187 => x"84989a18",
          5188 => x"34608105",
          5189 => x"7081ff06",
          5190 => x"5b587e7a",
          5191 => x"2681ac38",
          5192 => x"84b7bd33",
          5193 => x"587792fb",
          5194 => x"38ff1956",
          5195 => x"7583f8f9",
          5196 => x"34811c70",
          5197 => x"81ff065d",
          5198 => x"597b8326",
          5199 => x"f7a73883",
          5200 => x"f8f83384",
          5201 => x"b7bc3383",
          5202 => x"f8f93372",
          5203 => x"81ff0672",
          5204 => x"81ff0672",
          5205 => x"81ff0672",
          5206 => x"72290554",
          5207 => x"5b435b5b",
          5208 => x"5b84b7e4",
          5209 => x"3386a7a0",
          5210 => x"801b3484",
          5211 => x"b7bc3383",
          5212 => x"f8f93383",
          5213 => x"f8f62272",
          5214 => x"7129125e",
          5215 => x"415e56a0",
          5216 => x"0b83f8fa",
          5217 => x"1c3483f8",
          5218 => x"f8337671",
          5219 => x"291e5a5e",
          5220 => x"83f8f433",
          5221 => x"86a7b080",
          5222 => x"1a3484b7",
          5223 => x"bc337081",
          5224 => x"ff0683f8",
          5225 => x"f62283f8",
          5226 => x"f9337272",
          5227 => x"29115b44",
          5228 => x"5a405983",
          5229 => x"f8f43384",
          5230 => x"989a1834",
          5231 => x"60810570",
          5232 => x"81ff065b",
          5233 => x"58797f27",
          5234 => x"fed63877",
          5235 => x"83f8f934",
          5236 => x"fedf3982",
          5237 => x"0b84b8c4",
          5238 => x"0c800b84",
          5239 => x"b9c80c9c",
          5240 => x"3d0d0483",
          5241 => x"f8fa1733",
          5242 => x"5984b7c4",
          5243 => x"19337a34",
          5244 => x"83f8f933",
          5245 => x"7081ff06",
          5246 => x"58ff0556",
          5247 => x"f9ca3981",
          5248 => x"0b84b8ca",
          5249 => x"34800b84",
          5250 => x"b9c80c9c",
          5251 => x"3d0d0483",
          5252 => x"f8fa1733",
          5253 => x"5b84b7c4",
          5254 => x"1b337c34",
          5255 => x"83f8f833",
          5256 => x"84b7bc33",
          5257 => x"83f8f933",
          5258 => x"5b5b5b80",
          5259 => x"5cfcf439",
          5260 => x"84b8cc42",
          5261 => x"9c3ddc11",
          5262 => x"53d80551",
          5263 => x"ff8ac73f",
          5264 => x"84b9c808",
          5265 => x"802efbf0",
          5266 => x"3884b8c9",
          5267 => x"33811157",
          5268 => x"5a7584b8",
          5269 => x"c9347910",
          5270 => x"83fe0641",
          5271 => x"0280ca05",
          5272 => x"226184b9",
          5273 => x"9c0523fb",
          5274 => x"cf3983f8",
          5275 => x"fa17335c",
          5276 => x"84b7c41c",
          5277 => x"337b3483",
          5278 => x"f8f83384",
          5279 => x"b7bc3383",
          5280 => x"f8f9335b",
          5281 => x"5b5cf9e5",
          5282 => x"3984b7bc",
          5283 => x"3383f8f8",
          5284 => x"3383f8f9",
          5285 => x"33727229",
          5286 => x"05415d5b",
          5287 => x"84b7c419",
          5288 => x"337f86a7",
          5289 => x"a0800534",
          5290 => x"84b7bc33",
          5291 => x"83f8f933",
          5292 => x"83f8f622",
          5293 => x"72712912",
          5294 => x"5a435b56",
          5295 => x"7883f8fa",
          5296 => x"183483f8",
          5297 => x"f8337671",
          5298 => x"291b415e",
          5299 => x"83f8f433",
          5300 => x"6086a7b0",
          5301 => x"80053484",
          5302 => x"b7bc3370",
          5303 => x"81ff0683",
          5304 => x"f8f62283",
          5305 => x"f8f93372",
          5306 => x"72291141",
          5307 => x"5f5a425a",
          5308 => x"83f8f433",
          5309 => x"84989a1e",
          5310 => x"34811c70",
          5311 => x"81ff065c",
          5312 => x"58607b26",
          5313 => x"90a23884",
          5314 => x"b7bd3358",
          5315 => x"7790e238",
          5316 => x"ff1a5675",
          5317 => x"83f8f934",
          5318 => x"800b84b8",
          5319 => x"c40c84b7",
          5320 => x"bf33407f",
          5321 => x"802ef3bd",
          5322 => x"3884b7c0",
          5323 => x"335675f3",
          5324 => x"b4387852",
          5325 => x"8151eae4",
          5326 => x"3f800b84",
          5327 => x"b9c80c9c",
          5328 => x"3d0d0484",
          5329 => x"b9b03383",
          5330 => x"f8f83484",
          5331 => x"b9b13383",
          5332 => x"f8f93484",
          5333 => x"b9b23357",
          5334 => x"7683f8f6",
          5335 => x"23ffb939",
          5336 => x"83f8f833",
          5337 => x"84b9b034",
          5338 => x"83f8f933",
          5339 => x"84b9b134",
          5340 => x"83f8f733",
          5341 => x"84b9b234",
          5342 => x"ff9e3984",
          5343 => x"b8c9335b",
          5344 => x"7a802eff",
          5345 => x"933884b9",
          5346 => x"9c225d7c",
          5347 => x"862e0981",
          5348 => x"06ff8538",
          5349 => x"83f8f933",
          5350 => x"81055583",
          5351 => x"f8f83381",
          5352 => x"05549b53",
          5353 => x"83e48452",
          5354 => x"943d7052",
          5355 => x"57feedf8",
          5356 => x"3f7651fe",
          5357 => x"fef23f84",
          5358 => x"b9c80881",
          5359 => x"ff0683f7",
          5360 => x"cc335776",
          5361 => x"054160a0",
          5362 => x"24fecd38",
          5363 => x"765283f7",
          5364 => x"ac51fefd",
          5365 => x"bd3ffec0",
          5366 => x"39800b84",
          5367 => x"b8c9335b",
          5368 => x"587981ff",
          5369 => x"065b777b",
          5370 => x"27fead38",
          5371 => x"771084b9",
          5372 => x"9c058111",
          5373 => x"33574175",
          5374 => x"b1268aa5",
          5375 => x"38751010",
          5376 => x"83c7a405",
          5377 => x"5f7e0804",
          5378 => x"84b8c933",
          5379 => x"5e7d802e",
          5380 => x"8fa43883",
          5381 => x"f8f83384",
          5382 => x"b99d3371",
          5383 => x"71317009",
          5384 => x"709f2c72",
          5385 => x"065a4259",
          5386 => x"5e5c7583",
          5387 => x"f8f834fd",
          5388 => x"e73984b8",
          5389 => x"c9335675",
          5390 => x"802e8ee7",
          5391 => x"3884b99d",
          5392 => x"33ff0570",
          5393 => x"81ff0684",
          5394 => x"b7bc335d",
          5395 => x"575f757b",
          5396 => x"27fdc538",
          5397 => x"7583f8f9",
          5398 => x"34fdbd39",
          5399 => x"800b83f8",
          5400 => x"f93483f8",
          5401 => x"f8337081",
          5402 => x"ff065d57",
          5403 => x"7b802efd",
          5404 => x"a738ff17",
          5405 => x"567583f8",
          5406 => x"f834fd9c",
          5407 => x"39800b83",
          5408 => x"f8f93483",
          5409 => x"f8f83384",
          5410 => x"b7bb33ff",
          5411 => x"05575776",
          5412 => x"7625fd84",
          5413 => x"38811756",
          5414 => x"7583f8f8",
          5415 => x"34fcf939",
          5416 => x"84b8c933",
          5417 => x"407f802e",
          5418 => x"8de03883",
          5419 => x"f8f93384",
          5420 => x"b99d3371",
          5421 => x"71317009",
          5422 => x"709f2c72",
          5423 => x"065a4159",
          5424 => x"425a7583",
          5425 => x"f8f934fc",
          5426 => x"cf3984b8",
          5427 => x"c9335b7a",
          5428 => x"802efcc4",
          5429 => x"3884b99c",
          5430 => x"22416099",
          5431 => x"2e098106",
          5432 => x"fcb63884",
          5433 => x"b7bc3383",
          5434 => x"f8f93383",
          5435 => x"f8f83372",
          5436 => x"71291286",
          5437 => x"a7a08011",
          5438 => x"83f8f622",
          5439 => x"43515a58",
          5440 => x"71602905",
          5441 => x"7083ffff",
          5442 => x"0683f7cc",
          5443 => x"0887fffe",
          5444 => x"8006425a",
          5445 => x"5d5d7e84",
          5446 => x"82802e92",
          5447 => x"bf38800b",
          5448 => x"83f7cd34",
          5449 => x"fbf23984",
          5450 => x"b8c9335a",
          5451 => x"79802efb",
          5452 => x"e73884b9",
          5453 => x"9c225877",
          5454 => x"992e0981",
          5455 => x"06fbd938",
          5456 => x"810b83f7",
          5457 => x"cd34fbd0",
          5458 => x"3984b8c9",
          5459 => x"33567580",
          5460 => x"2e90be38",
          5461 => x"84b99d33",
          5462 => x"83f8f933",
          5463 => x"5d7c0584",
          5464 => x"b7bc33ff",
          5465 => x"11595e56",
          5466 => x"757d2583",
          5467 => x"38755776",
          5468 => x"83f8f934",
          5469 => x"fba23984",
          5470 => x"b8c93357",
          5471 => x"76802e8c",
          5472 => x"c83884b9",
          5473 => x"9d3383f8",
          5474 => x"f8334261",
          5475 => x"0584b7bb",
          5476 => x"33ff1159",
          5477 => x"41567560",
          5478 => x"25833875",
          5479 => x"577683f8",
          5480 => x"f834faf4",
          5481 => x"3983e490",
          5482 => x"51fee8dc",
          5483 => x"3f800b84",
          5484 => x"b8c93357",
          5485 => x"57767627",
          5486 => x"8bc73876",
          5487 => x"1084b99c",
          5488 => x"05702253",
          5489 => x"5a83e3f0",
          5490 => x"51fee8bc",
          5491 => x"3f811770",
          5492 => x"81ff0684",
          5493 => x"b8c93358",
          5494 => x"5858da39",
          5495 => x"820b84b8",
          5496 => x"c9335f57",
          5497 => x"7d802e8d",
          5498 => x"3884b99c",
          5499 => x"22567583",
          5500 => x"26833875",
          5501 => x"57815276",
          5502 => x"81ff0651",
          5503 => x"d5f33ffa",
          5504 => x"973984b8",
          5505 => x"c9335781",
          5506 => x"77278eb7",
          5507 => x"3884b99f",
          5508 => x"33ff0570",
          5509 => x"81ff0684",
          5510 => x"b99d33ff",
          5511 => x"057081ff",
          5512 => x"0684b7bb",
          5513 => x"337081ff",
          5514 => x"06ff1140",
          5515 => x"43525b59",
          5516 => x"5c5c777e",
          5517 => x"27833877",
          5518 => x"5a7983f8",
          5519 => x"f6237681",
          5520 => x"ff06ff18",
          5521 => x"585f777f",
          5522 => x"27833877",
          5523 => x"577683f8",
          5524 => x"f83484b7",
          5525 => x"bc33ff11",
          5526 => x"57407a60",
          5527 => x"27f9b438",
          5528 => x"7a567583",
          5529 => x"f8f934f9",
          5530 => x"af3984b8",
          5531 => x"c9335f7e",
          5532 => x"802e8aef",
          5533 => x"3884b99d",
          5534 => x"3384b7bb",
          5535 => x"33405b7a",
          5536 => x"7f26f994",
          5537 => x"3883f8f8",
          5538 => x"3384b7bc",
          5539 => x"337081ff",
          5540 => x"0683f8f9",
          5541 => x"33717429",
          5542 => x"1186a7a0",
          5543 => x"800583f8",
          5544 => x"f6225f40",
          5545 => x"717e2905",
          5546 => x"7083ffff",
          5547 => x"0683f7ce",
          5548 => x"33465259",
          5549 => x"595f5d60",
          5550 => x"812e84f0",
          5551 => x"387983ff",
          5552 => x"ff06707c",
          5553 => x"315d5780",
          5554 => x"7c248efe",
          5555 => x"3884b7bb",
          5556 => x"33567676",
          5557 => x"278ed638",
          5558 => x"ff165675",
          5559 => x"83f8f623",
          5560 => x"7c81ff06",
          5561 => x"707c3141",
          5562 => x"57806024",
          5563 => x"8ee53884",
          5564 => x"b7bb3356",
          5565 => x"7676278d",
          5566 => x"ee38ff16",
          5567 => x"567583f8",
          5568 => x"f8347e81",
          5569 => x"ff0683f8",
          5570 => x"f6225757",
          5571 => x"805a7676",
          5572 => x"26903875",
          5573 => x"77318105",
          5574 => x"7e81ff06",
          5575 => x"7171295c",
          5576 => x"5e5b7958",
          5577 => x"86a7a080",
          5578 => x"5b86a7b0",
          5579 => x"807f81ff",
          5580 => x"067f81ff",
          5581 => x"06717129",
          5582 => x"1d425842",
          5583 => x"5c797f27",
          5584 => x"f7d63884",
          5585 => x"989a1a57",
          5586 => x"e0e01733",
          5587 => x"5f84b7c4",
          5588 => x"1f337b70",
          5589 => x"81055d34",
          5590 => x"76708105",
          5591 => x"58337c70",
          5592 => x"81055e34",
          5593 => x"811884b7",
          5594 => x"bc3384b7",
          5595 => x"bb337171",
          5596 => x"291d4340",
          5597 => x"5e587760",
          5598 => x"27f79d38",
          5599 => x"e0e01733",
          5600 => x"5f84b7c4",
          5601 => x"1f337b70",
          5602 => x"81055d34",
          5603 => x"76708105",
          5604 => x"58337c70",
          5605 => x"81055e34",
          5606 => x"811884b7",
          5607 => x"bc3384b7",
          5608 => x"bb337171",
          5609 => x"291d4340",
          5610 => x"5e587f78",
          5611 => x"26ff9938",
          5612 => x"f6e63984",
          5613 => x"b8c93356",
          5614 => x"75802e87",
          5615 => x"e0388052",
          5616 => x"84b99d33",
          5617 => x"51d8b13f",
          5618 => x"f6ce3980",
          5619 => x"0b84b7bc",
          5620 => x"33ff1184",
          5621 => x"b8c9335d",
          5622 => x"59405879",
          5623 => x"782e9438",
          5624 => x"84b99c22",
          5625 => x"5675782e",
          5626 => x"0981068b",
          5627 => x"be3883f8",
          5628 => x"f9335876",
          5629 => x"81ff0683",
          5630 => x"f8f83379",
          5631 => x"435c5c76",
          5632 => x"ff2e81ed",
          5633 => x"3884b7bb",
          5634 => x"33407a60",
          5635 => x"26f68938",
          5636 => x"7e81ff06",
          5637 => x"56607626",
          5638 => x"f5fe387b",
          5639 => x"7626617d",
          5640 => x"27075776",
          5641 => x"f5f2387a",
          5642 => x"10101b70",
          5643 => x"90296205",
          5644 => x"86a7a080",
          5645 => x"11701f5d",
          5646 => x"5a86a7b0",
          5647 => x"80057983",
          5648 => x"0658515d",
          5649 => x"758bac38",
          5650 => x"79830657",
          5651 => x"768ba438",
          5652 => x"83f8f433",
          5653 => x"70982b71",
          5654 => x"902b0771",
          5655 => x"882b0771",
          5656 => x"07797f59",
          5657 => x"525f5777",
          5658 => x"7a279e38",
          5659 => x"80777084",
          5660 => x"05590c7d",
          5661 => x"76708405",
          5662 => x"580c7977",
          5663 => x"26ee3884",
          5664 => x"b7bc3384",
          5665 => x"b7bb3341",
          5666 => x"5f7e81ff",
          5667 => x"066081ff",
          5668 => x"0683f8f6",
          5669 => x"227d7329",
          5670 => x"64055959",
          5671 => x"595a7777",
          5672 => x"268c3876",
          5673 => x"78311b70",
          5674 => x"7b296205",
          5675 => x"57407576",
          5676 => x"1d575776",
          5677 => x"7626f4e0",
          5678 => x"3883f8f4",
          5679 => x"3384989a",
          5680 => x"18595aa0",
          5681 => x"0be0e019",
          5682 => x"34797870",
          5683 => x"81055a34",
          5684 => x"81175776",
          5685 => x"7626f4c0",
          5686 => x"38a00be0",
          5687 => x"e0193479",
          5688 => x"78708105",
          5689 => x"5a348117",
          5690 => x"57757727",
          5691 => x"d638f4a8",
          5692 => x"39ff1f70",
          5693 => x"81ff065d",
          5694 => x"58fe8a39",
          5695 => x"83f8f433",
          5696 => x"7080f006",
          5697 => x"71842b80",
          5698 => x"f0067184",
          5699 => x"2a07585d",
          5700 => x"577b80f0",
          5701 => x"2e098106",
          5702 => x"be3880f2",
          5703 => x"0b83f8f4",
          5704 => x"34811870",
          5705 => x"81ff0659",
          5706 => x"56f5b639",
          5707 => x"83f8fa17",
          5708 => x"335e84b7",
          5709 => x"c41e337c",
          5710 => x"3483f8f8",
          5711 => x"3384b7bc",
          5712 => x"3383f8f6",
          5713 => x"2284b7bb",
          5714 => x"33425c5f",
          5715 => x"5dfaee39",
          5716 => x"83f8f433",
          5717 => x"87075675",
          5718 => x"83f8f434",
          5719 => x"81187081",
          5720 => x"ff065956",
          5721 => x"f4fb3983",
          5722 => x"f8f43381",
          5723 => x"fd068507",
          5724 => x"567583f8",
          5725 => x"f434e539",
          5726 => x"83f8f433",
          5727 => x"81fb0683",
          5728 => x"07567583",
          5729 => x"f8f434d4",
          5730 => x"3983f8f4",
          5731 => x"3381f906",
          5732 => x"81075675",
          5733 => x"83f8f434",
          5734 => x"c33983f8",
          5735 => x"f433819f",
          5736 => x"06900756",
          5737 => x"7583f8f4",
          5738 => x"34ffb139",
          5739 => x"80f10b83",
          5740 => x"f8f43481",
          5741 => x"187081ff",
          5742 => x"065956f4",
          5743 => x"a43983f8",
          5744 => x"f433818f",
          5745 => x"06567583",
          5746 => x"f8f434ff",
          5747 => x"8f3983f8",
          5748 => x"f433819f",
          5749 => x"06900756",
          5750 => x"7583f8f4",
          5751 => x"34fefd39",
          5752 => x"83f8f433",
          5753 => x"81ef0680",
          5754 => x"e0075675",
          5755 => x"83f8f434",
          5756 => x"feea3983",
          5757 => x"f8f43381",
          5758 => x"cf0680c0",
          5759 => x"07567583",
          5760 => x"f8f434fe",
          5761 => x"d73983f8",
          5762 => x"f43381af",
          5763 => x"06a00756",
          5764 => x"7583f8f4",
          5765 => x"34fec539",
          5766 => x"83f8f433",
          5767 => x"81fe0686",
          5768 => x"07567583",
          5769 => x"f8f434fe",
          5770 => x"b33983f8",
          5771 => x"f43381fc",
          5772 => x"06840756",
          5773 => x"7583f8f4",
          5774 => x"34fea139",
          5775 => x"83f8f433",
          5776 => x"81fa0682",
          5777 => x"07567583",
          5778 => x"f8f434fe",
          5779 => x"8f3983f8",
          5780 => x"f43381f8",
          5781 => x"06567583",
          5782 => x"f8f434fd",
          5783 => x"ff3983f8",
          5784 => x"f43380f0",
          5785 => x"07567583",
          5786 => x"f8f434fd",
          5787 => x"ef3983f8",
          5788 => x"f43380f0",
          5789 => x"07567583",
          5790 => x"f8f434fd",
          5791 => x"df3983f8",
          5792 => x"f43381df",
          5793 => x"0680d007",
          5794 => x"567583f8",
          5795 => x"f434fdcc",
          5796 => x"3983f8f4",
          5797 => x"3381bf06",
          5798 => x"b0075675",
          5799 => x"83f8f434",
          5800 => x"fdba3980",
          5801 => x"0b83f8f9",
          5802 => x"34805281",
          5803 => x"51d2c93f",
          5804 => x"ecff3984",
          5805 => x"b9b03383",
          5806 => x"f8f83484",
          5807 => x"b9b13383",
          5808 => x"f8f93484",
          5809 => x"b9b23359",
          5810 => x"7883f8f6",
          5811 => x"23800b84",
          5812 => x"b8c40ce8",
          5813 => x"c739810b",
          5814 => x"84b8cb34",
          5815 => x"800b84b9",
          5816 => x"c80c9c3d",
          5817 => x"0d047783",
          5818 => x"f8f93483",
          5819 => x"f8f93370",
          5820 => x"81ff0658",
          5821 => x"ff0556e7",
          5822 => x"cf3984b8",
          5823 => x"cc429c3d",
          5824 => x"dc1153d8",
          5825 => x"0551fef8",
          5826 => x"fd3f84b9",
          5827 => x"c808a138",
          5828 => x"84b9c808",
          5829 => x"84b8c40c",
          5830 => x"800b84b8",
          5831 => x"c834800b",
          5832 => x"84b9c80c",
          5833 => x"9c3d0d04",
          5834 => x"7783f8f9",
          5835 => x"34efe939",
          5836 => x"84b8c933",
          5837 => x"81115c5c",
          5838 => x"7a84b8c9",
          5839 => x"347b1083",
          5840 => x"fe065d02",
          5841 => x"80ca0522",
          5842 => x"84b99c1e",
          5843 => x"23800b84",
          5844 => x"b8c834ca",
          5845 => x"39800b83",
          5846 => x"f8f93480",
          5847 => x"528151d1",
          5848 => x"973f83f8",
          5849 => x"f9337081",
          5850 => x"ff0658ff",
          5851 => x"0556e6d8",
          5852 => x"39800b83",
          5853 => x"f8f93480",
          5854 => x"528151d0",
          5855 => x"fb3fef98",
          5856 => x"398a51fe",
          5857 => x"ebd83fef",
          5858 => x"8f3983f8",
          5859 => x"f933ff05",
          5860 => x"7009709f",
          5861 => x"2c720658",
          5862 => x"5f57f2a6",
          5863 => x"39755281",
          5864 => x"51d93984",
          5865 => x"b7bc3340",
          5866 => x"756027ee",
          5867 => x"eb387583",
          5868 => x"f8f934ee",
          5869 => x"e33983f8",
          5870 => x"f833ff05",
          5871 => x"7009709f",
          5872 => x"2c720658",
          5873 => x"4057f0e2",
          5874 => x"3983f8f8",
          5875 => x"33810584",
          5876 => x"b7bb33ff",
          5877 => x"11595956",
          5878 => x"757825f3",
          5879 => x"c0387557",
          5880 => x"f3bb3984",
          5881 => x"b7bb3370",
          5882 => x"81ff0658",
          5883 => x"5c817726",
          5884 => x"eea63883",
          5885 => x"f8f83384",
          5886 => x"b7bc3370",
          5887 => x"81ff0683",
          5888 => x"f8f93371",
          5889 => x"74291186",
          5890 => x"a7a08005",
          5891 => x"83f8f622",
          5892 => x"5f5f717e",
          5893 => x"29057083",
          5894 => x"ffff0683",
          5895 => x"f7ce335d",
          5896 => x"5b44425f",
          5897 => x"5d77812e",
          5898 => x"81f53879",
          5899 => x"83ffff06",
          5900 => x"ff115c57",
          5901 => x"807b2484",
          5902 => x"893884b7",
          5903 => x"bb335676",
          5904 => x"76278398",
          5905 => x"38ff1656",
          5906 => x"7583f8f6",
          5907 => x"237c81ff",
          5908 => x"06ff1157",
          5909 => x"57807624",
          5910 => x"83df3884",
          5911 => x"b7bb3356",
          5912 => x"76762782",
          5913 => x"ec38ff16",
          5914 => x"567583f8",
          5915 => x"f8347b81",
          5916 => x"ff0683f8",
          5917 => x"f6225757",
          5918 => x"805a7676",
          5919 => x"26903875",
          5920 => x"77318105",
          5921 => x"7e81ff06",
          5922 => x"7171295c",
          5923 => x"5e5f7958",
          5924 => x"86a7a080",
          5925 => x"5b86a7b0",
          5926 => x"807c81ff",
          5927 => x"067f81ff",
          5928 => x"06717129",
          5929 => x"1d414242",
          5930 => x"5d797e27",
          5931 => x"ecea3884",
          5932 => x"989a1a57",
          5933 => x"e0e01733",
          5934 => x"5e84b7c4",
          5935 => x"1e337b70",
          5936 => x"81055d34",
          5937 => x"76708105",
          5938 => x"58337d70",
          5939 => x"81055f34",
          5940 => x"811884b7",
          5941 => x"bc3384b7",
          5942 => x"bb337171",
          5943 => x"291d5941",
          5944 => x"5d587776",
          5945 => x"27ecb138",
          5946 => x"e0e01733",
          5947 => x"5e84b7c4",
          5948 => x"1e337b70",
          5949 => x"81055d34",
          5950 => x"76708105",
          5951 => x"58337d70",
          5952 => x"81055f34",
          5953 => x"811884b7",
          5954 => x"bc3384b7",
          5955 => x"bb337171",
          5956 => x"291d5941",
          5957 => x"5d587578",
          5958 => x"26ff9938",
          5959 => x"ebfa3983",
          5960 => x"f8fa1733",
          5961 => x"5c84b7c4",
          5962 => x"1c337b34",
          5963 => x"83f8f833",
          5964 => x"84b7bc33",
          5965 => x"83f8f622",
          5966 => x"84b7bb33",
          5967 => x"5f5c5f5d",
          5968 => x"fde93976",
          5969 => x"ebd23884",
          5970 => x"b7bb3370",
          5971 => x"81ff06ff",
          5972 => x"115c4258",
          5973 => x"76612783",
          5974 => x"38765a79",
          5975 => x"83f8f623",
          5976 => x"7781ff06",
          5977 => x"ff19585a",
          5978 => x"807a2783",
          5979 => x"38805776",
          5980 => x"83f8f834",
          5981 => x"84b7bc33",
          5982 => x"7081ff06",
          5983 => x"ff125259",
          5984 => x"56807827",
          5985 => x"eb8d3880",
          5986 => x"567583f8",
          5987 => x"f934eb88",
          5988 => x"3983f8f9",
          5989 => x"33810584",
          5990 => x"b7bc33ff",
          5991 => x"11594056",
          5992 => x"757f25ef",
          5993 => x"ca387557",
          5994 => x"efc53975",
          5995 => x"812e0981",
          5996 => x"06f4c038",
          5997 => x"83f8f933",
          5998 => x"7081ff06",
          5999 => x"83f8f833",
          6000 => x"7a445d5d",
          6001 => x"5776ff2e",
          6002 => x"098106f4",
          6003 => x"b838f6a1",
          6004 => x"39ff1d56",
          6005 => x"7583f8f8",
          6006 => x"34fd9339",
          6007 => x"ff1a5675",
          6008 => x"83f8f623",
          6009 => x"fce7397c",
          6010 => x"7b315675",
          6011 => x"83f8f834",
          6012 => x"f2903977",
          6013 => x"7d585677",
          6014 => x"7a26f58d",
          6015 => x"38807670",
          6016 => x"81055834",
          6017 => x"83f8f433",
          6018 => x"77708105",
          6019 => x"5934757a",
          6020 => x"26f4ec38",
          6021 => x"80767081",
          6022 => x"05583483",
          6023 => x"f8f43377",
          6024 => x"70810559",
          6025 => x"34797627",
          6026 => x"d438f4d3",
          6027 => x"39797b31",
          6028 => x"567583f8",
          6029 => x"f623f1a8",
          6030 => x"39800b83",
          6031 => x"f8f834fc",
          6032 => x"ad397e83",
          6033 => x"f8f623fc",
          6034 => x"8439800b",
          6035 => x"83f8f623",
          6036 => x"f18e3980",
          6037 => x"0b83f8f8",
          6038 => x"34f1a739",
          6039 => x"83f8fa18",
          6040 => x"335a84b7",
          6041 => x"c41a3377",
          6042 => x"34800b83",
          6043 => x"f7cd34e9",
          6044 => x"a739fd3d",
          6045 => x"0d029705",
          6046 => x"3384b7be",
          6047 => x"33545472",
          6048 => x"802e9038",
          6049 => x"7351db9c",
          6050 => x"3f800b84",
          6051 => x"b9c80c85",
          6052 => x"3d0d0476",
          6053 => x"527351d7",
          6054 => x"ab3f800b",
          6055 => x"84b9c80c",
          6056 => x"853d0d04",
          6057 => x"f33d0d02",
          6058 => x"bf05335c",
          6059 => x"ff0b83f7",
          6060 => x"cc337081",
          6061 => x"ff0683f7",
          6062 => x"ac113358",
          6063 => x"55555974",
          6064 => x"802e80d6",
          6065 => x"38811456",
          6066 => x"7583f7cc",
          6067 => x"34745978",
          6068 => x"84b9c80c",
          6069 => x"8f3d0d04",
          6070 => x"83f7a808",
          6071 => x"54825373",
          6072 => x"802e9138",
          6073 => x"73733270",
          6074 => x"30710770",
          6075 => x"09709f2a",
          6076 => x"565d5e58",
          6077 => x"7283f7a8",
          6078 => x"0cff5980",
          6079 => x"547b812e",
          6080 => x"09810683",
          6081 => x"387b547b",
          6082 => x"83327030",
          6083 => x"70802576",
          6084 => x"075c5c5d",
          6085 => x"79802e85",
          6086 => x"c43884b7",
          6087 => x"bc3383f8",
          6088 => x"f93383f8",
          6089 => x"f8337271",
          6090 => x"291286a7",
          6091 => x"a0800583",
          6092 => x"f8f6225b",
          6093 => x"595d7179",
          6094 => x"29057083",
          6095 => x"ffff0683",
          6096 => x"f7cd3358",
          6097 => x"59555874",
          6098 => x"812e838c",
          6099 => x"3881f054",
          6100 => x"73878e80",
          6101 => x"8034800b",
          6102 => x"87c09888",
          6103 => x"0c87c098",
          6104 => x"88085675",
          6105 => x"802ef638",
          6106 => x"878e8084",
          6107 => x"08577683",
          6108 => x"f4f81534",
          6109 => x"81147081",
          6110 => x"ff065555",
          6111 => x"81f97427",
          6112 => x"cf388054",
          6113 => x"83f6e814",
          6114 => x"337081ff",
          6115 => x"0683f6f2",
          6116 => x"16335854",
          6117 => x"5572762e",
          6118 => x"85c13872",
          6119 => x"81ff2e86",
          6120 => x"b4387483",
          6121 => x"f6fc1534",
          6122 => x"7581ff06",
          6123 => x"5a7981ff",
          6124 => x"2e85cd38",
          6125 => x"7583f786",
          6126 => x"153483f6",
          6127 => x"e8143383",
          6128 => x"f6f21534",
          6129 => x"81147081",
          6130 => x"ff06555e",
          6131 => x"897427ff",
          6132 => x"b33883f6",
          6133 => x"f0337098",
          6134 => x"2b708025",
          6135 => x"58565475",
          6136 => x"83f7a034",
          6137 => x"7381ff06",
          6138 => x"70862a81",
          6139 => x"32708106",
          6140 => x"51545872",
          6141 => x"802e85e7",
          6142 => x"38810b83",
          6143 => x"f7a13473",
          6144 => x"09810653",
          6145 => x"72802e85",
          6146 => x"e438810b",
          6147 => x"83f7a234",
          6148 => x"800b83f7",
          6149 => x"a13383f7",
          6150 => x"a80883f7",
          6151 => x"a2337083",
          6152 => x"f7a43383",
          6153 => x"f7a3335d",
          6154 => x"5d425e5c",
          6155 => x"5e5683f6",
          6156 => x"fc163355",
          6157 => x"7481ff2e",
          6158 => x"8d3883f7",
          6159 => x"90163354",
          6160 => x"73802e82",
          6161 => x"823883f7",
          6162 => x"86163353",
          6163 => x"7281ff2e",
          6164 => x"8b3883f7",
          6165 => x"90163354",
          6166 => x"7381ec38",
          6167 => x"7481ff06",
          6168 => x"547381ff",
          6169 => x"2e8d3883",
          6170 => x"f7901633",
          6171 => x"5372812e",
          6172 => x"81da3874",
          6173 => x"81ff0653",
          6174 => x"7281ff2e",
          6175 => x"848c3883",
          6176 => x"f7901633",
          6177 => x"54817427",
          6178 => x"84803883",
          6179 => x"f79c0887",
          6180 => x"e80587c0",
          6181 => x"989c0854",
          6182 => x"54737327",
          6183 => x"83ec3881",
          6184 => x"0b87c098",
          6185 => x"9c0883f7",
          6186 => x"9c0c5881",
          6187 => x"167081ff",
          6188 => x"06575489",
          6189 => x"7627fef6",
          6190 => x"387683f7",
          6191 => x"a3347783",
          6192 => x"f7a434fe",
          6193 => x"9e195372",
          6194 => x"9c26828b",
          6195 => x"38721010",
          6196 => x"83c8ec05",
          6197 => x"5a790804",
          6198 => x"83f7d008",
          6199 => x"5473802e",
          6200 => x"913883f4",
          6201 => x"1487c098",
          6202 => x"9c085e5e",
          6203 => x"7d7d27fc",
          6204 => x"dc38800b",
          6205 => x"83f7ce33",
          6206 => x"54547281",
          6207 => x"2e833874",
          6208 => x"547383f7",
          6209 => x"ce3487c0",
          6210 => x"989c0883",
          6211 => x"f7d00c73",
          6212 => x"81ff0658",
          6213 => x"77812e94",
          6214 => x"3883f8fa",
          6215 => x"17335484",
          6216 => x"b7c41433",
          6217 => x"763481f0",
          6218 => x"54fca539",
          6219 => x"83f7a808",
          6220 => x"5372802e",
          6221 => x"829c3872",
          6222 => x"812e83f4",
          6223 => x"3880c376",
          6224 => x"3481f054",
          6225 => x"fc8a3980",
          6226 => x"58fee039",
          6227 => x"80745657",
          6228 => x"83597c81",
          6229 => x"2e9b3879",
          6230 => x"772e0981",
          6231 => x"0683b438",
          6232 => x"7d812e80",
          6233 => x"ed387981",
          6234 => x"2e80d738",
          6235 => x"7981ff06",
          6236 => x"59877727",
          6237 => x"75982b54",
          6238 => x"54728025",
          6239 => x"a1387380",
          6240 => x"2e9c3881",
          6241 => x"177081ff",
          6242 => x"06761081",
          6243 => x"fe068772",
          6244 => x"2771982b",
          6245 => x"57535758",
          6246 => x"54807324",
          6247 => x"e1387810",
          6248 => x"10107910",
          6249 => x"05761183",
          6250 => x"2b780583",
          6251 => x"f3d80570",
          6252 => x"335b5654",
          6253 => x"7887c098",
          6254 => x"9c0883f7",
          6255 => x"9c0c57fd",
          6256 => x"ea398059",
          6257 => x"7d812eff",
          6258 => x"a8387981",
          6259 => x"ff0659ff",
          6260 => x"a0398259",
          6261 => x"ff9b3978",
          6262 => x"ff2efa9f",
          6263 => x"38800b84",
          6264 => x"b7be3354",
          6265 => x"5472812e",
          6266 => x"83e8387b",
          6267 => x"82327030",
          6268 => x"70802576",
          6269 => x"07405956",
          6270 => x"7d8a387b",
          6271 => x"832e0981",
          6272 => x"06f9cc38",
          6273 => x"78ff2ef9",
          6274 => x"c6388053",
          6275 => x"72101010",
          6276 => x"83f7d405",
          6277 => x"70335d54",
          6278 => x"787c2e83",
          6279 => x"ba388113",
          6280 => x"7081ff06",
          6281 => x"54579373",
          6282 => x"27e23884",
          6283 => x"b7bf3353",
          6284 => x"72802ef9",
          6285 => x"9a3884b7",
          6286 => x"c0335574",
          6287 => x"f9913878",
          6288 => x"81ff0652",
          6289 => x"8251ccd4",
          6290 => x"3f7884b9",
          6291 => x"c80c8f3d",
          6292 => x"0d04be76",
          6293 => x"3481f054",
          6294 => x"f9f63972",
          6295 => x"81ff2e92",
          6296 => x"3883f790",
          6297 => x"14338105",
          6298 => x"5b7a83f7",
          6299 => x"901534fa",
          6300 => x"c939800b",
          6301 => x"83f79015",
          6302 => x"34ff0b83",
          6303 => x"f6fc1534",
          6304 => x"ff0b83f7",
          6305 => x"861534fa",
          6306 => x"b1397481",
          6307 => x"ff065372",
          6308 => x"81ff2efc",
          6309 => x"963883f7",
          6310 => x"90163355",
          6311 => x"817527fc",
          6312 => x"8a387781",
          6313 => x"ff065473",
          6314 => x"812e0981",
          6315 => x"06fbfc38",
          6316 => x"83f79c08",
          6317 => x"81fa0587",
          6318 => x"c0989c08",
          6319 => x"54557473",
          6320 => x"27fbe838",
          6321 => x"87c0989c",
          6322 => x"0883f79c",
          6323 => x"0c7681ff",
          6324 => x"0659fbd7",
          6325 => x"39ff0b83",
          6326 => x"f6fc1534",
          6327 => x"f9ca3972",
          6328 => x"83f7a134",
          6329 => x"73098106",
          6330 => x"5372fa9e",
          6331 => x"387283f7",
          6332 => x"a234800b",
          6333 => x"83f7a133",
          6334 => x"83f7a808",
          6335 => x"83f7a233",
          6336 => x"7083f7a4",
          6337 => x"3383f7a3",
          6338 => x"335d5d42",
          6339 => x"5e5c5e56",
          6340 => x"fa9c3979",
          6341 => x"822e0981",
          6342 => x"06fccb38",
          6343 => x"7a597a81",
          6344 => x"2efcce38",
          6345 => x"79812e09",
          6346 => x"8106fcc0",
          6347 => x"38fd9339",
          6348 => x"ef763481",
          6349 => x"f054f898",
          6350 => x"39800b84",
          6351 => x"b7bf3357",
          6352 => x"54758338",
          6353 => x"81547384",
          6354 => x"b7bf34ff",
          6355 => x"59f7ac39",
          6356 => x"800b84b7",
          6357 => x"be335854",
          6358 => x"76833881",
          6359 => x"547384b7",
          6360 => x"be34ff59",
          6361 => x"f7953981",
          6362 => x"5383f7a8",
          6363 => x"08842ef7",
          6364 => x"8338840b",
          6365 => x"83f7a80c",
          6366 => x"f6ff3984",
          6367 => x"b7bb3370",
          6368 => x"81ff06ff",
          6369 => x"11575a54",
          6370 => x"80792783",
          6371 => x"38805574",
          6372 => x"83f8f623",
          6373 => x"7381ff06",
          6374 => x"ff155553",
          6375 => x"80732783",
          6376 => x"38805473",
          6377 => x"83f8f834",
          6378 => x"84b7bc33",
          6379 => x"7081ff06",
          6380 => x"56ff0553",
          6381 => x"80752783",
          6382 => x"38805372",
          6383 => x"83f8f934",
          6384 => x"ff59f6b7",
          6385 => x"39815283",
          6386 => x"51ffbaa5",
          6387 => x"3fff59f6",
          6388 => x"aa397254",
          6389 => x"fc953984",
          6390 => x"14085283",
          6391 => x"f7ac51fe",
          6392 => x"dee53f81",
          6393 => x"0b83f7cc",
          6394 => x"3483f7ac",
          6395 => x"3359fcbb",
          6396 => x"39803d0d",
          6397 => x"8151f5ac",
          6398 => x"3f823d0d",
          6399 => x"04fa3d0d",
          6400 => x"800b83f3",
          6401 => x"d4085357",
          6402 => x"02a30533",
          6403 => x"82133483",
          6404 => x"f3d40851",
          6405 => x"80e07134",
          6406 => x"850b83f3",
          6407 => x"d4085556",
          6408 => x"fe0b8115",
          6409 => x"34800b87",
          6410 => x"9080e834",
          6411 => x"87c0989c",
          6412 => x"0883f3d4",
          6413 => x"085580ce",
          6414 => x"90055387",
          6415 => x"c0989c08",
          6416 => x"5287c098",
          6417 => x"9c085170",
          6418 => x"722ef638",
          6419 => x"81143387",
          6420 => x"c0989c08",
          6421 => x"56527473",
          6422 => x"27873871",
          6423 => x"81fe2edb",
          6424 => x"3887c098",
          6425 => x"a40851ff",
          6426 => x"55707327",
          6427 => x"80c83871",
          6428 => x"5571ff2e",
          6429 => x"80c03887",
          6430 => x"c0989c08",
          6431 => x"80ce9005",
          6432 => x"5387c098",
          6433 => x"9c085287",
          6434 => x"c0989c08",
          6435 => x"5574722e",
          6436 => x"f6388114",
          6437 => x"3387c098",
          6438 => x"9c085252",
          6439 => x"70732787",
          6440 => x"387181ff",
          6441 => x"2edb3887",
          6442 => x"c098a408",
          6443 => x"55727526",
          6444 => x"8338ff52",
          6445 => x"7155ff16",
          6446 => x"7081ff06",
          6447 => x"57537580",
          6448 => x"2e983874",
          6449 => x"81ff0652",
          6450 => x"71fed538",
          6451 => x"74ff2e8a",
          6452 => x"387684b9",
          6453 => x"c80c883d",
          6454 => x"0d04810b",
          6455 => x"84b9c80c",
          6456 => x"883d0d04",
          6457 => x"fa3d0d79",
          6458 => x"028405a3",
          6459 => x"05335652",
          6460 => x"800b83f3",
          6461 => x"d4087388",
          6462 => x"2b87fc80",
          6463 => x"80067075",
          6464 => x"982a0751",
          6465 => x"55555771",
          6466 => x"83153472",
          6467 => x"902a5170",
          6468 => x"84153471",
          6469 => x"902a5675",
          6470 => x"85153472",
          6471 => x"86153483",
          6472 => x"f3d40852",
          6473 => x"74821334",
          6474 => x"83f3d408",
          6475 => x"5180e171",
          6476 => x"34850b83",
          6477 => x"f3d40855",
          6478 => x"56fe0b81",
          6479 => x"1534800b",
          6480 => x"879080e8",
          6481 => x"3487c098",
          6482 => x"9c0883f3",
          6483 => x"d4085580",
          6484 => x"ce900553",
          6485 => x"87c0989c",
          6486 => x"085287c0",
          6487 => x"989c0851",
          6488 => x"70722ef6",
          6489 => x"38811433",
          6490 => x"87c0989c",
          6491 => x"08565274",
          6492 => x"73278738",
          6493 => x"7181fe2e",
          6494 => x"db3887c0",
          6495 => x"98a40851",
          6496 => x"ff557073",
          6497 => x"2780c838",
          6498 => x"715571ff",
          6499 => x"2e80c038",
          6500 => x"87c0989c",
          6501 => x"0880ce90",
          6502 => x"055387c0",
          6503 => x"989c0852",
          6504 => x"87c0989c",
          6505 => x"08557472",
          6506 => x"2ef63881",
          6507 => x"143387c0",
          6508 => x"989c0852",
          6509 => x"52707327",
          6510 => x"87387181",
          6511 => x"ff2edb38",
          6512 => x"87c098a4",
          6513 => x"08557275",
          6514 => x"268338ff",
          6515 => x"527155ff",
          6516 => x"167081ff",
          6517 => x"06575375",
          6518 => x"802e80c7",
          6519 => x"387481ff",
          6520 => x"065271fe",
          6521 => x"d4387451",
          6522 => x"7081ff06",
          6523 => x"5675aa38",
          6524 => x"80c6147b",
          6525 => x"84801155",
          6526 => x"52527073",
          6527 => x"27923871",
          6528 => x"70810553",
          6529 => x"33717081",
          6530 => x"05533472",
          6531 => x"7126f038",
          6532 => x"7684b9c8",
          6533 => x"0c883d0d",
          6534 => x"04810b84",
          6535 => x"b9c80c88",
          6536 => x"3d0d04ff",
          6537 => x"51c239fa",
          6538 => x"3d0d7902",
          6539 => x"8405a305",
          6540 => x"33565680",
          6541 => x"0b83f3d4",
          6542 => x"0877882b",
          6543 => x"87fc8080",
          6544 => x"06707998",
          6545 => x"2a075155",
          6546 => x"55577583",
          6547 => x"15347290",
          6548 => x"2a517084",
          6549 => x"15347590",
          6550 => x"2a527185",
          6551 => x"15347286",
          6552 => x"15347a83",
          6553 => x"f3d40880",
          6554 => x"c6118480",
          6555 => x"13565455",
          6556 => x"51707327",
          6557 => x"97387070",
          6558 => x"81055233",
          6559 => x"72708105",
          6560 => x"54347271",
          6561 => x"26f03883",
          6562 => x"f3d40854",
          6563 => x"74821534",
          6564 => x"83f3d408",
          6565 => x"5580e275",
          6566 => x"34850b83",
          6567 => x"f3d40855",
          6568 => x"56fe0b81",
          6569 => x"1534800b",
          6570 => x"879080e8",
          6571 => x"3487c098",
          6572 => x"9c0883f3",
          6573 => x"d4085580",
          6574 => x"ce900553",
          6575 => x"87c0989c",
          6576 => x"085287c0",
          6577 => x"989c0851",
          6578 => x"70722ef6",
          6579 => x"38811433",
          6580 => x"87c0989c",
          6581 => x"08565274",
          6582 => x"73278738",
          6583 => x"7181fe2e",
          6584 => x"db3887c0",
          6585 => x"98a40851",
          6586 => x"ff557073",
          6587 => x"2780c838",
          6588 => x"715571ff",
          6589 => x"2e80c038",
          6590 => x"87c0989c",
          6591 => x"0880ce90",
          6592 => x"055387c0",
          6593 => x"989c0852",
          6594 => x"87c0989c",
          6595 => x"08557472",
          6596 => x"2ef63881",
          6597 => x"143387c0",
          6598 => x"989c0852",
          6599 => x"52707327",
          6600 => x"87387181",
          6601 => x"ff2edb38",
          6602 => x"87c098a4",
          6603 => x"08557275",
          6604 => x"268338ff",
          6605 => x"527155ff",
          6606 => x"167081ff",
          6607 => x"06575375",
          6608 => x"802ea138",
          6609 => x"7481ff06",
          6610 => x"5271fed5",
          6611 => x"38745170",
          6612 => x"81ff0654",
          6613 => x"73802e83",
          6614 => x"38815776",
          6615 => x"84b9c80c",
          6616 => x"883d0d04",
          6617 => x"ff51e839",
          6618 => x"fb3d0d83",
          6619 => x"f3d40851",
          6620 => x"80d07134",
          6621 => x"850b83f3",
          6622 => x"d4085656",
          6623 => x"fe0b8116",
          6624 => x"34800b87",
          6625 => x"9080e834",
          6626 => x"87c0989c",
          6627 => x"0883f3d4",
          6628 => x"085680ce",
          6629 => x"90055487",
          6630 => x"c0989c08",
          6631 => x"5287c098",
          6632 => x"9c085372",
          6633 => x"722ef638",
          6634 => x"81153387",
          6635 => x"c0989c08",
          6636 => x"52527074",
          6637 => x"27873871",
          6638 => x"81fe2edb",
          6639 => x"3887c098",
          6640 => x"a40851ff",
          6641 => x"53707427",
          6642 => x"80c83871",
          6643 => x"5371ff2e",
          6644 => x"80c03887",
          6645 => x"c0989c08",
          6646 => x"80ce9005",
          6647 => x"5387c098",
          6648 => x"9c085287",
          6649 => x"c0989c08",
          6650 => x"5170722e",
          6651 => x"f6388115",
          6652 => x"3387c098",
          6653 => x"9c085552",
          6654 => x"73732787",
          6655 => x"387181ff",
          6656 => x"2edb3887",
          6657 => x"c098a408",
          6658 => x"51727126",
          6659 => x"8338ff52",
          6660 => x"7153ff16",
          6661 => x"7081ff06",
          6662 => x"57527580",
          6663 => x"2e8a3872",
          6664 => x"81ff0654",
          6665 => x"73fed538",
          6666 => x"ff39803d",
          6667 => x"0d83e4cc",
          6668 => x"51fed0bf",
          6669 => x"3f823d0d",
          6670 => x"04f93d0d",
          6671 => x"84b9b808",
          6672 => x"7a713183",
          6673 => x"2a7083ff",
          6674 => x"ff067083",
          6675 => x"2b731170",
          6676 => x"33811233",
          6677 => x"718b2b71",
          6678 => x"832b0777",
          6679 => x"11703381",
          6680 => x"12337198",
          6681 => x"2b71902b",
          6682 => x"075c5441",
          6683 => x"53535d57",
          6684 => x"59525657",
          6685 => x"53807124",
          6686 => x"81af3872",
          6687 => x"16821133",
          6688 => x"83123371",
          6689 => x"8b2b7183",
          6690 => x"2b077605",
          6691 => x"70338112",
          6692 => x"3371982b",
          6693 => x"71902b07",
          6694 => x"57535c52",
          6695 => x"59565280",
          6696 => x"7124839e",
          6697 => x"38841333",
          6698 => x"85143371",
          6699 => x"8b2b7183",
          6700 => x"2b077505",
          6701 => x"76882a52",
          6702 => x"54565774",
          6703 => x"86133473",
          6704 => x"81ff0654",
          6705 => x"73871334",
          6706 => x"84b9b808",
          6707 => x"70178412",
          6708 => x"33851333",
          6709 => x"71882b07",
          6710 => x"70882a5c",
          6711 => x"55595451",
          6712 => x"77841434",
          6713 => x"71851434",
          6714 => x"84b9b808",
          6715 => x"1652800b",
          6716 => x"86133480",
          6717 => x"0b871334",
          6718 => x"84b9b808",
          6719 => x"53748414",
          6720 => x"34738514",
          6721 => x"3484b9b8",
          6722 => x"08167033",
          6723 => x"81123371",
          6724 => x"882b0782",
          6725 => x"80800770",
          6726 => x"882a5858",
          6727 => x"52527472",
          6728 => x"34758113",
          6729 => x"34893d0d",
          6730 => x"04861233",
          6731 => x"87133371",
          6732 => x"8b2b7183",
          6733 => x"2b077511",
          6734 => x"84163385",
          6735 => x"17337188",
          6736 => x"2b077088",
          6737 => x"2a585854",
          6738 => x"51535858",
          6739 => x"71841234",
          6740 => x"72851234",
          6741 => x"84b9b808",
          6742 => x"70168411",
          6743 => x"33851233",
          6744 => x"718b2b71",
          6745 => x"832b0756",
          6746 => x"5a5a5272",
          6747 => x"05861233",
          6748 => x"87133371",
          6749 => x"882b0770",
          6750 => x"882a5255",
          6751 => x"59527786",
          6752 => x"13347287",
          6753 => x"133484b9",
          6754 => x"b8081570",
          6755 => x"33811233",
          6756 => x"71882b07",
          6757 => x"81ffff06",
          6758 => x"70882a5a",
          6759 => x"5a545276",
          6760 => x"72347781",
          6761 => x"133484b9",
          6762 => x"b8087017",
          6763 => x"70338112",
          6764 => x"33718b2b",
          6765 => x"71832b07",
          6766 => x"74057033",
          6767 => x"81123371",
          6768 => x"882b0770",
          6769 => x"832b8fff",
          6770 => x"f8067705",
          6771 => x"7b882a54",
          6772 => x"5253545c",
          6773 => x"5a575452",
          6774 => x"77821434",
          6775 => x"73831434",
          6776 => x"84b9b808",
          6777 => x"70177033",
          6778 => x"81123371",
          6779 => x"8b2b7183",
          6780 => x"2b077405",
          6781 => x"70338112",
          6782 => x"3371882b",
          6783 => x"0781ffff",
          6784 => x"0670882a",
          6785 => x"5f525355",
          6786 => x"5a575452",
          6787 => x"77733470",
          6788 => x"81143484",
          6789 => x"b9b80870",
          6790 => x"17821133",
          6791 => x"83123371",
          6792 => x"8b2b7183",
          6793 => x"2b077405",
          6794 => x"70338112",
          6795 => x"3371982b",
          6796 => x"71902b07",
          6797 => x"58535d52",
          6798 => x"5a575353",
          6799 => x"708025fc",
          6800 => x"e4387133",
          6801 => x"81133371",
          6802 => x"882b0782",
          6803 => x"80800770",
          6804 => x"882a5959",
          6805 => x"54767534",
          6806 => x"77811634",
          6807 => x"84b9b808",
          6808 => x"70177033",
          6809 => x"81123371",
          6810 => x"8b2b7183",
          6811 => x"2b077405",
          6812 => x"82143383",
          6813 => x"15337188",
          6814 => x"2b077088",
          6815 => x"2a575c5c",
          6816 => x"52585652",
          6817 => x"53728215",
          6818 => x"34758315",
          6819 => x"34893d0d",
          6820 => x"04f93d0d",
          6821 => x"7984b9b8",
          6822 => x"08585876",
          6823 => x"802e8f38",
          6824 => x"77802e86",
          6825 => x"387751fb",
          6826 => x"903f893d",
          6827 => x"0d0484ff",
          6828 => x"f40b84b9",
          6829 => x"b80ca080",
          6830 => x"0b84b9b4",
          6831 => x"23828080",
          6832 => x"53765284",
          6833 => x"fff451fe",
          6834 => x"d3b53f84",
          6835 => x"b9b80855",
          6836 => x"76753481",
          6837 => x"0b811634",
          6838 => x"84b9b808",
          6839 => x"54768415",
          6840 => x"34810b85",
          6841 => x"153484b9",
          6842 => x"b8085676",
          6843 => x"86173481",
          6844 => x"0b871734",
          6845 => x"84b9b808",
          6846 => x"84b9b422",
          6847 => x"ff05fe80",
          6848 => x"80077083",
          6849 => x"ffff0670",
          6850 => x"882a5851",
          6851 => x"55567488",
          6852 => x"17347389",
          6853 => x"173484b9",
          6854 => x"b4227010",
          6855 => x"101084b9",
          6856 => x"b80805f8",
          6857 => x"05555576",
          6858 => x"82153481",
          6859 => x"0b831534",
          6860 => x"feee39f7",
          6861 => x"3d0d7b52",
          6862 => x"80538151",
          6863 => x"8472278e",
          6864 => x"38fb1283",
          6865 => x"2a820570",
          6866 => x"83ffff06",
          6867 => x"51517083",
          6868 => x"ffff0684",
          6869 => x"b9b80884",
          6870 => x"11338512",
          6871 => x"3371882b",
          6872 => x"07705259",
          6873 => x"5a585581",
          6874 => x"ffff5475",
          6875 => x"802e80cc",
          6876 => x"38751010",
          6877 => x"10177033",
          6878 => x"81123371",
          6879 => x"882b0770",
          6880 => x"81ffff06",
          6881 => x"79317083",
          6882 => x"ffff0670",
          6883 => x"7a275653",
          6884 => x"5c5c5452",
          6885 => x"7274278a",
          6886 => x"3870802e",
          6887 => x"85387573",
          6888 => x"55588412",
          6889 => x"33851333",
          6890 => x"71882b07",
          6891 => x"575a75c1",
          6892 => x"387381ff",
          6893 => x"ff2e8538",
          6894 => x"77745456",
          6895 => x"8076832b",
          6896 => x"78117033",
          6897 => x"81123371",
          6898 => x"882b0770",
          6899 => x"81ffff06",
          6900 => x"56565d56",
          6901 => x"59597079",
          6902 => x"2e833881",
          6903 => x"59805174",
          6904 => x"7326828d",
          6905 => x"38785178",
          6906 => x"802e8285",
          6907 => x"3872752e",
          6908 => x"82883874",
          6909 => x"1670832b",
          6910 => x"78117482",
          6911 => x"80800770",
          6912 => x"882a5b5c",
          6913 => x"56565a76",
          6914 => x"74347881",
          6915 => x"153484b9",
          6916 => x"b8081576",
          6917 => x"882a5353",
          6918 => x"71821434",
          6919 => x"75831434",
          6920 => x"84b9b808",
          6921 => x"70197033",
          6922 => x"81123371",
          6923 => x"882b0770",
          6924 => x"832b8fff",
          6925 => x"f8067405",
          6926 => x"7e83ffff",
          6927 => x"0670882a",
          6928 => x"5c585357",
          6929 => x"59525275",
          6930 => x"82123472",
          6931 => x"81ff0653",
          6932 => x"72831234",
          6933 => x"84b9b808",
          6934 => x"18547574",
          6935 => x"34728115",
          6936 => x"3484b9b8",
          6937 => x"08701986",
          6938 => x"11338712",
          6939 => x"33718b2b",
          6940 => x"71832b07",
          6941 => x"7405585c",
          6942 => x"5c535775",
          6943 => x"84153472",
          6944 => x"85153484",
          6945 => x"b9b80870",
          6946 => x"16557805",
          6947 => x"86113387",
          6948 => x"12337188",
          6949 => x"2b077088",
          6950 => x"2a545458",
          6951 => x"59708615",
          6952 => x"34718715",
          6953 => x"3484b9b8",
          6954 => x"08701984",
          6955 => x"11338512",
          6956 => x"33718b2b",
          6957 => x"71832b07",
          6958 => x"7405585a",
          6959 => x"5c5a5275",
          6960 => x"86153472",
          6961 => x"87153484",
          6962 => x"b9b80870",
          6963 => x"16557805",
          6964 => x"84113385",
          6965 => x"12337188",
          6966 => x"2b077088",
          6967 => x"2a545c57",
          6968 => x"59708415",
          6969 => x"34798515",
          6970 => x"3484b9b8",
          6971 => x"08188405",
          6972 => x"517084b9",
          6973 => x"c80c8b3d",
          6974 => x"0d048614",
          6975 => x"33871533",
          6976 => x"718b2b71",
          6977 => x"832b0779",
          6978 => x"05841733",
          6979 => x"85183371",
          6980 => x"882b0770",
          6981 => x"882a5a5b",
          6982 => x"59535452",
          6983 => x"74841234",
          6984 => x"76851234",
          6985 => x"84b9b808",
          6986 => x"70198411",
          6987 => x"33851233",
          6988 => x"718b2b71",
          6989 => x"832b0774",
          6990 => x"05861433",
          6991 => x"87153371",
          6992 => x"882b0770",
          6993 => x"882a585d",
          6994 => x"5f52565b",
          6995 => x"57527086",
          6996 => x"1a347687",
          6997 => x"1a3484b9",
          6998 => x"b8081870",
          6999 => x"33811233",
          7000 => x"71882b07",
          7001 => x"81ffff06",
          7002 => x"70882a59",
          7003 => x"57545775",
          7004 => x"77347481",
          7005 => x"183484b9",
          7006 => x"b8081884",
          7007 => x"0551fef1",
          7008 => x"39f93d0d",
          7009 => x"7984b9b8",
          7010 => x"08585876",
          7011 => x"802ea038",
          7012 => x"7754778a",
          7013 => x"387384b9",
          7014 => x"c80c893d",
          7015 => x"0d047751",
          7016 => x"fb913f84",
          7017 => x"b9c80884",
          7018 => x"b9c80c89",
          7019 => x"3d0d0484",
          7020 => x"fff40b84",
          7021 => x"b9b80ca0",
          7022 => x"800b84b9",
          7023 => x"b4238280",
          7024 => x"80537652",
          7025 => x"84fff451",
          7026 => x"fecdb43f",
          7027 => x"84b9b808",
          7028 => x"55767534",
          7029 => x"810b8116",
          7030 => x"3484b9b8",
          7031 => x"08547684",
          7032 => x"1534810b",
          7033 => x"85153484",
          7034 => x"b9b80856",
          7035 => x"76861734",
          7036 => x"810b8717",
          7037 => x"3484b9b8",
          7038 => x"0884b9b4",
          7039 => x"22ff05fe",
          7040 => x"80800770",
          7041 => x"83ffff06",
          7042 => x"70882a58",
          7043 => x"51555674",
          7044 => x"88173473",
          7045 => x"89173484",
          7046 => x"b9b42270",
          7047 => x"10101084",
          7048 => x"b9b80805",
          7049 => x"f8055555",
          7050 => x"76821534",
          7051 => x"810b8315",
          7052 => x"34775477",
          7053 => x"802efedd",
          7054 => x"38fee339",
          7055 => x"ed3d0d65",
          7056 => x"67415f80",
          7057 => x"7084b9b8",
          7058 => x"08594541",
          7059 => x"76612e84",
          7060 => x"aa387e80",
          7061 => x"2e85af38",
          7062 => x"7f802e88",
          7063 => x"d7388154",
          7064 => x"8460278f",
          7065 => x"387ffb05",
          7066 => x"832a8205",
          7067 => x"7083ffff",
          7068 => x"06555873",
          7069 => x"83ffff06",
          7070 => x"7f783183",
          7071 => x"2a7083ff",
          7072 => x"ff067083",
          7073 => x"2b7a1170",
          7074 => x"33811233",
          7075 => x"71882b07",
          7076 => x"70753170",
          7077 => x"83ffff06",
          7078 => x"70101010",
          7079 => x"fc057383",
          7080 => x"2b611170",
          7081 => x"33811233",
          7082 => x"71882b07",
          7083 => x"70902b70",
          7084 => x"902c5342",
          7085 => x"45464453",
          7086 => x"5443445c",
          7087 => x"4859525e",
          7088 => x"5f42807a",
          7089 => x"2485fd38",
          7090 => x"82153383",
          7091 => x"16337188",
          7092 => x"2b077010",
          7093 => x"10101970",
          7094 => x"33811233",
          7095 => x"71982b71",
          7096 => x"902b0753",
          7097 => x"5c535656",
          7098 => x"56807424",
          7099 => x"85c9387a",
          7100 => x"622782f6",
          7101 => x"38631b58",
          7102 => x"77622e87",
          7103 => x"a2386080",
          7104 => x"2e85f938",
          7105 => x"601b5877",
          7106 => x"622587be",
          7107 => x"38631859",
          7108 => x"61792492",
          7109 => x"f738761e",
          7110 => x"70338112",
          7111 => x"33718b2b",
          7112 => x"71832b07",
          7113 => x"7a117033",
          7114 => x"81123371",
          7115 => x"982b7190",
          7116 => x"2b074743",
          7117 => x"59525357",
          7118 => x"5b588060",
          7119 => x"248cba38",
          7120 => x"761e8211",
          7121 => x"33831233",
          7122 => x"718b2b71",
          7123 => x"832b077a",
          7124 => x"11861133",
          7125 => x"87123371",
          7126 => x"8b2b7183",
          7127 => x"2b077e05",
          7128 => x"84143385",
          7129 => x"15337188",
          7130 => x"2b077088",
          7131 => x"2a595748",
          7132 => x"525b4158",
          7133 => x"535c5956",
          7134 => x"77841d34",
          7135 => x"79851d34",
          7136 => x"84b9b808",
          7137 => x"70178411",
          7138 => x"33851233",
          7139 => x"718b2b71",
          7140 => x"832b0774",
          7141 => x"05861433",
          7142 => x"87153371",
          7143 => x"882b0770",
          7144 => x"882a5f42",
          7145 => x"5e524057",
          7146 => x"41577786",
          7147 => x"16347b87",
          7148 => x"163484b9",
          7149 => x"b8081670",
          7150 => x"33811233",
          7151 => x"71882b07",
          7152 => x"81ffff06",
          7153 => x"70882a5a",
          7154 => x"5c5e5976",
          7155 => x"79347981",
          7156 => x"1a3484b9",
          7157 => x"b808701f",
          7158 => x"82113383",
          7159 => x"1233718b",
          7160 => x"2b71832b",
          7161 => x"07740573",
          7162 => x"33811533",
          7163 => x"71882b07",
          7164 => x"70882a41",
          7165 => x"5c455d5f",
          7166 => x"5a555579",
          7167 => x"79347581",
          7168 => x"1a3484b9",
          7169 => x"b808701f",
          7170 => x"70338112",
          7171 => x"33718b2b",
          7172 => x"71832b07",
          7173 => x"74058214",
          7174 => x"33831533",
          7175 => x"71882b07",
          7176 => x"70882a41",
          7177 => x"5c455d5f",
          7178 => x"5a555579",
          7179 => x"821a3475",
          7180 => x"831a3484",
          7181 => x"b9b80870",
          7182 => x"1f821133",
          7183 => x"83123371",
          7184 => x"882b0766",
          7185 => x"57625670",
          7186 => x"832b4252",
          7187 => x"5a5d7e05",
          7188 => x"840551fe",
          7189 => x"c4ec3f84",
          7190 => x"b9b8081e",
          7191 => x"84056165",
          7192 => x"051c7083",
          7193 => x"ffff065d",
          7194 => x"445f7a62",
          7195 => x"2681b638",
          7196 => x"7e547384",
          7197 => x"b9c80c95",
          7198 => x"3d0d0484",
          7199 => x"fff40b84",
          7200 => x"b9b80ca0",
          7201 => x"800b84b9",
          7202 => x"b4238280",
          7203 => x"80536052",
          7204 => x"84fff451",
          7205 => x"fec7e83f",
          7206 => x"84b9b808",
          7207 => x"5e607e34",
          7208 => x"810b811f",
          7209 => x"3484b9b8",
          7210 => x"085d6084",
          7211 => x"1e34810b",
          7212 => x"851e3484",
          7213 => x"b9b8085c",
          7214 => x"60861d34",
          7215 => x"810b871d",
          7216 => x"3484b9b8",
          7217 => x"0884b9b4",
          7218 => x"22ff05fe",
          7219 => x"80800770",
          7220 => x"83ffff06",
          7221 => x"70882a5c",
          7222 => x"5a5b5778",
          7223 => x"88183477",
          7224 => x"89183484",
          7225 => x"b9b42270",
          7226 => x"10101084",
          7227 => x"b9b80805",
          7228 => x"f8055556",
          7229 => x"60821534",
          7230 => x"810b8315",
          7231 => x"3484b9b8",
          7232 => x"08577efa",
          7233 => x"d3387680",
          7234 => x"2e828c38",
          7235 => x"7e547f80",
          7236 => x"2efedf38",
          7237 => x"7f51f49b",
          7238 => x"3f84b9c8",
          7239 => x"0884b9c8",
          7240 => x"0c953d0d",
          7241 => x"04611c84",
          7242 => x"b9b80871",
          7243 => x"832b7111",
          7244 => x"5e447f05",
          7245 => x"70338112",
          7246 => x"3371882b",
          7247 => x"0781ffff",
          7248 => x"0670882a",
          7249 => x"48445b5e",
          7250 => x"40637b34",
          7251 => x"60811c34",
          7252 => x"6184b9b8",
          7253 => x"08057c88",
          7254 => x"2a575875",
          7255 => x"8219347b",
          7256 => x"83193484",
          7257 => x"b9b80870",
          7258 => x"1f703381",
          7259 => x"12337188",
          7260 => x"2b077083",
          7261 => x"2b8ffff8",
          7262 => x"06740564",
          7263 => x"83ffff06",
          7264 => x"70882a4a",
          7265 => x"5c47575e",
          7266 => x"5b5d6363",
          7267 => x"82053476",
          7268 => x"81ff0641",
          7269 => x"60638305",
          7270 => x"3484b9b8",
          7271 => x"081e5b63",
          7272 => x"7b346081",
          7273 => x"1c346184",
          7274 => x"b9b80805",
          7275 => x"840551ed",
          7276 => x"883f7e54",
          7277 => x"fdbc397b",
          7278 => x"75317083",
          7279 => x"ffff0642",
          7280 => x"54faac39",
          7281 => x"7781ffff",
          7282 => x"06763170",
          7283 => x"83ffff06",
          7284 => x"82173383",
          7285 => x"18337188",
          7286 => x"2b077010",
          7287 => x"10101b70",
          7288 => x"33811233",
          7289 => x"71982b71",
          7290 => x"902b0753",
          7291 => x"5e535458",
          7292 => x"58455473",
          7293 => x"8025f9f7",
          7294 => x"38ffbc39",
          7295 => x"617824fa",
          7296 => x"8338807a",
          7297 => x"248b8f38",
          7298 => x"7783ffff",
          7299 => x"065b617b",
          7300 => x"27fcdd38",
          7301 => x"fe8f3984",
          7302 => x"fff40b84",
          7303 => x"b9b80ca0",
          7304 => x"800b84b9",
          7305 => x"b4238280",
          7306 => x"80537e52",
          7307 => x"84fff451",
          7308 => x"fec4cc3f",
          7309 => x"84b9b808",
          7310 => x"5a7e7a34",
          7311 => x"810b811b",
          7312 => x"3484b9b8",
          7313 => x"08597e84",
          7314 => x"1a34810b",
          7315 => x"851a3484",
          7316 => x"b9b80858",
          7317 => x"7e861934",
          7318 => x"810b8719",
          7319 => x"3484b9b8",
          7320 => x"0884b9b4",
          7321 => x"22ff05fe",
          7322 => x"80800770",
          7323 => x"83ffff06",
          7324 => x"70882a58",
          7325 => x"56574474",
          7326 => x"64880534",
          7327 => x"73648905",
          7328 => x"3484b9b4",
          7329 => x"22701010",
          7330 => x"1084b9b8",
          7331 => x"0805f805",
          7332 => x"42437e61",
          7333 => x"82053481",
          7334 => x"61830534",
          7335 => x"fcee3980",
          7336 => x"7a2483de",
          7337 => x"386183ff",
          7338 => x"ff065b61",
          7339 => x"7b27fbc0",
          7340 => x"38fcf239",
          7341 => x"76802e82",
          7342 => x"bd387e51",
          7343 => x"eafb3f7f",
          7344 => x"547384b9",
          7345 => x"c80c953d",
          7346 => x"0d04761e",
          7347 => x"82113383",
          7348 => x"1233718b",
          7349 => x"2b71832b",
          7350 => x"077a1186",
          7351 => x"11338712",
          7352 => x"33718b2b",
          7353 => x"71832b07",
          7354 => x"7e058414",
          7355 => x"33851533",
          7356 => x"71882b07",
          7357 => x"70882a43",
          7358 => x"4445565b",
          7359 => x"4658535c",
          7360 => x"45567864",
          7361 => x"8405347a",
          7362 => x"64850534",
          7363 => x"84b9b808",
          7364 => x"70178411",
          7365 => x"33851233",
          7366 => x"718b2b71",
          7367 => x"832b0774",
          7368 => x"05861433",
          7369 => x"87153371",
          7370 => x"882b0770",
          7371 => x"882a5b41",
          7372 => x"42485d59",
          7373 => x"5d417364",
          7374 => x"8605347a",
          7375 => x"64870534",
          7376 => x"84b9b808",
          7377 => x"16703381",
          7378 => x"12337188",
          7379 => x"2b0781ff",
          7380 => x"ff067088",
          7381 => x"2a5f5c5a",
          7382 => x"5d7b7d34",
          7383 => x"79811e34",
          7384 => x"84b9b808",
          7385 => x"701f8211",
          7386 => x"33831233",
          7387 => x"718b2b71",
          7388 => x"832b0774",
          7389 => x"05733381",
          7390 => x"15337188",
          7391 => x"2b077088",
          7392 => x"2a5e5c5e",
          7393 => x"40435745",
          7394 => x"54767c34",
          7395 => x"75811d34",
          7396 => x"84b9b808",
          7397 => x"701f7033",
          7398 => x"81123371",
          7399 => x"8b2b7183",
          7400 => x"2b077405",
          7401 => x"82143383",
          7402 => x"15337188",
          7403 => x"2b077088",
          7404 => x"2a404740",
          7405 => x"5b405c55",
          7406 => x"55788218",
          7407 => x"34608318",
          7408 => x"3484b9b8",
          7409 => x"08701f82",
          7410 => x"11338312",
          7411 => x"3371882b",
          7412 => x"07665762",
          7413 => x"5670832b",
          7414 => x"4252585d",
          7415 => x"7e058405",
          7416 => x"51febdde",
          7417 => x"3f84b9b8",
          7418 => x"081e8405",
          7419 => x"7883ffff",
          7420 => x"065c5ffc",
          7421 => x"993984ff",
          7422 => x"f40b84b9",
          7423 => x"b80ca080",
          7424 => x"0b84b9b4",
          7425 => x"23828080",
          7426 => x"537f5284",
          7427 => x"fff451fe",
          7428 => x"c0ed3f84",
          7429 => x"b9b80856",
          7430 => x"7f763481",
          7431 => x"0b811734",
          7432 => x"84b9b808",
          7433 => x"557f8416",
          7434 => x"34810b85",
          7435 => x"163484b9",
          7436 => x"b808547f",
          7437 => x"86153481",
          7438 => x"0b871534",
          7439 => x"84b9b808",
          7440 => x"84b9b422",
          7441 => x"ff05fe80",
          7442 => x"80077083",
          7443 => x"ffff0670",
          7444 => x"882a4543",
          7445 => x"445e6188",
          7446 => x"1f346089",
          7447 => x"1f3484b9",
          7448 => x"b4227010",
          7449 => x"101084b9",
          7450 => x"b80805f8",
          7451 => x"055c5d7f",
          7452 => x"821c3481",
          7453 => x"0b831c34",
          7454 => x"7e51e7bd",
          7455 => x"3f7f54fc",
          7456 => x"c0398619",
          7457 => x"33871a33",
          7458 => x"718b2b71",
          7459 => x"832b0779",
          7460 => x"05841c33",
          7461 => x"851d3371",
          7462 => x"882b0770",
          7463 => x"882a5c48",
          7464 => x"5e435955",
          7465 => x"76618405",
          7466 => x"34636185",
          7467 => x"053484b9",
          7468 => x"b808701e",
          7469 => x"84113385",
          7470 => x"1233718b",
          7471 => x"2b71832b",
          7472 => x"07740586",
          7473 => x"14338715",
          7474 => x"3371882b",
          7475 => x"0770882a",
          7476 => x"415f4848",
          7477 => x"59565940",
          7478 => x"79648605",
          7479 => x"34786487",
          7480 => x"053484b9",
          7481 => x"b8081d70",
          7482 => x"33811233",
          7483 => x"71882b07",
          7484 => x"81ffff06",
          7485 => x"70882a59",
          7486 => x"42585875",
          7487 => x"78347f81",
          7488 => x"193484b9",
          7489 => x"b808701f",
          7490 => x"70338112",
          7491 => x"33718b2b",
          7492 => x"71832b07",
          7493 => x"74057033",
          7494 => x"81123371",
          7495 => x"882b0770",
          7496 => x"832b8fff",
          7497 => x"f8067705",
          7498 => x"63882a48",
          7499 => x"5d5d5a5d",
          7500 => x"405d4441",
          7501 => x"7f821734",
          7502 => x"7b831734",
          7503 => x"84b9b808",
          7504 => x"701f7033",
          7505 => x"81123371",
          7506 => x"8b2b7183",
          7507 => x"2b077405",
          7508 => x"70338112",
          7509 => x"3371882b",
          7510 => x"0781ffff",
          7511 => x"0670882a",
          7512 => x"485d5e5e",
          7513 => x"465a415b",
          7514 => x"60603476",
          7515 => x"60810534",
          7516 => x"6183ffff",
          7517 => x"065bfab3",
          7518 => x"39861533",
          7519 => x"87163371",
          7520 => x"8b2b7183",
          7521 => x"2b077905",
          7522 => x"84183385",
          7523 => x"19337188",
          7524 => x"2b077088",
          7525 => x"2a5e5e5a",
          7526 => x"52415d78",
          7527 => x"841e3479",
          7528 => x"851e3484",
          7529 => x"b9b80870",
          7530 => x"19841133",
          7531 => x"85123371",
          7532 => x"8b2b7183",
          7533 => x"2b077405",
          7534 => x"86143387",
          7535 => x"15337188",
          7536 => x"2b077088",
          7537 => x"2a44565e",
          7538 => x"525a4255",
          7539 => x"567c6086",
          7540 => x"05347560",
          7541 => x"87053484",
          7542 => x"b9b80818",
          7543 => x"70338112",
          7544 => x"3371882b",
          7545 => x"0781ffff",
          7546 => x"0670882a",
          7547 => x"5b5b5855",
          7548 => x"77753478",
          7549 => x"81163484",
          7550 => x"b9b80870",
          7551 => x"1f703381",
          7552 => x"1233718b",
          7553 => x"2b71832b",
          7554 => x"07740570",
          7555 => x"33811233",
          7556 => x"71882b07",
          7557 => x"70832b8f",
          7558 => x"fff80677",
          7559 => x"0563882a",
          7560 => x"56545f5f",
          7561 => x"5859425e",
          7562 => x"557f8217",
          7563 => x"347b8317",
          7564 => x"3484b9b8",
          7565 => x"08701f70",
          7566 => x"33811233",
          7567 => x"718b2b71",
          7568 => x"832b0774",
          7569 => x"05703381",
          7570 => x"12337188",
          7571 => x"2b0781ff",
          7572 => x"ff067088",
          7573 => x"2a5d545e",
          7574 => x"585b595d",
          7575 => x"55757c34",
          7576 => x"76811d34",
          7577 => x"84b9b808",
          7578 => x"701f8211",
          7579 => x"33831233",
          7580 => x"718b2b71",
          7581 => x"832b0774",
          7582 => x"11861133",
          7583 => x"87123371",
          7584 => x"8b2b7183",
          7585 => x"2b077805",
          7586 => x"84143385",
          7587 => x"15337188",
          7588 => x"2b077088",
          7589 => x"2a595749",
          7590 => x"525c4259",
          7591 => x"535d5a57",
          7592 => x"5777841d",
          7593 => x"3479851d",
          7594 => x"3484b9b8",
          7595 => x"08701784",
          7596 => x"11338512",
          7597 => x"33718b2b",
          7598 => x"71832b07",
          7599 => x"74058614",
          7600 => x"33871533",
          7601 => x"71882b07",
          7602 => x"70882a5f",
          7603 => x"425e5240",
          7604 => x"57415777",
          7605 => x"8616347b",
          7606 => x"87163484",
          7607 => x"b9b80816",
          7608 => x"70338112",
          7609 => x"3371882b",
          7610 => x"0781ffff",
          7611 => x"0670882a",
          7612 => x"5a5c5e59",
          7613 => x"76793479",
          7614 => x"811a3484",
          7615 => x"b9b80870",
          7616 => x"1f821133",
          7617 => x"83123371",
          7618 => x"8b2b7183",
          7619 => x"2b077405",
          7620 => x"73338115",
          7621 => x"3371882b",
          7622 => x"0770882a",
          7623 => x"415c455d",
          7624 => x"5f5a5555",
          7625 => x"79793475",
          7626 => x"811a3484",
          7627 => x"b9b80870",
          7628 => x"1f703381",
          7629 => x"1233718b",
          7630 => x"2b71832b",
          7631 => x"07740582",
          7632 => x"14338315",
          7633 => x"3371882b",
          7634 => x"0770882a",
          7635 => x"415c455d",
          7636 => x"5f5a5555",
          7637 => x"79821a34",
          7638 => x"75831a34",
          7639 => x"84b9b808",
          7640 => x"701f8211",
          7641 => x"33831233",
          7642 => x"71882b07",
          7643 => x"66576256",
          7644 => x"70832b42",
          7645 => x"525a5d7e",
          7646 => x"05840551",
          7647 => x"feb6c33f",
          7648 => x"84b9b808",
          7649 => x"1e840561",
          7650 => x"65051c70",
          7651 => x"83ffff06",
          7652 => x"5d445ff1",
          7653 => x"d5398619",
          7654 => x"33871a33",
          7655 => x"718b2b71",
          7656 => x"832b0779",
          7657 => x"05841c33",
          7658 => x"851d3371",
          7659 => x"882b0770",
          7660 => x"882a4048",
          7661 => x"5d434155",
          7662 => x"7a618405",
          7663 => x"34636185",
          7664 => x"053484b9",
          7665 => x"b808701e",
          7666 => x"84113385",
          7667 => x"1233718b",
          7668 => x"2b71832b",
          7669 => x"07740586",
          7670 => x"14338715",
          7671 => x"3371882b",
          7672 => x"0770882a",
          7673 => x"5b415f48",
          7674 => x"5c594156",
          7675 => x"73648605",
          7676 => x"347a6487",
          7677 => x"053484b9",
          7678 => x"b8081d70",
          7679 => x"33811233",
          7680 => x"71882b07",
          7681 => x"81ffff06",
          7682 => x"70882a5c",
          7683 => x"5f425578",
          7684 => x"75347c81",
          7685 => x"163484b9",
          7686 => x"b808701f",
          7687 => x"70338112",
          7688 => x"33718b2b",
          7689 => x"71832b07",
          7690 => x"74057033",
          7691 => x"81123371",
          7692 => x"882b0770",
          7693 => x"832b8fff",
          7694 => x"f8067705",
          7695 => x"63882a5d",
          7696 => x"445c4958",
          7697 => x"5e455840",
          7698 => x"74821e34",
          7699 => x"7b831e34",
          7700 => x"84b9b808",
          7701 => x"701f7033",
          7702 => x"81123371",
          7703 => x"8b2b7183",
          7704 => x"2b077405",
          7705 => x"70338112",
          7706 => x"3371882b",
          7707 => x"0781ffff",
          7708 => x"0670882a",
          7709 => x"475f4958",
          7710 => x"46595e5b",
          7711 => x"7f7d3478",
          7712 => x"811e3477",
          7713 => x"83ffff06",
          7714 => x"5bf38339",
          7715 => x"7e605254",
          7716 => x"e5a13f84",
          7717 => x"b9c8085f",
          7718 => x"84b9c808",
          7719 => x"802e9338",
          7720 => x"62537352",
          7721 => x"84b9c808",
          7722 => x"51feb5be",
          7723 => x"3f7351df",
          7724 => x"883f615b",
          7725 => x"617b27ef",
          7726 => x"b738f0e9",
          7727 => x"39f93d0d",
          7728 => x"7a7a2984",
          7729 => x"b9b80858",
          7730 => x"5876802e",
          7731 => x"b7387754",
          7732 => x"778a3873",
          7733 => x"84b9c80c",
          7734 => x"893d0d04",
          7735 => x"7751e4d3",
          7736 => x"3f84b9c8",
          7737 => x"085484b9",
          7738 => x"c808802e",
          7739 => x"e6387753",
          7740 => x"805284b9",
          7741 => x"c80851fe",
          7742 => x"b7853f73",
          7743 => x"84b9c80c",
          7744 => x"893d0d04",
          7745 => x"84fff40b",
          7746 => x"84b9b80c",
          7747 => x"a0800b84",
          7748 => x"b9b42382",
          7749 => x"80805376",
          7750 => x"5284fff4",
          7751 => x"51feb6df",
          7752 => x"3f84b9b8",
          7753 => x"08557675",
          7754 => x"34810b81",
          7755 => x"163484b9",
          7756 => x"b8085476",
          7757 => x"84153481",
          7758 => x"0b851534",
          7759 => x"84b9b808",
          7760 => x"56768617",
          7761 => x"34810b87",
          7762 => x"173484b9",
          7763 => x"b80884b9",
          7764 => x"b422ff05",
          7765 => x"fe808007",
          7766 => x"7083ffff",
          7767 => x"0670882a",
          7768 => x"58515556",
          7769 => x"74881734",
          7770 => x"73891734",
          7771 => x"84b9b422",
          7772 => x"70101010",
          7773 => x"84b9b808",
          7774 => x"05f80555",
          7775 => x"55768215",
          7776 => x"34810b83",
          7777 => x"15347754",
          7778 => x"77802efe",
          7779 => x"c638fecc",
          7780 => x"39ff3d0d",
          7781 => x"028f0533",
          7782 => x"51815270",
          7783 => x"72268738",
          7784 => x"84b9c411",
          7785 => x"33527184",
          7786 => x"b9c80c83",
          7787 => x"3d0d04fe",
          7788 => x"3d0d0293",
          7789 => x"05335283",
          7790 => x"53718126",
          7791 => x"9d387151",
          7792 => x"d4bb3f84",
          7793 => x"b9c80881",
          7794 => x"ff065372",
          7795 => x"87387284",
          7796 => x"b9c41334",
          7797 => x"84b9c412",
          7798 => x"33537284",
          7799 => x"b9c80c84",
          7800 => x"3d0d04f7",
          7801 => x"3d0d7c7e",
          7802 => x"60028c05",
          7803 => x"af05335a",
          7804 => x"5c575981",
          7805 => x"54767426",
          7806 => x"873884b9",
          7807 => x"c4173354",
          7808 => x"73810654",
          7809 => x"835573bd",
          7810 => x"38735885",
          7811 => x"0b87c098",
          7812 => x"8c0c7853",
          7813 => x"75527651",
          7814 => x"d5ca3f84",
          7815 => x"b9c80881",
          7816 => x"ff065574",
          7817 => x"802ea738",
          7818 => x"87c0988c",
          7819 => x"085473e2",
          7820 => x"38797826",
          7821 => x"d63874fc",
          7822 => x"80800654",
          7823 => x"73802e83",
          7824 => x"38815473",
          7825 => x"557484b9",
          7826 => x"c80c8b3d",
          7827 => x"0d048480",
          7828 => x"16811970",
          7829 => x"81ff065a",
          7830 => x"55567978",
          7831 => x"26ffac38",
          7832 => x"d539f73d",
          7833 => x"0d7c7e60",
          7834 => x"028c05af",
          7835 => x"05335a5c",
          7836 => x"57598154",
          7837 => x"76742687",
          7838 => x"3884b9c4",
          7839 => x"17335473",
          7840 => x"81065483",
          7841 => x"5573bd38",
          7842 => x"7358850b",
          7843 => x"87c0988c",
          7844 => x"0c785375",
          7845 => x"527651d7",
          7846 => x"8e3f84b9",
          7847 => x"c80881ff",
          7848 => x"06557480",
          7849 => x"2ea73887",
          7850 => x"c0988c08",
          7851 => x"5473e238",
          7852 => x"797826d6",
          7853 => x"3874fc80",
          7854 => x"80065473",
          7855 => x"802e8338",
          7856 => x"81547355",
          7857 => x"7484b9c8",
          7858 => x"0c8b3d0d",
          7859 => x"04848016",
          7860 => x"81197081",
          7861 => x"ff065a55",
          7862 => x"56797826",
          7863 => x"ffac38d5",
          7864 => x"39fc3d0d",
          7865 => x"78028405",
          7866 => x"9b053302",
          7867 => x"88059f05",
          7868 => x"33535355",
          7869 => x"81537173",
          7870 => x"26873884",
          7871 => x"b9c41233",
          7872 => x"53728106",
          7873 => x"54835373",
          7874 => x"9b38850b",
          7875 => x"87c0988c",
          7876 => x"0c815370",
          7877 => x"732e9638",
          7878 => x"727125ad",
          7879 => x"3870832e",
          7880 => x"9a388453",
          7881 => x"7284b9c8",
          7882 => x"0c863d0d",
          7883 => x"0488800a",
          7884 => x"750c7384",
          7885 => x"b9c80c86",
          7886 => x"3d0d0481",
          7887 => x"80750c80",
          7888 => x"0b84b9c8",
          7889 => x"0c863d0d",
          7890 => x"0471842b",
          7891 => x"87c0928c",
          7892 => x"11535470",
          7893 => x"cd387108",
          7894 => x"70812a81",
          7895 => x"06515170",
          7896 => x"802e8a38",
          7897 => x"87c0988c",
          7898 => x"085574ea",
          7899 => x"3887c098",
          7900 => x"8c085170",
          7901 => x"ca388172",
          7902 => x"0c87c092",
          7903 => x"8c145271",
          7904 => x"08820654",
          7905 => x"73802eff",
          7906 => x"9b387108",
          7907 => x"82065473",
          7908 => x"ee38ff90",
          7909 => x"39f63d0d",
          7910 => x"7c58800b",
          7911 => x"83193371",
          7912 => x"5b565774",
          7913 => x"772e0981",
          7914 => x"06a83877",
          7915 => x"33567583",
          7916 => x"2e818738",
          7917 => x"80538052",
          7918 => x"81183351",
          7919 => x"fea33f84",
          7920 => x"b9c80880",
          7921 => x"2e833881",
          7922 => x"597884b9",
          7923 => x"c80c8c3d",
          7924 => x"0d048154",
          7925 => x"b4180853",
          7926 => x"b8187053",
          7927 => x"81193352",
          7928 => x"5afcff3f",
          7929 => x"815984b9",
          7930 => x"c808772e",
          7931 => x"098106d9",
          7932 => x"3884b9c8",
          7933 => x"08831934",
          7934 => x"b4180870",
          7935 => x"a81a0831",
          7936 => x"a01a0884",
          7937 => x"b9c8085c",
          7938 => x"58565b74",
          7939 => x"7627ff9b",
          7940 => x"38821833",
          7941 => x"5574822e",
          7942 => x"098106ff",
          7943 => x"8e388154",
          7944 => x"751b5379",
          7945 => x"52811833",
          7946 => x"51fcb73f",
          7947 => x"76783357",
          7948 => x"5975832e",
          7949 => x"098106fe",
          7950 => x"fb388418",
          7951 => x"33577681",
          7952 => x"2e098106",
          7953 => x"feee38b8",
          7954 => x"185a8480",
          7955 => x"7a565780",
          7956 => x"75708105",
          7957 => x"5734ff17",
          7958 => x"5776f438",
          7959 => x"80d50b84",
          7960 => x"b61934ff",
          7961 => x"aa0b84b7",
          7962 => x"193480d2",
          7963 => x"7a3480d2",
          7964 => x"0bb91934",
          7965 => x"80e10bba",
          7966 => x"193480c1",
          7967 => x"0bbb1934",
          7968 => x"80f20b84",
          7969 => x"9c193480",
          7970 => x"f20b849d",
          7971 => x"193480c1",
          7972 => x"0b849e19",
          7973 => x"3480e10b",
          7974 => x"849f1934",
          7975 => x"94180855",
          7976 => x"7484a019",
          7977 => x"3474882a",
          7978 => x"5b7a84a1",
          7979 => x"19347490",
          7980 => x"2a567584",
          7981 => x"a2193474",
          7982 => x"982a5b7a",
          7983 => x"84a31934",
          7984 => x"9018085b",
          7985 => x"7a84a419",
          7986 => x"347a882a",
          7987 => x"557484a5",
          7988 => x"19347a90",
          7989 => x"2a567584",
          7990 => x"a619347a",
          7991 => x"982a5574",
          7992 => x"84a71934",
          7993 => x"a4180881",
          7994 => x"0570b41a",
          7995 => x"0c5b8154",
          7996 => x"7a537952",
          7997 => x"81183351",
          7998 => x"fae83f76",
          7999 => x"84193480",
          8000 => x"53805281",
          8001 => x"183351fb",
          8002 => x"d83f84b9",
          8003 => x"c808802e",
          8004 => x"fdb738fd",
          8005 => x"b239f33d",
          8006 => x"0d606070",
          8007 => x"08595656",
          8008 => x"81762788",
          8009 => x"389c1708",
          8010 => x"76268c38",
          8011 => x"81587784",
          8012 => x"b9c80c8f",
          8013 => x"3d0d04ff",
          8014 => x"77335658",
          8015 => x"74822e81",
          8016 => x"cc387482",
          8017 => x"2482a538",
          8018 => x"74812e09",
          8019 => x"8106dd38",
          8020 => x"75812a16",
          8021 => x"70892aa8",
          8022 => x"1908055a",
          8023 => x"5a805bb4",
          8024 => x"1708792e",
          8025 => x"b0388317",
          8026 => x"335c7b7b",
          8027 => x"2e098106",
          8028 => x"83de3881",
          8029 => x"547853b8",
          8030 => x"17528117",
          8031 => x"3351f8e3",
          8032 => x"3f84b9c8",
          8033 => x"08802e85",
          8034 => x"38ff5981",
          8035 => x"5b78b418",
          8036 => x"0c7aff9a",
          8037 => x"387983ff",
          8038 => x"0617b811",
          8039 => x"33811c70",
          8040 => x"892aa81b",
          8041 => x"0805535d",
          8042 => x"5d59b417",
          8043 => x"08792eb5",
          8044 => x"38800b83",
          8045 => x"1833715c",
          8046 => x"565d747d",
          8047 => x"2e098106",
          8048 => x"84b53881",
          8049 => x"547853b8",
          8050 => x"17528117",
          8051 => x"3351f893",
          8052 => x"3f84b9c8",
          8053 => x"08802e85",
          8054 => x"38ff5981",
          8055 => x"5a78b418",
          8056 => x"0c79feca",
          8057 => x"387a83ff",
          8058 => x"0617b811",
          8059 => x"3370882b",
          8060 => x"7e077881",
          8061 => x"0671842a",
          8062 => x"535d5959",
          8063 => x"5d79feae",
          8064 => x"38769fff",
          8065 => x"0684b9c8",
          8066 => x"0c8f3d0d",
          8067 => x"0475882a",
          8068 => x"a8180805",
          8069 => x"59b41708",
          8070 => x"792eb538",
          8071 => x"800b8318",
          8072 => x"33715c5d",
          8073 => x"5b7b7b2e",
          8074 => x"09810681",
          8075 => x"c2388154",
          8076 => x"7853b817",
          8077 => x"52811733",
          8078 => x"51f7a83f",
          8079 => x"84b9c808",
          8080 => x"802e8538",
          8081 => x"ff59815a",
          8082 => x"78b4180c",
          8083 => x"79fddf38",
          8084 => x"751083fe",
          8085 => x"067705b8",
          8086 => x"05811133",
          8087 => x"71337188",
          8088 => x"2b0784b9",
          8089 => x"c80c575b",
          8090 => x"8f3d0d04",
          8091 => x"74832e09",
          8092 => x"8106fdb8",
          8093 => x"3875872a",
          8094 => x"a8180805",
          8095 => x"59b41708",
          8096 => x"792eb538",
          8097 => x"800b8318",
          8098 => x"33715c5e",
          8099 => x"5b7c7b2e",
          8100 => x"09810682",
          8101 => x"81388154",
          8102 => x"7853b817",
          8103 => x"52811733",
          8104 => x"51f6c03f",
          8105 => x"84b9c808",
          8106 => x"802e8538",
          8107 => x"ff59815a",
          8108 => x"78b4180c",
          8109 => x"79fcf738",
          8110 => x"75822b83",
          8111 => x"fc067705",
          8112 => x"b8058311",
          8113 => x"33821233",
          8114 => x"71902b71",
          8115 => x"882b0781",
          8116 => x"14337072",
          8117 => x"07882b75",
          8118 => x"337180ff",
          8119 => x"fffe8006",
          8120 => x"0784b9c8",
          8121 => x"0c415c5e",
          8122 => x"595a568f",
          8123 => x"3d0d0481",
          8124 => x"54b41708",
          8125 => x"53b81770",
          8126 => x"53811833",
          8127 => x"525cf6e2",
          8128 => x"3f815a84",
          8129 => x"b9c8087b",
          8130 => x"2e098106",
          8131 => x"febe3884",
          8132 => x"b9c80883",
          8133 => x"1834b417",
          8134 => x"08a81808",
          8135 => x"3184b9c8",
          8136 => x"085b5e7d",
          8137 => x"a0180827",
          8138 => x"fe843882",
          8139 => x"17335574",
          8140 => x"822e0981",
          8141 => x"06fdf738",
          8142 => x"8154b417",
          8143 => x"08a01808",
          8144 => x"05537b52",
          8145 => x"81173351",
          8146 => x"f6983f7a",
          8147 => x"5afddf39",
          8148 => x"8154b417",
          8149 => x"0853b817",
          8150 => x"70538118",
          8151 => x"33525cf6",
          8152 => x"813f84b9",
          8153 => x"c8087b2e",
          8154 => x"09810682",
          8155 => x"813884b9",
          8156 => x"c8088318",
          8157 => x"34b41708",
          8158 => x"a8180831",
          8159 => x"5d7ca018",
          8160 => x"08278b38",
          8161 => x"8217335e",
          8162 => x"7d822e81",
          8163 => x"cb3884b9",
          8164 => x"c8085bfb",
          8165 => x"de398154",
          8166 => x"b4170853",
          8167 => x"b8177053",
          8168 => x"81183352",
          8169 => x"5cf5bb3f",
          8170 => x"815a84b9",
          8171 => x"c8087b2e",
          8172 => x"098106fd",
          8173 => x"ff3884b9",
          8174 => x"c8088318",
          8175 => x"34b41708",
          8176 => x"a8180831",
          8177 => x"84b9c808",
          8178 => x"5b5e7da0",
          8179 => x"180827fd",
          8180 => x"c5388217",
          8181 => x"33557482",
          8182 => x"2e098106",
          8183 => x"fdb83881",
          8184 => x"54b41708",
          8185 => x"a0180805",
          8186 => x"537b5281",
          8187 => x"173351f4",
          8188 => x"f13f7a5a",
          8189 => x"fda03981",
          8190 => x"54b41708",
          8191 => x"53b81770",
          8192 => x"53811833",
          8193 => x"525ef4da",
          8194 => x"3f815a84",
          8195 => x"b9c8087d",
          8196 => x"2e098106",
          8197 => x"fbcb3884",
          8198 => x"b9c80883",
          8199 => x"1834b417",
          8200 => x"08a81808",
          8201 => x"3184b9c8",
          8202 => x"085b5574",
          8203 => x"a0180827",
          8204 => x"fb913882",
          8205 => x"17335574",
          8206 => x"822e0981",
          8207 => x"06fb8438",
          8208 => x"8154b417",
          8209 => x"08a01808",
          8210 => x"05537d52",
          8211 => x"81173351",
          8212 => x"f4903f7c",
          8213 => x"5afaec39",
          8214 => x"8154b417",
          8215 => x"08a01808",
          8216 => x"05537b52",
          8217 => x"81173351",
          8218 => x"f3f83ffa",
          8219 => x"8639815b",
          8220 => x"7af9bb38",
          8221 => x"fa9f39f2",
          8222 => x"3d0d6062",
          8223 => x"645d5759",
          8224 => x"82588176",
          8225 => x"279c3875",
          8226 => x"9c1a0827",
          8227 => x"95387833",
          8228 => x"5574782e",
          8229 => x"96387478",
          8230 => x"24818038",
          8231 => x"74812e82",
          8232 => x"8a387784",
          8233 => x"b9c80c90",
          8234 => x"3d0d0475",
          8235 => x"882aa81a",
          8236 => x"08055880",
          8237 => x"0bb41a08",
          8238 => x"585c7678",
          8239 => x"2e86b638",
          8240 => x"8319337c",
          8241 => x"5b5d7c7c",
          8242 => x"2e098106",
          8243 => x"83fa3881",
          8244 => x"547753b8",
          8245 => x"19528119",
          8246 => x"3351f287",
          8247 => x"3f84b9c8",
          8248 => x"08802e85",
          8249 => x"38ff5881",
          8250 => x"5a77b41a",
          8251 => x"0c795879",
          8252 => x"ffb03875",
          8253 => x"1083fe06",
          8254 => x"79057b83",
          8255 => x"ffff0658",
          8256 => x"5e76b81f",
          8257 => x"3476882a",
          8258 => x"5a79b91f",
          8259 => x"34810b83",
          8260 => x"1a347784",
          8261 => x"b9c80c90",
          8262 => x"3d0d0474",
          8263 => x"832e0981",
          8264 => x"06feff38",
          8265 => x"75872aa8",
          8266 => x"1a080558",
          8267 => x"800bb41a",
          8268 => x"08585c76",
          8269 => x"782e85e1",
          8270 => x"38831933",
          8271 => x"7c5b5d7c",
          8272 => x"7c2e0981",
          8273 => x"0684bd38",
          8274 => x"81547753",
          8275 => x"b8195281",
          8276 => x"193351f1",
          8277 => x"8e3f84b9",
          8278 => x"c808802e",
          8279 => x"8538ff58",
          8280 => x"815a77b4",
          8281 => x"1a0c7958",
          8282 => x"79feb738",
          8283 => x"75822b83",
          8284 => x"fc067905",
          8285 => x"b8118311",
          8286 => x"3370982b",
          8287 => x"8f0a067e",
          8288 => x"f00a0607",
          8289 => x"41575e5c",
          8290 => x"7d7d347d",
          8291 => x"882a5675",
          8292 => x"b91d347d",
          8293 => x"902a5a79",
          8294 => x"ba1d347d",
          8295 => x"982a5b7a",
          8296 => x"bb1d3481",
          8297 => x"0b831a34",
          8298 => x"fee83975",
          8299 => x"812a1670",
          8300 => x"892aa81b",
          8301 => x"0805b41b",
          8302 => x"0859595a",
          8303 => x"76782eb7",
          8304 => x"38800b83",
          8305 => x"1a33715e",
          8306 => x"565d747d",
          8307 => x"2e098106",
          8308 => x"82d43881",
          8309 => x"547753b8",
          8310 => x"19528119",
          8311 => x"3351f083",
          8312 => x"3f84b9c8",
          8313 => x"08802e85",
          8314 => x"38ff5881",
          8315 => x"5c77b41a",
          8316 => x"0c7b587b",
          8317 => x"fdac3879",
          8318 => x"83ff0619",
          8319 => x"b805811b",
          8320 => x"7781065f",
          8321 => x"5f577a55",
          8322 => x"7c802e8f",
          8323 => x"387a842b",
          8324 => x"9ff00677",
          8325 => x"338f0671",
          8326 => x"07565a74",
          8327 => x"7734810b",
          8328 => x"831a347d",
          8329 => x"892aa81a",
          8330 => x"08055680",
          8331 => x"0bb41a08",
          8332 => x"565f7476",
          8333 => x"2e83dd38",
          8334 => x"81547453",
          8335 => x"b8197053",
          8336 => x"811a3352",
          8337 => x"57f09b3f",
          8338 => x"815884b9",
          8339 => x"c8087f2e",
          8340 => x"09810680",
          8341 => x"c73884b9",
          8342 => x"c808831a",
          8343 => x"34b41908",
          8344 => x"70a81b08",
          8345 => x"31a01b08",
          8346 => x"84b9c808",
          8347 => x"5b5c565c",
          8348 => x"747a278b",
          8349 => x"38821933",
          8350 => x"5574822e",
          8351 => x"82e43881",
          8352 => x"54755376",
          8353 => x"52811933",
          8354 => x"51eed83f",
          8355 => x"84b9c808",
          8356 => x"802e8538",
          8357 => x"ff568158",
          8358 => x"75b41a0c",
          8359 => x"77fc8338",
          8360 => x"7d83ff06",
          8361 => x"19b8057b",
          8362 => x"842a5656",
          8363 => x"7c8f387a",
          8364 => x"882a7633",
          8365 => x"81f00671",
          8366 => x"8f060756",
          8367 => x"5c747634",
          8368 => x"810b831a",
          8369 => x"34fccb39",
          8370 => x"81547653",
          8371 => x"b8197053",
          8372 => x"811a3352",
          8373 => x"5def8b3f",
          8374 => x"815a84b9",
          8375 => x"c8087c2e",
          8376 => x"098106fc",
          8377 => x"883884b9",
          8378 => x"c808831a",
          8379 => x"34b41908",
          8380 => x"70a81b08",
          8381 => x"31a01b08",
          8382 => x"84b9c808",
          8383 => x"5d59405e",
          8384 => x"7e7727fb",
          8385 => x"ca388219",
          8386 => x"33557482",
          8387 => x"2e098106",
          8388 => x"fbbd3881",
          8389 => x"54761e53",
          8390 => x"7c528119",
          8391 => x"3351eec2",
          8392 => x"3f7b5afb",
          8393 => x"aa398154",
          8394 => x"7653b819",
          8395 => x"7053811a",
          8396 => x"335257ee",
          8397 => x"ad3f815c",
          8398 => x"84b9c808",
          8399 => x"7d2e0981",
          8400 => x"06fdae38",
          8401 => x"84b9c808",
          8402 => x"831a34b4",
          8403 => x"190870a8",
          8404 => x"1b0831a0",
          8405 => x"1b0884b9",
          8406 => x"c8085f40",
          8407 => x"565f747e",
          8408 => x"27fcf038",
          8409 => x"82193355",
          8410 => x"74822e09",
          8411 => x"8106fce3",
          8412 => x"3881547d",
          8413 => x"1f537652",
          8414 => x"81193351",
          8415 => x"ede43f7c",
          8416 => x"5cfcd039",
          8417 => x"81547653",
          8418 => x"b8197053",
          8419 => x"811a3352",
          8420 => x"57edcf3f",
          8421 => x"815a84b9",
          8422 => x"c8087c2e",
          8423 => x"098106fb",
          8424 => x"c53884b9",
          8425 => x"c808831a",
          8426 => x"34b41908",
          8427 => x"70a81b08",
          8428 => x"31a01b08",
          8429 => x"84b9c808",
          8430 => x"5d5f405e",
          8431 => x"7e7d27fb",
          8432 => x"87388219",
          8433 => x"33557482",
          8434 => x"2e098106",
          8435 => x"fafa3881",
          8436 => x"547c1e53",
          8437 => x"76528119",
          8438 => x"3351ed86",
          8439 => x"3f7b5afa",
          8440 => x"e7398154",
          8441 => x"791c5376",
          8442 => x"52811933",
          8443 => x"51ecf33f",
          8444 => x"7e58fd8b",
          8445 => x"397b7610",
          8446 => x"83fe067a",
          8447 => x"057c83ff",
          8448 => x"ff06595f",
          8449 => x"5876b81f",
          8450 => x"3476882a",
          8451 => x"5a79b91f",
          8452 => x"34f9fa39",
          8453 => x"7e58fd88",
          8454 => x"397b7682",
          8455 => x"2b83fc06",
          8456 => x"7a05b811",
          8457 => x"83113370",
          8458 => x"982b8f0a",
          8459 => x"067ff00a",
          8460 => x"06074258",
          8461 => x"5f5d587d",
          8462 => x"7d347d88",
          8463 => x"2a5675b9",
          8464 => x"1d347d90",
          8465 => x"2a5a79ba",
          8466 => x"1d347d98",
          8467 => x"2a5b7abb",
          8468 => x"1d34facf",
          8469 => x"39f63d0d",
          8470 => x"7c7e7108",
          8471 => x"5b5c5a7a",
          8472 => x"818a3890",
          8473 => x"19085776",
          8474 => x"802e80f4",
          8475 => x"38769c1a",
          8476 => x"082780ec",
          8477 => x"38941908",
          8478 => x"70565473",
          8479 => x"802e80d7",
          8480 => x"38767b2e",
          8481 => x"81933876",
          8482 => x"56811656",
          8483 => x"9c190876",
          8484 => x"26893882",
          8485 => x"56757726",
          8486 => x"82b23875",
          8487 => x"527951f0",
          8488 => x"f53f84b9",
          8489 => x"c808802e",
          8490 => x"81d03880",
          8491 => x"5884b9c8",
          8492 => x"08812eb1",
          8493 => x"3884b9c8",
          8494 => x"08097030",
          8495 => x"70720780",
          8496 => x"25707b07",
          8497 => x"51515555",
          8498 => x"7382aa38",
          8499 => x"75772e09",
          8500 => x"8106ffb5",
          8501 => x"38735574",
          8502 => x"84b9c80c",
          8503 => x"8c3d0d04",
          8504 => x"8157ff91",
          8505 => x"3984b9c8",
          8506 => x"0858ca39",
          8507 => x"7a527951",
          8508 => x"f0a43f81",
          8509 => x"557484b9",
          8510 => x"c80827db",
          8511 => x"3884b9c8",
          8512 => x"085584b9",
          8513 => x"c808ff2e",
          8514 => x"ce389c19",
          8515 => x"0884b9c8",
          8516 => x"0826c438",
          8517 => x"7a57fedd",
          8518 => x"39811b56",
          8519 => x"9c190876",
          8520 => x"26833882",
          8521 => x"56755279",
          8522 => x"51efeb3f",
          8523 => x"805884b9",
          8524 => x"c808812e",
          8525 => x"81a03884",
          8526 => x"b9c80809",
          8527 => x"70307072",
          8528 => x"07802570",
          8529 => x"7b0784b9",
          8530 => x"c8085451",
          8531 => x"51555573",
          8532 => x"ff853884",
          8533 => x"b9c80880",
          8534 => x"2e9a3890",
          8535 => x"19085481",
          8536 => x"7427fea3",
          8537 => x"38739c1a",
          8538 => x"0827fe9b",
          8539 => x"38737057",
          8540 => x"57fe9639",
          8541 => x"75802efe",
          8542 => x"8e38ff53",
          8543 => x"75527851",
          8544 => x"f5f53f84",
          8545 => x"b9c80884",
          8546 => x"b9c80830",
          8547 => x"7084b9c8",
          8548 => x"08078025",
          8549 => x"5658557a",
          8550 => x"80c43874",
          8551 => x"80e33875",
          8552 => x"901a0c9c",
          8553 => x"1908fe05",
          8554 => x"941a0856",
          8555 => x"58747826",
          8556 => x"8638ff15",
          8557 => x"941a0c84",
          8558 => x"19338107",
          8559 => x"5a79841a",
          8560 => x"34755574",
          8561 => x"84b9c80c",
          8562 => x"8c3d0d04",
          8563 => x"800b84b9",
          8564 => x"c80c8c3d",
          8565 => x"0d0484b9",
          8566 => x"c80858fe",
          8567 => x"da397380",
          8568 => x"2effb838",
          8569 => x"75537a52",
          8570 => x"7851f58b",
          8571 => x"3f84b9c8",
          8572 => x"0855ffa7",
          8573 => x"3984b9c8",
          8574 => x"0884b9c8",
          8575 => x"0c8c3d0d",
          8576 => x"04ff5674",
          8577 => x"812effb9",
          8578 => x"388155ff",
          8579 => x"b639f83d",
          8580 => x"0d7a7c71",
          8581 => x"08595558",
          8582 => x"73f0800a",
          8583 => x"2680df38",
          8584 => x"739f0653",
          8585 => x"7280d738",
          8586 => x"7390190c",
          8587 => x"88180855",
          8588 => x"7480df38",
          8589 => x"76335675",
          8590 => x"822680cc",
          8591 => x"3873852a",
          8592 => x"53820b88",
          8593 => x"18225a56",
          8594 => x"727927a9",
          8595 => x"38ac1708",
          8596 => x"98190c74",
          8597 => x"94190c98",
          8598 => x"18085382",
          8599 => x"5672802e",
          8600 => x"94387389",
          8601 => x"2a139819",
          8602 => x"0c7383ff",
          8603 => x"0617b805",
          8604 => x"9c190c80",
          8605 => x"567584b9",
          8606 => x"c80c8a3d",
          8607 => x"0d04820b",
          8608 => x"84b9c80c",
          8609 => x"8a3d0d04",
          8610 => x"ac170855",
          8611 => x"74802eff",
          8612 => x"ac388a17",
          8613 => x"2270892b",
          8614 => x"57597376",
          8615 => x"27a5389c",
          8616 => x"170853fe",
          8617 => x"15fe1454",
          8618 => x"56805975",
          8619 => x"73278d38",
          8620 => x"8a172276",
          8621 => x"7129b019",
          8622 => x"08055a53",
          8623 => x"7898190c",
          8624 => x"ff913974",
          8625 => x"527751ec",
          8626 => x"cd3f84b9",
          8627 => x"c8085584",
          8628 => x"b9c808ff",
          8629 => x"2ea43881",
          8630 => x"0b84b9c8",
          8631 => x"0827ff9e",
          8632 => x"389c1708",
          8633 => x"5384b9c8",
          8634 => x"087327ff",
          8635 => x"91387376",
          8636 => x"31547376",
          8637 => x"27cd38ff",
          8638 => x"aa39810b",
          8639 => x"84b9c80c",
          8640 => x"8a3d0d04",
          8641 => x"f33d0d7f",
          8642 => x"70089012",
          8643 => x"08a0055c",
          8644 => x"5a57f080",
          8645 => x"0a7a2786",
          8646 => x"38800b98",
          8647 => x"180c9817",
          8648 => x"08558456",
          8649 => x"74802eb2",
          8650 => x"387983ff",
          8651 => x"065b7a9d",
          8652 => x"38811594",
          8653 => x"18085758",
          8654 => x"75a93879",
          8655 => x"852a881a",
          8656 => x"22575574",
          8657 => x"762781f5",
          8658 => x"38779818",
          8659 => x"0c799018",
          8660 => x"0c781bb8",
          8661 => x"059c180c",
          8662 => x"80567584",
          8663 => x"b9c80c8f",
          8664 => x"3d0d0477",
          8665 => x"98180c8a",
          8666 => x"1922ff05",
          8667 => x"7a892a06",
          8668 => x"5c7bda38",
          8669 => x"75527651",
          8670 => x"eb9c3f84",
          8671 => x"b9c8085d",
          8672 => x"8256810b",
          8673 => x"84b9c808",
          8674 => x"27d03881",
          8675 => x"5684b9c8",
          8676 => x"08ff2ec6",
          8677 => x"389c1908",
          8678 => x"84b9c808",
          8679 => x"26829138",
          8680 => x"60802e81",
          8681 => x"98389417",
          8682 => x"08527651",
          8683 => x"f9a73f84",
          8684 => x"b9c8085d",
          8685 => x"875684b9",
          8686 => x"c808802e",
          8687 => x"ff9c3882",
          8688 => x"5684b9c8",
          8689 => x"08812eff",
          8690 => x"91388156",
          8691 => x"84b9c808",
          8692 => x"ff2eff86",
          8693 => x"3884b9c8",
          8694 => x"08831a33",
          8695 => x"5f587d80",
          8696 => x"ea38fe18",
          8697 => x"9c1a08fe",
          8698 => x"05595680",
          8699 => x"5c757827",
          8700 => x"8d388a19",
          8701 => x"22767129",
          8702 => x"b01b0805",
          8703 => x"5d5e7bb4",
          8704 => x"1a0cb819",
          8705 => x"58848078",
          8706 => x"57558076",
          8707 => x"70810558",
          8708 => x"34ff1555",
          8709 => x"74f43874",
          8710 => x"568a1922",
          8711 => x"55757527",
          8712 => x"81803881",
          8713 => x"54751c53",
          8714 => x"77528119",
          8715 => x"3351e4b2",
          8716 => x"3f84b9c8",
          8717 => x"0880e738",
          8718 => x"811656dd",
          8719 => x"397a9818",
          8720 => x"0c840b84",
          8721 => x"b9c80c8f",
          8722 => x"3d0d0475",
          8723 => x"54b41908",
          8724 => x"53b81970",
          8725 => x"53811a33",
          8726 => x"5256e486",
          8727 => x"3f84b9c8",
          8728 => x"0880f338",
          8729 => x"84b9c808",
          8730 => x"831a34b4",
          8731 => x"1908a81a",
          8732 => x"08315574",
          8733 => x"a01a0827",
          8734 => x"fee83882",
          8735 => x"19335c7b",
          8736 => x"822e0981",
          8737 => x"06fedb38",
          8738 => x"8154b419",
          8739 => x"08a01a08",
          8740 => x"05537552",
          8741 => x"81193351",
          8742 => x"e3c83ffe",
          8743 => x"c5398a19",
          8744 => x"22557483",
          8745 => x"ffff0655",
          8746 => x"74762e09",
          8747 => x"8106a738",
          8748 => x"7c94180c",
          8749 => x"fe1d9c1a",
          8750 => x"08fe055e",
          8751 => x"56805875",
          8752 => x"7d27fd85",
          8753 => x"388a1922",
          8754 => x"767129b0",
          8755 => x"1b080598",
          8756 => x"190c5cfc",
          8757 => x"f839810b",
          8758 => x"84b9c80c",
          8759 => x"8f3d0d04",
          8760 => x"ee3d0d64",
          8761 => x"66415c84",
          8762 => x"7c085a5b",
          8763 => x"81ff7098",
          8764 => x"1e08585e",
          8765 => x"5e75802e",
          8766 => x"82d238b8",
          8767 => x"195f755a",
          8768 => x"8058b419",
          8769 => x"08762e82",
          8770 => x"d1388319",
          8771 => x"33785855",
          8772 => x"74782e09",
          8773 => x"81068194",
          8774 => x"38815475",
          8775 => x"53b81952",
          8776 => x"81193351",
          8777 => x"e1bd3f84",
          8778 => x"b9c80880",
          8779 => x"2e8538ff",
          8780 => x"5a815779",
          8781 => x"b41a0c76",
          8782 => x"5b768290",
          8783 => x"389c1c08",
          8784 => x"70335858",
          8785 => x"76802e82",
          8786 => x"81388b18",
          8787 => x"33bf0670",
          8788 => x"81ff065b",
          8789 => x"4160861d",
          8790 => x"347681e5",
          8791 => x"32703078",
          8792 => x"ae327030",
          8793 => x"72802571",
          8794 => x"80250754",
          8795 => x"45455755",
          8796 => x"74933874",
          8797 => x"7adf0643",
          8798 => x"5661882e",
          8799 => x"81bf3875",
          8800 => x"602e8186",
          8801 => x"3881ff5d",
          8802 => x"80527b51",
          8803 => x"faf63f84",
          8804 => x"b9c8085b",
          8805 => x"84b9c808",
          8806 => x"81b23898",
          8807 => x"1c085675",
          8808 => x"fedc387a",
          8809 => x"84b9c80c",
          8810 => x"943d0d04",
          8811 => x"8154b419",
          8812 => x"08537e52",
          8813 => x"81193351",
          8814 => x"e1a83f81",
          8815 => x"5784b9c8",
          8816 => x"08782e09",
          8817 => x"8106feef",
          8818 => x"3884b9c8",
          8819 => x"08831a34",
          8820 => x"b41908a8",
          8821 => x"1a083184",
          8822 => x"b9c80858",
          8823 => x"5b7aa01a",
          8824 => x"0827feb5",
          8825 => x"38821933",
          8826 => x"4160822e",
          8827 => x"098106fe",
          8828 => x"a8388154",
          8829 => x"b41908a0",
          8830 => x"1a080553",
          8831 => x"7e528119",
          8832 => x"3351e0de",
          8833 => x"3f7757fe",
          8834 => x"9039798f",
          8835 => x"2e098106",
          8836 => x"81e73876",
          8837 => x"862a8106",
          8838 => x"5b7a802e",
          8839 => x"93388d18",
          8840 => x"337781bf",
          8841 => x"0670901f",
          8842 => x"087fac05",
          8843 => x"0c595e5e",
          8844 => x"767d2eab",
          8845 => x"3881ff55",
          8846 => x"745dfecc",
          8847 => x"39815675",
          8848 => x"602e0981",
          8849 => x"06febe38",
          8850 => x"c139845b",
          8851 => x"800b981d",
          8852 => x"0c7a84b9",
          8853 => x"c80c943d",
          8854 => x"0d04775b",
          8855 => x"fddf398d",
          8856 => x"1833577d",
          8857 => x"772e0981",
          8858 => x"06cb388c",
          8859 => x"19089b19",
          8860 => x"339a1a33",
          8861 => x"71882b07",
          8862 => x"58564175",
          8863 => x"ffb73877",
          8864 => x"337081bf",
          8865 => x"068d29f3",
          8866 => x"05515a81",
          8867 => x"76585b83",
          8868 => x"e5c81733",
          8869 => x"78058111",
          8870 => x"33713371",
          8871 => x"882b0752",
          8872 => x"44567a80",
          8873 => x"2e80c538",
          8874 => x"7981fe26",
          8875 => x"ff873879",
          8876 => x"10610576",
          8877 => x"5c427562",
          8878 => x"23811a5a",
          8879 => x"8117578c",
          8880 => x"7727cc38",
          8881 => x"77337086",
          8882 => x"2a810659",
          8883 => x"5777802e",
          8884 => x"90387981",
          8885 => x"fe26fedd",
          8886 => x"38791061",
          8887 => x"05438063",
          8888 => x"23ff1d70",
          8889 => x"81ff065e",
          8890 => x"41fd9d39",
          8891 => x"7583ffff",
          8892 => x"2eca3881",
          8893 => x"ff55fec0",
          8894 => x"397ca838",
          8895 => x"7c558b57",
          8896 => x"74812a75",
          8897 => x"81802905",
          8898 => x"78708105",
          8899 => x"5a33407f",
          8900 => x"057081ff",
          8901 => x"06ff1959",
          8902 => x"565976e4",
          8903 => x"38747e2e",
          8904 => x"fd8138ff",
          8905 => x"0bac1d0c",
          8906 => x"7a84b9c8",
          8907 => x"0c943d0d",
          8908 => x"04ef3d0d",
          8909 => x"6370085c",
          8910 => x"5c80527b",
          8911 => x"51f5cf3f",
          8912 => x"84b9c808",
          8913 => x"5a84b9c8",
          8914 => x"08828038",
          8915 => x"81ff7040",
          8916 => x"5dff0bac",
          8917 => x"1d0cb81b",
          8918 => x"5e981c08",
          8919 => x"568058b4",
          8920 => x"1b08762e",
          8921 => x"82cc3883",
          8922 => x"1b337858",
          8923 => x"5574782e",
          8924 => x"09810681",
          8925 => x"df388154",
          8926 => x"7553b81b",
          8927 => x"52811b33",
          8928 => x"51dce03f",
          8929 => x"84b9c808",
          8930 => x"802e8538",
          8931 => x"ff568157",
          8932 => x"75b41c0c",
          8933 => x"765a7681",
          8934 => x"b2389c1c",
          8935 => x"08703358",
          8936 => x"5976802e",
          8937 => x"8499388b",
          8938 => x"1933bf06",
          8939 => x"7081ff06",
          8940 => x"57587786",
          8941 => x"1d347681",
          8942 => x"e52e80f2",
          8943 => x"3875832a",
          8944 => x"81065575",
          8945 => x"8f2e81ef",
          8946 => x"387480e2",
          8947 => x"38758f2e",
          8948 => x"81e5387c",
          8949 => x"aa38787d",
          8950 => x"56588b57",
          8951 => x"74812a75",
          8952 => x"81802905",
          8953 => x"78708105",
          8954 => x"5a335776",
          8955 => x"057081ff",
          8956 => x"06ff1959",
          8957 => x"565d76e4",
          8958 => x"38747f2e",
          8959 => x"80cd38ab",
          8960 => x"1c338106",
          8961 => x"5776a738",
          8962 => x"8b0ba01d",
          8963 => x"59577870",
          8964 => x"81055a33",
          8965 => x"78708105",
          8966 => x"5a337171",
          8967 => x"31ff1a5a",
          8968 => x"58424076",
          8969 => x"802e81dc",
          8970 => x"3875802e",
          8971 => x"e13881ff",
          8972 => x"5dff0bac",
          8973 => x"1d0c8052",
          8974 => x"7b51f5c8",
          8975 => x"3f84b9c8",
          8976 => x"085a84b9",
          8977 => x"c808802e",
          8978 => x"fe8f3879",
          8979 => x"84b9c80c",
          8980 => x"933d0d04",
          8981 => x"8154b41b",
          8982 => x"08537d52",
          8983 => x"811b3351",
          8984 => x"dc803f81",
          8985 => x"5784b9c8",
          8986 => x"08782e09",
          8987 => x"8106fea4",
          8988 => x"3884b9c8",
          8989 => x"08831c34",
          8990 => x"b41b08a8",
          8991 => x"1c083184",
          8992 => x"b9c80858",
          8993 => x"5978a01c",
          8994 => x"0827fdea",
          8995 => x"38821b33",
          8996 => x"5a79822e",
          8997 => x"098106fd",
          8998 => x"dd388154",
          8999 => x"b41b08a0",
          9000 => x"1c080553",
          9001 => x"7d52811b",
          9002 => x"3351dbb6",
          9003 => x"3f7757fd",
          9004 => x"c539775a",
          9005 => x"fde439ab",
          9006 => x"1c337086",
          9007 => x"2a810642",
          9008 => x"5560fef2",
          9009 => x"3876862a",
          9010 => x"81065a79",
          9011 => x"802e9338",
          9012 => x"8d193377",
          9013 => x"81bf0670",
          9014 => x"901f087f",
          9015 => x"ac050c59",
          9016 => x"5e5f767d",
          9017 => x"2eaf3881",
          9018 => x"ff55745d",
          9019 => x"80527b51",
          9020 => x"f4923f84",
          9021 => x"b9c8085a",
          9022 => x"84b9c808",
          9023 => x"802efcd9",
          9024 => x"38fec839",
          9025 => x"75802efe",
          9026 => x"c23881ff",
          9027 => x"5dff0bac",
          9028 => x"1d0cfea2",
          9029 => x"398d1933",
          9030 => x"577e772e",
          9031 => x"098106c7",
          9032 => x"388c1b08",
          9033 => x"9b1a339a",
          9034 => x"1b337188",
          9035 => x"2b075942",
          9036 => x"4076ffb3",
          9037 => x"38783370",
          9038 => x"bf068d29",
          9039 => x"f3055b55",
          9040 => x"81775956",
          9041 => x"83e5c818",
          9042 => x"33790581",
          9043 => x"11337133",
          9044 => x"71882b07",
          9045 => x"52425775",
          9046 => x"802e80ed",
          9047 => x"387981fe",
          9048 => x"26ff8438",
          9049 => x"765181a1",
          9050 => x"8a3f84b9",
          9051 => x"c8087a10",
          9052 => x"61057022",
          9053 => x"5343811b",
          9054 => x"5b5681a0",
          9055 => x"f63f7584",
          9056 => x"b9c8082e",
          9057 => x"098106fe",
          9058 => x"de387656",
          9059 => x"8118588c",
          9060 => x"7827ffb0",
          9061 => x"38783370",
          9062 => x"862a8106",
          9063 => x"56597580",
          9064 => x"2e923874",
          9065 => x"802e8d38",
          9066 => x"79106005",
          9067 => x"70224141",
          9068 => x"7ffeb438",
          9069 => x"ff1d7081",
          9070 => x"ff065e5a",
          9071 => x"feae3984",
          9072 => x"0b84b9c8",
          9073 => x"0c933d0d",
          9074 => x"047683ff",
          9075 => x"ff2effbc",
          9076 => x"3881ff55",
          9077 => x"fe9439ea",
          9078 => x"3d0d6870",
          9079 => x"0870ab13",
          9080 => x"3381a006",
          9081 => x"585a5d5e",
          9082 => x"86567485",
          9083 => x"b538748c",
          9084 => x"1d087022",
          9085 => x"57575d74",
          9086 => x"802e8e38",
          9087 => x"811d7010",
          9088 => x"17702251",
          9089 => x"565d74f4",
          9090 => x"38953da0",
          9091 => x"1f5b408c",
          9092 => x"607b5858",
          9093 => x"55757081",
          9094 => x"05573377",
          9095 => x"70810559",
          9096 => x"34ff1555",
          9097 => x"74ef3802",
          9098 => x"80db0533",
          9099 => x"70810658",
          9100 => x"5676802e",
          9101 => x"82aa3880",
          9102 => x"c00bab1f",
          9103 => x"34810b94",
          9104 => x"3d405b8c",
          9105 => x"1c087b58",
          9106 => x"598b7a61",
          9107 => x"5a575577",
          9108 => x"70810559",
          9109 => x"33767081",
          9110 => x"055834ff",
          9111 => x"155574ef",
          9112 => x"38857b27",
          9113 => x"80c2387a",
          9114 => x"79225657",
          9115 => x"74802eb8",
          9116 => x"3874821a",
          9117 => x"5a568f58",
          9118 => x"75810677",
          9119 => x"10077681",
          9120 => x"2a7083ff",
          9121 => x"ff067290",
          9122 => x"2a810644",
          9123 => x"58565760",
          9124 => x"802e8738",
          9125 => x"7684a0a1",
          9126 => x"3257ff18",
          9127 => x"58778025",
          9128 => x"d7387822",
          9129 => x"5574ca38",
          9130 => x"87028405",
          9131 => x"80cf0557",
          9132 => x"5876b007",
          9133 => x"bf0655b9",
          9134 => x"75278438",
          9135 => x"87155574",
          9136 => x"7634ff16",
          9137 => x"ff197884",
          9138 => x"2a595956",
          9139 => x"76e33877",
          9140 => x"1f5980fe",
          9141 => x"7934767a",
          9142 => x"58568078",
          9143 => x"27a03879",
          9144 => x"335574a0",
          9145 => x"2e983881",
          9146 => x"16567578",
          9147 => x"2788a238",
          9148 => x"751a7033",
          9149 => x"565774a0",
          9150 => x"2e098106",
          9151 => x"ea388116",
          9152 => x"56a05577",
          9153 => x"87268e38",
          9154 => x"983d7805",
          9155 => x"ec058119",
          9156 => x"71335759",
          9157 => x"41747734",
          9158 => x"87762787",
          9159 => x"f4387d51",
          9160 => x"f88f3f84",
          9161 => x"b9c8088b",
          9162 => x"38811b5b",
          9163 => x"80e37b27",
          9164 => x"fe913887",
          9165 => x"567a80e4",
          9166 => x"2e82e738",
          9167 => x"84b9c808",
          9168 => x"5684b9c8",
          9169 => x"08842e09",
          9170 => x"810682d6",
          9171 => x"380280db",
          9172 => x"0533ab1f",
          9173 => x"347d0802",
          9174 => x"840580db",
          9175 => x"05335758",
          9176 => x"75812a81",
          9177 => x"065f815b",
          9178 => x"7e802e90",
          9179 => x"388d528c",
          9180 => x"1d51fe8a",
          9181 => x"b03f84b9",
          9182 => x"c8081b5b",
          9183 => x"80527d51",
          9184 => x"ed8c3f84",
          9185 => x"b9c80856",
          9186 => x"84b9c808",
          9187 => x"81823884",
          9188 => x"b9c808b8",
          9189 => x"195e5998",
          9190 => x"1e085680",
          9191 => x"57b41808",
          9192 => x"762e85f3",
          9193 => x"38831833",
          9194 => x"407f772e",
          9195 => x"09810682",
          9196 => x"a3388154",
          9197 => x"7553b818",
          9198 => x"52811833",
          9199 => x"51d4a43f",
          9200 => x"84b9c808",
          9201 => x"802e8538",
          9202 => x"ff568157",
          9203 => x"75b4190c",
          9204 => x"765676bc",
          9205 => x"389c1e08",
          9206 => x"70335642",
          9207 => x"7481e52e",
          9208 => x"81c93874",
          9209 => x"30708025",
          9210 => x"7807565f",
          9211 => x"74802e81",
          9212 => x"c9388119",
          9213 => x"59787b2e",
          9214 => x"86893881",
          9215 => x"527d51ee",
          9216 => x"833f84b9",
          9217 => x"c8085684",
          9218 => x"b9c80880",
          9219 => x"2eff8838",
          9220 => x"87587584",
          9221 => x"2e818938",
          9222 => x"75587581",
          9223 => x"8338ff1b",
          9224 => x"407f81f3",
          9225 => x"38981e08",
          9226 => x"57b41c08",
          9227 => x"772eaf38",
          9228 => x"831c3378",
          9229 => x"57407f84",
          9230 => x"82388154",
          9231 => x"7653b81c",
          9232 => x"52811c33",
          9233 => x"51d39c3f",
          9234 => x"84b9c808",
          9235 => x"802e8538",
          9236 => x"ff578156",
          9237 => x"76b41d0c",
          9238 => x"75587580",
          9239 => x"c338a00b",
          9240 => x"9c1f0857",
          9241 => x"55807670",
          9242 => x"81055834",
          9243 => x"ff155574",
          9244 => x"f4388b0b",
          9245 => x"9c1f087b",
          9246 => x"58585575",
          9247 => x"70810557",
          9248 => x"33777081",
          9249 => x"055934ff",
          9250 => x"155574ef",
          9251 => x"389c1e08",
          9252 => x"ab1f3398",
          9253 => x"065e5a7c",
          9254 => x"8c1b3481",
          9255 => x"0b831d34",
          9256 => x"77567584",
          9257 => x"b9c80c98",
          9258 => x"3d0d0481",
          9259 => x"75307080",
          9260 => x"25720757",
          9261 => x"405774fe",
          9262 => x"b9387459",
          9263 => x"81527d51",
          9264 => x"ecc23f84",
          9265 => x"b9c80856",
          9266 => x"84b9c808",
          9267 => x"802efdc7",
          9268 => x"38febd39",
          9269 => x"8154b418",
          9270 => x"08537c52",
          9271 => x"81183351",
          9272 => x"d3803f84",
          9273 => x"b9c80877",
          9274 => x"2e098106",
          9275 => x"83bf3884",
          9276 => x"b9c80883",
          9277 => x"1934b418",
          9278 => x"08a81908",
          9279 => x"315574a0",
          9280 => x"1908278b",
          9281 => x"38821833",
          9282 => x"4160822e",
          9283 => x"84ac3884",
          9284 => x"b9c80857",
          9285 => x"fd9c397f",
          9286 => x"852b901f",
          9287 => x"08713153",
          9288 => x"587d51e9",
          9289 => x"e93f84b9",
          9290 => x"c8085884",
          9291 => x"b9c808fe",
          9292 => x"ef387984",
          9293 => x"b9c80856",
          9294 => x"588b5774",
          9295 => x"812a7581",
          9296 => x"80290578",
          9297 => x"7081055a",
          9298 => x"33577605",
          9299 => x"7081ff06",
          9300 => x"ff195956",
          9301 => x"5d76e438",
          9302 => x"7481ff06",
          9303 => x"b81d4341",
          9304 => x"981e0857",
          9305 => x"8056b41c",
          9306 => x"08772eb2",
          9307 => x"38831c33",
          9308 => x"5b7a762e",
          9309 => x"09810682",
          9310 => x"c9388154",
          9311 => x"7653b81c",
          9312 => x"52811c33",
          9313 => x"51d0dc3f",
          9314 => x"84b9c808",
          9315 => x"802e8538",
          9316 => x"ff578156",
          9317 => x"76b41d0c",
          9318 => x"755875fe",
          9319 => x"83388c1c",
          9320 => x"089c1f08",
          9321 => x"6181ff06",
          9322 => x"5f5c5f60",
          9323 => x"8d1c348f",
          9324 => x"0b8b1c34",
          9325 => x"758c1c34",
          9326 => x"759a1c34",
          9327 => x"759b1c34",
          9328 => x"7c8d29f3",
          9329 => x"0576775a",
          9330 => x"58597683",
          9331 => x"ffff2e8b",
          9332 => x"3878101f",
          9333 => x"7022811b",
          9334 => x"5b585683",
          9335 => x"e5c81833",
          9336 => x"7b055576",
          9337 => x"75708105",
          9338 => x"57347688",
          9339 => x"2a567575",
          9340 => x"34768538",
          9341 => x"83ffff57",
          9342 => x"8118588c",
          9343 => x"7827cb38",
          9344 => x"7683ffff",
          9345 => x"2e81b338",
          9346 => x"78101f70",
          9347 => x"22585876",
          9348 => x"802e81a6",
          9349 => x"387c7b34",
          9350 => x"810b831d",
          9351 => x"3480527d",
          9352 => x"51e9e13f",
          9353 => x"84b9c808",
          9354 => x"5884b9c8",
          9355 => x"08fcf138",
          9356 => x"7fff0540",
          9357 => x"7ffea938",
          9358 => x"fbeb3981",
          9359 => x"54b41c08",
          9360 => x"53b81c70",
          9361 => x"53811d33",
          9362 => x"5259d096",
          9363 => x"3f815684",
          9364 => x"b9c808fc",
          9365 => x"833884b9",
          9366 => x"c808831d",
          9367 => x"34b41c08",
          9368 => x"a81d0831",
          9369 => x"84b9c808",
          9370 => x"574160a0",
          9371 => x"1d0827fb",
          9372 => x"c938821c",
          9373 => x"33426182",
          9374 => x"2e098106",
          9375 => x"fbbc3881",
          9376 => x"54b41c08",
          9377 => x"a01d0805",
          9378 => x"53785281",
          9379 => x"1c3351cf",
          9380 => x"d13f7756",
          9381 => x"fba43976",
          9382 => x"9c1f0870",
          9383 => x"33574356",
          9384 => x"7481e52e",
          9385 => x"098106fa",
          9386 => x"ba38fbff",
          9387 => x"39817057",
          9388 => x"5776802e",
          9389 => x"fa9f38fa",
          9390 => x"d7397c80",
          9391 => x"c0075dfe",
          9392 => x"d4398154",
          9393 => x"b41c0853",
          9394 => x"6152811c",
          9395 => x"3351cf92",
          9396 => x"3f84b9c8",
          9397 => x"08762e09",
          9398 => x"8106bc38",
          9399 => x"84b9c808",
          9400 => x"831d34b4",
          9401 => x"1c08a81d",
          9402 => x"08315574",
          9403 => x"a01d0827",
          9404 => x"8a38821c",
          9405 => x"335f7e82",
          9406 => x"2eaa3884",
          9407 => x"b9c80856",
          9408 => x"fcf83975",
          9409 => x"ff1c4158",
          9410 => x"7f802efa",
          9411 => x"9838fc87",
          9412 => x"39751a57",
          9413 => x"f7e83981",
          9414 => x"70595675",
          9415 => x"802efcfe",
          9416 => x"38fafd39",
          9417 => x"8154b41c",
          9418 => x"08a01d08",
          9419 => x"05536152",
          9420 => x"811c3351",
          9421 => x"ceac3ffc",
          9422 => x"c1398154",
          9423 => x"b41808a0",
          9424 => x"19080553",
          9425 => x"7c528118",
          9426 => x"3351ce96",
          9427 => x"3ff8e339",
          9428 => x"f33d0d7f",
          9429 => x"61710840",
          9430 => x"5e5c800b",
          9431 => x"961e3498",
          9432 => x"1c08802e",
          9433 => x"82b538ac",
          9434 => x"1c08ff2e",
          9435 => x"80d93880",
          9436 => x"7071608c",
          9437 => x"05087022",
          9438 => x"57585b5c",
          9439 => x"5872782e",
          9440 => x"bc387754",
          9441 => x"74147022",
          9442 => x"811b5b55",
          9443 => x"567a8295",
          9444 => x"3880d080",
          9445 => x"147083ff",
          9446 => x"ff06585a",
          9447 => x"768fff26",
          9448 => x"82833873",
          9449 => x"791a7611",
          9450 => x"70225d58",
          9451 => x"555b79d4",
          9452 => x"387a3070",
          9453 => x"80257030",
          9454 => x"7a065a5c",
          9455 => x"5e7c1894",
          9456 => x"0557800b",
          9457 => x"82183480",
          9458 => x"70891f59",
          9459 => x"57589c1c",
          9460 => x"08167033",
          9461 => x"81185856",
          9462 => x"5374a02e",
          9463 => x"b2387485",
          9464 => x"2e81bc38",
          9465 => x"75893270",
          9466 => x"30707207",
          9467 => x"8025555b",
          9468 => x"54778b26",
          9469 => x"90387280",
          9470 => x"2e8b38ae",
          9471 => x"77708105",
          9472 => x"59348118",
          9473 => x"58747770",
          9474 => x"81055934",
          9475 => x"8118588a",
          9476 => x"7627ffba",
          9477 => x"387c1888",
          9478 => x"0555800b",
          9479 => x"81163496",
          9480 => x"1d335372",
          9481 => x"a5387781",
          9482 => x"f338bf0b",
          9483 => x"961e3481",
          9484 => x"577c1794",
          9485 => x"0556800b",
          9486 => x"8217349c",
          9487 => x"1c088c11",
          9488 => x"33555373",
          9489 => x"89387389",
          9490 => x"1e349c1c",
          9491 => x"08538b13",
          9492 => x"33881e34",
          9493 => x"9c1c089c",
          9494 => x"11831133",
          9495 => x"82123371",
          9496 => x"902b7188",
          9497 => x"2b078114",
          9498 => x"33707207",
          9499 => x"882b7533",
          9500 => x"7107640c",
          9501 => x"59971633",
          9502 => x"96173371",
          9503 => x"882b075f",
          9504 => x"415b405a",
          9505 => x"565b5577",
          9506 => x"861e2399",
          9507 => x"15339816",
          9508 => x"3371882b",
          9509 => x"075d547b",
          9510 => x"841e238f",
          9511 => x"3d0d0481",
          9512 => x"e555fec0",
          9513 => x"39771d96",
          9514 => x"1181ff7a",
          9515 => x"31585b57",
          9516 => x"83b5527a",
          9517 => x"902b7407",
          9518 => x"51819189",
          9519 => x"3f84b9c8",
          9520 => x"0883ffff",
          9521 => x"065581ff",
          9522 => x"7527ad38",
          9523 => x"81762781",
          9524 => x"b3387488",
          9525 => x"2a54737a",
          9526 => x"34749718",
          9527 => x"34827805",
          9528 => x"58800b8c",
          9529 => x"1f08565b",
          9530 => x"78197511",
          9531 => x"70225c57",
          9532 => x"5479fd90",
          9533 => x"38fdba39",
          9534 => x"74307630",
          9535 => x"70780780",
          9536 => x"25728025",
          9537 => x"07585557",
          9538 => x"7580f938",
          9539 => x"747a3481",
          9540 => x"78055880",
          9541 => x"0b8c1f08",
          9542 => x"565bcd39",
          9543 => x"7273891f",
          9544 => x"335a5757",
          9545 => x"77802efe",
          9546 => x"88387c96",
          9547 => x"1e7e5759",
          9548 => x"54891433",
          9549 => x"ffbf115a",
          9550 => x"54789926",
          9551 => x"a4389c1c",
          9552 => x"088c1133",
          9553 => x"545b8876",
          9554 => x"27b43872",
          9555 => x"842a5372",
          9556 => x"81065e7d",
          9557 => x"802e8a38",
          9558 => x"a0147083",
          9559 => x"ffff0655",
          9560 => x"53737870",
          9561 => x"81055a34",
          9562 => x"81168116",
          9563 => x"81197189",
          9564 => x"13335e57",
          9565 => x"59565679",
          9566 => x"ffb738fd",
          9567 => x"b4397283",
          9568 => x"2a53cc39",
          9569 => x"807b3070",
          9570 => x"80257030",
          9571 => x"7306535d",
          9572 => x"5f58fca9",
          9573 => x"39ef3d0d",
          9574 => x"63700870",
          9575 => x"42575c80",
          9576 => x"65703357",
          9577 => x"555374af",
          9578 => x"2e833881",
          9579 => x"537480dc",
          9580 => x"2e81df38",
          9581 => x"72802e81",
          9582 => x"d9389816",
          9583 => x"08881d0c",
          9584 => x"7333963d",
          9585 => x"943d4142",
          9586 => x"559f7527",
          9587 => x"82a73873",
          9588 => x"428c1608",
          9589 => x"58805761",
          9590 => x"70708105",
          9591 => x"52335553",
          9592 => x"7381df38",
          9593 => x"727f0c73",
          9594 => x"ff2e81ec",
          9595 => x"3883ffff",
          9596 => x"74278b38",
          9597 => x"76101856",
          9598 => x"80762381",
          9599 => x"17577383",
          9600 => x"ffff0670",
          9601 => x"af327030",
          9602 => x"9f732771",
          9603 => x"80250757",
          9604 => x"5b5b5573",
          9605 => x"82903874",
          9606 => x"80dc2e82",
          9607 => x"89387480",
          9608 => x"ff26b238",
          9609 => x"83e4e40b",
          9610 => x"83e4e433",
          9611 => x"7081ff06",
          9612 => x"56545673",
          9613 => x"802e81ab",
          9614 => x"3873752e",
          9615 => x"8f388116",
          9616 => x"70337081",
          9617 => x"ff065654",
          9618 => x"5673ee38",
          9619 => x"7281ff06",
          9620 => x"5b7a8184",
          9621 => x"387681fe",
          9622 => x"2680fd38",
          9623 => x"7610185d",
          9624 => x"747d2381",
          9625 => x"17627070",
          9626 => x"81055233",
          9627 => x"56545773",
          9628 => x"802efef0",
          9629 => x"3880cb39",
          9630 => x"817380dc",
          9631 => x"32703070",
          9632 => x"80257307",
          9633 => x"51555855",
          9634 => x"72802ea1",
          9635 => x"38811470",
          9636 => x"46548074",
          9637 => x"33545572",
          9638 => x"af2edd38",
          9639 => x"7280dc32",
          9640 => x"70307080",
          9641 => x"25770751",
          9642 => x"545772e1",
          9643 => x"3872881d",
          9644 => x"0c733396",
          9645 => x"3d943d41",
          9646 => x"4255749f",
          9647 => x"26fe9038",
          9648 => x"b43983b5",
          9649 => x"52735181",
          9650 => x"8de73f84",
          9651 => x"b9c80883",
          9652 => x"ffff0654",
          9653 => x"73fe8d38",
          9654 => x"86547384",
          9655 => x"b9c80c93",
          9656 => x"3d0d0483",
          9657 => x"e4e43370",
          9658 => x"81ff065c",
          9659 => x"537a802e",
          9660 => x"fee338e4",
          9661 => x"39ff800b",
          9662 => x"ab1d3480",
          9663 => x"527b51de",
          9664 => x"8d3f84b9",
          9665 => x"c80884b9",
          9666 => x"c80c933d",
          9667 => x"0d048173",
          9668 => x"80dc3270",
          9669 => x"30708025",
          9670 => x"73074155",
          9671 => x"5a567d80",
          9672 => x"2ea13881",
          9673 => x"14428062",
          9674 => x"70335555",
          9675 => x"5672af2e",
          9676 => x"dd387280",
          9677 => x"dc327030",
          9678 => x"70802578",
          9679 => x"07405459",
          9680 => x"7de13873",
          9681 => x"610c9f75",
          9682 => x"27822b5a",
          9683 => x"76812e84",
          9684 => x"f8387682",
          9685 => x"2e83d138",
          9686 => x"76175976",
          9687 => x"802ea738",
          9688 => x"76177811",
          9689 => x"fe057022",
          9690 => x"70a03270",
          9691 => x"30709f2a",
          9692 => x"5242565f",
          9693 => x"56597cae",
          9694 => x"2e843872",
          9695 => x"8938ff17",
          9696 => x"5776dd38",
          9697 => x"76597719",
          9698 => x"56807623",
          9699 => x"76802efe",
          9700 => x"c7388078",
          9701 => x"227083ff",
          9702 => x"ff067258",
          9703 => x"5d55567a",
          9704 => x"a02e82e6",
          9705 => x"387383ff",
          9706 => x"ff065372",
          9707 => x"ae2e82f1",
          9708 => x"3876802e",
          9709 => x"aa387719",
          9710 => x"fe057022",
          9711 => x"5a5478ae",
          9712 => x"2e9d3876",
          9713 => x"1018fe05",
          9714 => x"54ff1757",
          9715 => x"76802e8f",
          9716 => x"38fe1470",
          9717 => x"225e547c",
          9718 => x"ae2e0981",
          9719 => x"06eb388b",
          9720 => x"0ba01d55",
          9721 => x"53a07470",
          9722 => x"81055634",
          9723 => x"ff135372",
          9724 => x"f4387273",
          9725 => x"5c5e8878",
          9726 => x"16702281",
          9727 => x"19595754",
          9728 => x"5d74802e",
          9729 => x"80ed3874",
          9730 => x"a02e83d0",
          9731 => x"3874ae32",
          9732 => x"70307080",
          9733 => x"25555a54",
          9734 => x"75772e85",
          9735 => x"ce387283",
          9736 => x"bb387259",
          9737 => x"7c7b2683",
          9738 => x"38815975",
          9739 => x"77327030",
          9740 => x"70720780",
          9741 => x"25707c07",
          9742 => x"51515454",
          9743 => x"72802e83",
          9744 => x"e0387c8b",
          9745 => x"2e868338",
          9746 => x"75772e8a",
          9747 => x"38798307",
          9748 => x"5a757726",
          9749 => x"9e387656",
          9750 => x"885b8b7e",
          9751 => x"822b81fc",
          9752 => x"06771857",
          9753 => x"5f5d7715",
          9754 => x"70228118",
          9755 => x"58565374",
          9756 => x"ff9538a0",
          9757 => x"1c335776",
          9758 => x"81e52e83",
          9759 => x"84387c88",
          9760 => x"2e82e338",
          9761 => x"7d8c0658",
          9762 => x"778c2e82",
          9763 => x"ed387d83",
          9764 => x"06557483",
          9765 => x"2e82e338",
          9766 => x"79812a81",
          9767 => x"0656759d",
          9768 => x"387d8106",
          9769 => x"5d7c802e",
          9770 => x"85387990",
          9771 => x"075a7d82",
          9772 => x"2a81065e",
          9773 => x"7d802e85",
          9774 => x"38798807",
          9775 => x"5a79ab1d",
          9776 => x"347b51e4",
          9777 => x"ec3f84b9",
          9778 => x"c808ab1d",
          9779 => x"33565484",
          9780 => x"b9c80880",
          9781 => x"2e81ac38",
          9782 => x"84b9c808",
          9783 => x"842e0981",
          9784 => x"06fbf738",
          9785 => x"74852a81",
          9786 => x"065a7980",
          9787 => x"2e84f038",
          9788 => x"74822a81",
          9789 => x"06597882",
          9790 => x"98387b08",
          9791 => x"65555673",
          9792 => x"428c1608",
          9793 => x"588057f9",
          9794 => x"ce398116",
          9795 => x"70117911",
          9796 => x"70224040",
          9797 => x"56567ca0",
          9798 => x"2ef03875",
          9799 => x"802efd85",
          9800 => x"38798307",
          9801 => x"5afd8a39",
          9802 => x"82182256",
          9803 => x"75ae2e09",
          9804 => x"8106fcac",
          9805 => x"38772254",
          9806 => x"73ae2e09",
          9807 => x"8106fca0",
          9808 => x"38761018",
          9809 => x"5b807b23",
          9810 => x"800ba01d",
          9811 => x"5653ae54",
          9812 => x"76732683",
          9813 => x"38a05473",
          9814 => x"75708105",
          9815 => x"57348113",
          9816 => x"538a7327",
          9817 => x"e93879a0",
          9818 => x"075877ab",
          9819 => x"1d347b51",
          9820 => x"e3bf3f84",
          9821 => x"b9c808ab",
          9822 => x"1d335654",
          9823 => x"84b9c808",
          9824 => x"fed63874",
          9825 => x"822a8106",
          9826 => x"5877face",
          9827 => x"38861c33",
          9828 => x"70842a81",
          9829 => x"06565d74",
          9830 => x"802e83cd",
          9831 => x"38901c08",
          9832 => x"83ff0660",
          9833 => x"0580d311",
          9834 => x"3380d212",
          9835 => x"3371882b",
          9836 => x"07623341",
          9837 => x"5754547d",
          9838 => x"832e82d8",
          9839 => x"3874881d",
          9840 => x"0c7b0865",
          9841 => x"5556feb7",
          9842 => x"39772255",
          9843 => x"74ae2efe",
          9844 => x"f0387617",
          9845 => x"5976fb88",
          9846 => x"38fbab39",
          9847 => x"79830776",
          9848 => x"17565afd",
          9849 => x"81397d82",
          9850 => x"2b81fc06",
          9851 => x"708c0659",
          9852 => x"5e778c2e",
          9853 => x"098106fd",
          9854 => x"95387982",
          9855 => x"075afd98",
          9856 => x"39850ba0",
          9857 => x"1d347c88",
          9858 => x"2e098106",
          9859 => x"fcf638d6",
          9860 => x"39ff800b",
          9861 => x"ab1d3480",
          9862 => x"0b84b9c8",
          9863 => x"0c933d0d",
          9864 => x"047480ff",
          9865 => x"269d3881",
          9866 => x"ff752780",
          9867 => x"c938ff1d",
          9868 => x"59787b26",
          9869 => x"81f73879",
          9870 => x"83077d77",
          9871 => x"18575c5a",
          9872 => x"fca43979",
          9873 => x"82075a83",
          9874 => x"b5527451",
          9875 => x"8185f63f",
          9876 => x"84b9c808",
          9877 => x"83ffff06",
          9878 => x"70872a81",
          9879 => x"065a5578",
          9880 => x"802ec438",
          9881 => x"7480ff06",
          9882 => x"83e5d811",
          9883 => x"33565474",
          9884 => x"81ff26ff",
          9885 => x"b9387480",
          9886 => x"2e818538",
          9887 => x"83e4f00b",
          9888 => x"83e4f033",
          9889 => x"7081ff06",
          9890 => x"56545973",
          9891 => x"802e80e0",
          9892 => x"3873752e",
          9893 => x"8f388119",
          9894 => x"70337081",
          9895 => x"ff065654",
          9896 => x"5973ee38",
          9897 => x"7281ff06",
          9898 => x"597880d4",
          9899 => x"38ffbf15",
          9900 => x"54739926",
          9901 => x"8a387d82",
          9902 => x"077081ff",
          9903 => x"065f53ff",
          9904 => x"9f155978",
          9905 => x"99269338",
          9906 => x"7d810770",
          9907 => x"81ff06e0",
          9908 => x"177083ff",
          9909 => x"ff065856",
          9910 => x"5f537b1b",
          9911 => x"a0055974",
          9912 => x"7934811b",
          9913 => x"5b751655",
          9914 => x"fafc3980",
          9915 => x"53fab339",
          9916 => x"83e4f033",
          9917 => x"7081ff06",
          9918 => x"5a537880",
          9919 => x"2effae38",
          9920 => x"80df7a83",
          9921 => x"077d1da0",
          9922 => x"055b5b55",
          9923 => x"74793481",
          9924 => x"1b5bd239",
          9925 => x"80cd1433",
          9926 => x"80cc1533",
          9927 => x"71982b71",
          9928 => x"902b0777",
          9929 => x"07881f0c",
          9930 => x"5a57fd95",
          9931 => x"397b1ba0",
          9932 => x"0575882a",
          9933 => x"54547274",
          9934 => x"34811b7c",
          9935 => x"11a0055a",
          9936 => x"5b747934",
          9937 => x"811b5bff",
          9938 => x"9c397983",
          9939 => x"07a01d33",
          9940 => x"585a7681",
          9941 => x"e52e0981",
          9942 => x"06faa338",
          9943 => x"fda33974",
          9944 => x"822a8106",
          9945 => x"5c7bf6f2",
          9946 => x"38850b84",
          9947 => x"b9c80c93",
          9948 => x"3d0d04eb",
          9949 => x"3d0d6769",
          9950 => x"02880580",
          9951 => x"e7053342",
          9952 => x"425e8061",
          9953 => x"0cff7e08",
          9954 => x"70595b42",
          9955 => x"79802e85",
          9956 => x"d7387970",
          9957 => x"81055b33",
          9958 => x"709f2656",
          9959 => x"5675ba2e",
          9960 => x"85d03874",
          9961 => x"ed3875ba",
          9962 => x"2e85c738",
          9963 => x"84d1a433",
          9964 => x"56807624",
          9965 => x"85b23875",
          9966 => x"101084d1",
          9967 => x"90057008",
          9968 => x"585a8c58",
          9969 => x"76802e85",
          9970 => x"96387661",
          9971 => x"0c7f81fe",
          9972 => x"0677335d",
          9973 => x"597b802e",
          9974 => x"9b388117",
          9975 => x"3351ffbb",
          9976 => x"b03f84b9",
          9977 => x"c80881ff",
          9978 => x"06708106",
          9979 => x"5e587c80",
          9980 => x"2e869638",
          9981 => x"80773475",
          9982 => x"165d84b9",
          9983 => x"bc1d3381",
          9984 => x"18348152",
          9985 => x"81173351",
          9986 => x"ffbba43f",
          9987 => x"84b9c808",
          9988 => x"81ff0670",
          9989 => x"81064156",
          9990 => x"83587f84",
          9991 => x"c2387880",
          9992 => x"2e8d3875",
          9993 => x"822a8106",
          9994 => x"418a5860",
          9995 => x"84b13880",
          9996 => x"5b7a8318",
          9997 => x"34ff0bb4",
          9998 => x"180c7a7b",
          9999 => x"5a558154",
         10000 => x"7a53b817",
         10001 => x"70538118",
         10002 => x"335258ff",
         10003 => x"bb953f84",
         10004 => x"b9c8087b",
         10005 => x"2e8538ff",
         10006 => x"55815974",
         10007 => x"b4180c84",
         10008 => x"56789938",
         10009 => x"84b71733",
         10010 => x"84b61833",
         10011 => x"71882b07",
         10012 => x"56568356",
         10013 => x"7482d4d5",
         10014 => x"2e85a538",
         10015 => x"7581268b",
         10016 => x"3884b9bd",
         10017 => x"1d334261",
         10018 => x"85bf3881",
         10019 => x"5875842e",
         10020 => x"83cd388d",
         10021 => x"58758126",
         10022 => x"83c53880",
         10023 => x"c4173380",
         10024 => x"c3183371",
         10025 => x"882b075e",
         10026 => x"597c8480",
         10027 => x"2e098106",
         10028 => x"83ad3880",
         10029 => x"cf173380",
         10030 => x"ce183371",
         10031 => x"882b0757",
         10032 => x"5a75a438",
         10033 => x"80dc1783",
         10034 => x"11338212",
         10035 => x"3371902b",
         10036 => x"71882b07",
         10037 => x"81143370",
         10038 => x"7207882b",
         10039 => x"75337107",
         10040 => x"565a4543",
         10041 => x"5e5f5675",
         10042 => x"a0180c80",
         10043 => x"c8173382",
         10044 => x"183480c8",
         10045 => x"1733ff11",
         10046 => x"7081ff06",
         10047 => x"5f40598d",
         10048 => x"587c8126",
         10049 => x"82d93878",
         10050 => x"81ff0676",
         10051 => x"712980c5",
         10052 => x"19335a5f",
         10053 => x"5a778a18",
         10054 => x"23775977",
         10055 => x"802e87c4",
         10056 => x"38ff1878",
         10057 => x"06426187",
         10058 => x"bb3880ca",
         10059 => x"173380c9",
         10060 => x"18337188",
         10061 => x"2b075640",
         10062 => x"74881823",
         10063 => x"74758f06",
         10064 => x"5e5a8d58",
         10065 => x"7c829838",
         10066 => x"80cc1733",
         10067 => x"80cb1833",
         10068 => x"71882b07",
         10069 => x"565c74a4",
         10070 => x"3880d817",
         10071 => x"83113382",
         10072 => x"12337190",
         10073 => x"2b71882b",
         10074 => x"07811433",
         10075 => x"70720788",
         10076 => x"2b753371",
         10077 => x"0753445a",
         10078 => x"58424242",
         10079 => x"80c71733",
         10080 => x"80c61833",
         10081 => x"71882b07",
         10082 => x"5d588d58",
         10083 => x"7b802e81",
         10084 => x"ce387d1c",
         10085 => x"7a842a05",
         10086 => x"5a797526",
         10087 => x"81c13878",
         10088 => x"52747a31",
         10089 => x"51fdedfd",
         10090 => x"3f84b9c8",
         10091 => x"085684b9",
         10092 => x"c808802e",
         10093 => x"81a93884",
         10094 => x"b9c80880",
         10095 => x"fffffff5",
         10096 => x"26833883",
         10097 => x"5d7583ff",
         10098 => x"f5268338",
         10099 => x"825d759f",
         10100 => x"f52685eb",
         10101 => x"38815d82",
         10102 => x"16709c19",
         10103 => x"0c7ba419",
         10104 => x"0c7b1d70",
         10105 => x"a81a0c7b",
         10106 => x"1db01a0c",
         10107 => x"57597c83",
         10108 => x"2e8a8738",
         10109 => x"8817225c",
         10110 => x"8d587b80",
         10111 => x"2e80e038",
         10112 => x"7d16ac18",
         10113 => x"0c781955",
         10114 => x"7c822e8d",
         10115 => x"38781019",
         10116 => x"70812a7a",
         10117 => x"81060556",
         10118 => x"5a83ff15",
         10119 => x"892a598d",
         10120 => x"5878a018",
         10121 => x"0826b838",
         10122 => x"ff0b9418",
         10123 => x"0cff0b90",
         10124 => x"180cff80",
         10125 => x"0b841834",
         10126 => x"7c832e86",
         10127 => x"96387c77",
         10128 => x"3484d1a0",
         10129 => x"2281055d",
         10130 => x"7c84d1a0",
         10131 => x"237c8618",
         10132 => x"2384d1a8",
         10133 => x"0b8c180c",
         10134 => x"800b9818",
         10135 => x"0c805877",
         10136 => x"84b9c80c",
         10137 => x"973d0d04",
         10138 => x"8b0b84b9",
         10139 => x"c80c973d",
         10140 => x"0d047633",
         10141 => x"d0117081",
         10142 => x"ff065757",
         10143 => x"58748926",
         10144 => x"91388217",
         10145 => x"7881ff06",
         10146 => x"d0055d59",
         10147 => x"787a2e87",
         10148 => x"fe38807e",
         10149 => x"0883e5b8",
         10150 => x"5f405c7c",
         10151 => x"087f5a5b",
         10152 => x"7a708105",
         10153 => x"5c337970",
         10154 => x"81055b33",
         10155 => x"ff9f125a",
         10156 => x"58567799",
         10157 => x"268938e0",
         10158 => x"167081ff",
         10159 => x"065755ff",
         10160 => x"9f175877",
         10161 => x"99268938",
         10162 => x"e0177081",
         10163 => x"ff065855",
         10164 => x"7530709f",
         10165 => x"2a595575",
         10166 => x"772e0981",
         10167 => x"06853877",
         10168 => x"ffbe3878",
         10169 => x"7a327030",
         10170 => x"7072079f",
         10171 => x"2a7a075d",
         10172 => x"58557a80",
         10173 => x"2e879838",
         10174 => x"811c841e",
         10175 => x"5e5c837c",
         10176 => x"25ff9838",
         10177 => x"6156f9a9",
         10178 => x"3978802e",
         10179 => x"fecf3877",
         10180 => x"822a8106",
         10181 => x"5e8a587d",
         10182 => x"fec53880",
         10183 => x"58fec039",
         10184 => x"7a783357",
         10185 => x"597581e9",
         10186 => x"2e098106",
         10187 => x"83388159",
         10188 => x"7581eb32",
         10189 => x"70307080",
         10190 => x"257b075a",
         10191 => x"5b5c7783",
         10192 => x"ad387581",
         10193 => x"e82e83a6",
         10194 => x"38933d77",
         10195 => x"575a8359",
         10196 => x"83fa1633",
         10197 => x"70595b7a",
         10198 => x"802ea538",
         10199 => x"84811633",
         10200 => x"84801733",
         10201 => x"71902b71",
         10202 => x"882b0783",
         10203 => x"ff193370",
         10204 => x"7207882b",
         10205 => x"83fe1b33",
         10206 => x"71075259",
         10207 => x"5b404040",
         10208 => x"777a7084",
         10209 => x"055c0cff",
         10210 => x"19901757",
         10211 => x"59788025",
         10212 => x"ffbe3884",
         10213 => x"b9bd1d33",
         10214 => x"7030709f",
         10215 => x"2a727131",
         10216 => x"9b3d7110",
         10217 => x"1005f005",
         10218 => x"84b61c44",
         10219 => x"5d52435b",
         10220 => x"4278085b",
         10221 => x"83567a80",
         10222 => x"2e80fb38",
         10223 => x"800b8318",
         10224 => x"34ff0bb4",
         10225 => x"180c7a55",
         10226 => x"80567aff",
         10227 => x"2ea53881",
         10228 => x"547a53b8",
         10229 => x"17528117",
         10230 => x"3351ffb4",
         10231 => x"863f84b9",
         10232 => x"c808762e",
         10233 => x"8538ff55",
         10234 => x"815674b4",
         10235 => x"180c8458",
         10236 => x"75bf3881",
         10237 => x"1f337f33",
         10238 => x"71882b07",
         10239 => x"5d5e8358",
         10240 => x"7b82d4d5",
         10241 => x"2e098106",
         10242 => x"a838800b",
         10243 => x"b8183357",
         10244 => x"587581e9",
         10245 => x"2e82b738",
         10246 => x"7581eb32",
         10247 => x"70307080",
         10248 => x"257a0742",
         10249 => x"42427fbc",
         10250 => x"387581e8",
         10251 => x"2eb63882",
         10252 => x"587781ff",
         10253 => x"0656800b",
         10254 => x"84b9bd1e",
         10255 => x"335d587b",
         10256 => x"782e0981",
         10257 => x"06833881",
         10258 => x"58817627",
         10259 => x"f8bd3877",
         10260 => x"802ef8b7",
         10261 => x"38811a84",
         10262 => x"1a5a5a83",
         10263 => x"7a27fed1",
         10264 => x"38f8a839",
         10265 => x"830b80ee",
         10266 => x"1883e4f8",
         10267 => x"405d587b",
         10268 => x"7081055d",
         10269 => x"337e7081",
         10270 => x"05403371",
         10271 => x"7131ff1b",
         10272 => x"5b525656",
         10273 => x"77802e80",
         10274 => x"c5387580",
         10275 => x"2ee13885",
         10276 => x"0b818a18",
         10277 => x"83e4fc40",
         10278 => x"5d587b70",
         10279 => x"81055d33",
         10280 => x"7e708105",
         10281 => x"40337171",
         10282 => x"31ff1b5b",
         10283 => x"58424077",
         10284 => x"802e858e",
         10285 => x"3875802e",
         10286 => x"e1388258",
         10287 => x"fef3398d",
         10288 => x"587cfa93",
         10289 => x"387784b9",
         10290 => x"c80c973d",
         10291 => x"0d047558",
         10292 => x"75802efe",
         10293 => x"dc38850b",
         10294 => x"818a1883",
         10295 => x"e4fc405d",
         10296 => x"58ffb739",
         10297 => x"8d0b84b9",
         10298 => x"c80c973d",
         10299 => x"0d04830b",
         10300 => x"80ee1883",
         10301 => x"e4f85c5a",
         10302 => x"58787081",
         10303 => x"055a337a",
         10304 => x"7081055c",
         10305 => x"33717131",
         10306 => x"ff1b5b57",
         10307 => x"5f5f7780",
         10308 => x"2e83d138",
         10309 => x"74802ee1",
         10310 => x"38850b81",
         10311 => x"8a1883e4",
         10312 => x"fc5c5a58",
         10313 => x"78708105",
         10314 => x"5a337a70",
         10315 => x"81055c33",
         10316 => x"717131ff",
         10317 => x"1b5b5842",
         10318 => x"4077802e",
         10319 => x"84913875",
         10320 => x"802ee138",
         10321 => x"933d7757",
         10322 => x"5a8359fc",
         10323 => x"83398158",
         10324 => x"fdc63980",
         10325 => x"e9173380",
         10326 => x"e8183371",
         10327 => x"882b0757",
         10328 => x"5575812e",
         10329 => x"098106f9",
         10330 => x"d538811b",
         10331 => x"58805ab4",
         10332 => x"1708782e",
         10333 => x"b1388317",
         10334 => x"335b7a7a",
         10335 => x"2e098106",
         10336 => x"829b3881",
         10337 => x"547753b8",
         10338 => x"17528117",
         10339 => x"3351ffb0",
         10340 => x"d23f84b9",
         10341 => x"c808802e",
         10342 => x"8538ff58",
         10343 => x"815a77b4",
         10344 => x"180c79f9",
         10345 => x"99387984",
         10346 => x"183484b7",
         10347 => x"173384b6",
         10348 => x"18337188",
         10349 => x"2b07575e",
         10350 => x"7582d4d5",
         10351 => x"2e098106",
         10352 => x"f8fc38b8",
         10353 => x"17831133",
         10354 => x"82123371",
         10355 => x"902b7188",
         10356 => x"2b078114",
         10357 => x"33707207",
         10358 => x"882b7533",
         10359 => x"71075e41",
         10360 => x"5945425c",
         10361 => x"5977848b",
         10362 => x"85a4d22e",
         10363 => x"098106f8",
         10364 => x"cd38849c",
         10365 => x"17831133",
         10366 => x"82123371",
         10367 => x"902b7188",
         10368 => x"2b078114",
         10369 => x"33707207",
         10370 => x"882b7533",
         10371 => x"71074744",
         10372 => x"405b5c5a",
         10373 => x"5e60868a",
         10374 => x"85e4f22e",
         10375 => x"098106f8",
         10376 => x"9d3884a0",
         10377 => x"17831133",
         10378 => x"82123371",
         10379 => x"902b7188",
         10380 => x"2b078114",
         10381 => x"33707207",
         10382 => x"882b7533",
         10383 => x"7107941e",
         10384 => x"0c5d84a4",
         10385 => x"1c831133",
         10386 => x"82123371",
         10387 => x"902b7188",
         10388 => x"2b078114",
         10389 => x"33707207",
         10390 => x"882b7533",
         10391 => x"71076290",
         10392 => x"050c5944",
         10393 => x"49465c45",
         10394 => x"40455b56",
         10395 => x"5a7c7734",
         10396 => x"84d1a022",
         10397 => x"81055d7c",
         10398 => x"84d1a023",
         10399 => x"7c861823",
         10400 => x"84d1a80b",
         10401 => x"8c180c80",
         10402 => x"0b98180c",
         10403 => x"f7cf397b",
         10404 => x"8324f8f0",
         10405 => x"387b7a7f",
         10406 => x"0c56f295",
         10407 => x"397554b4",
         10408 => x"170853b8",
         10409 => x"17705381",
         10410 => x"18335259",
         10411 => x"ffafb33f",
         10412 => x"84b9c808",
         10413 => x"7a2e0981",
         10414 => x"0681a438",
         10415 => x"84b9c808",
         10416 => x"831834b4",
         10417 => x"1708a818",
         10418 => x"0831407f",
         10419 => x"a0180827",
         10420 => x"8b388217",
         10421 => x"33416082",
         10422 => x"2e818d38",
         10423 => x"84b9c808",
         10424 => x"5afda039",
         10425 => x"74567480",
         10426 => x"2ef39138",
         10427 => x"850b818a",
         10428 => x"1883e4fc",
         10429 => x"5c5a58fc",
         10430 => x"ab3980e3",
         10431 => x"173380e2",
         10432 => x"18337188",
         10433 => x"2b075f5a",
         10434 => x"8d587df6",
         10435 => x"d2388817",
         10436 => x"224261f6",
         10437 => x"ca3880e4",
         10438 => x"17831133",
         10439 => x"82123371",
         10440 => x"902b7188",
         10441 => x"2b078114",
         10442 => x"33707207",
         10443 => x"882b7533",
         10444 => x"7107ac1e",
         10445 => x"0c5a7d82",
         10446 => x"2b5a4344",
         10447 => x"405940f5",
         10448 => x"d8397558",
         10449 => x"75802ef9",
         10450 => x"e8388258",
         10451 => x"f9e33975",
         10452 => x"802ef2a8",
         10453 => x"38933d77",
         10454 => x"575a8359",
         10455 => x"f7f23975",
         10456 => x"5a79f5da",
         10457 => x"38fcbf39",
         10458 => x"7554b417",
         10459 => x"08a01808",
         10460 => x"05537852",
         10461 => x"81173351",
         10462 => x"ffade73f",
         10463 => x"fc8539f0",
         10464 => x"3d0d0280",
         10465 => x"d3053364",
         10466 => x"7043933d",
         10467 => x"41575dff",
         10468 => x"765a4075",
         10469 => x"802e80e9",
         10470 => x"38787081",
         10471 => x"055a3370",
         10472 => x"9f265555",
         10473 => x"74ba2e80",
         10474 => x"e23873ed",
         10475 => x"3874ba2e",
         10476 => x"80d93884",
         10477 => x"d1a43354",
         10478 => x"80742480",
         10479 => x"c4387310",
         10480 => x"1084d190",
         10481 => x"05700855",
         10482 => x"5573802e",
         10483 => x"84388074",
         10484 => x"34625473",
         10485 => x"802e8638",
         10486 => x"80743462",
         10487 => x"5473750c",
         10488 => x"7c547c80",
         10489 => x"2e923880",
         10490 => x"53933d70",
         10491 => x"53840551",
         10492 => x"ef813f84",
         10493 => x"b9c80854",
         10494 => x"7384b9c8",
         10495 => x"0c923d0d",
         10496 => x"048b0b84",
         10497 => x"b9c80c92",
         10498 => x"3d0d0475",
         10499 => x"33d01170",
         10500 => x"81ff0656",
         10501 => x"56577389",
         10502 => x"26913882",
         10503 => x"167781ff",
         10504 => x"06d0055c",
         10505 => x"5877792e",
         10506 => x"80f73880",
         10507 => x"7f0883e5",
         10508 => x"b85e5f5b",
         10509 => x"7b087e59",
         10510 => x"5a797081",
         10511 => x"055b3378",
         10512 => x"7081055a",
         10513 => x"33ff9f12",
         10514 => x"59575576",
         10515 => x"99268938",
         10516 => x"e0157081",
         10517 => x"ff065654",
         10518 => x"ff9f1657",
         10519 => x"76992689",
         10520 => x"38e01670",
         10521 => x"81ff0657",
         10522 => x"54743070",
         10523 => x"9f2a5854",
         10524 => x"74762e09",
         10525 => x"81068538",
         10526 => x"76ffbe38",
         10527 => x"77793270",
         10528 => x"30707207",
         10529 => x"9f2a7907",
         10530 => x"5c575479",
         10531 => x"802e9238",
         10532 => x"811b841d",
         10533 => x"5d5b837b",
         10534 => x"25ff9938",
         10535 => x"7f54fe98",
         10536 => x"397a8324",
         10537 => x"f7387a79",
         10538 => x"600c54fe",
         10539 => x"8b39e63d",
         10540 => x"0d6c0284",
         10541 => x"0580fb05",
         10542 => x"33565989",
         10543 => x"5678802e",
         10544 => x"a63874bf",
         10545 => x"0670549d",
         10546 => x"3dcc0553",
         10547 => x"9e3d8405",
         10548 => x"5258ed9f",
         10549 => x"3f84b9c8",
         10550 => x"085784b9",
         10551 => x"c808802e",
         10552 => x"8f388079",
         10553 => x"0c765675",
         10554 => x"84b9c80c",
         10555 => x"9c3d0d04",
         10556 => x"7e406d52",
         10557 => x"903d7052",
         10558 => x"5ae19a3f",
         10559 => x"84b9c808",
         10560 => x"5784b9c8",
         10561 => x"08802e81",
         10562 => x"ba38779c",
         10563 => x"065d7c80",
         10564 => x"2e81ca38",
         10565 => x"76802e83",
         10566 => x"c1387684",
         10567 => x"2e83ea38",
         10568 => x"77880758",
         10569 => x"76ffbb38",
         10570 => x"77832a81",
         10571 => x"065b7a80",
         10572 => x"2e81d138",
         10573 => x"669b1133",
         10574 => x"9a123371",
         10575 => x"882b0761",
         10576 => x"70334258",
         10577 => x"5e5e567d",
         10578 => x"832e84e9",
         10579 => x"38800b8e",
         10580 => x"1734800b",
         10581 => x"8f1734a1",
         10582 => x"0b901734",
         10583 => x"80cc0b91",
         10584 => x"17346656",
         10585 => x"a00b8b17",
         10586 => x"347e6757",
         10587 => x"5e800b9a",
         10588 => x"1734800b",
         10589 => x"9b17347d",
         10590 => x"335d7c83",
         10591 => x"2e84a938",
         10592 => x"665b800b",
         10593 => x"9c1c3480",
         10594 => x"0b9d1c34",
         10595 => x"800b9e1c",
         10596 => x"34800b9f",
         10597 => x"1c347e55",
         10598 => x"810b8316",
         10599 => x"347b802e",
         10600 => x"80e2387e",
         10601 => x"b411087d",
         10602 => x"7c085357",
         10603 => x"5f57817c",
         10604 => x"2789389c",
         10605 => x"17087c26",
         10606 => x"838a3882",
         10607 => x"5780790c",
         10608 => x"fea33902",
         10609 => x"80e70533",
         10610 => x"70982b5d",
         10611 => x"5b7b8025",
         10612 => x"feb83886",
         10613 => x"789c065e",
         10614 => x"577cfeb8",
         10615 => x"3876fe82",
         10616 => x"380280c2",
         10617 => x"05337084",
         10618 => x"2a81065d",
         10619 => x"567b8291",
         10620 => x"3877812a",
         10621 => x"81065e7d",
         10622 => x"802e8938",
         10623 => x"7581065a",
         10624 => x"7981f638",
         10625 => x"77832a81",
         10626 => x"06567580",
         10627 => x"2e863877",
         10628 => x"80c00758",
         10629 => x"7eb41108",
         10630 => x"a01b0c67",
         10631 => x"a41b0c67",
         10632 => x"9b11339a",
         10633 => x"12337188",
         10634 => x"2b077333",
         10635 => x"405e4057",
         10636 => x"5a7b832e",
         10637 => x"81f1387a",
         10638 => x"881a0c9c",
         10639 => x"16831133",
         10640 => x"82123371",
         10641 => x"902b7188",
         10642 => x"2b078114",
         10643 => x"33707207",
         10644 => x"882b7533",
         10645 => x"71077060",
         10646 => x"8c050c60",
         10647 => x"600c5152",
         10648 => x"4159575d",
         10649 => x"5e861a22",
         10650 => x"841a2377",
         10651 => x"901a3480",
         10652 => x"0b911a34",
         10653 => x"800b9c1a",
         10654 => x"0c77852a",
         10655 => x"81065574",
         10656 => x"802e84ac",
         10657 => x"3875802e",
         10658 => x"84f13875",
         10659 => x"941a0c8a",
         10660 => x"1a227089",
         10661 => x"2b7c525b",
         10662 => x"58763070",
         10663 => x"78078025",
         10664 => x"565b7976",
         10665 => x"27849238",
         10666 => x"81707606",
         10667 => x"5f5b7d80",
         10668 => x"2e848638",
         10669 => x"77527851",
         10670 => x"ffacdb3f",
         10671 => x"84b9c808",
         10672 => x"5884b9c8",
         10673 => x"08812683",
         10674 => x"38825784",
         10675 => x"b9c808ff",
         10676 => x"2e80cb38",
         10677 => x"757a3156",
         10678 => x"c0390280",
         10679 => x"c2053391",
         10680 => x"065e7d95",
         10681 => x"3877822a",
         10682 => x"81065574",
         10683 => x"802efcb8",
         10684 => x"38885780",
         10685 => x"790cfbed",
         10686 => x"39875780",
         10687 => x"790cfbe5",
         10688 => x"39845780",
         10689 => x"790cfbdd",
         10690 => x"397951cd",
         10691 => x"ca3f84b9",
         10692 => x"c8087888",
         10693 => x"07595776",
         10694 => x"fbc838fc",
         10695 => x"8b397a76",
         10696 => x"7b315757",
         10697 => x"fef33995",
         10698 => x"16339417",
         10699 => x"3371982b",
         10700 => x"71902b07",
         10701 => x"7d075d5e",
         10702 => x"5cfdfc39",
         10703 => x"7c557c7b",
         10704 => x"2781bd38",
         10705 => x"74527951",
         10706 => x"ffabcb3f",
         10707 => x"84b9c808",
         10708 => x"5d84b9c8",
         10709 => x"08802e81",
         10710 => x"a73884b9",
         10711 => x"c808812e",
         10712 => x"fcd93884",
         10713 => x"b9c808ff",
         10714 => x"2e839938",
         10715 => x"80537452",
         10716 => x"7651ffb2",
         10717 => x"823f84b9",
         10718 => x"c8088390",
         10719 => x"389c1708",
         10720 => x"fe119419",
         10721 => x"0858565b",
         10722 => x"757527ff",
         10723 => x"af388116",
         10724 => x"94180c84",
         10725 => x"17338107",
         10726 => x"55748418",
         10727 => x"347c557a",
         10728 => x"7d26ffa0",
         10729 => x"3880d939",
         10730 => x"800b9417",
         10731 => x"34800b95",
         10732 => x"1734fbcc",
         10733 => x"39951633",
         10734 => x"94173371",
         10735 => x"982b7190",
         10736 => x"2b077e07",
         10737 => x"5e565b80",
         10738 => x"0b8e1734",
         10739 => x"800b8f17",
         10740 => x"34a10b90",
         10741 => x"173480cc",
         10742 => x"0b911734",
         10743 => x"6656a00b",
         10744 => x"8b17347e",
         10745 => x"67575e80",
         10746 => x"0b9a1734",
         10747 => x"800b9b17",
         10748 => x"347d335d",
         10749 => x"7c832e09",
         10750 => x"8106fb84",
         10751 => x"38ffa939",
         10752 => x"807f7f72",
         10753 => x"5e59575d",
         10754 => x"b416087e",
         10755 => x"2eae3883",
         10756 => x"16335a79",
         10757 => x"7d2e0981",
         10758 => x"06b53881",
         10759 => x"547d53b8",
         10760 => x"16528116",
         10761 => x"3351ffa3",
         10762 => x"ba3f84b9",
         10763 => x"c808802e",
         10764 => x"8538ff57",
         10765 => x"815b76b4",
         10766 => x"170c7e56",
         10767 => x"7aff1d90",
         10768 => x"180c577a",
         10769 => x"802efbbc",
         10770 => x"3880790c",
         10771 => x"f9973981",
         10772 => x"54b41608",
         10773 => x"53b81670",
         10774 => x"53811733",
         10775 => x"525affa4",
         10776 => x"813f84b9",
         10777 => x"c8087d2e",
         10778 => x"09810681",
         10779 => x"aa3884b9",
         10780 => x"c8088317",
         10781 => x"34b41608",
         10782 => x"a8170831",
         10783 => x"84b9c808",
         10784 => x"5c5574a0",
         10785 => x"170827ff",
         10786 => x"92388216",
         10787 => x"33557482",
         10788 => x"2e098106",
         10789 => x"ff853881",
         10790 => x"54b41608",
         10791 => x"a0170805",
         10792 => x"53795281",
         10793 => x"163351ff",
         10794 => x"a3b83f7c",
         10795 => x"5bfeec39",
         10796 => x"74941a0c",
         10797 => x"7656f8af",
         10798 => x"3977981a",
         10799 => x"0c76f8a2",
         10800 => x"387583ff",
         10801 => x"065a7980",
         10802 => x"2ef89a38",
         10803 => x"7efe199c",
         10804 => x"1208fe05",
         10805 => x"5f595a77",
         10806 => x"7d27f9df",
         10807 => x"388a1a22",
         10808 => x"787129b0",
         10809 => x"1c080556",
         10810 => x"5c74802e",
         10811 => x"f9cd3875",
         10812 => x"892a159c",
         10813 => x"1a0c7656",
         10814 => x"f7ed3975",
         10815 => x"941a0c76",
         10816 => x"56f7e439",
         10817 => x"81578079",
         10818 => x"0cf7da39",
         10819 => x"84b9c808",
         10820 => x"5780790c",
         10821 => x"f7cf3981",
         10822 => x"7f575bfe",
         10823 => x"9f39f03d",
         10824 => x"0d626567",
         10825 => x"6640405d",
         10826 => x"5a807e0c",
         10827 => x"89577980",
         10828 => x"2e9f3879",
         10829 => x"08567580",
         10830 => x"2e973875",
         10831 => x"33557480",
         10832 => x"2e8f3886",
         10833 => x"1622841b",
         10834 => x"22595978",
         10835 => x"782e84b7",
         10836 => x"38805574",
         10837 => x"41765576",
         10838 => x"828c3891",
         10839 => x"1a335574",
         10840 => x"82843890",
         10841 => x"1a338106",
         10842 => x"57875676",
         10843 => x"802e81ed",
         10844 => x"38941a08",
         10845 => x"8c1b0871",
         10846 => x"3156567b",
         10847 => x"752681ef",
         10848 => x"387b802e",
         10849 => x"81d53860",
         10850 => x"597583ff",
         10851 => x"065b7a81",
         10852 => x"e3388a19",
         10853 => x"22ff0576",
         10854 => x"892a065b",
         10855 => x"7a9b3875",
         10856 => x"83d33888",
         10857 => x"1a085581",
         10858 => x"75278485",
         10859 => x"3874ff2e",
         10860 => x"83f03874",
         10861 => x"981b0c60",
         10862 => x"59981a08",
         10863 => x"fe059c1a",
         10864 => x"08fe0541",
         10865 => x"57766027",
         10866 => x"83e7388a",
         10867 => x"19227078",
         10868 => x"29b01b08",
         10869 => x"05565674",
         10870 => x"802e83d5",
         10871 => x"387a157c",
         10872 => x"892a5957",
         10873 => x"77802e83",
         10874 => x"8138771b",
         10875 => x"55757527",
         10876 => x"8538757b",
         10877 => x"31587754",
         10878 => x"76537c52",
         10879 => x"81193351",
         10880 => x"ff9fe03f",
         10881 => x"84b9c808",
         10882 => x"83983860",
         10883 => x"83113357",
         10884 => x"5975802e",
         10885 => x"a938b419",
         10886 => x"08773156",
         10887 => x"7578279e",
         10888 => x"38848076",
         10889 => x"71291eb8",
         10890 => x"1b585855",
         10891 => x"75708105",
         10892 => x"57337770",
         10893 => x"81055934",
         10894 => x"ff155574",
         10895 => x"ef387789",
         10896 => x"2b587b78",
         10897 => x"317e0819",
         10898 => x"7f0c781e",
         10899 => x"941c081a",
         10900 => x"7059941d",
         10901 => x"0c5e5c7b",
         10902 => x"feaf3880",
         10903 => x"567584b9",
         10904 => x"c80c923d",
         10905 => x"0d047484",
         10906 => x"b9c80c92",
         10907 => x"3d0d0474",
         10908 => x"5cfe8e39",
         10909 => x"9c1a0857",
         10910 => x"7583ff06",
         10911 => x"84807131",
         10912 => x"595b7b78",
         10913 => x"2783387b",
         10914 => x"587656b4",
         10915 => x"1908772e",
         10916 => x"b638800b",
         10917 => x"831a3371",
         10918 => x"5d415f7f",
         10919 => x"7f2e0981",
         10920 => x"0680e438",
         10921 => x"81547653",
         10922 => x"b8195281",
         10923 => x"193351ff",
         10924 => x"9eb13f84",
         10925 => x"b9c80880",
         10926 => x"2e8538ff",
         10927 => x"56815b75",
         10928 => x"b41a0c7a",
         10929 => x"81dc3860",
         10930 => x"941b0883",
         10931 => x"ff061179",
         10932 => x"7f5a58b8",
         10933 => x"05565977",
         10934 => x"802efee6",
         10935 => x"38747081",
         10936 => x"05563377",
         10937 => x"70810559",
         10938 => x"34ff1656",
         10939 => x"75802efe",
         10940 => x"d1387470",
         10941 => x"81055633",
         10942 => x"77708105",
         10943 => x"5934ff16",
         10944 => x"5675da38",
         10945 => x"febc3981",
         10946 => x"54b41908",
         10947 => x"53b81970",
         10948 => x"53811a33",
         10949 => x"5240ff9e",
         10950 => x"c93f815b",
         10951 => x"84b9c808",
         10952 => x"7f2e0981",
         10953 => x"06ff9c38",
         10954 => x"84b9c808",
         10955 => x"831a34b4",
         10956 => x"1908a81a",
         10957 => x"083184b9",
         10958 => x"c8085c55",
         10959 => x"74a01a08",
         10960 => x"27fee138",
         10961 => x"82193355",
         10962 => x"74822e09",
         10963 => x"8106fed4",
         10964 => x"388154b4",
         10965 => x"1908a01a",
         10966 => x"0805537f",
         10967 => x"52811933",
         10968 => x"51ff9dfe",
         10969 => x"3f7e5bfe",
         10970 => x"bb39769c",
         10971 => x"1b0c941a",
         10972 => x"0856fe84",
         10973 => x"39981a08",
         10974 => x"527951ff",
         10975 => x"a3983f84",
         10976 => x"b9c80855",
         10977 => x"fca13981",
         10978 => x"163351ff",
         10979 => x"9c833f84",
         10980 => x"b9c80881",
         10981 => x"065574fb",
         10982 => x"b838747a",
         10983 => x"085657fb",
         10984 => x"b239810b",
         10985 => x"911b3481",
         10986 => x"0b84b9c8",
         10987 => x"0c923d0d",
         10988 => x"04820b91",
         10989 => x"1b34820b",
         10990 => x"84b9c80c",
         10991 => x"923d0d04",
         10992 => x"f03d0d62",
         10993 => x"65676640",
         10994 => x"405c5a80",
         10995 => x"7e0c8957",
         10996 => x"79802e9f",
         10997 => x"38790856",
         10998 => x"75802e97",
         10999 => x"38753355",
         11000 => x"74802e8f",
         11001 => x"38861622",
         11002 => x"841b2259",
         11003 => x"5978782e",
         11004 => x"85fd3880",
         11005 => x"55744176",
         11006 => x"557682c4",
         11007 => x"38911a33",
         11008 => x"557482bc",
         11009 => x"38901a33",
         11010 => x"70812a81",
         11011 => x"06585887",
         11012 => x"5676802e",
         11013 => x"82a13894",
         11014 => x"1a087b11",
         11015 => x"5d577b77",
         11016 => x"27843876",
         11017 => x"095b7a80",
         11018 => x"2e828138",
         11019 => x"7683ff06",
         11020 => x"5f7e82a2",
         11021 => x"38608a11",
         11022 => x"22ff0578",
         11023 => x"892a065a",
         11024 => x"5678aa38",
         11025 => x"76849e38",
         11026 => x"881a0855",
         11027 => x"74802e84",
         11028 => x"b1387481",
         11029 => x"2e86a138",
         11030 => x"74ff2e86",
         11031 => x"8c387498",
         11032 => x"1b0c881a",
         11033 => x"08853874",
         11034 => x"881b0c60",
         11035 => x"56b41608",
         11036 => x"9c1b082e",
         11037 => x"81d33898",
         11038 => x"1a08fe05",
         11039 => x"9c1708fe",
         11040 => x"05585877",
         11041 => x"772785f0",
         11042 => x"388a1622",
         11043 => x"707929b0",
         11044 => x"18080556",
         11045 => x"5774802e",
         11046 => x"85de3878",
         11047 => x"157b892a",
         11048 => x"595c7780",
         11049 => x"2e839838",
         11050 => x"77195f76",
         11051 => x"7f278538",
         11052 => x"76793158",
         11053 => x"77547b53",
         11054 => x"7c528116",
         11055 => x"3351ff9b",
         11056 => x"a13f84b9",
         11057 => x"c80885a1",
         11058 => x"3860b411",
         11059 => x"087d3156",
         11060 => x"57747827",
         11061 => x"a5388480",
         11062 => x"0bb81876",
         11063 => x"72291f57",
         11064 => x"58567470",
         11065 => x"81055633",
         11066 => x"77708105",
         11067 => x"5934ff16",
         11068 => x"5675ef38",
         11069 => x"60597583",
         11070 => x"1a347789",
         11071 => x"2b597a79",
         11072 => x"317e081a",
         11073 => x"7f0c791e",
         11074 => x"941c081b",
         11075 => x"7071941f",
         11076 => x"0c8c1e08",
         11077 => x"5a5a575e",
         11078 => x"5b757527",
         11079 => x"83387456",
         11080 => x"758c1b0c",
         11081 => x"7afe8538",
         11082 => x"901a3358",
         11083 => x"7780c007",
         11084 => x"5b7a901b",
         11085 => x"34805675",
         11086 => x"84b9c80c",
         11087 => x"923d0d04",
         11088 => x"7484b9c8",
         11089 => x"0c923d0d",
         11090 => x"04831633",
         11091 => x"557482c8",
         11092 => x"386056fe",
         11093 => x"a239609c",
         11094 => x"1b085956",
         11095 => x"7683ff06",
         11096 => x"84807131",
         11097 => x"5a5c7a79",
         11098 => x"2783387a",
         11099 => x"597757b4",
         11100 => x"1608782e",
         11101 => x"b638800b",
         11102 => x"83173371",
         11103 => x"5e415f7f",
         11104 => x"7f2e0981",
         11105 => x"0680d538",
         11106 => x"81547753",
         11107 => x"b8165281",
         11108 => x"163351ff",
         11109 => x"98cd3f84",
         11110 => x"b9c80880",
         11111 => x"2e8538ff",
         11112 => x"57815c76",
         11113 => x"b4170c7b",
         11114 => x"83bf3860",
         11115 => x"941b0883",
         11116 => x"ff06117a",
         11117 => x"58b8057e",
         11118 => x"59565878",
         11119 => x"802e9538",
         11120 => x"76708105",
         11121 => x"58337570",
         11122 => x"81055734",
         11123 => x"ff165675",
         11124 => x"ef386058",
         11125 => x"810b8319",
         11126 => x"34fea339",
         11127 => x"8154b416",
         11128 => x"0853b816",
         11129 => x"70538117",
         11130 => x"335240ff",
         11131 => x"98f43f81",
         11132 => x"5c84b9c8",
         11133 => x"087f2e09",
         11134 => x"8106ffab",
         11135 => x"3884b9c8",
         11136 => x"08831734",
         11137 => x"b41608a8",
         11138 => x"17083184",
         11139 => x"b9c8085d",
         11140 => x"5574a017",
         11141 => x"0827fef0",
         11142 => x"38821633",
         11143 => x"5574822e",
         11144 => x"098106fe",
         11145 => x"e3388154",
         11146 => x"b41608a0",
         11147 => x"17080553",
         11148 => x"7f528116",
         11149 => x"3351ff98",
         11150 => x"a93f7e5c",
         11151 => x"feca3994",
         11152 => x"1a08578c",
         11153 => x"1a087726",
         11154 => x"93388316",
         11155 => x"33407f81",
         11156 => x"b938607c",
         11157 => x"b4120c94",
         11158 => x"1b085856",
         11159 => x"7b7c9c1c",
         11160 => x"0c58fdf8",
         11161 => x"39981a08",
         11162 => x"527951ff",
         11163 => x"abe73f84",
         11164 => x"b9c80855",
         11165 => x"84b9c808",
         11166 => x"fbd83890",
         11167 => x"1a3358fd",
         11168 => x"ab397652",
         11169 => x"7951ffab",
         11170 => x"cc3f84b9",
         11171 => x"c8085584",
         11172 => x"b9c808fb",
         11173 => x"bd38e439",
         11174 => x"8154b416",
         11175 => x"0853b816",
         11176 => x"70538117",
         11177 => x"335257ff",
         11178 => x"97b83f84",
         11179 => x"b9c80881",
         11180 => x"b83884b9",
         11181 => x"c8088317",
         11182 => x"34b41608",
         11183 => x"a8170831",
         11184 => x"5877a017",
         11185 => x"0827fd89",
         11186 => x"38821633",
         11187 => x"5c7b822e",
         11188 => x"098106fc",
         11189 => x"fc388154",
         11190 => x"b41608a0",
         11191 => x"17080553",
         11192 => x"76528116",
         11193 => x"3351ff96",
         11194 => x"f93f6056",
         11195 => x"fb893981",
         11196 => x"163351ff",
         11197 => x"959b3f84",
         11198 => x"b9c80881",
         11199 => x"065574f9",
         11200 => x"f238747a",
         11201 => x"085657f9",
         11202 => x"ec398154",
         11203 => x"b4160853",
         11204 => x"b8167053",
         11205 => x"81173352",
         11206 => x"57ff96c6",
         11207 => x"3f84b9c8",
         11208 => x"0880c638",
         11209 => x"84b9c808",
         11210 => x"831734b4",
         11211 => x"1608a817",
         11212 => x"08315574",
         11213 => x"a0170827",
         11214 => x"fe983882",
         11215 => x"16335877",
         11216 => x"822e0981",
         11217 => x"06fe8b38",
         11218 => x"8154b416",
         11219 => x"08a01708",
         11220 => x"05537652",
         11221 => x"81163351",
         11222 => x"ff96873f",
         11223 => x"607cb412",
         11224 => x"0c941b08",
         11225 => x"5856fdf4",
         11226 => x"39810b91",
         11227 => x"1b34810b",
         11228 => x"84b9c80c",
         11229 => x"923d0d04",
         11230 => x"820b911b",
         11231 => x"34820b84",
         11232 => x"b9c80c92",
         11233 => x"3d0d04f5",
         11234 => x"3d0d7d58",
         11235 => x"895a7780",
         11236 => x"2e9f3877",
         11237 => x"08567580",
         11238 => x"2e973875",
         11239 => x"33557480",
         11240 => x"2e8f3886",
         11241 => x"16228419",
         11242 => x"22585978",
         11243 => x"772e83b5",
         11244 => x"38805574",
         11245 => x"5c795679",
         11246 => x"81d83890",
         11247 => x"18337086",
         11248 => x"2a81065c",
         11249 => x"577a802e",
         11250 => x"81c8387b",
         11251 => x"a019085a",
         11252 => x"57b41708",
         11253 => x"792eac38",
         11254 => x"8317335b",
         11255 => x"7a81bc38",
         11256 => x"81547853",
         11257 => x"b8175281",
         11258 => x"173351ff",
         11259 => x"93f53f84",
         11260 => x"b9c80880",
         11261 => x"2e8538ff",
         11262 => x"59815678",
         11263 => x"b4180c75",
         11264 => x"819038a4",
         11265 => x"18088b11",
         11266 => x"33a0075a",
         11267 => x"57788b18",
         11268 => x"34770888",
         11269 => x"19087083",
         11270 => x"ffff065d",
         11271 => x"5a567a9a",
         11272 => x"18347a88",
         11273 => x"2a5a799b",
         11274 => x"18349c17",
         11275 => x"76339619",
         11276 => x"5c565b74",
         11277 => x"832e81c1",
         11278 => x"388c1808",
         11279 => x"55747b34",
         11280 => x"74882a5b",
         11281 => x"7a9d1834",
         11282 => x"74902a56",
         11283 => x"759e1834",
         11284 => x"74982a59",
         11285 => x"789f1834",
         11286 => x"807a3480",
         11287 => x"0b971834",
         11288 => x"a10b9818",
         11289 => x"3480cc0b",
         11290 => x"99183480",
         11291 => x"0b921834",
         11292 => x"800b9318",
         11293 => x"347b5b81",
         11294 => x"0b831c34",
         11295 => x"7b51ff96",
         11296 => x"943f84b9",
         11297 => x"c8089019",
         11298 => x"3381bf06",
         11299 => x"5b567990",
         11300 => x"19347584",
         11301 => x"b9c80c8d",
         11302 => x"3d0d0481",
         11303 => x"54b41708",
         11304 => x"53b81770",
         11305 => x"53811833",
         11306 => x"525bff93",
         11307 => x"b53f8156",
         11308 => x"84b9c808",
         11309 => x"fec93884",
         11310 => x"b9c80883",
         11311 => x"1834b417",
         11312 => x"08a81808",
         11313 => x"3184b9c8",
         11314 => x"08575574",
         11315 => x"a0180827",
         11316 => x"fe8e3882",
         11317 => x"17335574",
         11318 => x"822e0981",
         11319 => x"06fe8138",
         11320 => x"8154b417",
         11321 => x"08a01808",
         11322 => x"05537a52",
         11323 => x"81173351",
         11324 => x"ff92ef3f",
         11325 => x"7956fde8",
         11326 => x"3978902a",
         11327 => x"55749418",
         11328 => x"3474882a",
         11329 => x"56759518",
         11330 => x"348c1808",
         11331 => x"55747b34",
         11332 => x"74882a5b",
         11333 => x"7a9d1834",
         11334 => x"74902a56",
         11335 => x"759e1834",
         11336 => x"74982a59",
         11337 => x"789f1834",
         11338 => x"807a3480",
         11339 => x"0b971834",
         11340 => x"a10b9818",
         11341 => x"3480cc0b",
         11342 => x"99183480",
         11343 => x"0b921834",
         11344 => x"800b9318",
         11345 => x"347b5b81",
         11346 => x"0b831c34",
         11347 => x"7b51ff94",
         11348 => x"c43f84b9",
         11349 => x"c8089019",
         11350 => x"3381bf06",
         11351 => x"5b567990",
         11352 => x"1934feae",
         11353 => x"39811633",
         11354 => x"51ff90a5",
         11355 => x"3f84b9c8",
         11356 => x"08810655",
         11357 => x"74fcba38",
         11358 => x"74780856",
         11359 => x"5afcb439",
         11360 => x"f93d0d79",
         11361 => x"705255fb",
         11362 => x"fe3f84b9",
         11363 => x"c8085484",
         11364 => x"b9c808b1",
         11365 => x"38895674",
         11366 => x"802e9e38",
         11367 => x"74085372",
         11368 => x"802e9638",
         11369 => x"72335271",
         11370 => x"802e8e38",
         11371 => x"86132284",
         11372 => x"16225852",
         11373 => x"71772e96",
         11374 => x"38805271",
         11375 => x"58755475",
         11376 => x"84387575",
         11377 => x"0c7384b9",
         11378 => x"c80c893d",
         11379 => x"0d048113",
         11380 => x"3351ff8f",
         11381 => x"bc3f84b9",
         11382 => x"c8088106",
         11383 => x"5372da38",
         11384 => x"73750853",
         11385 => x"56d539f6",
         11386 => x"3d0dff7d",
         11387 => x"705b575b",
         11388 => x"75802eb2",
         11389 => x"38757081",
         11390 => x"05573370",
         11391 => x"9f265252",
         11392 => x"71ba2eac",
         11393 => x"3870ee38",
         11394 => x"71ba2ea4",
         11395 => x"3884d1a4",
         11396 => x"33518071",
         11397 => x"24903870",
         11398 => x"84d1a434",
         11399 => x"800b84b9",
         11400 => x"c80c8c3d",
         11401 => x"0d048b0b",
         11402 => x"84b9c80c",
         11403 => x"8c3d0d04",
         11404 => x"7833d011",
         11405 => x"7081ff06",
         11406 => x"53535370",
         11407 => x"89269138",
         11408 => x"82197381",
         11409 => x"ff06d005",
         11410 => x"59547376",
         11411 => x"2e80f538",
         11412 => x"800b83e5",
         11413 => x"b85b5879",
         11414 => x"08795657",
         11415 => x"76708105",
         11416 => x"58337570",
         11417 => x"81055733",
         11418 => x"ff9f1253",
         11419 => x"54527099",
         11420 => x"268938e0",
         11421 => x"127081ff",
         11422 => x"065354ff",
         11423 => x"9f135170",
         11424 => x"99268938",
         11425 => x"e0137081",
         11426 => x"ff065454",
         11427 => x"7130709f",
         11428 => x"2a555171",
         11429 => x"732e0981",
         11430 => x"06853873",
         11431 => x"ffbe3874",
         11432 => x"76327030",
         11433 => x"7072079f",
         11434 => x"2a760759",
         11435 => x"52527680",
         11436 => x"2e923881",
         11437 => x"18841b5b",
         11438 => x"58837825",
         11439 => x"ff99387a",
         11440 => x"51fecf39",
         11441 => x"778324f7",
         11442 => x"3877765e",
         11443 => x"51fec339",
         11444 => x"ea3d0d80",
         11445 => x"53983dcc",
         11446 => x"0552993d",
         11447 => x"51d1943f",
         11448 => x"84b9c808",
         11449 => x"5584b9c8",
         11450 => x"08802e8a",
         11451 => x"387484b9",
         11452 => x"c80c983d",
         11453 => x"0d047a5c",
         11454 => x"6852983d",
         11455 => x"d00551c5",
         11456 => x"943f84b9",
         11457 => x"c8085584",
         11458 => x"b9c80880",
         11459 => x"c6380280",
         11460 => x"d7053370",
         11461 => x"982b585a",
         11462 => x"80772480",
         11463 => x"e23802b2",
         11464 => x"05337084",
         11465 => x"2a810657",
         11466 => x"5975802e",
         11467 => x"b2387a63",
         11468 => x"9b11339a",
         11469 => x"12337188",
         11470 => x"2b077333",
         11471 => x"5e5a5b57",
         11472 => x"5879832e",
         11473 => x"a4387698",
         11474 => x"190c7484",
         11475 => x"b9c80c98",
         11476 => x"3d0d0484",
         11477 => x"b9c80884",
         11478 => x"2e098106",
         11479 => x"ff8f3885",
         11480 => x"0b84b9c8",
         11481 => x"0c983d0d",
         11482 => x"04951633",
         11483 => x"94173371",
         11484 => x"982b7190",
         11485 => x"2b077907",
         11486 => x"981b0c5b",
         11487 => x"54cc397a",
         11488 => x"7e98120c",
         11489 => x"587484b9",
         11490 => x"c80c983d",
         11491 => x"0d04ff9e",
         11492 => x"3d0d80e6",
         11493 => x"3d0880e6",
         11494 => x"3d085d40",
         11495 => x"807c3480",
         11496 => x"5380e43d",
         11497 => x"fdb40552",
         11498 => x"80e53d51",
         11499 => x"cfc53f84",
         11500 => x"b9c80859",
         11501 => x"84b9c808",
         11502 => x"83c83860",
         11503 => x"80d93d0c",
         11504 => x"7f619811",
         11505 => x"0880dd3d",
         11506 => x"0c5880db",
         11507 => x"3d085b58",
         11508 => x"79802e82",
         11509 => x"cc3880d8",
         11510 => x"3d983d40",
         11511 => x"5ba0527a",
         11512 => x"51ffa4aa",
         11513 => x"3f84b9c8",
         11514 => x"085984b9",
         11515 => x"c8088392",
         11516 => x"386080df",
         11517 => x"3d085856",
         11518 => x"b4160877",
         11519 => x"2eb13884",
         11520 => x"b9c80883",
         11521 => x"17335f5d",
         11522 => x"7d83c738",
         11523 => x"81547653",
         11524 => x"b8165281",
         11525 => x"163351ff",
         11526 => x"8bc93f84",
         11527 => x"b9c80880",
         11528 => x"2e8538ff",
         11529 => x"57815976",
         11530 => x"b4170c78",
         11531 => x"82d43880",
         11532 => x"df3d089b",
         11533 => x"11339a12",
         11534 => x"3371882b",
         11535 => x"07637033",
         11536 => x"5d405956",
         11537 => x"5678832e",
         11538 => x"82da3876",
         11539 => x"80db3d0c",
         11540 => x"80527a51",
         11541 => x"ffa3b73f",
         11542 => x"84b9c808",
         11543 => x"5984b9c8",
         11544 => x"08829f38",
         11545 => x"80527a51",
         11546 => x"ffa8f53f",
         11547 => x"84b9c808",
         11548 => x"5984b9c8",
         11549 => x"08bb3880",
         11550 => x"df3d089b",
         11551 => x"11339a12",
         11552 => x"3371882b",
         11553 => x"07637033",
         11554 => x"4258595e",
         11555 => x"567d832e",
         11556 => x"81fd3876",
         11557 => x"7a2ea438",
         11558 => x"84b9c808",
         11559 => x"527a51ff",
         11560 => x"a4e23f84",
         11561 => x"b9c80859",
         11562 => x"84b9c808",
         11563 => x"802effb4",
         11564 => x"3878842e",
         11565 => x"83d83878",
         11566 => x"81c83880",
         11567 => x"e43dfdb8",
         11568 => x"05527a51",
         11569 => x"ffbd893f",
         11570 => x"787f8205",
         11571 => x"335b5779",
         11572 => x"802e9038",
         11573 => x"821f5681",
         11574 => x"17811770",
         11575 => x"335f5757",
         11576 => x"7cf53881",
         11577 => x"17567578",
         11578 => x"26819538",
         11579 => x"76802e9c",
         11580 => x"387e1782",
         11581 => x"0556ff18",
         11582 => x"80e63d08",
         11583 => x"11ff19ff",
         11584 => x"19595956",
         11585 => x"58753375",
         11586 => x"3476eb38",
         11587 => x"ff1880e6",
         11588 => x"3d08115f",
         11589 => x"58af7e34",
         11590 => x"80da3d08",
         11591 => x"5a79fdbd",
         11592 => x"3877602e",
         11593 => x"828a3880",
         11594 => x"0b84d1a4",
         11595 => x"33701010",
         11596 => x"83e5b805",
         11597 => x"70087033",
         11598 => x"4359595e",
         11599 => x"5a7e7a2e",
         11600 => x"8d38811a",
         11601 => x"70177033",
         11602 => x"575f5a74",
         11603 => x"f538821a",
         11604 => x"5b7a7826",
         11605 => x"ab388057",
         11606 => x"767a2794",
         11607 => x"3876165f",
         11608 => x"7e337c70",
         11609 => x"81055e34",
         11610 => x"81175779",
         11611 => x"7726ee38",
         11612 => x"ba7c7081",
         11613 => x"055e3476",
         11614 => x"ff2e0981",
         11615 => x"0681df38",
         11616 => x"9159807c",
         11617 => x"347884b9",
         11618 => x"c80c80e4",
         11619 => x"3d0d0495",
         11620 => x"16339417",
         11621 => x"3371982b",
         11622 => x"71902b07",
         11623 => x"79075956",
         11624 => x"5efdf039",
         11625 => x"95163394",
         11626 => x"17337198",
         11627 => x"2b71902b",
         11628 => x"07790780",
         11629 => x"dd3d0c5a",
         11630 => x"5d80527a",
         11631 => x"51ffa0ce",
         11632 => x"3f84b9c8",
         11633 => x"085984b9",
         11634 => x"c808802e",
         11635 => x"fd9638ff",
         11636 => x"b1398154",
         11637 => x"b4160853",
         11638 => x"b8167053",
         11639 => x"81173352",
         11640 => x"5eff88fe",
         11641 => x"3f815984",
         11642 => x"b9c808fc",
         11643 => x"be3884b9",
         11644 => x"c8088317",
         11645 => x"34b41608",
         11646 => x"a8170831",
         11647 => x"84b9c808",
         11648 => x"5a5574a0",
         11649 => x"170827fc",
         11650 => x"83388216",
         11651 => x"33557482",
         11652 => x"2e098106",
         11653 => x"fbf63881",
         11654 => x"54b41608",
         11655 => x"a0170805",
         11656 => x"537d5281",
         11657 => x"163351ff",
         11658 => x"88b83f7c",
         11659 => x"59fbdd39",
         11660 => x"ff1880e6",
         11661 => x"3d08115c",
         11662 => x"58af7b34",
         11663 => x"800b84d1",
         11664 => x"a4337010",
         11665 => x"1083e5b8",
         11666 => x"05700870",
         11667 => x"33435959",
         11668 => x"5e5a7e7a",
         11669 => x"2e098106",
         11670 => x"fde838fd",
         11671 => x"f13980e5",
         11672 => x"3d081881",
         11673 => x"19595a79",
         11674 => x"337c7081",
         11675 => x"055e3477",
         11676 => x"6027fe8e",
         11677 => x"3880e53d",
         11678 => x"08188119",
         11679 => x"595a7933",
         11680 => x"7c708105",
         11681 => x"5e347f78",
         11682 => x"26d438fd",
         11683 => x"f5398259",
         11684 => x"807c3478",
         11685 => x"84b9c80c",
         11686 => x"80e43d0d",
         11687 => x"04f73d0d",
         11688 => x"7b7d5855",
         11689 => x"89567480",
         11690 => x"2e9f3874",
         11691 => x"08547380",
         11692 => x"2e973873",
         11693 => x"33537280",
         11694 => x"2e8f3886",
         11695 => x"14228416",
         11696 => x"22595978",
         11697 => x"782e83a0",
         11698 => x"38805372",
         11699 => x"5a755375",
         11700 => x"81c23891",
         11701 => x"15335372",
         11702 => x"81ba388c",
         11703 => x"15085676",
         11704 => x"762681b9",
         11705 => x"38941508",
         11706 => x"54805876",
         11707 => x"782e81cc",
         11708 => x"38798a11",
         11709 => x"2270892b",
         11710 => x"525a5673",
         11711 => x"782e81f7",
         11712 => x"387552ff",
         11713 => x"1751fdbb",
         11714 => x"9c3f84b9",
         11715 => x"c808ff15",
         11716 => x"77547053",
         11717 => x"5553fdbb",
         11718 => x"8c3f84b9",
         11719 => x"c8087326",
         11720 => x"81d53875",
         11721 => x"30740670",
         11722 => x"94170c77",
         11723 => x"71319817",
         11724 => x"08565859",
         11725 => x"73802e82",
         11726 => x"98387577",
         11727 => x"2781d938",
         11728 => x"76763194",
         11729 => x"16081794",
         11730 => x"170c9016",
         11731 => x"3370812a",
         11732 => x"8106515a",
         11733 => x"5778802e",
         11734 => x"81fe3873",
         11735 => x"527451ff",
         11736 => x"99f33f84",
         11737 => x"b9c80854",
         11738 => x"84b9c808",
         11739 => x"802e81a3",
         11740 => x"3873ff2e",
         11741 => x"98388174",
         11742 => x"2782b438",
         11743 => x"7953739c",
         11744 => x"14082782",
         11745 => x"aa387398",
         11746 => x"160cffae",
         11747 => x"39810b91",
         11748 => x"16348153",
         11749 => x"7284b9c8",
         11750 => x"0c8b3d0d",
         11751 => x"04901533",
         11752 => x"70812a81",
         11753 => x"06555873",
         11754 => x"febb3875",
         11755 => x"94160855",
         11756 => x"57805876",
         11757 => x"782e0981",
         11758 => x"06feb638",
         11759 => x"7794160c",
         11760 => x"94150854",
         11761 => x"75742790",
         11762 => x"38738c16",
         11763 => x"0c901533",
         11764 => x"80c00757",
         11765 => x"76901634",
         11766 => x"7383ff06",
         11767 => x"5978802e",
         11768 => x"8c389c15",
         11769 => x"08782e85",
         11770 => x"38779c16",
         11771 => x"0c800b84",
         11772 => x"b9c80c8b",
         11773 => x"3d0d0480",
         11774 => x"0b94160c",
         11775 => x"88150854",
         11776 => x"73802e80",
         11777 => x"fe387398",
         11778 => x"160c7380",
         11779 => x"2e80c238",
         11780 => x"fea83984",
         11781 => x"b9c80857",
         11782 => x"94150817",
         11783 => x"94160c76",
         11784 => x"83ff0656",
         11785 => x"75802ea9",
         11786 => x"3879fe15",
         11787 => x"9c1208fe",
         11788 => x"055a5556",
         11789 => x"73782780",
         11790 => x"f6388a16",
         11791 => x"22747129",
         11792 => x"b0180805",
         11793 => x"78892a11",
         11794 => x"5a5a5378",
         11795 => x"802e80df",
         11796 => x"388c1508",
         11797 => x"56fee939",
         11798 => x"73527451",
         11799 => x"ff89b73f",
         11800 => x"84b9c808",
         11801 => x"54fe8a39",
         11802 => x"81143351",
         11803 => x"ff82a23f",
         11804 => x"84b9c808",
         11805 => x"81065372",
         11806 => x"fccf3872",
         11807 => x"75085456",
         11808 => x"fcc93973",
         11809 => x"527451ff",
         11810 => x"97cb3f84",
         11811 => x"b9c80854",
         11812 => x"84b9c808",
         11813 => x"812e9838",
         11814 => x"84b9c808",
         11815 => x"ff2efded",
         11816 => x"3884b9c8",
         11817 => x"0888160c",
         11818 => x"7398160c",
         11819 => x"fedc3982",
         11820 => x"0b911634",
         11821 => x"820b84b9",
         11822 => x"c80c8b3d",
         11823 => x"0d04f63d",
         11824 => x"0d7c5689",
         11825 => x"5475802e",
         11826 => x"a2388053",
         11827 => x"8c3dfc05",
         11828 => x"528d3d84",
         11829 => x"0551c59b",
         11830 => x"3f84b9c8",
         11831 => x"085584b9",
         11832 => x"c808802e",
         11833 => x"8f388076",
         11834 => x"0c745473",
         11835 => x"84b9c80c",
         11836 => x"8c3d0d04",
         11837 => x"7a760c7d",
         11838 => x"527551ff",
         11839 => x"b9973f84",
         11840 => x"b9c80855",
         11841 => x"84b9c808",
         11842 => x"80d138ab",
         11843 => x"16337098",
         11844 => x"2b595980",
         11845 => x"7824af38",
         11846 => x"86163370",
         11847 => x"842a8106",
         11848 => x"5b547980",
         11849 => x"2e80c538",
         11850 => x"9c16089b",
         11851 => x"11339a12",
         11852 => x"3371882b",
         11853 => x"077d7033",
         11854 => x"5d5d5a55",
         11855 => x"5778832e",
         11856 => x"b3387788",
         11857 => x"170c7a58",
         11858 => x"86182284",
         11859 => x"17237452",
         11860 => x"7551ff99",
         11861 => x"b93f84b9",
         11862 => x"c8085574",
         11863 => x"842e8d38",
         11864 => x"74802eff",
         11865 => x"84388076",
         11866 => x"0cfefe39",
         11867 => x"85558076",
         11868 => x"0cfef639",
         11869 => x"95173394",
         11870 => x"18337198",
         11871 => x"2b71902b",
         11872 => x"077a0788",
         11873 => x"190c5a5a",
         11874 => x"ffbc39fa",
         11875 => x"3d0d7855",
         11876 => x"89547480",
         11877 => x"2e9e3874",
         11878 => x"08537280",
         11879 => x"2e963872",
         11880 => x"33527180",
         11881 => x"2e8e3886",
         11882 => x"13228416",
         11883 => x"22575271",
         11884 => x"762e9438",
         11885 => x"80527157",
         11886 => x"73843873",
         11887 => x"750c7384",
         11888 => x"b9c80c88",
         11889 => x"3d0d0481",
         11890 => x"133351fe",
         11891 => x"ffc33f84",
         11892 => x"b9c80881",
         11893 => x"065271dc",
         11894 => x"38717508",
         11895 => x"5354d739",
         11896 => x"f83d0d7a",
         11897 => x"7c585589",
         11898 => x"5674802e",
         11899 => x"9f387408",
         11900 => x"5473802e",
         11901 => x"97387333",
         11902 => x"5372802e",
         11903 => x"8f388614",
         11904 => x"22841622",
         11905 => x"59537278",
         11906 => x"2e819738",
         11907 => x"80537259",
         11908 => x"75537580",
         11909 => x"c7387680",
         11910 => x"2e80f338",
         11911 => x"75527451",
         11912 => x"ff9dbd3f",
         11913 => x"84b9c808",
         11914 => x"5384b9c8",
         11915 => x"08842eb5",
         11916 => x"3884b9c8",
         11917 => x"08a63876",
         11918 => x"527451ff",
         11919 => x"b2923f72",
         11920 => x"527451ff",
         11921 => x"99be3f84",
         11922 => x"b9c80884",
         11923 => x"32703070",
         11924 => x"72079f2c",
         11925 => x"84b9c808",
         11926 => x"06555754",
         11927 => x"7284b9c8",
         11928 => x"0c8a3d0d",
         11929 => x"04757753",
         11930 => x"755253ff",
         11931 => x"b1e23f72",
         11932 => x"527451ff",
         11933 => x"998e3f84",
         11934 => x"b9c80884",
         11935 => x"32703070",
         11936 => x"72079f2c",
         11937 => x"84b9c808",
         11938 => x"06555754",
         11939 => x"cf397552",
         11940 => x"7451ff96",
         11941 => x"f93f84b9",
         11942 => x"c80884b9",
         11943 => x"c80c8a3d",
         11944 => x"0d048114",
         11945 => x"3351fefd",
         11946 => x"e83f84b9",
         11947 => x"c8088106",
         11948 => x"5372fed8",
         11949 => x"38727508",
         11950 => x"5456fed2",
         11951 => x"39ed3d0d",
         11952 => x"66578053",
         11953 => x"893d7053",
         11954 => x"973d5256",
         11955 => x"c1a53f84",
         11956 => x"b9c80855",
         11957 => x"84b9c808",
         11958 => x"802e8a38",
         11959 => x"7484b9c8",
         11960 => x"0c953d0d",
         11961 => x"04655275",
         11962 => x"51ffb5a9",
         11963 => x"3f84b9c8",
         11964 => x"085584b9",
         11965 => x"c808e538",
         11966 => x"0280cb05",
         11967 => x"3370982b",
         11968 => x"55588074",
         11969 => x"24973876",
         11970 => x"802ed138",
         11971 => x"76527551",
         11972 => x"ffb0bd3f",
         11973 => x"7484b9c8",
         11974 => x"0c953d0d",
         11975 => x"04860b84",
         11976 => x"b9c80c95",
         11977 => x"3d0d04ed",
         11978 => x"3d0d6668",
         11979 => x"565f8053",
         11980 => x"953dec05",
         11981 => x"52963d51",
         11982 => x"c0b93f84",
         11983 => x"b9c8085a",
         11984 => x"84b9c808",
         11985 => x"9a387f75",
         11986 => x"0c74089c",
         11987 => x"1108fe11",
         11988 => x"94130859",
         11989 => x"57595775",
         11990 => x"75268d38",
         11991 => x"757f0c79",
         11992 => x"84b9c80c",
         11993 => x"953d0d04",
         11994 => x"84b9c808",
         11995 => x"77335a5b",
         11996 => x"78812e82",
         11997 => x"933877a8",
         11998 => x"180884b9",
         11999 => x"c8085a5d",
         12000 => x"597780c1",
         12001 => x"387b811d",
         12002 => x"715c5d56",
         12003 => x"b4170876",
         12004 => x"2e82ef38",
         12005 => x"83173378",
         12006 => x"5f5d7c81",
         12007 => x"8d388154",
         12008 => x"7553b817",
         12009 => x"52811733",
         12010 => x"51fefcb7",
         12011 => x"3f84b9c8",
         12012 => x"08802e85",
         12013 => x"38ff5a81",
         12014 => x"5e79b418",
         12015 => x"0c7f7e5b",
         12016 => x"577d80cc",
         12017 => x"3876335e",
         12018 => x"7d822e82",
         12019 => x"8d387717",
         12020 => x"b8058311",
         12021 => x"33821233",
         12022 => x"71902b71",
         12023 => x"882b0781",
         12024 => x"14337072",
         12025 => x"07882b75",
         12026 => x"337180ff",
         12027 => x"fffe8006",
         12028 => x"07703070",
         12029 => x"80256305",
         12030 => x"60840583",
         12031 => x"ff0662ff",
         12032 => x"05434143",
         12033 => x"53545253",
         12034 => x"58405e56",
         12035 => x"78fef238",
         12036 => x"7a7f0c7a",
         12037 => x"94180c84",
         12038 => x"17338107",
         12039 => x"58778418",
         12040 => x"347984b9",
         12041 => x"c80c953d",
         12042 => x"0d048154",
         12043 => x"b4170853",
         12044 => x"b8177053",
         12045 => x"81183352",
         12046 => x"5dfefca6",
         12047 => x"3f815e84",
         12048 => x"b9c808fe",
         12049 => x"f83884b9",
         12050 => x"c8088318",
         12051 => x"34b41708",
         12052 => x"a8180831",
         12053 => x"84b9c808",
         12054 => x"5f5574a0",
         12055 => x"180827fe",
         12056 => x"bd388217",
         12057 => x"33557482",
         12058 => x"2e098106",
         12059 => x"feb03881",
         12060 => x"54b41708",
         12061 => x"a0180805",
         12062 => x"537c5281",
         12063 => x"173351fe",
         12064 => x"fbe03f77",
         12065 => x"5efe9739",
         12066 => x"82774292",
         12067 => x"3d595675",
         12068 => x"527751ff",
         12069 => x"81803f84",
         12070 => x"b9c808ff",
         12071 => x"2e80e838",
         12072 => x"84b9c808",
         12073 => x"812e80f7",
         12074 => x"3884b9c8",
         12075 => x"08307084",
         12076 => x"b9c80807",
         12077 => x"80257c05",
         12078 => x"8118625a",
         12079 => x"585c5c9c",
         12080 => x"17087626",
         12081 => x"ca387a7f",
         12082 => x"0c7a9418",
         12083 => x"0c841733",
         12084 => x"81075877",
         12085 => x"841834fe",
         12086 => x"c8397717",
         12087 => x"b8058111",
         12088 => x"33713371",
         12089 => x"882b0770",
         12090 => x"30708025",
         12091 => x"1f821d83",
         12092 => x"ff06ff1f",
         12093 => x"5f5d5f59",
         12094 => x"5f5f5578",
         12095 => x"fd8338fe",
         12096 => x"8f39775a",
         12097 => x"fdbf3981",
         12098 => x"60585a7a",
         12099 => x"7f0c7a94",
         12100 => x"180c8417",
         12101 => x"33810758",
         12102 => x"77841834",
         12103 => x"fe833982",
         12104 => x"60585ae7",
         12105 => x"39f73d0d",
         12106 => x"7b578956",
         12107 => x"76802e9f",
         12108 => x"38760855",
         12109 => x"74802e97",
         12110 => x"38743354",
         12111 => x"73802e8f",
         12112 => x"38861522",
         12113 => x"84182259",
         12114 => x"5978782e",
         12115 => x"81da3880",
         12116 => x"54735a75",
         12117 => x"80dc3891",
         12118 => x"17335675",
         12119 => x"80d43890",
         12120 => x"17337081",
         12121 => x"2a810655",
         12122 => x"58875573",
         12123 => x"802e80c4",
         12124 => x"38941708",
         12125 => x"54738c18",
         12126 => x"0827b738",
         12127 => x"7381d538",
         12128 => x"88170877",
         12129 => x"08575481",
         12130 => x"74278838",
         12131 => x"9c160874",
         12132 => x"26b33882",
         12133 => x"56800b88",
         12134 => x"180c9417",
         12135 => x"088c180c",
         12136 => x"7780c007",
         12137 => x"59789018",
         12138 => x"3475802e",
         12139 => x"85387591",
         12140 => x"18347555",
         12141 => x"7484b9c8",
         12142 => x"0c8b3d0d",
         12143 => x"04785478",
         12144 => x"782780ff",
         12145 => x"38735276",
         12146 => x"51fefeca",
         12147 => x"3f84b9c8",
         12148 => x"085984b9",
         12149 => x"c808802e",
         12150 => x"80e93884",
         12151 => x"b9c80881",
         12152 => x"2e82d838",
         12153 => x"84b9c808",
         12154 => x"ff2e82e5",
         12155 => x"38805373",
         12156 => x"527551ff",
         12157 => x"85813f84",
         12158 => x"b9c80882",
         12159 => x"c8389c16",
         12160 => x"08fe1194",
         12161 => x"18085755",
         12162 => x"58747427",
         12163 => x"ffaf3881",
         12164 => x"1594170c",
         12165 => x"84163381",
         12166 => x"07547384",
         12167 => x"17347854",
         12168 => x"777926ff",
         12169 => x"a0389c39",
         12170 => x"81153351",
         12171 => x"fef6e23f",
         12172 => x"84b9c808",
         12173 => x"81065473",
         12174 => x"fe953873",
         12175 => x"77085556",
         12176 => x"fe8f3980",
         12177 => x"0b901833",
         12178 => x"59547356",
         12179 => x"800b8818",
         12180 => x"0cfec739",
         12181 => x"98170852",
         12182 => x"7651fefd",
         12183 => x"b93f84b9",
         12184 => x"c808ff2e",
         12185 => x"81c23884",
         12186 => x"b9c80881",
         12187 => x"2e81be38",
         12188 => x"7581ae38",
         12189 => x"795884b9",
         12190 => x"c8089c19",
         12191 => x"082781a1",
         12192 => x"3884b9c8",
         12193 => x"08981808",
         12194 => x"78085856",
         12195 => x"54810b84",
         12196 => x"b9c80827",
         12197 => x"81a13884",
         12198 => x"b9c8089c",
         12199 => x"17082781",
         12200 => x"96387480",
         12201 => x"2e9738ff",
         12202 => x"53745275",
         12203 => x"51ff83c7",
         12204 => x"3f84b9c8",
         12205 => x"085584b9",
         12206 => x"c80880e3",
         12207 => x"38735276",
         12208 => x"51fefcd2",
         12209 => x"3f84b9c8",
         12210 => x"085984b9",
         12211 => x"c808802e",
         12212 => x"80cb3884",
         12213 => x"b9c80881",
         12214 => x"2e80dc38",
         12215 => x"84b9c808",
         12216 => x"ff2e80fe",
         12217 => x"38805373",
         12218 => x"527551ff",
         12219 => x"83893f84",
         12220 => x"b9c80880",
         12221 => x"e6389c16",
         12222 => x"08fe1194",
         12223 => x"18085755",
         12224 => x"58747427",
         12225 => x"90388115",
         12226 => x"94170c84",
         12227 => x"16338107",
         12228 => x"54738417",
         12229 => x"34785477",
         12230 => x"7926ffa1",
         12231 => x"38805574",
         12232 => x"56901733",
         12233 => x"58fcf339",
         12234 => x"8156febb",
         12235 => x"39820b90",
         12236 => x"18335956",
         12237 => x"fce43982",
         12238 => x"56e73982",
         12239 => x"0b901833",
         12240 => x"5954fe86",
         12241 => x"3984b9c8",
         12242 => x"08901833",
         12243 => x"5954fdfa",
         12244 => x"39810b90",
         12245 => x"18335954",
         12246 => x"fdf03984",
         12247 => x"b9c80856",
         12248 => x"c0398156",
         12249 => x"ffbb39db",
         12250 => x"3d0d8253",
         12251 => x"a73dff9c",
         12252 => x"0552a83d",
         12253 => x"51ffb7fb",
         12254 => x"3f84b9c8",
         12255 => x"085684b9",
         12256 => x"c808802e",
         12257 => x"8a387584",
         12258 => x"b9c80ca7",
         12259 => x"3d0d047d",
         12260 => x"4ba83d08",
         12261 => x"529b3d70",
         12262 => x"5259ffab",
         12263 => x"f83f84b9",
         12264 => x"c8085684",
         12265 => x"b9c808de",
         12266 => x"38028193",
         12267 => x"05337085",
         12268 => x"2a810659",
         12269 => x"57865677",
         12270 => x"cd387698",
         12271 => x"2b5b807b",
         12272 => x"24c43802",
         12273 => x"80ee0533",
         12274 => x"7081065d",
         12275 => x"5787567b",
         12276 => x"ffb4387d",
         12277 => x"a33d089b",
         12278 => x"11339a12",
         12279 => x"3371882b",
         12280 => x"07733341",
         12281 => x"5e5c5758",
         12282 => x"7c832e80",
         12283 => x"d5387684",
         12284 => x"2a810657",
         12285 => x"76802e80",
         12286 => x"ed388756",
         12287 => x"9818087b",
         12288 => x"2eff8338",
         12289 => x"775f7a41",
         12290 => x"84b9c808",
         12291 => x"528f3d70",
         12292 => x"5255ff8b",
         12293 => x"f93f84b9",
         12294 => x"c8085684",
         12295 => x"b9c808fe",
         12296 => x"e53884b9",
         12297 => x"c8085274",
         12298 => x"51ff91b4",
         12299 => x"3f84b9c8",
         12300 => x"085684b9",
         12301 => x"c808a038",
         12302 => x"870b84b9",
         12303 => x"c80ca73d",
         12304 => x"0d049516",
         12305 => x"33941733",
         12306 => x"71982b71",
         12307 => x"902b077d",
         12308 => x"075d5d5d",
         12309 => x"ff983984",
         12310 => x"b9c80884",
         12311 => x"2e883884",
         12312 => x"b9c808fe",
         12313 => x"a1387808",
         12314 => x"6fa83d08",
         12315 => x"575d5774",
         12316 => x"ff2e80d3",
         12317 => x"38745278",
         12318 => x"51ff8b92",
         12319 => x"3f84b9c8",
         12320 => x"085684b9",
         12321 => x"c808802e",
         12322 => x"be387530",
         12323 => x"70770780",
         12324 => x"25565a7a",
         12325 => x"802e9a38",
         12326 => x"74802e95",
         12327 => x"387a7908",
         12328 => x"5855817b",
         12329 => x"2789389c",
         12330 => x"17087b26",
         12331 => x"81fd3882",
         12332 => x"5675fdd2",
         12333 => x"387d51fe",
         12334 => x"f5db3f84",
         12335 => x"b9c80884",
         12336 => x"b9c80ca7",
         12337 => x"3d0d04b8",
         12338 => x"175d9819",
         12339 => x"0856805a",
         12340 => x"b4170876",
         12341 => x"2e82b938",
         12342 => x"8317337a",
         12343 => x"5955747a",
         12344 => x"2e098106",
         12345 => x"80dd3881",
         12346 => x"547553b8",
         12347 => x"17528117",
         12348 => x"3351fef1",
         12349 => x"ee3f84b9",
         12350 => x"c808802e",
         12351 => x"8538ff56",
         12352 => x"815875b4",
         12353 => x"180c7756",
         12354 => x"77ab389c",
         12355 => x"190858e5",
         12356 => x"7834810b",
         12357 => x"83183490",
         12358 => x"19087c27",
         12359 => x"feec3880",
         12360 => x"527851ff",
         12361 => x"8bde3f84",
         12362 => x"b9c80856",
         12363 => x"84b9c808",
         12364 => x"802eff96",
         12365 => x"3875842e",
         12366 => x"098106fe",
         12367 => x"cd388256",
         12368 => x"fec83981",
         12369 => x"54b41708",
         12370 => x"537c5281",
         12371 => x"173351fe",
         12372 => x"f2903f81",
         12373 => x"5884b9c8",
         12374 => x"087a2e09",
         12375 => x"8106ffa6",
         12376 => x"3884b9c8",
         12377 => x"08831834",
         12378 => x"b41708a8",
         12379 => x"18083184",
         12380 => x"b9c80859",
         12381 => x"5574a018",
         12382 => x"0827feeb",
         12383 => x"38821733",
         12384 => x"5574822e",
         12385 => x"098106fe",
         12386 => x"de388154",
         12387 => x"b41708a0",
         12388 => x"18080553",
         12389 => x"7c528117",
         12390 => x"3351fef1",
         12391 => x"c53f7958",
         12392 => x"fec53979",
         12393 => x"55797827",
         12394 => x"80e13874",
         12395 => x"527851fe",
         12396 => x"f6e43f84",
         12397 => x"b9c8085a",
         12398 => x"84b9c808",
         12399 => x"802e80cb",
         12400 => x"3884b9c8",
         12401 => x"08812efd",
         12402 => x"e63884b9",
         12403 => x"c808ff2e",
         12404 => x"80cb3880",
         12405 => x"53745276",
         12406 => x"51fefd9b",
         12407 => x"3f84b9c8",
         12408 => x"08b3389c",
         12409 => x"1708fe11",
         12410 => x"94190858",
         12411 => x"5c58757b",
         12412 => x"27ffb038",
         12413 => x"81169418",
         12414 => x"0c841733",
         12415 => x"81075c7b",
         12416 => x"84183479",
         12417 => x"55777a26",
         12418 => x"ffa13880",
         12419 => x"56fda239",
         12420 => x"7956fdf7",
         12421 => x"3984b9c8",
         12422 => x"0856fd95",
         12423 => x"398156fd",
         12424 => x"9039e33d",
         12425 => x"0d82539f",
         12426 => x"3dffbc05",
         12427 => x"52a03d51",
         12428 => x"ffb2c03f",
         12429 => x"84b9c808",
         12430 => x"5684b9c8",
         12431 => x"08802e8a",
         12432 => x"387584b9",
         12433 => x"c80c9f3d",
         12434 => x"0d047d43",
         12435 => x"6f52933d",
         12436 => x"70525aff",
         12437 => x"a6bf3f84",
         12438 => x"b9c80856",
         12439 => x"84b9c808",
         12440 => x"8b38880b",
         12441 => x"84b9c80c",
         12442 => x"9f3d0d04",
         12443 => x"84b9c808",
         12444 => x"842e0981",
         12445 => x"06cb3802",
         12446 => x"80f30533",
         12447 => x"70852a81",
         12448 => x"06565886",
         12449 => x"5674ffb9",
         12450 => x"387d5f74",
         12451 => x"528f3d70",
         12452 => x"525dff83",
         12453 => x"c03f84b9",
         12454 => x"c8087557",
         12455 => x"5c84b9c8",
         12456 => x"08833887",
         12457 => x"5684b9c8",
         12458 => x"08812e80",
         12459 => x"f93884b9",
         12460 => x"c808ff2e",
         12461 => x"81cb3875",
         12462 => x"81c9387d",
         12463 => x"84b9c808",
         12464 => x"8312335d",
         12465 => x"5a577a80",
         12466 => x"e238fe19",
         12467 => x"9c1808fe",
         12468 => x"055a5680",
         12469 => x"5b757927",
         12470 => x"8d388a17",
         12471 => x"22767129",
         12472 => x"b0190805",
         12473 => x"5c587ab4",
         12474 => x"180cb817",
         12475 => x"59848079",
         12476 => x"57558076",
         12477 => x"70810558",
         12478 => x"34ff1555",
         12479 => x"74f43874",
         12480 => x"588a1722",
         12481 => x"55777527",
         12482 => x"81f93881",
         12483 => x"54771b53",
         12484 => x"78528117",
         12485 => x"3351feee",
         12486 => x"c93f84b9",
         12487 => x"c80881df",
         12488 => x"38811858",
         12489 => x"dc398256",
         12490 => x"ff843981",
         12491 => x"54b41708",
         12492 => x"53b81770",
         12493 => x"53811833",
         12494 => x"5258feee",
         12495 => x"a53f8156",
         12496 => x"84b9c808",
         12497 => x"be3884b9",
         12498 => x"c8088318",
         12499 => x"34b41708",
         12500 => x"a8180831",
         12501 => x"5574a018",
         12502 => x"0827feee",
         12503 => x"38821733",
         12504 => x"5b7a822e",
         12505 => x"098106fe",
         12506 => x"e1387554",
         12507 => x"b41708a0",
         12508 => x"18080553",
         12509 => x"77528117",
         12510 => x"3351feed",
         12511 => x"e53ffeca",
         12512 => x"3981567b",
         12513 => x"7d085855",
         12514 => x"817c27fd",
         12515 => x"b4387b9c",
         12516 => x"180827fd",
         12517 => x"ac387452",
         12518 => x"7c51fef2",
         12519 => x"f93f84b9",
         12520 => x"c8085a84",
         12521 => x"b9c80880",
         12522 => x"2efd9638",
         12523 => x"84b9c808",
         12524 => x"812efd8d",
         12525 => x"3884b9c8",
         12526 => x"08ff2efd",
         12527 => x"84388053",
         12528 => x"74527651",
         12529 => x"fef9b03f",
         12530 => x"84b9c808",
         12531 => x"fcf3389c",
         12532 => x"1708fe11",
         12533 => x"9419085a",
         12534 => x"5c59777b",
         12535 => x"27903881",
         12536 => x"1894180c",
         12537 => x"84173381",
         12538 => x"075c7b84",
         12539 => x"18347955",
         12540 => x"787a26ff",
         12541 => x"a1387584",
         12542 => x"b9c80c9f",
         12543 => x"3d0d048a",
         12544 => x"17225574",
         12545 => x"83ffff06",
         12546 => x"57815676",
         12547 => x"782e0981",
         12548 => x"06fef038",
         12549 => x"8b0bb81f",
         12550 => x"5656a075",
         12551 => x"70810557",
         12552 => x"34ff1656",
         12553 => x"75f4387d",
         12554 => x"57ae0bb8",
         12555 => x"18347d58",
         12556 => x"900b80c3",
         12557 => x"19347d59",
         12558 => x"7580ce1a",
         12559 => x"347580cf",
         12560 => x"1a34a10b",
         12561 => x"80d01a34",
         12562 => x"80cc0b80",
         12563 => x"d11a347d",
         12564 => x"7c83ffff",
         12565 => x"06595677",
         12566 => x"80d21734",
         12567 => x"77882a5b",
         12568 => x"7a80d317",
         12569 => x"34753355",
         12570 => x"74832e81",
         12571 => x"cc387d59",
         12572 => x"a00b80d8",
         12573 => x"1ab81b57",
         12574 => x"58567470",
         12575 => x"81055633",
         12576 => x"77708105",
         12577 => x"5934ff16",
         12578 => x"5675ef38",
         12579 => x"7d56ae0b",
         12580 => x"80d91734",
         12581 => x"647e7183",
         12582 => x"ffff065b",
         12583 => x"57577880",
         12584 => x"f2173478",
         12585 => x"882a5b7a",
         12586 => x"80f31734",
         12587 => x"75335574",
         12588 => x"832e80f0",
         12589 => x"387d5b81",
         12590 => x"0b831c34",
         12591 => x"7951ff92",
         12592 => x"963f84b9",
         12593 => x"c8085684",
         12594 => x"b9c808fd",
         12595 => x"b6386956",
         12596 => x"84b9c808",
         12597 => x"96173484",
         12598 => x"b9c80897",
         12599 => x"1734a10b",
         12600 => x"98173480",
         12601 => x"cc0b9917",
         12602 => x"347d6a58",
         12603 => x"5d779a18",
         12604 => x"3477882a",
         12605 => x"59789b18",
         12606 => x"347c335a",
         12607 => x"79832e80",
         12608 => x"d9386955",
         12609 => x"900b8b16",
         12610 => x"347d5781",
         12611 => x"0b831834",
         12612 => x"7d51feed",
         12613 => x"803f84b9",
         12614 => x"c8085675",
         12615 => x"84b9c80c",
         12616 => x"9f3d0d04",
         12617 => x"76902a55",
         12618 => x"7480ec17",
         12619 => x"3474882a",
         12620 => x"577680ed",
         12621 => x"1734fefd",
         12622 => x"397b902a",
         12623 => x"5b7a80cc",
         12624 => x"17347a88",
         12625 => x"2a557480",
         12626 => x"cd17347d",
         12627 => x"59a00b80",
         12628 => x"d81ab81b",
         12629 => x"575856fe",
         12630 => x"a1397b90",
         12631 => x"2a587794",
         12632 => x"18347788",
         12633 => x"2a5c7b95",
         12634 => x"18346955",
         12635 => x"900b8b16",
         12636 => x"347d5781",
         12637 => x"0b831834",
         12638 => x"7d51feec",
         12639 => x"983f84b9",
         12640 => x"c80856ff",
         12641 => x"9639d13d",
         12642 => x"0db33db4",
         12643 => x"3d087059",
         12644 => x"5b5f7980",
         12645 => x"2e9b3879",
         12646 => x"7081055b",
         12647 => x"33709f26",
         12648 => x"565675ba",
         12649 => x"2e81b838",
         12650 => x"74ed3875",
         12651 => x"ba2e81af",
         12652 => x"388253b1",
         12653 => x"3dfefc05",
         12654 => x"52b23d51",
         12655 => x"ffabb43f",
         12656 => x"84b9c808",
         12657 => x"5684b9c8",
         12658 => x"08802e8a",
         12659 => x"387584b9",
         12660 => x"c80cb13d",
         12661 => x"0d047fa6",
         12662 => x"3d0cb23d",
         12663 => x"0852a53d",
         12664 => x"705259ff",
         12665 => x"9faf3f84",
         12666 => x"b9c80856",
         12667 => x"84b9c808",
         12668 => x"dc380281",
         12669 => x"bb053381",
         12670 => x"a0065d86",
         12671 => x"567cce38",
         12672 => x"a00b923d",
         12673 => x"ae3d0858",
         12674 => x"58557570",
         12675 => x"81055733",
         12676 => x"77708105",
         12677 => x"5934ff15",
         12678 => x"5574ef38",
         12679 => x"993d58b0",
         12680 => x"787a5858",
         12681 => x"55757081",
         12682 => x"05573377",
         12683 => x"70810559",
         12684 => x"34ff1555",
         12685 => x"74ef38b3",
         12686 => x"3d085277",
         12687 => x"51ff9ed5",
         12688 => x"3f84b9c8",
         12689 => x"085684b9",
         12690 => x"c80885d8",
         12691 => x"386aa83d",
         12692 => x"082e81cb",
         12693 => x"38880b84",
         12694 => x"b9c80cb1",
         12695 => x"3d0d0476",
         12696 => x"33d01170",
         12697 => x"81ff0657",
         12698 => x"57587489",
         12699 => x"26913882",
         12700 => x"177881ff",
         12701 => x"06d0055d",
         12702 => x"59787a2e",
         12703 => x"80fa3880",
         12704 => x"7f0883e5",
         12705 => x"b8700872",
         12706 => x"5d5e5f5f",
         12707 => x"5c7a7081",
         12708 => x"055c3379",
         12709 => x"7081055b",
         12710 => x"33ff9f12",
         12711 => x"5a585677",
         12712 => x"99268938",
         12713 => x"e0167081",
         12714 => x"ff065755",
         12715 => x"ff9f1758",
         12716 => x"77992689",
         12717 => x"38e01770",
         12718 => x"81ff0658",
         12719 => x"55753070",
         12720 => x"9f2a5955",
         12721 => x"75772e09",
         12722 => x"81068538",
         12723 => x"77ffbe38",
         12724 => x"787a3270",
         12725 => x"30707207",
         12726 => x"9f2a7a07",
         12727 => x"5d58557a",
         12728 => x"802e9538",
         12729 => x"811c841e",
         12730 => x"5e5c7b83",
         12731 => x"24fdc238",
         12732 => x"7c087e5a",
         12733 => x"5bff9639",
         12734 => x"7b8324fd",
         12735 => x"b438797f",
         12736 => x"0c8253b1",
         12737 => x"3dfefc05",
         12738 => x"52b23d51",
         12739 => x"ffa8e43f",
         12740 => x"84b9c808",
         12741 => x"5684b9c8",
         12742 => x"08fdb238",
         12743 => x"fdb8396c",
         12744 => x"aa3d082e",
         12745 => x"098106fe",
         12746 => x"ac387751",
         12747 => x"ff8da83f",
         12748 => x"84b9c808",
         12749 => x"5684b9c8",
         12750 => x"08fd9238",
         12751 => x"6f58930b",
         12752 => x"8d190288",
         12753 => x"0580cd05",
         12754 => x"58565a75",
         12755 => x"70810557",
         12756 => x"33757081",
         12757 => x"055734ff",
         12758 => x"1a5a79ef",
         12759 => x"380280cb",
         12760 => x"05338b19",
         12761 => x"348b1833",
         12762 => x"70842a81",
         12763 => x"0640567e",
         12764 => x"893875a0",
         12765 => x"0757768b",
         12766 => x"19347f5d",
         12767 => x"810b831e",
         12768 => x"348b1833",
         12769 => x"70842a81",
         12770 => x"06575c75",
         12771 => x"802e81c5",
         12772 => x"38a73d08",
         12773 => x"6b2e81bd",
         12774 => x"387f9b19",
         12775 => x"339a1a33",
         12776 => x"71882b07",
         12777 => x"72334158",
         12778 => x"5c577d83",
         12779 => x"2e82e038",
         12780 => x"fe169c18",
         12781 => x"08fe055e",
         12782 => x"56757d27",
         12783 => x"82c7388a",
         12784 => x"17227671",
         12785 => x"29b01908",
         12786 => x"05575e75",
         12787 => x"802e82b5",
         12788 => x"38757a5d",
         12789 => x"58b41708",
         12790 => x"762eaa38",
         12791 => x"8317335f",
         12792 => x"7e83bc38",
         12793 => x"81547553",
         12794 => x"b8175281",
         12795 => x"173351fe",
         12796 => x"e3f13f84",
         12797 => x"b9c80880",
         12798 => x"2e8538ff",
         12799 => x"58815c77",
         12800 => x"b4180c7f",
         12801 => x"577b80d8",
         12802 => x"1856567b",
         12803 => x"fbbf3881",
         12804 => x"15335a79",
         12805 => x"ae2e0981",
         12806 => x"06bb386a",
         12807 => x"7083ffff",
         12808 => x"065d567b",
         12809 => x"80f21834",
         12810 => x"7b882a58",
         12811 => x"7780f318",
         12812 => x"3476335b",
         12813 => x"7a832e09",
         12814 => x"81069338",
         12815 => x"75902a5e",
         12816 => x"7d80ec18",
         12817 => x"347d882a",
         12818 => x"567580ed",
         12819 => x"18347f57",
         12820 => x"810b8318",
         12821 => x"347808aa",
         12822 => x"3d08b23d",
         12823 => x"08575c56",
         12824 => x"74ff2e95",
         12825 => x"38745278",
         12826 => x"51fefba2",
         12827 => x"3f84b9c8",
         12828 => x"085584b9",
         12829 => x"c80880f5",
         12830 => x"38b8165c",
         12831 => x"98190857",
         12832 => x"805ab416",
         12833 => x"08772eb4",
         12834 => x"38831633",
         12835 => x"7a595f7e",
         12836 => x"7a2e0981",
         12837 => x"0681a838",
         12838 => x"81547653",
         12839 => x"b8165281",
         12840 => x"163351fe",
         12841 => x"e2bd3f84",
         12842 => x"b9c80880",
         12843 => x"2e8538ff",
         12844 => x"57815876",
         12845 => x"b4170c77",
         12846 => x"5577aa38",
         12847 => x"9c19085a",
         12848 => x"e57a3481",
         12849 => x"0b831734",
         12850 => x"9019087b",
         12851 => x"27a53880",
         12852 => x"527851fe",
         12853 => x"fcae3f84",
         12854 => x"b9c80855",
         12855 => x"84b9c808",
         12856 => x"802eff98",
         12857 => x"38825674",
         12858 => x"842ef9e1",
         12859 => x"38745674",
         12860 => x"f9db387f",
         12861 => x"51fee59d",
         12862 => x"3f84b9c8",
         12863 => x"0884b9c8",
         12864 => x"0cb13d0d",
         12865 => x"04820b84",
         12866 => x"b9c80cb1",
         12867 => x"3d0d0495",
         12868 => x"18339419",
         12869 => x"3371982b",
         12870 => x"71902b07",
         12871 => x"78075856",
         12872 => x"5cfd8d39",
         12873 => x"84b9c808",
         12874 => x"842efbfe",
         12875 => x"3884b9c8",
         12876 => x"08802efe",
         12877 => x"a0387584",
         12878 => x"b9c80cb1",
         12879 => x"3d0d0481",
         12880 => x"54b41608",
         12881 => x"537b5281",
         12882 => x"163351fe",
         12883 => x"e2943f81",
         12884 => x"5884b9c8",
         12885 => x"087a2e09",
         12886 => x"8106fedb",
         12887 => x"3884b9c8",
         12888 => x"08831734",
         12889 => x"b41608a8",
         12890 => x"17083184",
         12891 => x"b9c80859",
         12892 => x"5574a017",
         12893 => x"0827fea0",
         12894 => x"38821633",
         12895 => x"5d7c822e",
         12896 => x"098106fe",
         12897 => x"93388154",
         12898 => x"b41608a0",
         12899 => x"17080553",
         12900 => x"7b528116",
         12901 => x"3351fee1",
         12902 => x"c93f7958",
         12903 => x"fdfa3981",
         12904 => x"54b41708",
         12905 => x"53b81770",
         12906 => x"53811833",
         12907 => x"525bfee1",
         12908 => x"b13f815c",
         12909 => x"84b9c808",
         12910 => x"fcc93884",
         12911 => x"b9c80883",
         12912 => x"1834b417",
         12913 => x"08a81808",
         12914 => x"3184b9c8",
         12915 => x"085d5574",
         12916 => x"a0180827",
         12917 => x"fc8e3882",
         12918 => x"17335d7c",
         12919 => x"822e0981",
         12920 => x"06fc8138",
         12921 => x"8154b417",
         12922 => x"08a01808",
         12923 => x"05537a52",
         12924 => x"81173351",
         12925 => x"fee0eb3f",
         12926 => x"795cfbe8",
         12927 => x"39ec3d0d",
         12928 => x"0280df05",
         12929 => x"33028405",
         12930 => x"80e30533",
         12931 => x"56578253",
         12932 => x"963dcc05",
         12933 => x"52973d51",
         12934 => x"ffa2d83f",
         12935 => x"84b9c808",
         12936 => x"5684b9c8",
         12937 => x"08802e8a",
         12938 => x"387584b9",
         12939 => x"c80c963d",
         12940 => x"0d04785a",
         12941 => x"6652963d",
         12942 => x"d00551ff",
         12943 => x"96d73f84",
         12944 => x"b9c80856",
         12945 => x"84b9c808",
         12946 => x"e0380280",
         12947 => x"cf053381",
         12948 => x"a0065486",
         12949 => x"5673d238",
         12950 => x"74a70661",
         12951 => x"71098b12",
         12952 => x"3371067a",
         12953 => x"74060751",
         12954 => x"56575573",
         12955 => x"8b173478",
         12956 => x"55810b83",
         12957 => x"16347851",
         12958 => x"fee29a3f",
         12959 => x"84b9c808",
         12960 => x"84b9c80c",
         12961 => x"963d0d04",
         12962 => x"ec3d0d67",
         12963 => x"57825396",
         12964 => x"3dcc0552",
         12965 => x"973d51ff",
         12966 => x"a1d93f84",
         12967 => x"b9c80855",
         12968 => x"84b9c808",
         12969 => x"802e8a38",
         12970 => x"7484b9c8",
         12971 => x"0c963d0d",
         12972 => x"04785a66",
         12973 => x"52963dd0",
         12974 => x"0551ff95",
         12975 => x"d83f84b9",
         12976 => x"c8085584",
         12977 => x"b9c808e0",
         12978 => x"380280cf",
         12979 => x"053381a0",
         12980 => x"06568655",
         12981 => x"75d23860",
         12982 => x"84182286",
         12983 => x"19227190",
         12984 => x"2b075959",
         12985 => x"56769617",
         12986 => x"3476882a",
         12987 => x"55749717",
         12988 => x"3476902a",
         12989 => x"58779817",
         12990 => x"3476982a",
         12991 => x"54739917",
         12992 => x"34785781",
         12993 => x"0b831834",
         12994 => x"7851fee1",
         12995 => x"883f84b9",
         12996 => x"c80884b9",
         12997 => x"c80c963d",
         12998 => x"0d04e83d",
         12999 => x"0d6b6d5d",
         13000 => x"5b80539a",
         13001 => x"3dcc0552",
         13002 => x"9b3d51ff",
         13003 => x"a0c53f84",
         13004 => x"b9c80884",
         13005 => x"b9c80830",
         13006 => x"7084b9c8",
         13007 => x"08078025",
         13008 => x"5156577a",
         13009 => x"802e8b38",
         13010 => x"81707606",
         13011 => x"5a567881",
         13012 => x"a4387630",
         13013 => x"70780780",
         13014 => x"25565b7b",
         13015 => x"802e818c",
         13016 => x"38817076",
         13017 => x"065a5878",
         13018 => x"802e8180",
         13019 => x"387ca411",
         13020 => x"08585680",
         13021 => x"5ab41608",
         13022 => x"772e82f6",
         13023 => x"38831633",
         13024 => x"7a5a5574",
         13025 => x"7a2e0981",
         13026 => x"06819838",
         13027 => x"81547653",
         13028 => x"b8165281",
         13029 => x"163351fe",
         13030 => x"dcc93f84",
         13031 => x"b9c80880",
         13032 => x"2e8538ff",
         13033 => x"57815976",
         13034 => x"b4170c78",
         13035 => x"5778bd38",
         13036 => x"7c703356",
         13037 => x"5880c356",
         13038 => x"74832e8b",
         13039 => x"3880e456",
         13040 => x"74842e83",
         13041 => x"38a75675",
         13042 => x"18b80583",
         13043 => x"11338212",
         13044 => x"3371902b",
         13045 => x"71882b07",
         13046 => x"81143370",
         13047 => x"7207882b",
         13048 => x"75337107",
         13049 => x"620c5f5d",
         13050 => x"5e575956",
         13051 => x"7684b9c8",
         13052 => x"0c9a3d0d",
         13053 => x"047c5e80",
         13054 => x"4080528e",
         13055 => x"3d705255",
         13056 => x"fef48b3f",
         13057 => x"84b9c808",
         13058 => x"5784b9c8",
         13059 => x"08802e81",
         13060 => x"8d387684",
         13061 => x"2e098106",
         13062 => x"feb83880",
         13063 => x"7b348057",
         13064 => x"feb03977",
         13065 => x"54b41608",
         13066 => x"53b81670",
         13067 => x"53811733",
         13068 => x"525bfedc",
         13069 => x"ad3f7759",
         13070 => x"84b9c808",
         13071 => x"7a2e0981",
         13072 => x"06fee838",
         13073 => x"84b9c808",
         13074 => x"831734b4",
         13075 => x"1608a817",
         13076 => x"083184b9",
         13077 => x"c8085a55",
         13078 => x"74a01708",
         13079 => x"27fead38",
         13080 => x"82163355",
         13081 => x"74822e09",
         13082 => x"8106fea0",
         13083 => x"387754b4",
         13084 => x"1608a017",
         13085 => x"0805537a",
         13086 => x"52811633",
         13087 => x"51fedbe2",
         13088 => x"3f795981",
         13089 => x"547653b8",
         13090 => x"16528116",
         13091 => x"3351feda",
         13092 => x"d23f84b9",
         13093 => x"c808802e",
         13094 => x"fe8d38fe",
         13095 => x"86397552",
         13096 => x"7451fef8",
         13097 => x"bb3f84b9",
         13098 => x"c8085784",
         13099 => x"b9c808fe",
         13100 => x"e13884b9",
         13101 => x"c80884b9",
         13102 => x"c808665c",
         13103 => x"59597918",
         13104 => x"81197c1b",
         13105 => x"57595675",
         13106 => x"33753481",
         13107 => x"19598a78",
         13108 => x"27ec388b",
         13109 => x"701c5758",
         13110 => x"80763477",
         13111 => x"802efcf2",
         13112 => x"38ff187b",
         13113 => x"1170335c",
         13114 => x"575879a0",
         13115 => x"2eea38fc",
         13116 => x"e1397957",
         13117 => x"fdba39e1",
         13118 => x"3d0d8253",
         13119 => x"a13dffb4",
         13120 => x"0552a23d",
         13121 => x"51ff9ceb",
         13122 => x"3f84b9c8",
         13123 => x"085684b9",
         13124 => x"c80882a6",
         13125 => x"388f3d5d",
         13126 => x"8b7d5755",
         13127 => x"a0767081",
         13128 => x"055834ff",
         13129 => x"155574f4",
         13130 => x"3874a33d",
         13131 => x"08703370",
         13132 => x"81ff065b",
         13133 => x"58585a9f",
         13134 => x"782781b7",
         13135 => x"38a23d90",
         13136 => x"3d5c5c75",
         13137 => x"81ff0681",
         13138 => x"18575574",
         13139 => x"81f53875",
         13140 => x"7c0c7483",
         13141 => x"ffff2681",
         13142 => x"ff387451",
         13143 => x"a1953f83",
         13144 => x"b55284b9",
         13145 => x"c808519f",
         13146 => x"dc3f84b9",
         13147 => x"c80883ff",
         13148 => x"ff065776",
         13149 => x"802e81e0",
         13150 => x"3883e6d8",
         13151 => x"0b83e6d8",
         13152 => x"337081ff",
         13153 => x"065b5658",
         13154 => x"78802e81",
         13155 => x"d6387456",
         13156 => x"78772e99",
         13157 => x"38811870",
         13158 => x"337081ff",
         13159 => x"06575758",
         13160 => x"74802e89",
         13161 => x"3874772e",
         13162 => x"098106e9",
         13163 => x"387581ff",
         13164 => x"06597881",
         13165 => x"a33881ff",
         13166 => x"772781f8",
         13167 => x"38798926",
         13168 => x"81963881",
         13169 => x"ff77278f",
         13170 => x"3876882a",
         13171 => x"55747b70",
         13172 => x"81055d34",
         13173 => x"811a5a76",
         13174 => x"7b708105",
         13175 => x"5d34811a",
         13176 => x"a33d0870",
         13177 => x"337081ff",
         13178 => x"065b5858",
         13179 => x"5a779f26",
         13180 => x"fed1388f",
         13181 => x"3d335786",
         13182 => x"567681e5",
         13183 => x"2ebc3879",
         13184 => x"802e9938",
         13185 => x"02b70556",
         13186 => x"79167033",
         13187 => x"5c5c7aa0",
         13188 => x"2e098106",
         13189 => x"8738ff1a",
         13190 => x"5a79ed38",
         13191 => x"7d458047",
         13192 => x"8052953d",
         13193 => x"705256fe",
         13194 => x"efe43f84",
         13195 => x"b9c80855",
         13196 => x"84b9c808",
         13197 => x"802eb438",
         13198 => x"74567584",
         13199 => x"b9c80ca1",
         13200 => x"3d0d0483",
         13201 => x"b5527451",
         13202 => x"9ee73f84",
         13203 => x"b9c80883",
         13204 => x"ffff0655",
         13205 => x"74fdf838",
         13206 => x"86567584",
         13207 => x"b9c80ca1",
         13208 => x"3d0d0483",
         13209 => x"e6d83356",
         13210 => x"fec33981",
         13211 => x"527551fe",
         13212 => x"f4ee3f84",
         13213 => x"b9c80855",
         13214 => x"84b9c808",
         13215 => x"80c13879",
         13216 => x"802e82c4",
         13217 => x"388b6c7e",
         13218 => x"59575576",
         13219 => x"70810558",
         13220 => x"33767081",
         13221 => x"055834ff",
         13222 => x"155574ef",
         13223 => x"387d5d81",
         13224 => x"0b831e34",
         13225 => x"7d51fed9",
         13226 => x"ec3f84b9",
         13227 => x"c8085574",
         13228 => x"56ff8739",
         13229 => x"8a7a27fe",
         13230 => x"8a388656",
         13231 => x"ff9c3984",
         13232 => x"b9c80884",
         13233 => x"2e098106",
         13234 => x"feee3880",
         13235 => x"5579752e",
         13236 => x"fee63875",
         13237 => x"08755376",
         13238 => x"5258feee",
         13239 => x"b13f84b9",
         13240 => x"c8085784",
         13241 => x"b9c80875",
         13242 => x"2e098106",
         13243 => x"81843884",
         13244 => x"b9c808b8",
         13245 => x"195c5a98",
         13246 => x"16085780",
         13247 => x"59b41808",
         13248 => x"772eb238",
         13249 => x"83183355",
         13250 => x"74792e09",
         13251 => x"810681d7",
         13252 => x"38815476",
         13253 => x"53b81852",
         13254 => x"81183351",
         13255 => x"fed5c43f",
         13256 => x"84b9c808",
         13257 => x"802e8538",
         13258 => x"ff578159",
         13259 => x"76b4190c",
         13260 => x"785778be",
         13261 => x"38789c17",
         13262 => x"08703357",
         13263 => x"5a577481",
         13264 => x"e52e819e",
         13265 => x"38743070",
         13266 => x"80257807",
         13267 => x"565c7480",
         13268 => x"2e81d738",
         13269 => x"811a5a79",
         13270 => x"812ea538",
         13271 => x"81527551",
         13272 => x"feefa13f",
         13273 => x"84b9c808",
         13274 => x"5784b9c8",
         13275 => x"08802eff",
         13276 => x"86388755",
         13277 => x"76842efd",
         13278 => x"bf387655",
         13279 => x"76fdb938",
         13280 => x"a06c5755",
         13281 => x"80767081",
         13282 => x"055834ff",
         13283 => x"155574f4",
         13284 => x"386b5688",
         13285 => x"0b8b1734",
         13286 => x"8b6c7e59",
         13287 => x"57557670",
         13288 => x"81055833",
         13289 => x"76708105",
         13290 => x"5834ff15",
         13291 => x"5574802e",
         13292 => x"fdeb3876",
         13293 => x"70810558",
         13294 => x"33767081",
         13295 => x"055834ff",
         13296 => x"155574da",
         13297 => x"38fdd639",
         13298 => x"6b5ae57a",
         13299 => x"347d5d81",
         13300 => x"0b831e34",
         13301 => x"7d51fed7",
         13302 => x"bc3f84b9",
         13303 => x"c80855fd",
         13304 => x"ce398157",
         13305 => x"fedf3981",
         13306 => x"54b41808",
         13307 => x"537a5281",
         13308 => x"183351fe",
         13309 => x"d4ec3f84",
         13310 => x"b9c80879",
         13311 => x"2e098106",
         13312 => x"80c33884",
         13313 => x"b9c80883",
         13314 => x"1934b418",
         13315 => x"08a81908",
         13316 => x"315c7ba0",
         13317 => x"1908278a",
         13318 => x"38821833",
         13319 => x"5574822e",
         13320 => x"b13884b9",
         13321 => x"c80859fd",
         13322 => x"e839745a",
         13323 => x"81527551",
         13324 => x"feedd13f",
         13325 => x"84b9c808",
         13326 => x"5784b9c8",
         13327 => x"08802efd",
         13328 => x"b638feae",
         13329 => x"39817058",
         13330 => x"5978802e",
         13331 => x"fde738fe",
         13332 => x"a1398154",
         13333 => x"b41808a0",
         13334 => x"19080553",
         13335 => x"7a528118",
         13336 => x"3351fed3",
         13337 => x"fd3ffda9",
         13338 => x"39f23d0d",
         13339 => x"60620288",
         13340 => x"0580cb05",
         13341 => x"335e5b57",
         13342 => x"89567680",
         13343 => x"2e9f3876",
         13344 => x"08557480",
         13345 => x"2e973874",
         13346 => x"33547380",
         13347 => x"2e8f3886",
         13348 => x"15228418",
         13349 => x"22595978",
         13350 => x"782e81c2",
         13351 => x"38805473",
         13352 => x"5f7581a5",
         13353 => x"38911733",
         13354 => x"5675819d",
         13355 => x"3879802e",
         13356 => x"81a2388c",
         13357 => x"1708819c",
         13358 => x"38901733",
         13359 => x"70812a81",
         13360 => x"06565d74",
         13361 => x"802e818c",
         13362 => x"387e8a11",
         13363 => x"2270892b",
         13364 => x"70557c54",
         13365 => x"575c59fd",
         13366 => x"87cb3fff",
         13367 => x"157a0670",
         13368 => x"30707207",
         13369 => x"9f2a84b9",
         13370 => x"c8080590",
         13371 => x"1c087942",
         13372 => x"535f5558",
         13373 => x"81782788",
         13374 => x"389c1908",
         13375 => x"78268338",
         13376 => x"82587778",
         13377 => x"565b8059",
         13378 => x"74527651",
         13379 => x"fed8873f",
         13380 => x"81157f55",
         13381 => x"559c1408",
         13382 => x"75268338",
         13383 => x"825584b9",
         13384 => x"c808812e",
         13385 => x"81dc3884",
         13386 => x"b9c808ff",
         13387 => x"2e81d838",
         13388 => x"84b9c808",
         13389 => x"81c53881",
         13390 => x"1959787d",
         13391 => x"2ebb3874",
         13392 => x"782e0981",
         13393 => x"06c23887",
         13394 => x"56755473",
         13395 => x"84b9c80c",
         13396 => x"903d0d04",
         13397 => x"870b84b9",
         13398 => x"c80c903d",
         13399 => x"0d048115",
         13400 => x"3351fed0",
         13401 => x"ac3f84b9",
         13402 => x"c8088106",
         13403 => x"5473fead",
         13404 => x"38737708",
         13405 => x"5556fea7",
         13406 => x"397b802e",
         13407 => x"818e387a",
         13408 => x"7d56587c",
         13409 => x"802eab38",
         13410 => x"81185474",
         13411 => x"812e80e6",
         13412 => x"38735377",
         13413 => x"527e51fe",
         13414 => x"dddd3f84",
         13415 => x"b9c80856",
         13416 => x"84b9c808",
         13417 => x"ffa33877",
         13418 => x"8119ff17",
         13419 => x"57595e74",
         13420 => x"d7387e7e",
         13421 => x"90120c55",
         13422 => x"7b802eff",
         13423 => x"8c387a88",
         13424 => x"180c798c",
         13425 => x"180c9017",
         13426 => x"3380c007",
         13427 => x"5c7b9018",
         13428 => x"349c1508",
         13429 => x"fe059416",
         13430 => x"08585a76",
         13431 => x"7a26fee9",
         13432 => x"38767d31",
         13433 => x"94160c84",
         13434 => x"15338107",
         13435 => x"5d7c8416",
         13436 => x"347554fe",
         13437 => x"d639ff54",
         13438 => x"ff973974",
         13439 => x"5b8059fe",
         13440 => x"be398254",
         13441 => x"fec53981",
         13442 => x"54fec039",
         13443 => x"ff1b5eff",
         13444 => x"a13984b9",
         13445 => x"d408e33d",
         13446 => x"0da33d08",
         13447 => x"a53d0802",
         13448 => x"88058187",
         13449 => x"05334442",
         13450 => x"5fff0ba2",
         13451 => x"3d08705f",
         13452 => x"5b407980",
         13453 => x"2e858a38",
         13454 => x"79708105",
         13455 => x"5b33709f",
         13456 => x"26565675",
         13457 => x"ba2e859b",
         13458 => x"3874ed38",
         13459 => x"75ba2e85",
         13460 => x"923884d1",
         13461 => x"a4335680",
         13462 => x"762484e5",
         13463 => x"38751010",
         13464 => x"84d19005",
         13465 => x"7008565a",
         13466 => x"74802e84",
         13467 => x"38807534",
         13468 => x"751684b9",
         13469 => x"bc113384",
         13470 => x"b9bd1233",
         13471 => x"405b5d81",
         13472 => x"527951fe",
         13473 => x"cea93f84",
         13474 => x"b9c80881",
         13475 => x"ff067081",
         13476 => x"065d5683",
         13477 => x"577b84ab",
         13478 => x"3875822a",
         13479 => x"8106408a",
         13480 => x"577f849f",
         13481 => x"389f3dfc",
         13482 => x"05538352",
         13483 => x"7951fed0",
         13484 => x"b03f84b9",
         13485 => x"c8088498",
         13486 => x"386d5574",
         13487 => x"802e8490",
         13488 => x"38748280",
         13489 => x"80268488",
         13490 => x"38ff1575",
         13491 => x"06557483",
         13492 => x"ff387e80",
         13493 => x"2e883884",
         13494 => x"807f2683",
         13495 => x"f8387e81",
         13496 => x"800a2683",
         13497 => x"f038ff1f",
         13498 => x"7f065574",
         13499 => x"83e7387e",
         13500 => x"892aa63d",
         13501 => x"08892a70",
         13502 => x"892b7759",
         13503 => x"4c475b60",
         13504 => x"802e85ab",
         13505 => x"38653070",
         13506 => x"80257707",
         13507 => x"565f9157",
         13508 => x"7483b038",
         13509 => x"7d802e84",
         13510 => x"df388154",
         13511 => x"74536052",
         13512 => x"7951fecd",
         13513 => x"be3f8157",
         13514 => x"84b9c808",
         13515 => x"83953860",
         13516 => x"83ff0533",
         13517 => x"6183fe05",
         13518 => x"3371882b",
         13519 => x"0759568e",
         13520 => x"577782d4",
         13521 => x"d52e0981",
         13522 => x"0682f838",
         13523 => x"7d902961",
         13524 => x"0583b211",
         13525 => x"33445862",
         13526 => x"802e82e7",
         13527 => x"3883b618",
         13528 => x"83113382",
         13529 => x"12337190",
         13530 => x"2b71882b",
         13531 => x"07811433",
         13532 => x"70720788",
         13533 => x"2b753371",
         13534 => x"0783ba1f",
         13535 => x"83113382",
         13536 => x"12337190",
         13537 => x"2b71882b",
         13538 => x"07811433",
         13539 => x"70720788",
         13540 => x"2b753371",
         13541 => x"075ca23d",
         13542 => x"0c42a33d",
         13543 => x"0ca33d0c",
         13544 => x"444e5445",
         13545 => x"594f415a",
         13546 => x"4b784d8e",
         13547 => x"5780ff79",
         13548 => x"27829038",
         13549 => x"93577a81",
         13550 => x"80268287",
         13551 => x"3861812a",
         13552 => x"70810645",
         13553 => x"4963802e",
         13554 => x"83f93861",
         13555 => x"87064564",
         13556 => x"822e8938",
         13557 => x"61810647",
         13558 => x"6683f438",
         13559 => x"836e7030",
         13560 => x"4a46437a",
         13561 => x"5862832e",
         13562 => x"8ac2387a",
         13563 => x"ae38788c",
         13564 => x"2a57810b",
         13565 => x"83e6ec22",
         13566 => x"56587480",
         13567 => x"2e9d3874",
         13568 => x"77269838",
         13569 => x"83e6ec56",
         13570 => x"77108217",
         13571 => x"70225757",
         13572 => x"5874802e",
         13573 => x"86387675",
         13574 => x"27ee3877",
         13575 => x"527851fd",
         13576 => x"81833f84",
         13577 => x"b9c80810",
         13578 => x"84055584",
         13579 => x"b9c8089f",
         13580 => x"f5269638",
         13581 => x"810b84b9",
         13582 => x"c8081084",
         13583 => x"b9c80805",
         13584 => x"7111722a",
         13585 => x"8305574c",
         13586 => x"4383ff15",
         13587 => x"892a5d81",
         13588 => x"5ca0477b",
         13589 => x"1f7d1168",
         13590 => x"056611ff",
         13591 => x"05706b06",
         13592 => x"7231584e",
         13593 => x"57446283",
         13594 => x"2e89b838",
         13595 => x"741d5d77",
         13596 => x"90291670",
         13597 => x"60315657",
         13598 => x"74792682",
         13599 => x"f238787c",
         13600 => x"317d3178",
         13601 => x"53706831",
         13602 => x"5256fd80",
         13603 => x"983f84b9",
         13604 => x"c8084062",
         13605 => x"832e89f6",
         13606 => x"3862822e",
         13607 => x"09810682",
         13608 => x"dd3883ff",
         13609 => x"f50b84b9",
         13610 => x"c8082782",
         13611 => x"ac387a89",
         13612 => x"f9387718",
         13613 => x"557480c0",
         13614 => x"2689ef38",
         13615 => x"745bfea3",
         13616 => x"398b5776",
         13617 => x"84b9c80c",
         13618 => x"9f3d0d84",
         13619 => x"b9d40c04",
         13620 => x"814efbfe",
         13621 => x"39930b84",
         13622 => x"b9c80c9f",
         13623 => x"3d0d84b9",
         13624 => x"d40c047c",
         13625 => x"33d01170",
         13626 => x"81ff0657",
         13627 => x"57577489",
         13628 => x"26913882",
         13629 => x"1d7781ff",
         13630 => x"06d0055d",
         13631 => x"58777a2e",
         13632 => x"81b23880",
         13633 => x"0b83e5b8",
         13634 => x"5f5c7d08",
         13635 => x"7d575b7a",
         13636 => x"7081055c",
         13637 => x"33767081",
         13638 => x"055833ff",
         13639 => x"9f124559",
         13640 => x"57629926",
         13641 => x"8938e017",
         13642 => x"7081ff06",
         13643 => x"5844ff9f",
         13644 => x"18456499",
         13645 => x"268938e0",
         13646 => x"187081ff",
         13647 => x"06594676",
         13648 => x"30709f2a",
         13649 => x"5a477678",
         13650 => x"2e098106",
         13651 => x"853878ff",
         13652 => x"be38757a",
         13653 => x"32703070",
         13654 => x"72079f2a",
         13655 => x"7b075d4a",
         13656 => x"4a7a802e",
         13657 => x"80ce3881",
         13658 => x"1c841f5f",
         13659 => x"5c837c25",
         13660 => x"ff98387f",
         13661 => x"56f9e039",
         13662 => x"9f3df805",
         13663 => x"53815279",
         13664 => x"51fecadd",
         13665 => x"3f815784",
         13666 => x"b9c808fe",
         13667 => x"b6386183",
         13668 => x"2a770684",
         13669 => x"b9c80840",
         13670 => x"56758338",
         13671 => x"bf5f6c55",
         13672 => x"8e577e75",
         13673 => x"26fe9c38",
         13674 => x"747f3159",
         13675 => x"fbfb3981",
         13676 => x"56fad239",
         13677 => x"7b8324ff",
         13678 => x"ba387b7a",
         13679 => x"a33d0c56",
         13680 => x"f9953961",
         13681 => x"81064893",
         13682 => x"5767802e",
         13683 => x"fdf53882",
         13684 => x"6e70304a",
         13685 => x"4643fc8b",
         13686 => x"3984b9c8",
         13687 => x"089ff526",
         13688 => x"9d387a8b",
         13689 => x"3877185b",
         13690 => x"81807b27",
         13691 => x"fbf5388e",
         13692 => x"577684b9",
         13693 => x"c80c9f3d",
         13694 => x"0d84b9d4",
         13695 => x"0c048055",
         13696 => x"62812e86",
         13697 => x"99389ff5",
         13698 => x"60278b38",
         13699 => x"7481065b",
         13700 => x"8e577afd",
         13701 => x"ae388480",
         13702 => x"61575580",
         13703 => x"76708105",
         13704 => x"5834ff15",
         13705 => x"5574f438",
         13706 => x"8b6183e5",
         13707 => x"84595755",
         13708 => x"76708105",
         13709 => x"58337670",
         13710 => x"81055834",
         13711 => x"ff155574",
         13712 => x"ef38608b",
         13713 => x"05457465",
         13714 => x"3482618c",
         13715 => x"05347761",
         13716 => x"8d05347b",
         13717 => x"83ffff06",
         13718 => x"4b6a618e",
         13719 => x"05346a88",
         13720 => x"2a5c7b61",
         13721 => x"8f053481",
         13722 => x"61900534",
         13723 => x"62833270",
         13724 => x"305a4880",
         13725 => x"61910534",
         13726 => x"789e2a82",
         13727 => x"06496861",
         13728 => x"9205346c",
         13729 => x"567583ff",
         13730 => x"ff2686ad",
         13731 => x"387583ff",
         13732 => x"ff065574",
         13733 => x"61930534",
         13734 => x"74882a4c",
         13735 => x"6b619405",
         13736 => x"34f86195",
         13737 => x"0534bf61",
         13738 => x"98053480",
         13739 => x"61990534",
         13740 => x"ff619a05",
         13741 => x"3480619b",
         13742 => x"05347e61",
         13743 => x"9c05347e",
         13744 => x"882a4867",
         13745 => x"619d0534",
         13746 => x"7e902a4c",
         13747 => x"6b619e05",
         13748 => x"347e982a",
         13749 => x"84b9d40c",
         13750 => x"84b9d408",
         13751 => x"619f0534",
         13752 => x"62832e85",
         13753 => x"f7388061",
         13754 => x"a7053480",
         13755 => x"61a80534",
         13756 => x"a161a905",
         13757 => x"3480cc61",
         13758 => x"aa05347c",
         13759 => x"83ffff06",
         13760 => x"55746196",
         13761 => x"05347488",
         13762 => x"2a4b6a61",
         13763 => x"970534ff",
         13764 => x"8061a405",
         13765 => x"34a961a6",
         13766 => x"05349361",
         13767 => x"ab0583e5",
         13768 => x"90595755",
         13769 => x"76708105",
         13770 => x"58337670",
         13771 => x"81055834",
         13772 => x"ff155574",
         13773 => x"ef386083",
         13774 => x"fe054980",
         13775 => x"d5693460",
         13776 => x"83ff054b",
         13777 => x"ffaa6b34",
         13778 => x"81547e53",
         13779 => x"60527951",
         13780 => x"fec68f3f",
         13781 => x"815784b9",
         13782 => x"c808fae7",
         13783 => x"3860175c",
         13784 => x"62832e87",
         13785 => x"9c386961",
         13786 => x"57558076",
         13787 => x"70810558",
         13788 => x"34ff1555",
         13789 => x"74f43863",
         13790 => x"75415b62",
         13791 => x"832e86c0",
         13792 => x"3887ffff",
         13793 => x"f8576281",
         13794 => x"2e8338f8",
         13795 => x"57766134",
         13796 => x"76882a7c",
         13797 => x"45557464",
         13798 => x"70810546",
         13799 => x"3476902a",
         13800 => x"59786470",
         13801 => x"81054634",
         13802 => x"76982a56",
         13803 => x"7564347c",
         13804 => x"57655976",
         13805 => x"66268338",
         13806 => x"76597854",
         13807 => x"7a536052",
         13808 => x"7951fec5",
         13809 => x"9d3f84b9",
         13810 => x"c80885e6",
         13811 => x"38848061",
         13812 => x"57558076",
         13813 => x"70810558",
         13814 => x"34ff1555",
         13815 => x"74f43878",
         13816 => x"1b777a31",
         13817 => x"585b76c9",
         13818 => x"387f8105",
         13819 => x"407f802e",
         13820 => x"ff893877",
         13821 => x"5662832e",
         13822 => x"83386656",
         13823 => x"65557566",
         13824 => x"26833875",
         13825 => x"5574547a",
         13826 => x"53605279",
         13827 => x"51fec4d2",
         13828 => x"3f84b9c8",
         13829 => x"08859b38",
         13830 => x"741b7676",
         13831 => x"31575b75",
         13832 => x"db388c58",
         13833 => x"62832e93",
         13834 => x"3886586c",
         13835 => x"83ffff26",
         13836 => x"8a388458",
         13837 => x"62822e83",
         13838 => x"3881587d",
         13839 => x"84c13861",
         13840 => x"832a8106",
         13841 => x"5e7d81b3",
         13842 => x"38848061",
         13843 => x"56598075",
         13844 => x"70810557",
         13845 => x"34ff1959",
         13846 => x"78f43880",
         13847 => x"d56934ff",
         13848 => x"aa6b3460",
         13849 => x"83be0547",
         13850 => x"78673481",
         13851 => x"67810534",
         13852 => x"81678205",
         13853 => x"34786783",
         13854 => x"05347767",
         13855 => x"8405346c",
         13856 => x"4380fdc1",
         13857 => x"52621f51",
         13858 => x"fcf89a3f",
         13859 => x"fe678505",
         13860 => x"3484b9c8",
         13861 => x"08822abf",
         13862 => x"07577667",
         13863 => x"86053484",
         13864 => x"b9c80867",
         13865 => x"8705347e",
         13866 => x"6183c605",
         13867 => x"34676183",
         13868 => x"c705346b",
         13869 => x"6183c805",
         13870 => x"3484b9d4",
         13871 => x"086183c9",
         13872 => x"05346261",
         13873 => x"83ca0534",
         13874 => x"62882a45",
         13875 => x"646183cb",
         13876 => x"05346290",
         13877 => x"2a587761",
         13878 => x"83cc0534",
         13879 => x"62982a5f",
         13880 => x"7e6183cd",
         13881 => x"05348154",
         13882 => x"78536052",
         13883 => x"7951fec2",
         13884 => x"f13f8157",
         13885 => x"84b9c808",
         13886 => x"f7c93880",
         13887 => x"53805279",
         13888 => x"51fec3dd",
         13889 => x"3f815784",
         13890 => x"b9c808f7",
         13891 => x"b63884b9",
         13892 => x"c80884b9",
         13893 => x"c80c9f3d",
         13894 => x"0d84b9d4",
         13895 => x"0c046255",
         13896 => x"f9e43974",
         13897 => x"1c641645",
         13898 => x"5cf6c439",
         13899 => x"7aae3878",
         13900 => x"912a5781",
         13901 => x"0b83e6fc",
         13902 => x"22565874",
         13903 => x"802e9d38",
         13904 => x"74772698",
         13905 => x"3883e6fc",
         13906 => x"56771082",
         13907 => x"17702257",
         13908 => x"57587480",
         13909 => x"2e863876",
         13910 => x"7527ee38",
         13911 => x"77527851",
         13912 => x"fcf6c23f",
         13913 => x"84b9c808",
         13914 => x"10108487",
         13915 => x"0570892a",
         13916 => x"5e5ca05c",
         13917 => x"800b84b9",
         13918 => x"c808fc80",
         13919 => x"8a055847",
         13920 => x"fdfff00a",
         13921 => x"7727f5cb",
         13922 => x"388e57f8",
         13923 => x"e43984b9",
         13924 => x"c80883ff",
         13925 => x"f526f8e6",
         13926 => x"387af8d3",
         13927 => x"3877812a",
         13928 => x"5b7af4bf",
         13929 => x"388e57f8",
         13930 => x"c8396881",
         13931 => x"06446380",
         13932 => x"2ef8af38",
         13933 => x"8343f4ab",
         13934 => x"397561a0",
         13935 => x"05347588",
         13936 => x"2a496861",
         13937 => x"a1053475",
         13938 => x"902a5b7a",
         13939 => x"61a20534",
         13940 => x"75982a57",
         13941 => x"7661a305",
         13942 => x"34f9c639",
         13943 => x"806180c3",
         13944 => x"05348061",
         13945 => x"80c40534",
         13946 => x"a16180c5",
         13947 => x"053480cc",
         13948 => x"6180c605",
         13949 => x"347c61a4",
         13950 => x"05347c88",
         13951 => x"2a5c7b61",
         13952 => x"a505347c",
         13953 => x"902a5978",
         13954 => x"61a60534",
         13955 => x"7c982a56",
         13956 => x"7561a705",
         13957 => x"348261ac",
         13958 => x"05348061",
         13959 => x"ad053480",
         13960 => x"61ae0534",
         13961 => x"8061af05",
         13962 => x"348161b0",
         13963 => x"05348061",
         13964 => x"b1053486",
         13965 => x"61b20534",
         13966 => x"8061b305",
         13967 => x"34ff8061",
         13968 => x"80c00534",
         13969 => x"a96180c2",
         13970 => x"05349361",
         13971 => x"80c70583",
         13972 => x"e5a45957",
         13973 => x"55767081",
         13974 => x"05583376",
         13975 => x"70810558",
         13976 => x"34ff1555",
         13977 => x"74802ef9",
         13978 => x"cd387670",
         13979 => x"81055833",
         13980 => x"76708105",
         13981 => x"5834ff15",
         13982 => x"5574da38",
         13983 => x"f9b83981",
         13984 => x"54805360",
         13985 => x"527951fe",
         13986 => x"bed93f81",
         13987 => x"5784b9c8",
         13988 => x"08f4b038",
         13989 => x"7d902961",
         13990 => x"05427762",
         13991 => x"83b20534",
         13992 => x"765484b9",
         13993 => x"c8085360",
         13994 => x"527951fe",
         13995 => x"bfb43ffc",
         13996 => x"c339810b",
         13997 => x"84b9c80c",
         13998 => x"9f3d0d84",
         13999 => x"b9d40c04",
         14000 => x"f861347b",
         14001 => x"4aff6a70",
         14002 => x"81054c34",
         14003 => x"ff6a7081",
         14004 => x"054c34ff",
         14005 => x"6a34ff61",
         14006 => x"840534ff",
         14007 => x"61850534",
         14008 => x"ff618605",
         14009 => x"34ff6187",
         14010 => x"0534ff61",
         14011 => x"880534ff",
         14012 => x"61890534",
         14013 => x"ff618a05",
         14014 => x"348f6534",
         14015 => x"7c57f9b1",
         14016 => x"39765486",
         14017 => x"1f536052",
         14018 => x"7951febe",
         14019 => x"d53f8480",
         14020 => x"61565780",
         14021 => x"75708105",
         14022 => x"5734ff17",
         14023 => x"5776f438",
         14024 => x"605c80d2",
         14025 => x"7c708105",
         14026 => x"5e347b55",
         14027 => x"80d27570",
         14028 => x"81055734",
         14029 => x"80e17570",
         14030 => x"81055734",
         14031 => x"80c17534",
         14032 => x"80f26183",
         14033 => x"e4053480",
         14034 => x"f26183e5",
         14035 => x"053480c1",
         14036 => x"6183e605",
         14037 => x"3480e161",
         14038 => x"83e70534",
         14039 => x"7fff055b",
         14040 => x"7a6183e8",
         14041 => x"05347a88",
         14042 => x"2a597861",
         14043 => x"83e90534",
         14044 => x"7a902a56",
         14045 => x"756183ea",
         14046 => x"05347a98",
         14047 => x"2a407f61",
         14048 => x"83eb0534",
         14049 => x"826183ec",
         14050 => x"05347661",
         14051 => x"83ed0534",
         14052 => x"766183ee",
         14053 => x"05347661",
         14054 => x"83ef0534",
         14055 => x"80d56934",
         14056 => x"ffaa6b34",
         14057 => x"8154871f",
         14058 => x"53605279",
         14059 => x"51febdb2",
         14060 => x"3f815481",
         14061 => x"1f536052",
         14062 => x"7951febd",
         14063 => x"a53f6961",
         14064 => x"5755f7a6",
         14065 => x"39f43d0d",
         14066 => x"7e615b5b",
         14067 => x"807b61ff",
         14068 => x"055a5757",
         14069 => x"767825b8",
         14070 => x"388d3d59",
         14071 => x"8e3df805",
         14072 => x"54815378",
         14073 => x"527951ff",
         14074 => x"9ab43f7b",
         14075 => x"812e0981",
         14076 => x"069e388d",
         14077 => x"3d335574",
         14078 => x"8d2e9038",
         14079 => x"74767081",
         14080 => x"05583481",
         14081 => x"1757748a",
         14082 => x"2e863877",
         14083 => x"7724cd38",
         14084 => x"8076347a",
         14085 => x"55768338",
         14086 => x"76557484",
         14087 => x"b9c80c8e",
         14088 => x"3d0d04f7",
         14089 => x"3d0d7b02",
         14090 => x"8405b305",
         14091 => x"33595777",
         14092 => x"8a2e80d5",
         14093 => x"38841708",
         14094 => x"56807624",
         14095 => x"9e388817",
         14096 => x"0877178c",
         14097 => x"05565977",
         14098 => x"75348116",
         14099 => x"5574bb24",
         14100 => x"8e387484",
         14101 => x"180c8119",
         14102 => x"88180c8b",
         14103 => x"3d0d048b",
         14104 => x"3dfc0554",
         14105 => x"74538c17",
         14106 => x"52760851",
         14107 => x"ff9ed13f",
         14108 => x"747a3270",
         14109 => x"30707207",
         14110 => x"9f2a7030",
         14111 => x"841b0c81",
         14112 => x"1c881b0c",
         14113 => x"5a5656d3",
         14114 => x"398d5276",
         14115 => x"51ff943f",
         14116 => x"ffa339e3",
         14117 => x"3d0d0280",
         14118 => x"ff05338d",
         14119 => x"3d585880",
         14120 => x"cc775755",
         14121 => x"80767081",
         14122 => x"055834ff",
         14123 => x"155574f4",
         14124 => x"38a13d08",
         14125 => x"770c778a",
         14126 => x"2e80f738",
         14127 => x"7c568076",
         14128 => x"2480c038",
         14129 => x"7d77178c",
         14130 => x"05565977",
         14131 => x"75348116",
         14132 => x"5574bb24",
         14133 => x"b8387484",
         14134 => x"180c8119",
         14135 => x"88180c7c",
         14136 => x"55807524",
         14137 => x"9e389f3d",
         14138 => x"ffac1155",
         14139 => x"7554c005",
         14140 => x"52760851",
         14141 => x"ff9dc93f",
         14142 => x"84b9c808",
         14143 => x"86387c7a",
         14144 => x"2eba38ff",
         14145 => x"0b84b9c8",
         14146 => x"0c9f3d0d",
         14147 => x"049f3dff",
         14148 => x"b0115575",
         14149 => x"54c00552",
         14150 => x"760851ff",
         14151 => x"9da23f74",
         14152 => x"7b327030",
         14153 => x"7072079f",
         14154 => x"2a703052",
         14155 => x"5a5656ff",
         14156 => x"a5398d52",
         14157 => x"7651fdeb",
         14158 => x"3fff8139",
         14159 => x"7d84b9c8",
         14160 => x"0c9f3d0d",
         14161 => x"04fd3d0d",
         14162 => x"75028405",
         14163 => x"9a052252",
         14164 => x"53805272",
         14165 => x"80ff2690",
         14166 => x"387283ff",
         14167 => x"ff065271",
         14168 => x"84b9c80c",
         14169 => x"853d0d04",
         14170 => x"83ffff73",
         14171 => x"27547083",
         14172 => x"b52e0981",
         14173 => x"06e93873",
         14174 => x"802ee438",
         14175 => x"83e78c22",
         14176 => x"5172712e",
         14177 => x"9c388112",
         14178 => x"7083ffff",
         14179 => x"06535471",
         14180 => x"80ff268d",
         14181 => x"38711083",
         14182 => x"e78c0570",
         14183 => x"225151e1",
         14184 => x"39818012",
         14185 => x"7081ff06",
         14186 => x"84b9c80c",
         14187 => x"53853d0d",
         14188 => x"04fe3d0d",
         14189 => x"02920522",
         14190 => x"02840596",
         14191 => x"05225351",
         14192 => x"80537080",
         14193 => x"ff268c38",
         14194 => x"70537284",
         14195 => x"b9c80c84",
         14196 => x"3d0d0471",
         14197 => x"83b52e09",
         14198 => x"8106ef38",
         14199 => x"7081ff26",
         14200 => x"e9387010",
         14201 => x"83e58c05",
         14202 => x"702284b9",
         14203 => x"c80c5184",
         14204 => x"3d0d04fb",
         14205 => x"3d0d7751",
         14206 => x"7083ffff",
         14207 => x"2680e138",
         14208 => x"7083ffff",
         14209 => x"0683e98c",
         14210 => x"5656759f",
         14211 => x"ff2680d9",
         14212 => x"38747082",
         14213 => x"05562275",
         14214 => x"71307080",
         14215 => x"25737a26",
         14216 => x"07545653",
         14217 => x"5370b738",
         14218 => x"71708205",
         14219 => x"53227271",
         14220 => x"882a5456",
         14221 => x"81ff0670",
         14222 => x"14525470",
         14223 => x"7624b138",
         14224 => x"71cf3873",
         14225 => x"10157070",
         14226 => x"82055222",
         14227 => x"54733070",
         14228 => x"80257579",
         14229 => x"26075355",
         14230 => x"5270802e",
         14231 => x"cb387551",
         14232 => x"7084b9c8",
         14233 => x"0c873d0d",
         14234 => x"0483ed80",
         14235 => x"55ffa239",
         14236 => x"718826ea",
         14237 => x"38711010",
         14238 => x"83c9e005",
         14239 => x"54730804",
         14240 => x"c7a01670",
         14241 => x"83ffff06",
         14242 => x"57517551",
         14243 => x"d339ffb0",
         14244 => x"167083ff",
         14245 => x"ff065751",
         14246 => x"f1398816",
         14247 => x"7083ffff",
         14248 => x"065751e6",
         14249 => x"39e61670",
         14250 => x"83ffff06",
         14251 => x"5751db39",
         14252 => x"d0167083",
         14253 => x"ffff0657",
         14254 => x"51d039e0",
         14255 => x"167083ff",
         14256 => x"ff065751",
         14257 => x"c539f016",
         14258 => x"7083ffff",
         14259 => x"065751ff",
         14260 => x"b9397573",
         14261 => x"31810676",
         14262 => x"71317083",
         14263 => x"ffff0658",
         14264 => x"5255ffa6",
         14265 => x"39757331",
         14266 => x"10750570",
         14267 => x"225252fe",
         14268 => x"ef390000",
         14269 => x"00ffffff",
         14270 => x"ff00ffff",
         14271 => x"ffff00ff",
         14272 => x"ffffff00",
         14273 => x"0000198b",
         14274 => x"00001980",
         14275 => x"00001975",
         14276 => x"0000196a",
         14277 => x"0000195f",
         14278 => x"00001954",
         14279 => x"00001949",
         14280 => x"0000193e",
         14281 => x"00001933",
         14282 => x"00001928",
         14283 => x"0000191d",
         14284 => x"00001912",
         14285 => x"00001907",
         14286 => x"000018fc",
         14287 => x"000018f1",
         14288 => x"000018e6",
         14289 => x"000018db",
         14290 => x"000018d0",
         14291 => x"000018c5",
         14292 => x"000018ba",
         14293 => x"00001ebf",
         14294 => x"00001f59",
         14295 => x"00001f59",
         14296 => x"00001f59",
         14297 => x"00001f59",
         14298 => x"00001f59",
         14299 => x"00001f59",
         14300 => x"00001f59",
         14301 => x"00001f59",
         14302 => x"00001f59",
         14303 => x"00001f59",
         14304 => x"00001f59",
         14305 => x"00001f59",
         14306 => x"00001f59",
         14307 => x"00001f59",
         14308 => x"00001f59",
         14309 => x"00001f59",
         14310 => x"00001f59",
         14311 => x"00001f59",
         14312 => x"00001f59",
         14313 => x"00001f59",
         14314 => x"00001f59",
         14315 => x"00001f59",
         14316 => x"00001f59",
         14317 => x"00001f59",
         14318 => x"00001f59",
         14319 => x"00001f59",
         14320 => x"00001f59",
         14321 => x"00001f59",
         14322 => x"00001f59",
         14323 => x"00001f59",
         14324 => x"00001f59",
         14325 => x"00001f59",
         14326 => x"00001f59",
         14327 => x"00001f59",
         14328 => x"00001f59",
         14329 => x"00001f59",
         14330 => x"00001f59",
         14331 => x"00001f59",
         14332 => x"00001f59",
         14333 => x"00001f59",
         14334 => x"00001f59",
         14335 => x"00001f59",
         14336 => x"00002471",
         14337 => x"00001f59",
         14338 => x"00001f59",
         14339 => x"00001f59",
         14340 => x"00001f59",
         14341 => x"00001f59",
         14342 => x"00001f59",
         14343 => x"00001f59",
         14344 => x"00001f59",
         14345 => x"00001f59",
         14346 => x"00001f59",
         14347 => x"00001f59",
         14348 => x"00001f59",
         14349 => x"00001f59",
         14350 => x"00001f59",
         14351 => x"00001f59",
         14352 => x"00001f59",
         14353 => x"00002407",
         14354 => x"00002306",
         14355 => x"00001f59",
         14356 => x"0000228a",
         14357 => x"000024a8",
         14358 => x"00002367",
         14359 => x"0000222c",
         14360 => x"000021ce",
         14361 => x"00001f59",
         14362 => x"00001f59",
         14363 => x"00001f59",
         14364 => x"00001f59",
         14365 => x"00001f59",
         14366 => x"00001f59",
         14367 => x"00001f59",
         14368 => x"00001f59",
         14369 => x"00001f59",
         14370 => x"00001f59",
         14371 => x"00001f59",
         14372 => x"00001f59",
         14373 => x"00001f59",
         14374 => x"00001f59",
         14375 => x"00001f59",
         14376 => x"00001f59",
         14377 => x"00001f59",
         14378 => x"00001f59",
         14379 => x"00001f59",
         14380 => x"00001f59",
         14381 => x"00001f59",
         14382 => x"00001f59",
         14383 => x"00001f59",
         14384 => x"00001f59",
         14385 => x"00001f59",
         14386 => x"00001f59",
         14387 => x"00001f59",
         14388 => x"00001f59",
         14389 => x"00001f59",
         14390 => x"00001f59",
         14391 => x"00001f59",
         14392 => x"00001f59",
         14393 => x"00001f59",
         14394 => x"00001f59",
         14395 => x"00001f59",
         14396 => x"00001f59",
         14397 => x"00001f59",
         14398 => x"00001f59",
         14399 => x"00001f59",
         14400 => x"00001f59",
         14401 => x"00001f59",
         14402 => x"00001f59",
         14403 => x"00001f59",
         14404 => x"00001f59",
         14405 => x"00001f59",
         14406 => x"00001f59",
         14407 => x"00001f59",
         14408 => x"00001f59",
         14409 => x"00001f59",
         14410 => x"00001f59",
         14411 => x"00001f59",
         14412 => x"00001f59",
         14413 => x"000021ab",
         14414 => x"00002170",
         14415 => x"00001f59",
         14416 => x"00001f59",
         14417 => x"00001f59",
         14418 => x"00001f59",
         14419 => x"00001f59",
         14420 => x"00001f59",
         14421 => x"00001f59",
         14422 => x"00001f59",
         14423 => x"00002163",
         14424 => x"00002158",
         14425 => x"00001f59",
         14426 => x"00002141",
         14427 => x"00001f59",
         14428 => x"00002151",
         14429 => x"00002147",
         14430 => x"0000213a",
         14431 => x"00003222",
         14432 => x"0000323a",
         14433 => x"00003246",
         14434 => x"00003252",
         14435 => x"0000325e",
         14436 => x"0000322e",
         14437 => x"00003b97",
         14438 => x"00003a85",
         14439 => x"00003901",
         14440 => x"0000364f",
         14441 => x"00003a21",
         14442 => x"000034de",
         14443 => x"0000379b",
         14444 => x"00003674",
         14445 => x"000039cb",
         14446 => x"000036a3",
         14447 => x"00003712",
         14448 => x"0000392a",
         14449 => x"000034de",
         14450 => x"00003901",
         14451 => x"0000380b",
         14452 => x"0000379b",
         14453 => x"000034de",
         14454 => x"000034de",
         14455 => x"00003712",
         14456 => x"000036a3",
         14457 => x"00003674",
         14458 => x"0000364f",
         14459 => x"0000467c",
         14460 => x"00004695",
         14461 => x"000046ba",
         14462 => x"000046db",
         14463 => x"0000463c",
         14464 => x"00004700",
         14465 => x"00004655",
         14466 => x"000047a5",
         14467 => x"00004762",
         14468 => x"00004762",
         14469 => x"00004762",
         14470 => x"00004762",
         14471 => x"00004762",
         14472 => x"00004762",
         14473 => x"0000473b",
         14474 => x"00004762",
         14475 => x"00004762",
         14476 => x"00004762",
         14477 => x"00004762",
         14478 => x"00004762",
         14479 => x"00004762",
         14480 => x"00004762",
         14481 => x"00004762",
         14482 => x"00004762",
         14483 => x"00004762",
         14484 => x"00004762",
         14485 => x"00004762",
         14486 => x"00004762",
         14487 => x"00004762",
         14488 => x"00004762",
         14489 => x"00004762",
         14490 => x"00004762",
         14491 => x"00004762",
         14492 => x"00004762",
         14493 => x"00004762",
         14494 => x"00004762",
         14495 => x"00004762",
         14496 => x"0000487a",
         14497 => x"00004868",
         14498 => x"00004855",
         14499 => x"00004842",
         14500 => x"0000476c",
         14501 => x"00004830",
         14502 => x"0000481d",
         14503 => x"00004785",
         14504 => x"00004762",
         14505 => x"00004785",
         14506 => x"0000480d",
         14507 => x"0000488a",
         14508 => x"000047b6",
         14509 => x"00004794",
         14510 => x"000047fb",
         14511 => x"000047e9",
         14512 => x"000047d7",
         14513 => x"000047c8",
         14514 => x"00004762",
         14515 => x"0000476c",
         14516 => x"00005408",
         14517 => x"00005577",
         14518 => x"00005549",
         14519 => x"000054a0",
         14520 => x"0000547d",
         14521 => x"0000545c",
         14522 => x"00005432",
         14523 => x"00005602",
         14524 => x"00005289",
         14525 => x"000055dc",
         14526 => x"000057cb",
         14527 => x"00005289",
         14528 => x"00005289",
         14529 => x"00005289",
         14530 => x"00005289",
         14531 => x"00005289",
         14532 => x"00005289",
         14533 => x"000055a5",
         14534 => x"000057b3",
         14535 => x"0000566a",
         14536 => x"00005289",
         14537 => x"00005289",
         14538 => x"00005289",
         14539 => x"00005289",
         14540 => x"00005289",
         14541 => x"00005289",
         14542 => x"00005289",
         14543 => x"00005289",
         14544 => x"00005289",
         14545 => x"00005289",
         14546 => x"00005289",
         14547 => x"00005289",
         14548 => x"00005289",
         14549 => x"00005289",
         14550 => x"00005289",
         14551 => x"00005289",
         14552 => x"00005289",
         14553 => x"00005289",
         14554 => x"00005289",
         14555 => x"00005527",
         14556 => x"00005289",
         14557 => x"00005289",
         14558 => x"00005289",
         14559 => x"000054ca",
         14560 => x"000053d9",
         14561 => x"0000537b",
         14562 => x"00005289",
         14563 => x"00005289",
         14564 => x"00005289",
         14565 => x"00005289",
         14566 => x"00005360",
         14567 => x"00005289",
         14568 => x"00005343",
         14569 => x"000059ac",
         14570 => x"00005921",
         14571 => x"00005921",
         14572 => x"00005921",
         14573 => x"00005921",
         14574 => x"00005921",
         14575 => x"00005921",
         14576 => x"000058fc",
         14577 => x"00005921",
         14578 => x"00005921",
         14579 => x"00005921",
         14580 => x"00005921",
         14581 => x"00005921",
         14582 => x"00005921",
         14583 => x"00005921",
         14584 => x"00005921",
         14585 => x"00005921",
         14586 => x"00005921",
         14587 => x"00005921",
         14588 => x"00005921",
         14589 => x"00005921",
         14590 => x"00005921",
         14591 => x"00005921",
         14592 => x"00005921",
         14593 => x"00005921",
         14594 => x"00005921",
         14595 => x"00005921",
         14596 => x"00005921",
         14597 => x"00005921",
         14598 => x"00005921",
         14599 => x"000059be",
         14600 => x"00005a06",
         14601 => x"000059f3",
         14602 => x"000059e0",
         14603 => x"000059ce",
         14604 => x"00005a91",
         14605 => x"00005a7e",
         14606 => x"00005a6e",
         14607 => x"00005921",
         14608 => x"00005a5e",
         14609 => x"00005a4e",
         14610 => x"00005a3c",
         14611 => x"00005a2a",
         14612 => x"00005a18",
         14613 => x"00005989",
         14614 => x"00005978",
         14615 => x"00005967",
         14616 => x"00005950",
         14617 => x"00005921",
         14618 => x"0000599a",
         14619 => x"0000637b",
         14620 => x"000061d7",
         14621 => x"000061d7",
         14622 => x"000061d7",
         14623 => x"000061d7",
         14624 => x"000061d7",
         14625 => x"000061d7",
         14626 => x"000061d7",
         14627 => x"000061d7",
         14628 => x"000061d7",
         14629 => x"000061d7",
         14630 => x"000061d7",
         14631 => x"000061d7",
         14632 => x"000061d7",
         14633 => x"00005ef9",
         14634 => x"000061d7",
         14635 => x"000061d7",
         14636 => x"000061d7",
         14637 => x"000061d7",
         14638 => x"000061d7",
         14639 => x"000061d7",
         14640 => x"000063c5",
         14641 => x"000061d7",
         14642 => x"000061d7",
         14643 => x"00006350",
         14644 => x"000061d7",
         14645 => x"00006367",
         14646 => x"00005ed8",
         14647 => x"00006339",
         14648 => x"0000dee5",
         14649 => x"0000ded2",
         14650 => x"0000dec6",
         14651 => x"0000debb",
         14652 => x"0000deb0",
         14653 => x"0000dea5",
         14654 => x"0000de9a",
         14655 => x"0000de8e",
         14656 => x"0000de80",
         14657 => x"00000e01",
         14658 => x"00000bfd",
         14659 => x"00000bfd",
         14660 => x"00000f49",
         14661 => x"00000bfd",
         14662 => x"00000bfd",
         14663 => x"00000bfd",
         14664 => x"00000bfd",
         14665 => x"00000bfd",
         14666 => x"00000bfd",
         14667 => x"00000bfd",
         14668 => x"00000dfd",
         14669 => x"00000bfd",
         14670 => x"00000f7f",
         14671 => x"00000f0d",
         14672 => x"00000bfd",
         14673 => x"00000bfd",
         14674 => x"00000bfd",
         14675 => x"00000bfd",
         14676 => x"00000bfd",
         14677 => x"00000bfd",
         14678 => x"00000bfd",
         14679 => x"00000bfd",
         14680 => x"00000bfd",
         14681 => x"00000bfd",
         14682 => x"00000bfd",
         14683 => x"00000bfd",
         14684 => x"00000bfd",
         14685 => x"00000bfd",
         14686 => x"00000bfd",
         14687 => x"00000bfd",
         14688 => x"00000bfd",
         14689 => x"00000bfd",
         14690 => x"00000bfd",
         14691 => x"00000bfd",
         14692 => x"00000bfd",
         14693 => x"00000bfd",
         14694 => x"00000bfd",
         14695 => x"00000bfd",
         14696 => x"00000bfd",
         14697 => x"00000bfd",
         14698 => x"00000bfd",
         14699 => x"00000bfd",
         14700 => x"00000bfd",
         14701 => x"00000bfd",
         14702 => x"00000bfd",
         14703 => x"00000bfd",
         14704 => x"00000bfd",
         14705 => x"00000bfd",
         14706 => x"00000bfd",
         14707 => x"00000bfd",
         14708 => x"00000f1d",
         14709 => x"00000bfd",
         14710 => x"00000bfd",
         14711 => x"00000bfd",
         14712 => x"00000bfd",
         14713 => x"00000e17",
         14714 => x"00000bfd",
         14715 => x"00000bfd",
         14716 => x"00000bfd",
         14717 => x"00000bfd",
         14718 => x"00000bfd",
         14719 => x"00000bfd",
         14720 => x"00000bfd",
         14721 => x"00000bfd",
         14722 => x"00000bfd",
         14723 => x"00000bfd",
         14724 => x"00000e2b",
         14725 => x"00000ee1",
         14726 => x"00000eb8",
         14727 => x"00000eb8",
         14728 => x"00000eb8",
         14729 => x"00000bfd",
         14730 => x"00000ee1",
         14731 => x"00000bfd",
         14732 => x"00000bfd",
         14733 => x"00000eff",
         14734 => x"00000bfd",
         14735 => x"00000bfd",
         14736 => x"00000c16",
         14737 => x"00000e0f",
         14738 => x"00000bfd",
         14739 => x"00000bfd",
         14740 => x"00000f58",
         14741 => x"00000bfd",
         14742 => x"00000c18",
         14743 => x"00000bfd",
         14744 => x"00000bfd",
         14745 => x"00000e17",
         14746 => x"64696e69",
         14747 => x"74000000",
         14748 => x"64696f63",
         14749 => x"746c0000",
         14750 => x"66696e69",
         14751 => x"74000000",
         14752 => x"666c6f61",
         14753 => x"64000000",
         14754 => x"66657865",
         14755 => x"63000000",
         14756 => x"6d636c65",
         14757 => x"61720000",
         14758 => x"6d636f70",
         14759 => x"79000000",
         14760 => x"6d646966",
         14761 => x"66000000",
         14762 => x"6d64756d",
         14763 => x"70000000",
         14764 => x"6d656200",
         14765 => x"6d656800",
         14766 => x"6d657700",
         14767 => x"68696400",
         14768 => x"68696500",
         14769 => x"68666400",
         14770 => x"68666500",
         14771 => x"63616c6c",
         14772 => x"00000000",
         14773 => x"6a6d7000",
         14774 => x"72657374",
         14775 => x"61727400",
         14776 => x"72657365",
         14777 => x"74000000",
         14778 => x"696e666f",
         14779 => x"00000000",
         14780 => x"74657374",
         14781 => x"00000000",
         14782 => x"636c7300",
         14783 => x"7a383000",
         14784 => x"74626173",
         14785 => x"69630000",
         14786 => x"6d626173",
         14787 => x"69630000",
         14788 => x"6b696c6f",
         14789 => x"00000000",
         14790 => x"65640000",
         14791 => x"556e6b6e",
         14792 => x"6f776e20",
         14793 => x"6572726f",
         14794 => x"722e0000",
         14795 => x"50617261",
         14796 => x"6d657465",
         14797 => x"72732069",
         14798 => x"6e636f72",
         14799 => x"72656374",
         14800 => x"2e000000",
         14801 => x"546f6f20",
         14802 => x"6d616e79",
         14803 => x"206f7065",
         14804 => x"6e206669",
         14805 => x"6c65732e",
         14806 => x"00000000",
         14807 => x"496e7375",
         14808 => x"66666963",
         14809 => x"69656e74",
         14810 => x"206d656d",
         14811 => x"6f72792e",
         14812 => x"00000000",
         14813 => x"46696c65",
         14814 => x"20697320",
         14815 => x"6c6f636b",
         14816 => x"65642e00",
         14817 => x"54696d65",
         14818 => x"6f75742c",
         14819 => x"206f7065",
         14820 => x"72617469",
         14821 => x"6f6e2063",
         14822 => x"616e6365",
         14823 => x"6c6c6564",
         14824 => x"2e000000",
         14825 => x"466f726d",
         14826 => x"61742061",
         14827 => x"626f7274",
         14828 => x"65642e00",
         14829 => x"4e6f2063",
         14830 => x"6f6d7061",
         14831 => x"7469626c",
         14832 => x"65206669",
         14833 => x"6c657379",
         14834 => x"7374656d",
         14835 => x"20666f75",
         14836 => x"6e64206f",
         14837 => x"6e206469",
         14838 => x"736b2e00",
         14839 => x"4469736b",
         14840 => x"206e6f74",
         14841 => x"20656e61",
         14842 => x"626c6564",
         14843 => x"2e000000",
         14844 => x"44726976",
         14845 => x"65206e75",
         14846 => x"6d626572",
         14847 => x"20697320",
         14848 => x"696e7661",
         14849 => x"6c69642e",
         14850 => x"00000000",
         14851 => x"53442069",
         14852 => x"73207772",
         14853 => x"69746520",
         14854 => x"70726f74",
         14855 => x"65637465",
         14856 => x"642e0000",
         14857 => x"46696c65",
         14858 => x"2068616e",
         14859 => x"646c6520",
         14860 => x"696e7661",
         14861 => x"6c69642e",
         14862 => x"00000000",
         14863 => x"46696c65",
         14864 => x"20616c72",
         14865 => x"65616479",
         14866 => x"20657869",
         14867 => x"7374732e",
         14868 => x"00000000",
         14869 => x"41636365",
         14870 => x"73732064",
         14871 => x"656e6965",
         14872 => x"642e0000",
         14873 => x"496e7661",
         14874 => x"6c696420",
         14875 => x"66696c65",
         14876 => x"6e616d65",
         14877 => x"2e000000",
         14878 => x"4e6f2070",
         14879 => x"61746820",
         14880 => x"666f756e",
         14881 => x"642e0000",
         14882 => x"4e6f2066",
         14883 => x"696c6520",
         14884 => x"666f756e",
         14885 => x"642e0000",
         14886 => x"4469736b",
         14887 => x"206e6f74",
         14888 => x"20726561",
         14889 => x"64792e00",
         14890 => x"496e7465",
         14891 => x"726e616c",
         14892 => x"20657272",
         14893 => x"6f722e00",
         14894 => x"4469736b",
         14895 => x"20457272",
         14896 => x"6f720000",
         14897 => x"53756363",
         14898 => x"6573732e",
         14899 => x"00000000",
         14900 => x"0a256c75",
         14901 => x"20627974",
         14902 => x"65732025",
         14903 => x"73206174",
         14904 => x"20256c75",
         14905 => x"20627974",
         14906 => x"65732f73",
         14907 => x"65632e0a",
         14908 => x"00000000",
         14909 => x"72656164",
         14910 => x"00000000",
         14911 => x"2530386c",
         14912 => x"58000000",
         14913 => x"3a202000",
         14914 => x"25303258",
         14915 => x"00000000",
         14916 => x"207c0000",
         14917 => x"7c000000",
         14918 => x"20200000",
         14919 => x"25303458",
         14920 => x"00000000",
         14921 => x"20202020",
         14922 => x"20202020",
         14923 => x"00000000",
         14924 => x"7a4f5300",
         14925 => x"2a2a2025",
         14926 => x"73202800",
         14927 => x"31312f30",
         14928 => x"352f3230",
         14929 => x"32310000",
         14930 => x"76312e33",
         14931 => x"62000000",
         14932 => x"205a5055",
         14933 => x"2c207265",
         14934 => x"76202530",
         14935 => x"32782920",
         14936 => x"25732025",
         14937 => x"73202a2a",
         14938 => x"0a0a0000",
         14939 => x"4f533a00",
         14940 => x"20202020",
         14941 => x"42617365",
         14942 => x"20416464",
         14943 => x"72657373",
         14944 => x"20202020",
         14945 => x"20202020",
         14946 => x"20202020",
         14947 => x"203d2025",
         14948 => x"30386c78",
         14949 => x"0a000000",
         14950 => x"20202020",
         14951 => x"41707020",
         14952 => x"41646472",
         14953 => x"65737320",
         14954 => x"20202020",
         14955 => x"20202020",
         14956 => x"20202020",
         14957 => x"203d2025",
         14958 => x"30386c78",
         14959 => x"0a000000",
         14960 => x"5a505520",
         14961 => x"496e7465",
         14962 => x"72727570",
         14963 => x"74204861",
         14964 => x"6e646c65",
         14965 => x"72000000",
         14966 => x"55415254",
         14967 => x"31205458",
         14968 => x"20696e74",
         14969 => x"65727275",
         14970 => x"70740000",
         14971 => x"55415254",
         14972 => x"31205258",
         14973 => x"20696e74",
         14974 => x"65727275",
         14975 => x"70740000",
         14976 => x"55415254",
         14977 => x"30205458",
         14978 => x"20696e74",
         14979 => x"65727275",
         14980 => x"70740000",
         14981 => x"55415254",
         14982 => x"30205258",
         14983 => x"20696e74",
         14984 => x"65727275",
         14985 => x"70740000",
         14986 => x"494f4354",
         14987 => x"4c205752",
         14988 => x"20696e74",
         14989 => x"65727275",
         14990 => x"70740000",
         14991 => x"494f4354",
         14992 => x"4c205244",
         14993 => x"20696e74",
         14994 => x"65727275",
         14995 => x"70740000",
         14996 => x"50533220",
         14997 => x"696e7465",
         14998 => x"72727570",
         14999 => x"74000000",
         15000 => x"54696d65",
         15001 => x"7220696e",
         15002 => x"74657272",
         15003 => x"75707400",
         15004 => x"53657474",
         15005 => x"696e6720",
         15006 => x"75702074",
         15007 => x"696d6572",
         15008 => x"2e2e2e00",
         15009 => x"456e6162",
         15010 => x"6c696e67",
         15011 => x"2074696d",
         15012 => x"65722e2e",
         15013 => x"2e000000",
         15014 => x"6175746f",
         15015 => x"65786563",
         15016 => x"2e626174",
         15017 => x"00000000",
         15018 => x"7a4f535f",
         15019 => x"7a70752e",
         15020 => x"68737400",
         15021 => x"4661696c",
         15022 => x"65642074",
         15023 => x"6f20696e",
         15024 => x"69746961",
         15025 => x"6c697365",
         15026 => x"20736420",
         15027 => x"63617264",
         15028 => x"20302c20",
         15029 => x"706c6561",
         15030 => x"73652069",
         15031 => x"6e697420",
         15032 => x"6d616e75",
         15033 => x"616c6c79",
         15034 => x"2e000000",
         15035 => x"2a200000",
         15036 => x"25643a5c",
         15037 => x"25730000",
         15038 => x"303a0000",
         15039 => x"42616420",
         15040 => x"636f6d6d",
         15041 => x"616e642e",
         15042 => x"00000000",
         15043 => x"5a505500",
         15044 => x"62696e00",
         15045 => x"25643a5c",
         15046 => x"25735c25",
         15047 => x"732e2573",
         15048 => x"00000000",
         15049 => x"436f6c64",
         15050 => x"20726562",
         15051 => x"6f6f7469",
         15052 => x"6e672e2e",
         15053 => x"2e000000",
         15054 => x"52657374",
         15055 => x"61727469",
         15056 => x"6e672061",
         15057 => x"70706c69",
         15058 => x"63617469",
         15059 => x"6f6e2e2e",
         15060 => x"2e000000",
         15061 => x"43616c6c",
         15062 => x"696e6720",
         15063 => x"636f6465",
         15064 => x"20402025",
         15065 => x"30386c78",
         15066 => x"202e2e2e",
         15067 => x"0a000000",
         15068 => x"43616c6c",
         15069 => x"20726574",
         15070 => x"75726e65",
         15071 => x"6420636f",
         15072 => x"64652028",
         15073 => x"2564292e",
         15074 => x"0a000000",
         15075 => x"45786563",
         15076 => x"7574696e",
         15077 => x"6720636f",
         15078 => x"64652040",
         15079 => x"20253038",
         15080 => x"6c78202e",
         15081 => x"2e2e0a00",
         15082 => x"2530386c",
         15083 => x"58202530",
         15084 => x"386c582d",
         15085 => x"00000000",
         15086 => x"2530386c",
         15087 => x"58202530",
         15088 => x"34582d00",
         15089 => x"436f6d70",
         15090 => x"6172696e",
         15091 => x"672e2e2e",
         15092 => x"00000000",
         15093 => x"2530386c",
         15094 => x"78282530",
         15095 => x"3878292d",
         15096 => x"3e253038",
         15097 => x"6c782825",
         15098 => x"30387829",
         15099 => x"0a000000",
         15100 => x"436f7079",
         15101 => x"696e672e",
         15102 => x"2e2e0000",
         15103 => x"2530386c",
         15104 => x"58202530",
         15105 => x"32582d00",
         15106 => x"436c6561",
         15107 => x"72696e67",
         15108 => x"2e2e2e2e",
         15109 => x"00000000",
         15110 => x"44756d70",
         15111 => x"204d656d",
         15112 => x"6f727900",
         15113 => x"0a436f6d",
         15114 => x"706c6574",
         15115 => x"652e0000",
         15116 => x"25643a5c",
         15117 => x"25735c25",
         15118 => x"73000000",
         15119 => x"4d656d6f",
         15120 => x"72792065",
         15121 => x"78686175",
         15122 => x"73746564",
         15123 => x"2c206361",
         15124 => x"6e6e6f74",
         15125 => x"2070726f",
         15126 => x"63657373",
         15127 => x"20636f6d",
         15128 => x"6d616e64",
         15129 => x"2e000000",
         15130 => x"3f3f3f00",
         15131 => x"25642f25",
         15132 => x"642f2564",
         15133 => x"2025643a",
         15134 => x"25643a25",
         15135 => x"642e2564",
         15136 => x"25640a00",
         15137 => x"536f4320",
         15138 => x"436f6e66",
         15139 => x"69677572",
         15140 => x"6174696f",
         15141 => x"6e000000",
         15142 => x"3a0a4465",
         15143 => x"76696365",
         15144 => x"7320696d",
         15145 => x"706c656d",
         15146 => x"656e7465",
         15147 => x"643a0000",
         15148 => x"41646472",
         15149 => x"65737365",
         15150 => x"733a0000",
         15151 => x"20202020",
         15152 => x"43505520",
         15153 => x"52657365",
         15154 => x"74205665",
         15155 => x"63746f72",
         15156 => x"20416464",
         15157 => x"72657373",
         15158 => x"203d2025",
         15159 => x"3038580a",
         15160 => x"00000000",
         15161 => x"20202020",
         15162 => x"43505520",
         15163 => x"4d656d6f",
         15164 => x"72792053",
         15165 => x"74617274",
         15166 => x"20416464",
         15167 => x"72657373",
         15168 => x"203d2025",
         15169 => x"3038580a",
         15170 => x"00000000",
         15171 => x"20202020",
         15172 => x"53746163",
         15173 => x"6b205374",
         15174 => x"61727420",
         15175 => x"41646472",
         15176 => x"65737320",
         15177 => x"20202020",
         15178 => x"203d2025",
         15179 => x"3038580a",
         15180 => x"00000000",
         15181 => x"4d697363",
         15182 => x"3a000000",
         15183 => x"20202020",
         15184 => x"5a505520",
         15185 => x"49642020",
         15186 => x"20202020",
         15187 => x"20202020",
         15188 => x"20202020",
         15189 => x"20202020",
         15190 => x"203d2025",
         15191 => x"3034580a",
         15192 => x"00000000",
         15193 => x"20202020",
         15194 => x"53797374",
         15195 => x"656d2043",
         15196 => x"6c6f636b",
         15197 => x"20467265",
         15198 => x"71202020",
         15199 => x"20202020",
         15200 => x"203d2025",
         15201 => x"642e2530",
         15202 => x"34644d48",
         15203 => x"7a0a0000",
         15204 => x"20202020",
         15205 => x"57697368",
         15206 => x"626f6e65",
         15207 => x"20534452",
         15208 => x"414d2043",
         15209 => x"6c6f636b",
         15210 => x"20467265",
         15211 => x"713d2025",
         15212 => x"642e2530",
         15213 => x"34644d48",
         15214 => x"7a0a0000",
         15215 => x"20202020",
         15216 => x"53445241",
         15217 => x"4d20436c",
         15218 => x"6f636b20",
         15219 => x"46726571",
         15220 => x"20202020",
         15221 => x"20202020",
         15222 => x"203d2025",
         15223 => x"642e2530",
         15224 => x"34644d48",
         15225 => x"7a0a0000",
         15226 => x"20202020",
         15227 => x"53504900",
         15228 => x"20202020",
         15229 => x"50533200",
         15230 => x"20202020",
         15231 => x"494f4354",
         15232 => x"4c000000",
         15233 => x"20202020",
         15234 => x"57422049",
         15235 => x"32430000",
         15236 => x"20202020",
         15237 => x"57495348",
         15238 => x"424f4e45",
         15239 => x"20425553",
         15240 => x"00000000",
         15241 => x"20202020",
         15242 => x"494e5452",
         15243 => x"20435452",
         15244 => x"4c202843",
         15245 => x"68616e6e",
         15246 => x"656c733d",
         15247 => x"25303264",
         15248 => x"292e0a00",
         15249 => x"20202020",
         15250 => x"54494d45",
         15251 => x"52312020",
         15252 => x"20202854",
         15253 => x"696d6572",
         15254 => x"7320203d",
         15255 => x"25303264",
         15256 => x"292e0a00",
         15257 => x"20202020",
         15258 => x"53442043",
         15259 => x"41524420",
         15260 => x"20202844",
         15261 => x"65766963",
         15262 => x"6573203d",
         15263 => x"25303264",
         15264 => x"292e0a00",
         15265 => x"20202020",
         15266 => x"52414d20",
         15267 => x"20202020",
         15268 => x"20202825",
         15269 => x"3038583a",
         15270 => x"25303858",
         15271 => x"292e0a00",
         15272 => x"20202020",
         15273 => x"4252414d",
         15274 => x"20202020",
         15275 => x"20202825",
         15276 => x"3038583a",
         15277 => x"25303858",
         15278 => x"292e0a00",
         15279 => x"20202020",
         15280 => x"494e534e",
         15281 => x"20425241",
         15282 => x"4d202825",
         15283 => x"3038583a",
         15284 => x"25303858",
         15285 => x"292e0a00",
         15286 => x"20202020",
         15287 => x"53445241",
         15288 => x"4d202020",
         15289 => x"20202825",
         15290 => x"3038583a",
         15291 => x"25303858",
         15292 => x"292e0a00",
         15293 => x"20202020",
         15294 => x"57422053",
         15295 => x"4452414d",
         15296 => x"20202825",
         15297 => x"3038583a",
         15298 => x"25303858",
         15299 => x"292e0a00",
         15300 => x"20286672",
         15301 => x"6f6d2053",
         15302 => x"6f432063",
         15303 => x"6f6e6669",
         15304 => x"67290000",
         15305 => x"556e6b6e",
         15306 => x"6f776e00",
         15307 => x"45564f6d",
         15308 => x"00000000",
         15309 => x"536d616c",
         15310 => x"6c000000",
         15311 => x"4d656469",
         15312 => x"756d0000",
         15313 => x"466c6578",
         15314 => x"00000000",
         15315 => x"45564f00",
         15316 => x"0000f0ac",
         15317 => x"01000000",
         15318 => x"00000002",
         15319 => x"0000f0a8",
         15320 => x"01000000",
         15321 => x"00000003",
         15322 => x"0000f0a4",
         15323 => x"01000000",
         15324 => x"00000004",
         15325 => x"0000f0a0",
         15326 => x"01000000",
         15327 => x"00000005",
         15328 => x"0000f09c",
         15329 => x"01000000",
         15330 => x"00000006",
         15331 => x"0000f098",
         15332 => x"01000000",
         15333 => x"00000007",
         15334 => x"0000f094",
         15335 => x"01000000",
         15336 => x"00000001",
         15337 => x"0000f090",
         15338 => x"01000000",
         15339 => x"00000008",
         15340 => x"0000f08c",
         15341 => x"01000000",
         15342 => x"0000000b",
         15343 => x"0000f088",
         15344 => x"01000000",
         15345 => x"00000009",
         15346 => x"0000f084",
         15347 => x"01000000",
         15348 => x"0000000a",
         15349 => x"0000f080",
         15350 => x"04000000",
         15351 => x"0000000d",
         15352 => x"0000f07c",
         15353 => x"04000000",
         15354 => x"0000000c",
         15355 => x"0000f078",
         15356 => x"04000000",
         15357 => x"0000000e",
         15358 => x"0000f074",
         15359 => x"03000000",
         15360 => x"0000000f",
         15361 => x"0000f070",
         15362 => x"04000000",
         15363 => x"0000000f",
         15364 => x"0000f06c",
         15365 => x"04000000",
         15366 => x"00000010",
         15367 => x"0000f068",
         15368 => x"04000000",
         15369 => x"00000011",
         15370 => x"0000f064",
         15371 => x"03000000",
         15372 => x"00000012",
         15373 => x"0000f060",
         15374 => x"03000000",
         15375 => x"00000013",
         15376 => x"0000f05c",
         15377 => x"03000000",
         15378 => x"00000014",
         15379 => x"0000f058",
         15380 => x"03000000",
         15381 => x"00000015",
         15382 => x"1b5b4400",
         15383 => x"1b5b4300",
         15384 => x"1b5b4200",
         15385 => x"1b5b4100",
         15386 => x"1b5b367e",
         15387 => x"1b5b357e",
         15388 => x"1b5b347e",
         15389 => x"1b304600",
         15390 => x"1b5b337e",
         15391 => x"1b5b327e",
         15392 => x"1b5b317e",
         15393 => x"10000000",
         15394 => x"0e000000",
         15395 => x"0d000000",
         15396 => x"0b000000",
         15397 => x"08000000",
         15398 => x"06000000",
         15399 => x"05000000",
         15400 => x"04000000",
         15401 => x"03000000",
         15402 => x"02000000",
         15403 => x"01000000",
         15404 => x"43616e6e",
         15405 => x"6f74206f",
         15406 => x"70656e2f",
         15407 => x"63726561",
         15408 => x"74652068",
         15409 => x"6973746f",
         15410 => x"72792066",
         15411 => x"696c652c",
         15412 => x"20646973",
         15413 => x"61626c69",
         15414 => x"6e672e00",
         15415 => x"68697374",
         15416 => x"6f727900",
         15417 => x"68697374",
         15418 => x"00000000",
         15419 => x"21000000",
         15420 => x"2530366c",
         15421 => x"75202025",
         15422 => x"730a0000",
         15423 => x"4661696c",
         15424 => x"65642074",
         15425 => x"6f207265",
         15426 => x"73657420",
         15427 => x"74686520",
         15428 => x"68697374",
         15429 => x"6f727920",
         15430 => x"66696c65",
         15431 => x"20746f20",
         15432 => x"454f462e",
         15433 => x"00000000",
         15434 => x"3e25730a",
         15435 => x"00000000",
         15436 => x"1b5b317e",
         15437 => x"00000000",
         15438 => x"1b5b4100",
         15439 => x"1b5b4200",
         15440 => x"1b5b4300",
         15441 => x"1b5b4400",
         15442 => x"1b5b3130",
         15443 => x"7e000000",
         15444 => x"1b5b3131",
         15445 => x"7e000000",
         15446 => x"1b5b3132",
         15447 => x"7e000000",
         15448 => x"1b5b3133",
         15449 => x"7e000000",
         15450 => x"1b5b3134",
         15451 => x"7e000000",
         15452 => x"1b5b3135",
         15453 => x"7e000000",
         15454 => x"1b5b3137",
         15455 => x"7e000000",
         15456 => x"1b5b3138",
         15457 => x"7e000000",
         15458 => x"1b5b3139",
         15459 => x"7e000000",
         15460 => x"1b5b3230",
         15461 => x"7e000000",
         15462 => x"1b5b327e",
         15463 => x"00000000",
         15464 => x"1b5b337e",
         15465 => x"00000000",
         15466 => x"1b5b4600",
         15467 => x"1b5b357e",
         15468 => x"00000000",
         15469 => x"1b5b367e",
         15470 => x"00000000",
         15471 => x"583a2564",
         15472 => x"2c25642c",
         15473 => x"25642c25",
         15474 => x"642c2564",
         15475 => x"2c25643a",
         15476 => x"25303278",
         15477 => x"00000000",
         15478 => x"443a2564",
         15479 => x"2d25642d",
         15480 => x"25643a25",
         15481 => x"633a2564",
         15482 => x"2c25642c",
         15483 => x"25643a00",
         15484 => x"25642c00",
         15485 => x"4b3a2564",
         15486 => x"3a000000",
         15487 => x"25303278",
         15488 => x"2c000000",
         15489 => x"25635b25",
         15490 => x"643b2564",
         15491 => x"52000000",
         15492 => x"5265706f",
         15493 => x"72742043",
         15494 => x"7572736f",
         15495 => x"723a0000",
         15496 => x"55703a25",
         15497 => x"30327820",
         15498 => x"25303278",
         15499 => x"00000000",
         15500 => x"44773a25",
         15501 => x"30327820",
         15502 => x"25303278",
         15503 => x"00000000",
         15504 => x"48643a25",
         15505 => x"30327820",
         15506 => x"00000000",
         15507 => x"4e6f2074",
         15508 => x"65737420",
         15509 => x"64656669",
         15510 => x"6e65642e",
         15511 => x"00000000",
         15512 => x"53440000",
         15513 => x"222a3a3c",
         15514 => x"3e3f7c7f",
         15515 => x"00000000",
         15516 => x"2b2c3b3d",
         15517 => x"5b5d0000",
         15518 => x"46415400",
         15519 => x"46415433",
         15520 => x"32000000",
         15521 => x"ebfe904d",
         15522 => x"53444f53",
         15523 => x"352e3000",
         15524 => x"4e4f204e",
         15525 => x"414d4520",
         15526 => x"20202046",
         15527 => x"41542020",
         15528 => x"20202000",
         15529 => x"4e4f204e",
         15530 => x"414d4520",
         15531 => x"20202046",
         15532 => x"41543332",
         15533 => x"20202000",
         15534 => x"0000f260",
         15535 => x"00000000",
         15536 => x"00000000",
         15537 => x"00000000",
         15538 => x"01030507",
         15539 => x"090e1012",
         15540 => x"1416181c",
         15541 => x"1e000000",
         15542 => x"809a4541",
         15543 => x"8e418f80",
         15544 => x"45454549",
         15545 => x"49498e8f",
         15546 => x"9092924f",
         15547 => x"994f5555",
         15548 => x"59999a9b",
         15549 => x"9c9d9e9f",
         15550 => x"41494f55",
         15551 => x"a5a5a6a7",
         15552 => x"a8a9aaab",
         15553 => x"acadaeaf",
         15554 => x"b0b1b2b3",
         15555 => x"b4b5b6b7",
         15556 => x"b8b9babb",
         15557 => x"bcbdbebf",
         15558 => x"c0c1c2c3",
         15559 => x"c4c5c6c7",
         15560 => x"c8c9cacb",
         15561 => x"cccdcecf",
         15562 => x"d0d1d2d3",
         15563 => x"d4d5d6d7",
         15564 => x"d8d9dadb",
         15565 => x"dcdddedf",
         15566 => x"e0e1e2e3",
         15567 => x"e4e5e6e7",
         15568 => x"e8e9eaeb",
         15569 => x"ecedeeef",
         15570 => x"f0f1f2f3",
         15571 => x"f4f5f6f7",
         15572 => x"f8f9fafb",
         15573 => x"fcfdfeff",
         15574 => x"2b2e2c3b",
         15575 => x"3d5b5d2f",
         15576 => x"5c222a3a",
         15577 => x"3c3e3f7c",
         15578 => x"7f000000",
         15579 => x"00010004",
         15580 => x"00100040",
         15581 => x"01000200",
         15582 => x"00000000",
         15583 => x"00010002",
         15584 => x"00040008",
         15585 => x"00100020",
         15586 => x"00000000",
         15587 => x"00c700fc",
         15588 => x"00e900e2",
         15589 => x"00e400e0",
         15590 => x"00e500e7",
         15591 => x"00ea00eb",
         15592 => x"00e800ef",
         15593 => x"00ee00ec",
         15594 => x"00c400c5",
         15595 => x"00c900e6",
         15596 => x"00c600f4",
         15597 => x"00f600f2",
         15598 => x"00fb00f9",
         15599 => x"00ff00d6",
         15600 => x"00dc00a2",
         15601 => x"00a300a5",
         15602 => x"20a70192",
         15603 => x"00e100ed",
         15604 => x"00f300fa",
         15605 => x"00f100d1",
         15606 => x"00aa00ba",
         15607 => x"00bf2310",
         15608 => x"00ac00bd",
         15609 => x"00bc00a1",
         15610 => x"00ab00bb",
         15611 => x"25912592",
         15612 => x"25932502",
         15613 => x"25242561",
         15614 => x"25622556",
         15615 => x"25552563",
         15616 => x"25512557",
         15617 => x"255d255c",
         15618 => x"255b2510",
         15619 => x"25142534",
         15620 => x"252c251c",
         15621 => x"2500253c",
         15622 => x"255e255f",
         15623 => x"255a2554",
         15624 => x"25692566",
         15625 => x"25602550",
         15626 => x"256c2567",
         15627 => x"25682564",
         15628 => x"25652559",
         15629 => x"25582552",
         15630 => x"2553256b",
         15631 => x"256a2518",
         15632 => x"250c2588",
         15633 => x"2584258c",
         15634 => x"25902580",
         15635 => x"03b100df",
         15636 => x"039303c0",
         15637 => x"03a303c3",
         15638 => x"00b503c4",
         15639 => x"03a60398",
         15640 => x"03a903b4",
         15641 => x"221e03c6",
         15642 => x"03b52229",
         15643 => x"226100b1",
         15644 => x"22652264",
         15645 => x"23202321",
         15646 => x"00f72248",
         15647 => x"00b02219",
         15648 => x"00b7221a",
         15649 => x"207f00b2",
         15650 => x"25a000a0",
         15651 => x"0061031a",
         15652 => x"00e00317",
         15653 => x"00f80307",
         15654 => x"00ff0001",
         15655 => x"01780100",
         15656 => x"01300132",
         15657 => x"01060139",
         15658 => x"0110014a",
         15659 => x"012e0179",
         15660 => x"01060180",
         15661 => x"004d0243",
         15662 => x"01810182",
         15663 => x"01820184",
         15664 => x"01840186",
         15665 => x"01870187",
         15666 => x"0189018a",
         15667 => x"018b018b",
         15668 => x"018d018e",
         15669 => x"018f0190",
         15670 => x"01910191",
         15671 => x"01930194",
         15672 => x"01f60196",
         15673 => x"01970198",
         15674 => x"0198023d",
         15675 => x"019b019c",
         15676 => x"019d0220",
         15677 => x"019f01a0",
         15678 => x"01a001a2",
         15679 => x"01a201a4",
         15680 => x"01a401a6",
         15681 => x"01a701a7",
         15682 => x"01a901aa",
         15683 => x"01ab01ac",
         15684 => x"01ac01ae",
         15685 => x"01af01af",
         15686 => x"01b101b2",
         15687 => x"01b301b3",
         15688 => x"01b501b5",
         15689 => x"01b701b8",
         15690 => x"01b801ba",
         15691 => x"01bb01bc",
         15692 => x"01bc01be",
         15693 => x"01f701c0",
         15694 => x"01c101c2",
         15695 => x"01c301c4",
         15696 => x"01c501c4",
         15697 => x"01c701c8",
         15698 => x"01c701ca",
         15699 => x"01cb01ca",
         15700 => x"01cd0110",
         15701 => x"01dd0001",
         15702 => x"018e01de",
         15703 => x"011201f3",
         15704 => x"000301f1",
         15705 => x"01f401f4",
         15706 => x"01f80128",
         15707 => x"02220112",
         15708 => x"023a0009",
         15709 => x"2c65023b",
         15710 => x"023b023d",
         15711 => x"2c66023f",
         15712 => x"02400241",
         15713 => x"02410246",
         15714 => x"010a0253",
         15715 => x"00400181",
         15716 => x"01860255",
         15717 => x"0189018a",
         15718 => x"0258018f",
         15719 => x"025a0190",
         15720 => x"025c025d",
         15721 => x"025e025f",
         15722 => x"01930261",
         15723 => x"02620194",
         15724 => x"02640265",
         15725 => x"02660267",
         15726 => x"01970196",
         15727 => x"026a2c62",
         15728 => x"026c026d",
         15729 => x"026e019c",
         15730 => x"02700271",
         15731 => x"019d0273",
         15732 => x"0274019f",
         15733 => x"02760277",
         15734 => x"02780279",
         15735 => x"027a027b",
         15736 => x"027c2c64",
         15737 => x"027e027f",
         15738 => x"01a60281",
         15739 => x"028201a9",
         15740 => x"02840285",
         15741 => x"02860287",
         15742 => x"01ae0244",
         15743 => x"01b101b2",
         15744 => x"0245028d",
         15745 => x"028e028f",
         15746 => x"02900291",
         15747 => x"01b7037b",
         15748 => x"000303fd",
         15749 => x"03fe03ff",
         15750 => x"03ac0004",
         15751 => x"03860388",
         15752 => x"0389038a",
         15753 => x"03b10311",
         15754 => x"03c20002",
         15755 => x"03a303a3",
         15756 => x"03c40308",
         15757 => x"03cc0003",
         15758 => x"038c038e",
         15759 => x"038f03d8",
         15760 => x"011803f2",
         15761 => x"000a03f9",
         15762 => x"03f303f4",
         15763 => x"03f503f6",
         15764 => x"03f703f7",
         15765 => x"03f903fa",
         15766 => x"03fa0430",
         15767 => x"03200450",
         15768 => x"07100460",
         15769 => x"0122048a",
         15770 => x"013604c1",
         15771 => x"010e04cf",
         15772 => x"000104c0",
         15773 => x"04d00144",
         15774 => x"05610426",
         15775 => x"00000000",
         15776 => x"1d7d0001",
         15777 => x"2c631e00",
         15778 => x"01961ea0",
         15779 => x"015a1f00",
         15780 => x"06081f10",
         15781 => x"06061f20",
         15782 => x"06081f30",
         15783 => x"06081f40",
         15784 => x"06061f51",
         15785 => x"00071f59",
         15786 => x"1f521f5b",
         15787 => x"1f541f5d",
         15788 => x"1f561f5f",
         15789 => x"1f600608",
         15790 => x"1f70000e",
         15791 => x"1fba1fbb",
         15792 => x"1fc81fc9",
         15793 => x"1fca1fcb",
         15794 => x"1fda1fdb",
         15795 => x"1ff81ff9",
         15796 => x"1fea1feb",
         15797 => x"1ffa1ffb",
         15798 => x"1f800608",
         15799 => x"1f900608",
         15800 => x"1fa00608",
         15801 => x"1fb00004",
         15802 => x"1fb81fb9",
         15803 => x"1fb21fbc",
         15804 => x"1fcc0001",
         15805 => x"1fc31fd0",
         15806 => x"06021fe0",
         15807 => x"06021fe5",
         15808 => x"00011fec",
         15809 => x"1ff30001",
         15810 => x"1ffc214e",
         15811 => x"00012132",
         15812 => x"21700210",
         15813 => x"21840001",
         15814 => x"218324d0",
         15815 => x"051a2c30",
         15816 => x"042f2c60",
         15817 => x"01022c67",
         15818 => x"01062c75",
         15819 => x"01022c80",
         15820 => x"01642d00",
         15821 => x"0826ff41",
         15822 => x"031a0000",
         15823 => x"00000000",
         15824 => x"0000e668",
         15825 => x"01020100",
         15826 => x"00000000",
         15827 => x"00000000",
         15828 => x"0000e670",
         15829 => x"01040100",
         15830 => x"00000000",
         15831 => x"00000000",
         15832 => x"0000e678",
         15833 => x"01140300",
         15834 => x"00000000",
         15835 => x"00000000",
         15836 => x"0000e680",
         15837 => x"012b0300",
         15838 => x"00000000",
         15839 => x"00000000",
         15840 => x"0000e688",
         15841 => x"01300300",
         15842 => x"00000000",
         15843 => x"00000000",
         15844 => x"0000e690",
         15845 => x"013c0400",
         15846 => x"00000000",
         15847 => x"00000000",
         15848 => x"0000e698",
         15849 => x"013d0400",
         15850 => x"00000000",
         15851 => x"00000000",
         15852 => x"0000e6a0",
         15853 => x"013f0400",
         15854 => x"00000000",
         15855 => x"00000000",
         15856 => x"0000e6a8",
         15857 => x"01400400",
         15858 => x"00000000",
         15859 => x"00000000",
         15860 => x"0000e6b0",
         15861 => x"01410400",
         15862 => x"00000000",
         15863 => x"00000000",
         15864 => x"0000e6b4",
         15865 => x"01420400",
         15866 => x"00000000",
         15867 => x"00000000",
         15868 => x"0000e6b8",
         15869 => x"01430400",
         15870 => x"00000000",
         15871 => x"00000000",
         15872 => x"0000e6bc",
         15873 => x"01500500",
         15874 => x"00000000",
         15875 => x"00000000",
         15876 => x"0000e6c0",
         15877 => x"01510500",
         15878 => x"00000000",
         15879 => x"00000000",
         15880 => x"0000e6c4",
         15881 => x"01540500",
         15882 => x"00000000",
         15883 => x"00000000",
         15884 => x"0000e6c8",
         15885 => x"01550500",
         15886 => x"00000000",
         15887 => x"00000000",
         15888 => x"0000e6cc",
         15889 => x"01790700",
         15890 => x"00000000",
         15891 => x"00000000",
         15892 => x"0000e6d4",
         15893 => x"01780700",
         15894 => x"00000000",
         15895 => x"00000000",
         15896 => x"0000e6d8",
         15897 => x"01820800",
         15898 => x"00000000",
         15899 => x"00000000",
         15900 => x"0000e6e0",
         15901 => x"01830800",
         15902 => x"00000000",
         15903 => x"00000000",
         15904 => x"0000e6e8",
         15905 => x"01850800",
         15906 => x"00000000",
         15907 => x"00000000",
         15908 => x"0000e6f0",
         15909 => x"01870800",
         15910 => x"00000000",
         15911 => x"00000000",
         15912 => x"0000e6f8",
         15913 => x"01880800",
         15914 => x"00000000",
         15915 => x"00000000",
         15916 => x"0000e6fc",
         15917 => x"01890800",
         15918 => x"00000000",
         15919 => x"00000000",
         15920 => x"0000e700",
         15921 => x"018c0900",
         15922 => x"00000000",
         15923 => x"00000000",
         15924 => x"0000e708",
         15925 => x"018d0900",
         15926 => x"00000000",
         15927 => x"00000000",
         15928 => x"0000e710",
         15929 => x"018e0900",
         15930 => x"00000000",
         15931 => x"00000000",
         15932 => x"0000e718",
         15933 => x"018f0900",
         15934 => x"00000000",
         15935 => x"00000000",
         15936 => x"00000000",
         15937 => x"00000000",
         15938 => x"00007fff",
         15939 => x"00000000",
         15940 => x"00007fff",
         15941 => x"00010000",
         15942 => x"00007fff",
         15943 => x"00010000",
         15944 => x"00810000",
         15945 => x"01000000",
         15946 => x"017fffff",
         15947 => x"00000000",
         15948 => x"00000000",
         15949 => x"00007800",
         15950 => x"00000000",
         15951 => x"05f5e100",
         15952 => x"05f5e100",
         15953 => x"05f5e100",
         15954 => x"00000000",
         15955 => x"01010101",
         15956 => x"01010101",
         15957 => x"01011001",
         15958 => x"01000000",
         15959 => x"00000000",
         15960 => x"00000000",
         15961 => x"00000000",
         15962 => x"00000000",
         15963 => x"00000000",
         15964 => x"00000000",
         15965 => x"00000000",
         15966 => x"00000000",
         15967 => x"00000000",
         15968 => x"00000000",
         15969 => x"00000000",
         15970 => x"00000000",
         15971 => x"00000000",
         15972 => x"00000000",
         15973 => x"00000000",
         15974 => x"00000000",
         15975 => x"00000000",
         15976 => x"00000000",
         15977 => x"00000000",
         15978 => x"00000000",
         15979 => x"00000000",
         15980 => x"00000000",
         15981 => x"00000000",
         15982 => x"00000000",
         15983 => x"0000f0dc",
         15984 => x"01000000",
         15985 => x"0000f0e4",
         15986 => x"01000000",
         15987 => x"0000f0ec",
         15988 => x"02000000",
         15989 => x"0001fd80",
         15990 => x"1bfc5ffd",
         15991 => x"f03b3a0d",
         15992 => x"797a405b",
         15993 => x"5df0f0f0",
         15994 => x"71727374",
         15995 => x"75767778",
         15996 => x"696a6b6c",
         15997 => x"6d6e6f70",
         15998 => x"61626364",
         15999 => x"65666768",
         16000 => x"31323334",
         16001 => x"35363738",
         16002 => x"5cf32d20",
         16003 => x"30392c2e",
         16004 => x"f67ff3f4",
         16005 => x"f1f23f2f",
         16006 => x"08f0f0f0",
         16007 => x"f0f0f0f0",
         16008 => x"80818283",
         16009 => x"84f0f0f0",
         16010 => x"1bfc58fd",
         16011 => x"f03a3b0d",
         16012 => x"595a405b",
         16013 => x"5df0f0f0",
         16014 => x"51525354",
         16015 => x"55565758",
         16016 => x"494a4b4c",
         16017 => x"4d4e4f50",
         16018 => x"41424344",
         16019 => x"45464748",
         16020 => x"31323334",
         16021 => x"35363738",
         16022 => x"5cf32d20",
         16023 => x"30392c2e",
         16024 => x"f67ff3f4",
         16025 => x"f1f23f2f",
         16026 => x"08f0f0f0",
         16027 => x"f0f0f0f0",
         16028 => x"80818283",
         16029 => x"84f0f0f0",
         16030 => x"1bfc58fd",
         16031 => x"f02b2a0d",
         16032 => x"595a607b",
         16033 => x"7df0f0f0",
         16034 => x"51525354",
         16035 => x"55565758",
         16036 => x"494a4b4c",
         16037 => x"4d4e4f50",
         16038 => x"41424344",
         16039 => x"45464748",
         16040 => x"21222324",
         16041 => x"25262728",
         16042 => x"7c7e3d20",
         16043 => x"20293c3e",
         16044 => x"f7e2e0e1",
         16045 => x"f9f83f2f",
         16046 => x"fbf0f0f0",
         16047 => x"f0f0f0f0",
         16048 => x"85868788",
         16049 => x"89f0f0f0",
         16050 => x"1bfe1efa",
         16051 => x"f0f0f0f0",
         16052 => x"191a001b",
         16053 => x"1df0f0f0",
         16054 => x"11121314",
         16055 => x"15161718",
         16056 => x"090a0b0c",
         16057 => x"0d0e0f10",
         16058 => x"01020304",
         16059 => x"05060708",
         16060 => x"f0f0f0f0",
         16061 => x"f0f0f0f0",
         16062 => x"f01ef0f0",
         16063 => x"f01ff0f0",
         16064 => x"f0f0f0f0",
         16065 => x"f0f0f01c",
         16066 => x"f0f0f0f0",
         16067 => x"f0f0f0f0",
         16068 => x"80818283",
         16069 => x"84f0f0f0",
         16070 => x"bff0cfc9",
         16071 => x"f0b54dcd",
         16072 => x"3577d7b3",
         16073 => x"b7f0f0f0",
         16074 => x"7c704131",
         16075 => x"39a678dd",
         16076 => x"3d5d6c56",
         16077 => x"1d33d5b1",
         16078 => x"466ed948",
         16079 => x"74434c73",
         16080 => x"3f367e3b",
         16081 => x"7a1e5fa2",
         16082 => x"d39fd100",
         16083 => x"9da3d0b9",
         16084 => x"c6c5c2c1",
         16085 => x"c3c4bbbe",
         16086 => x"f0f0f0f0",
         16087 => x"f0f0f0f0",
         16088 => x"80818283",
         16089 => x"84f0f0f0",
         16090 => x"00000000",
         16091 => x"00000000",
         16092 => x"00000000",
         16093 => x"00000000",
         16094 => x"00000000",
         16095 => x"00000000",
         16096 => x"00000000",
         16097 => x"00000000",
         16098 => x"00000000",
         16099 => x"00000000",
         16100 => x"00000000",
         16101 => x"00000000",
         16102 => x"00000000",
         16103 => x"00000000",
         16104 => x"00000000",
         16105 => x"00000000",
         16106 => x"00000000",
         16107 => x"00000000",
         16108 => x"00000000",
         16109 => x"00000000",
         16110 => x"00000000",
         16111 => x"00000000",
         16112 => x"00000000",
         16113 => x"00000000",
         16114 => x"00000000",
         16115 => x"00010000",
         16116 => x"00000000",
         16117 => x"f8000000",
         16118 => x"0000f130",
         16119 => x"f3000000",
         16120 => x"0000f138",
         16121 => x"f4000000",
         16122 => x"0000f13c",
         16123 => x"f1000000",
         16124 => x"0000f140",
         16125 => x"f2000000",
         16126 => x"0000f144",
         16127 => x"80000000",
         16128 => x"0000f148",
         16129 => x"81000000",
         16130 => x"0000f150",
         16131 => x"82000000",
         16132 => x"0000f158",
         16133 => x"83000000",
         16134 => x"0000f160",
         16135 => x"84000000",
         16136 => x"0000f168",
         16137 => x"85000000",
         16138 => x"0000f170",
         16139 => x"86000000",
         16140 => x"0000f178",
         16141 => x"87000000",
         16142 => x"0000f180",
         16143 => x"88000000",
         16144 => x"0000f188",
         16145 => x"89000000",
         16146 => x"0000f190",
         16147 => x"f6000000",
         16148 => x"0000f198",
         16149 => x"7f000000",
         16150 => x"0000f1a0",
         16151 => x"f9000000",
         16152 => x"0000f1a8",
         16153 => x"e0000000",
         16154 => x"0000f1ac",
         16155 => x"e1000000",
         16156 => x"0000f1b4",
         16157 => x"71000000",
         16158 => x"00000000",
         16159 => x"00000000",
         16160 => x"00000000",
         16161 => x"00000000",
         16162 => x"00000000",
         16163 => x"00000000",
         16164 => x"00000000",
         16165 => x"00000000",
         16166 => x"00000000",
         16167 => x"00000000",
         16168 => x"00000000",
         16169 => x"00000000",
         16170 => x"00000000",
         16171 => x"00000000",
         16172 => x"00000000",
         16173 => x"00000000",
         16174 => x"00000000",
         16175 => x"00000000",
         16176 => x"00000000",
         16177 => x"00000000",
         16178 => x"00000000",
         16179 => x"00000000",
         16180 => x"00000000",
         16181 => x"00000000",
         16182 => x"00000000",
         16183 => x"00000000",
         16184 => x"00000000",
         16185 => x"00000000",
         16186 => x"00000000",
         16187 => x"00000000",
         16188 => x"00000000",
         16189 => x"00000000",
         16190 => x"00000000",
         16191 => x"00000000",
         16192 => x"00000000",
         16193 => x"00000000",
         16194 => x"00000000",
         16195 => x"00000000",
         16196 => x"00000000",
         16197 => x"00000000",
         16198 => x"00000000",
         16199 => x"00000000",
         16200 => x"00000000",
         16201 => x"00000000",
         16202 => x"00000000",
         16203 => x"00000000",
         16204 => x"00000000",
         16205 => x"00000000",
         16206 => x"00000000",
         16207 => x"00000000",
         16208 => x"00000000",
         16209 => x"00000000",
         16210 => x"00000000",
         16211 => x"00000000",
         16212 => x"00000000",
         16213 => x"00000000",
         16214 => x"00000000",
         16215 => x"00000000",
         16216 => x"00000000",
         16217 => x"00000000",
         16218 => x"00000000",
         16219 => x"00000000",
         16220 => x"00000000",
         16221 => x"00000000",
         16222 => x"00000000",
         16223 => x"00000000",
         16224 => x"00000000",
         16225 => x"00000000",
         16226 => x"00000000",
         16227 => x"00000000",
         16228 => x"00000000",
         16229 => x"00000000",
         16230 => x"00000000",
         16231 => x"00000000",
         16232 => x"00000000",
         16233 => x"00000000",
         16234 => x"00000000",
         16235 => x"00000000",
         16236 => x"00000000",
         16237 => x"00000000",
         16238 => x"00000000",
         16239 => x"00000000",
         16240 => x"00000000",
         16241 => x"00000000",
         16242 => x"00000000",
         16243 => x"00000000",
         16244 => x"00000000",
         16245 => x"00000000",
         16246 => x"00000000",
         16247 => x"00000000",
         16248 => x"00000000",
         16249 => x"00000000",
         16250 => x"00000000",
         16251 => x"00000000",
         16252 => x"00000000",
         16253 => x"00000000",
         16254 => x"00000000",
         16255 => x"00000000",
         16256 => x"00000000",
         16257 => x"00000000",
         16258 => x"00000000",
         16259 => x"00000000",
         16260 => x"00000000",
         16261 => x"00000000",
         16262 => x"00000000",
         16263 => x"00000000",
         16264 => x"00000000",
         16265 => x"00000000",
         16266 => x"00000000",
         16267 => x"00000000",
         16268 => x"00000000",
         16269 => x"00000000",
         16270 => x"00000000",
         16271 => x"00000000",
         16272 => x"00000000",
         16273 => x"00000000",
         16274 => x"00000000",
         16275 => x"00000000",
         16276 => x"00000000",
         16277 => x"00000000",
         16278 => x"00000000",
         16279 => x"00000000",
         16280 => x"00000000",
         16281 => x"00000000",
         16282 => x"00000000",
         16283 => x"00000000",
         16284 => x"00000000",
         16285 => x"00000000",
         16286 => x"00000000",
         16287 => x"00000000",
         16288 => x"00000000",
         16289 => x"00000000",
         16290 => x"00000000",
         16291 => x"00000000",
         16292 => x"00000000",
         16293 => x"00000000",
         16294 => x"00000000",
         16295 => x"00000000",
         16296 => x"00000000",
         16297 => x"00000000",
         16298 => x"00000000",
         16299 => x"00000000",
         16300 => x"00000000",
         16301 => x"00000000",
         16302 => x"00000000",
         16303 => x"00000000",
         16304 => x"00000000",
         16305 => x"00000000",
         16306 => x"00000000",
         16307 => x"00000000",
         16308 => x"00000000",
         16309 => x"00000000",
         16310 => x"00000000",
         16311 => x"00000000",
         16312 => x"00000000",
         16313 => x"00000000",
         16314 => x"00000000",
         16315 => x"00000000",
         16316 => x"00000000",
         16317 => x"00000000",
         16318 => x"00000000",
         16319 => x"00000000",
         16320 => x"00000000",
         16321 => x"00000000",
         16322 => x"00000000",
         16323 => x"00000000",
         16324 => x"00000000",
         16325 => x"00000000",
         16326 => x"00000000",
         16327 => x"00000000",
         16328 => x"00000000",
         16329 => x"00000000",
         16330 => x"00000000",
         16331 => x"00000000",
         16332 => x"00000000",
         16333 => x"00000000",
         16334 => x"00000000",
         16335 => x"00000000",
         16336 => x"00000000",
         16337 => x"00000000",
         16338 => x"00000000",
         16339 => x"00000000",
         16340 => x"00000000",
         16341 => x"00000000",
         16342 => x"00000000",
         16343 => x"00000000",
         16344 => x"00000000",
         16345 => x"00000000",
         16346 => x"00000000",
         16347 => x"00000000",
         16348 => x"00000000",
         16349 => x"00000000",
         16350 => x"00000000",
         16351 => x"00000000",
         16352 => x"00000000",
         16353 => x"00000000",
         16354 => x"00000000",
         16355 => x"00000000",
         16356 => x"00000000",
         16357 => x"00000000",
         16358 => x"00000000",
         16359 => x"00000000",
         16360 => x"00000000",
         16361 => x"00000000",
         16362 => x"00000000",
         16363 => x"00000000",
         16364 => x"00000000",
         16365 => x"00000000",
         16366 => x"00000000",
         16367 => x"00000000",
         16368 => x"00000000",
         16369 => x"00000000",
         16370 => x"00000000",
         16371 => x"00000000",
         16372 => x"00000000",
         16373 => x"00000000",
         16374 => x"00000000",
         16375 => x"00000000",
         16376 => x"00000000",
         16377 => x"00000000",
         16378 => x"00000000",
         16379 => x"00000000",
         16380 => x"00000000",
         16381 => x"00000000",
         16382 => x"00000000",
         16383 => x"00000000",
         16384 => x"00000000",
         16385 => x"00000000",
         16386 => x"00000000",
         16387 => x"00000000",
         16388 => x"00000000",
         16389 => x"00000000",
         16390 => x"00000000",
         16391 => x"00000000",
         16392 => x"00000000",
         16393 => x"00000000",
         16394 => x"00000000",
         16395 => x"00000000",
         16396 => x"00000000",
         16397 => x"00000000",
         16398 => x"00000000",
         16399 => x"00000000",
         16400 => x"00000000",
         16401 => x"00000000",
         16402 => x"00000000",
         16403 => x"00000000",
         16404 => x"00000000",
         16405 => x"00000000",
         16406 => x"00000000",
         16407 => x"00000000",
         16408 => x"00000000",
         16409 => x"00000000",
         16410 => x"00000000",
         16411 => x"00000000",
         16412 => x"00000000",
         16413 => x"00000000",
         16414 => x"00000000",
         16415 => x"00000000",
         16416 => x"00000000",
         16417 => x"00000000",
         16418 => x"00000000",
         16419 => x"00000000",
         16420 => x"00000000",
         16421 => x"00000000",
         16422 => x"00000000",
         16423 => x"00000000",
         16424 => x"00000000",
         16425 => x"00000000",
         16426 => x"00000000",
         16427 => x"00000000",
         16428 => x"00000000",
         16429 => x"00000000",
         16430 => x"00000000",
         16431 => x"00000000",
         16432 => x"00000000",
         16433 => x"00000000",
         16434 => x"00000000",
         16435 => x"00000000",
         16436 => x"00000000",
         16437 => x"00000000",
         16438 => x"00000000",
         16439 => x"00000000",
         16440 => x"00000000",
         16441 => x"00000000",
         16442 => x"00000000",
         16443 => x"00000000",
         16444 => x"00000000",
         16445 => x"00000000",
         16446 => x"00000000",
         16447 => x"00000000",
         16448 => x"00000000",
         16449 => x"00000000",
         16450 => x"00000000",
         16451 => x"00000000",
         16452 => x"00000000",
         16453 => x"00000000",
         16454 => x"00000000",
         16455 => x"00000000",
         16456 => x"00000000",
         16457 => x"00000000",
         16458 => x"00000000",
         16459 => x"00000000",
         16460 => x"00000000",
         16461 => x"00000000",
         16462 => x"00000000",
         16463 => x"00000000",
         16464 => x"00000000",
         16465 => x"00000000",
         16466 => x"00000000",
         16467 => x"00000000",
         16468 => x"00000000",
         16469 => x"00000000",
         16470 => x"00000000",
         16471 => x"00000000",
         16472 => x"00000000",
         16473 => x"00000000",
         16474 => x"00000000",
         16475 => x"00000000",
         16476 => x"00000000",
         16477 => x"00000000",
         16478 => x"00000000",
         16479 => x"00000000",
         16480 => x"00000000",
         16481 => x"00000000",
         16482 => x"00000000",
         16483 => x"00000000",
         16484 => x"00000000",
         16485 => x"00000000",
         16486 => x"00000000",
         16487 => x"00000000",
         16488 => x"00000000",
         16489 => x"00000000",
         16490 => x"00000000",
         16491 => x"00000000",
         16492 => x"00000000",
         16493 => x"00000000",
         16494 => x"00000000",
         16495 => x"00000000",
         16496 => x"00000000",
         16497 => x"00000000",
         16498 => x"00000000",
         16499 => x"00000000",
         16500 => x"00000000",
         16501 => x"00000000",
         16502 => x"00000000",
         16503 => x"00000000",
         16504 => x"00000000",
         16505 => x"00000000",
         16506 => x"00000000",
         16507 => x"00000000",
         16508 => x"00000000",
         16509 => x"00000000",
         16510 => x"00000000",
         16511 => x"00000000",
         16512 => x"00000000",
         16513 => x"00000000",
         16514 => x"00000000",
         16515 => x"00000000",
         16516 => x"00000000",
         16517 => x"00000000",
         16518 => x"00000000",
         16519 => x"00000000",
         16520 => x"00000000",
         16521 => x"00000000",
         16522 => x"00000000",
         16523 => x"00000000",
         16524 => x"00000000",
         16525 => x"00000000",
         16526 => x"00000000",
         16527 => x"00000000",
         16528 => x"00000000",
         16529 => x"00000000",
         16530 => x"00000000",
         16531 => x"00000000",
         16532 => x"00000000",
         16533 => x"00000000",
         16534 => x"00000000",
         16535 => x"00000000",
         16536 => x"00000000",
         16537 => x"00000000",
         16538 => x"00000000",
         16539 => x"00000000",
         16540 => x"00000000",
         16541 => x"00000000",
         16542 => x"00000000",
         16543 => x"00000000",
         16544 => x"00000000",
         16545 => x"00000000",
         16546 => x"00000000",
         16547 => x"00000000",
         16548 => x"00000000",
         16549 => x"00000000",
         16550 => x"00000000",
         16551 => x"00000000",
         16552 => x"00000000",
         16553 => x"00000000",
         16554 => x"00000000",
         16555 => x"00000000",
         16556 => x"00000000",
         16557 => x"00000000",
         16558 => x"00000000",
         16559 => x"00000000",
         16560 => x"00000000",
         16561 => x"00000000",
         16562 => x"00000000",
         16563 => x"00000000",
         16564 => x"00000000",
         16565 => x"00000000",
         16566 => x"00000000",
         16567 => x"00000000",
         16568 => x"00000000",
         16569 => x"00000000",
         16570 => x"00000000",
         16571 => x"00000000",
         16572 => x"00000000",
         16573 => x"00000000",
         16574 => x"00000000",
         16575 => x"00000000",
         16576 => x"00000000",
         16577 => x"00000000",
         16578 => x"00000000",
         16579 => x"00000000",
         16580 => x"00000000",
         16581 => x"00000000",
         16582 => x"00000000",
         16583 => x"00000000",
         16584 => x"00000000",
         16585 => x"00000000",
         16586 => x"00000000",
         16587 => x"00000000",
         16588 => x"00000000",
         16589 => x"00000000",
         16590 => x"00000000",
         16591 => x"00000000",
         16592 => x"00000000",
         16593 => x"00000000",
         16594 => x"00000000",
         16595 => x"00000000",
         16596 => x"00000000",
         16597 => x"00000000",
         16598 => x"00000000",
         16599 => x"00000000",
         16600 => x"00000000",
         16601 => x"00000000",
         16602 => x"00000000",
         16603 => x"00000000",
         16604 => x"00000000",
         16605 => x"00000000",
         16606 => x"00000000",
         16607 => x"00000000",
         16608 => x"00000000",
         16609 => x"00000000",
         16610 => x"00000000",
         16611 => x"00000000",
         16612 => x"00000000",
         16613 => x"00000000",
         16614 => x"00000000",
         16615 => x"00000000",
         16616 => x"00000000",
         16617 => x"00000000",
         16618 => x"00000000",
         16619 => x"00000000",
         16620 => x"00000000",
         16621 => x"00000000",
         16622 => x"00000000",
         16623 => x"00000000",
         16624 => x"00000000",
         16625 => x"00000000",
         16626 => x"00000000",
         16627 => x"00000000",
         16628 => x"00000000",
         16629 => x"00000000",
         16630 => x"00000000",
         16631 => x"00000000",
         16632 => x"00000000",
         16633 => x"00000000",
         16634 => x"00000000",
         16635 => x"00000000",
         16636 => x"00000000",
         16637 => x"00000000",
         16638 => x"00000000",
         16639 => x"00000000",
         16640 => x"00000000",
         16641 => x"00000000",
         16642 => x"00000000",
         16643 => x"00000000",
         16644 => x"00000000",
         16645 => x"00000000",
         16646 => x"00000000",
         16647 => x"00000000",
         16648 => x"00000000",
         16649 => x"00000000",
         16650 => x"00000000",
         16651 => x"00000000",
         16652 => x"00000000",
         16653 => x"00000000",
         16654 => x"00000000",
         16655 => x"00000000",
         16656 => x"00000000",
         16657 => x"00000000",
         16658 => x"00000000",
         16659 => x"00000000",
         16660 => x"00000000",
         16661 => x"00000000",
         16662 => x"00000000",
         16663 => x"00000000",
         16664 => x"00000000",
         16665 => x"00000000",
         16666 => x"00000000",
         16667 => x"00000000",
         16668 => x"00000000",
         16669 => x"00000000",
         16670 => x"00000000",
         16671 => x"00000000",
         16672 => x"00000000",
         16673 => x"00000000",
         16674 => x"00000000",
         16675 => x"00000000",
         16676 => x"00000000",
         16677 => x"00000000",
         16678 => x"00000000",
         16679 => x"00000000",
         16680 => x"00000000",
         16681 => x"00000000",
         16682 => x"00000000",
         16683 => x"00000000",
         16684 => x"00000000",
         16685 => x"00000000",
         16686 => x"00000000",
         16687 => x"00000000",
         16688 => x"00000000",
         16689 => x"00000000",
         16690 => x"00000000",
         16691 => x"00000000",
         16692 => x"00000000",
         16693 => x"00000000",
         16694 => x"00000000",
         16695 => x"00000000",
         16696 => x"00000000",
         16697 => x"00000000",
         16698 => x"00000000",
         16699 => x"00000000",
         16700 => x"00000000",
         16701 => x"00000000",
         16702 => x"00000000",
         16703 => x"00000000",
         16704 => x"00000000",
         16705 => x"00000000",
         16706 => x"00000000",
         16707 => x"00000000",
         16708 => x"00000000",
         16709 => x"00000000",
         16710 => x"00000000",
         16711 => x"00000000",
         16712 => x"00000000",
         16713 => x"00000000",
         16714 => x"00000000",
         16715 => x"00000000",
         16716 => x"00000000",
         16717 => x"00000000",
         16718 => x"00000000",
         16719 => x"00000000",
         16720 => x"00000000",
         16721 => x"00000000",
         16722 => x"00000000",
         16723 => x"00000000",
         16724 => x"00000000",
         16725 => x"00000000",
         16726 => x"00000000",
         16727 => x"00000000",
         16728 => x"00000000",
         16729 => x"00000000",
         16730 => x"00000000",
         16731 => x"00000000",
         16732 => x"00000000",
         16733 => x"00000000",
         16734 => x"00000000",
         16735 => x"00000000",
         16736 => x"00000000",
         16737 => x"00000000",
         16738 => x"00000000",
         16739 => x"00000000",
         16740 => x"00000000",
         16741 => x"00000000",
         16742 => x"00000000",
         16743 => x"00000000",
         16744 => x"00000000",
         16745 => x"00000000",
         16746 => x"00000000",
         16747 => x"00000000",
         16748 => x"00000000",
         16749 => x"00000000",
         16750 => x"00000000",
         16751 => x"00000000",
         16752 => x"00000000",
         16753 => x"00000000",
         16754 => x"00000000",
         16755 => x"00000000",
         16756 => x"00000000",
         16757 => x"00000000",
         16758 => x"00000000",
         16759 => x"00000000",
         16760 => x"00000000",
         16761 => x"00000000",
         16762 => x"00000000",
         16763 => x"00000000",
         16764 => x"00000000",
         16765 => x"00000000",
         16766 => x"00000000",
         16767 => x"00000000",
         16768 => x"00000000",
         16769 => x"00000000",
         16770 => x"00000000",
         16771 => x"00000000",
         16772 => x"00000000",
         16773 => x"00000000",
         16774 => x"00000000",
         16775 => x"00000000",
         16776 => x"00000000",
         16777 => x"00000000",
         16778 => x"00000000",
         16779 => x"00000000",
         16780 => x"00000000",
         16781 => x"00000000",
         16782 => x"00000000",
         16783 => x"00000000",
         16784 => x"00000000",
         16785 => x"00000000",
         16786 => x"00000000",
         16787 => x"00000000",
         16788 => x"00000000",
         16789 => x"00000000",
         16790 => x"00000000",
         16791 => x"00000000",
         16792 => x"00000000",
         16793 => x"00000000",
         16794 => x"00000000",
         16795 => x"00000000",
         16796 => x"00000000",
         16797 => x"00000000",
         16798 => x"00000000",
         16799 => x"00000000",
         16800 => x"00000000",
         16801 => x"00000000",
         16802 => x"00000000",
         16803 => x"00000000",
         16804 => x"00000000",
         16805 => x"00000000",
         16806 => x"00000000",
         16807 => x"00000000",
         16808 => x"00000000",
         16809 => x"00000000",
         16810 => x"00000000",
         16811 => x"00000000",
         16812 => x"00000000",
         16813 => x"00000000",
         16814 => x"00000000",
         16815 => x"00000000",
         16816 => x"00000000",
         16817 => x"00000000",
         16818 => x"00000000",
         16819 => x"00000000",
         16820 => x"00000000",
         16821 => x"00000000",
         16822 => x"00000000",
         16823 => x"00000000",
         16824 => x"00000000",
         16825 => x"00000000",
         16826 => x"00000000",
         16827 => x"00000000",
         16828 => x"00000000",
         16829 => x"00000000",
         16830 => x"00000000",
         16831 => x"00000000",
         16832 => x"00000000",
         16833 => x"00000000",
         16834 => x"00000000",
         16835 => x"00000000",
         16836 => x"00000000",
         16837 => x"00000000",
         16838 => x"00000000",
         16839 => x"00000000",
         16840 => x"00000000",
         16841 => x"00000000",
         16842 => x"00000000",
         16843 => x"00000000",
         16844 => x"00000000",
         16845 => x"00000000",
         16846 => x"00000000",
         16847 => x"00000000",
         16848 => x"00000000",
         16849 => x"00000000",
         16850 => x"00000000",
         16851 => x"00000000",
         16852 => x"00000000",
         16853 => x"00000000",
         16854 => x"00000000",
         16855 => x"00000000",
         16856 => x"00000000",
         16857 => x"00000000",
         16858 => x"00000000",
         16859 => x"00000000",
         16860 => x"00000000",
         16861 => x"00000000",
         16862 => x"00000000",
         16863 => x"00000000",
         16864 => x"00000000",
         16865 => x"00000000",
         16866 => x"00000000",
         16867 => x"00000000",
         16868 => x"00000000",
         16869 => x"00000000",
         16870 => x"00000000",
         16871 => x"00000000",
         16872 => x"00000000",
         16873 => x"00000000",
         16874 => x"00000000",
         16875 => x"00000000",
         16876 => x"00000000",
         16877 => x"00000000",
         16878 => x"00000000",
         16879 => x"00000000",
         16880 => x"00000000",
         16881 => x"00000000",
         16882 => x"00000000",
         16883 => x"00000000",
         16884 => x"00000000",
         16885 => x"00000000",
         16886 => x"00000000",
         16887 => x"00000000",
         16888 => x"00000000",
         16889 => x"00000000",
         16890 => x"00000000",
         16891 => x"00000000",
         16892 => x"00000000",
         16893 => x"00000000",
         16894 => x"00000000",
         16895 => x"00000000",
         16896 => x"00000000",
         16897 => x"00000000",
         16898 => x"00000000",
         16899 => x"00000000",
         16900 => x"00000000",
         16901 => x"00000000",
         16902 => x"00000000",
         16903 => x"00000000",
         16904 => x"00000000",
         16905 => x"00000000",
         16906 => x"00000000",
         16907 => x"00000000",
         16908 => x"00000000",
         16909 => x"00000000",
         16910 => x"00000000",
         16911 => x"00000000",
         16912 => x"00000000",
         16913 => x"00000000",
         16914 => x"00000000",
         16915 => x"00000000",
         16916 => x"00000000",
         16917 => x"00000000",
         16918 => x"00000000",
         16919 => x"00000000",
         16920 => x"00000000",
         16921 => x"00000000",
         16922 => x"00000000",
         16923 => x"00000000",
         16924 => x"00000000",
         16925 => x"00000000",
         16926 => x"00000000",
         16927 => x"00000000",
         16928 => x"00000000",
         16929 => x"00000000",
         16930 => x"00000000",
         16931 => x"00000000",
         16932 => x"00000000",
         16933 => x"00000000",
         16934 => x"00000000",
         16935 => x"00000000",
         16936 => x"00000000",
         16937 => x"00000000",
         16938 => x"00000000",
         16939 => x"00000000",
         16940 => x"00000000",
         16941 => x"00000000",
         16942 => x"00000000",
         16943 => x"00000000",
         16944 => x"00000000",
         16945 => x"00000000",
         16946 => x"00000000",
         16947 => x"00000000",
         16948 => x"00000000",
         16949 => x"00000000",
         16950 => x"00000000",
         16951 => x"00000000",
         16952 => x"00000000",
         16953 => x"00000000",
         16954 => x"00000000",
         16955 => x"00000000",
         16956 => x"00000000",
         16957 => x"00000000",
         16958 => x"00000000",
         16959 => x"00000000",
         16960 => x"00000000",
         16961 => x"00000000",
         16962 => x"00000000",
         16963 => x"00000000",
         16964 => x"00000000",
         16965 => x"00000000",
         16966 => x"00000000",
         16967 => x"00000000",
         16968 => x"00000000",
         16969 => x"00000000",
         16970 => x"00000000",
         16971 => x"00000000",
         16972 => x"00000000",
         16973 => x"00000000",
         16974 => x"00000000",
         16975 => x"00000000",
         16976 => x"00000000",
         16977 => x"00000000",
         16978 => x"00000000",
         16979 => x"00000000",
         16980 => x"00000000",
         16981 => x"00000000",
         16982 => x"00000000",
         16983 => x"00000000",
         16984 => x"00000000",
         16985 => x"00000000",
         16986 => x"00000000",
         16987 => x"00000000",
         16988 => x"00000000",
         16989 => x"00000000",
         16990 => x"00000000",
         16991 => x"00000000",
         16992 => x"00000000",
         16993 => x"00000000",
         16994 => x"00000000",
         16995 => x"00000000",
         16996 => x"00000000",
         16997 => x"00000000",
         16998 => x"00000000",
         16999 => x"00000000",
         17000 => x"00000000",
         17001 => x"00000000",
         17002 => x"00000000",
         17003 => x"00000000",
         17004 => x"00000000",
         17005 => x"00000000",
         17006 => x"00000000",
         17007 => x"00000000",
         17008 => x"00000000",
         17009 => x"00000000",
         17010 => x"00000000",
         17011 => x"00000000",
         17012 => x"00000000",
         17013 => x"00000000",
         17014 => x"00000000",
         17015 => x"00000000",
         17016 => x"00000000",
         17017 => x"00000000",
         17018 => x"00000000",
         17019 => x"00000000",
         17020 => x"00000000",
         17021 => x"00000000",
         17022 => x"00000000",
         17023 => x"00000000",
         17024 => x"00000000",
         17025 => x"00000000",
         17026 => x"00000000",
         17027 => x"00000000",
         17028 => x"00000000",
         17029 => x"00000000",
         17030 => x"00000000",
         17031 => x"00000000",
         17032 => x"00000000",
         17033 => x"00000000",
         17034 => x"00000000",
         17035 => x"00000000",
         17036 => x"00000000",
         17037 => x"00000000",
         17038 => x"00000000",
         17039 => x"00000000",
         17040 => x"00000000",
         17041 => x"00000000",
         17042 => x"00000000",
         17043 => x"00000000",
         17044 => x"00000000",
         17045 => x"00000000",
         17046 => x"00000000",
         17047 => x"00000000",
         17048 => x"00000000",
         17049 => x"00000000",
         17050 => x"00000000",
         17051 => x"00000000",
         17052 => x"00000000",
         17053 => x"00000000",
         17054 => x"00000000",
         17055 => x"00000000",
         17056 => x"00000000",
         17057 => x"00000000",
         17058 => x"00000000",
         17059 => x"00000000",
         17060 => x"00000000",
         17061 => x"00000000",
         17062 => x"00000000",
         17063 => x"00000000",
         17064 => x"00000000",
         17065 => x"00000000",
         17066 => x"00000000",
         17067 => x"00000000",
         17068 => x"00000000",
         17069 => x"00000000",
         17070 => x"00000000",
         17071 => x"00000000",
         17072 => x"00000000",
         17073 => x"00000000",
         17074 => x"00000000",
         17075 => x"00000000",
         17076 => x"00000000",
         17077 => x"00000000",
         17078 => x"00000000",
         17079 => x"00000000",
         17080 => x"00000000",
         17081 => x"00000000",
         17082 => x"00000000",
         17083 => x"00000000",
         17084 => x"00000000",
         17085 => x"00000000",
         17086 => x"00000000",
         17087 => x"00000000",
         17088 => x"00000000",
         17089 => x"00000000",
         17090 => x"00000000",
         17091 => x"00000000",
         17092 => x"00000000",
         17093 => x"00000000",
         17094 => x"00000000",
         17095 => x"00000000",
         17096 => x"00000000",
         17097 => x"00000000",
         17098 => x"00000000",
         17099 => x"00000000",
         17100 => x"00000000",
         17101 => x"00000000",
         17102 => x"00000000",
         17103 => x"00000000",
         17104 => x"00000000",
         17105 => x"00000000",
         17106 => x"00000000",
         17107 => x"00000000",
         17108 => x"00000000",
         17109 => x"00000000",
         17110 => x"00000000",
         17111 => x"00000000",
         17112 => x"00000000",
         17113 => x"00000000",
         17114 => x"00000000",
         17115 => x"00000000",
         17116 => x"00000000",
         17117 => x"00000000",
         17118 => x"00000000",
         17119 => x"00000000",
         17120 => x"00000000",
         17121 => x"00000000",
         17122 => x"00000000",
         17123 => x"00000000",
         17124 => x"00000000",
         17125 => x"00000000",
         17126 => x"00000000",
         17127 => x"00000000",
         17128 => x"00000000",
         17129 => x"00000000",
         17130 => x"00000000",
         17131 => x"00000000",
         17132 => x"00000000",
         17133 => x"00000000",
         17134 => x"00000000",
         17135 => x"00000000",
         17136 => x"00000000",
         17137 => x"00000000",
         17138 => x"00000000",
         17139 => x"00000000",
         17140 => x"00000000",
         17141 => x"00000000",
         17142 => x"00000000",
         17143 => x"00000000",
         17144 => x"00000000",
         17145 => x"00000000",
         17146 => x"00000000",
         17147 => x"00000000",
         17148 => x"00000000",
         17149 => x"00000000",
         17150 => x"00000000",
         17151 => x"00000000",
         17152 => x"00000000",
         17153 => x"00000000",
         17154 => x"00000000",
         17155 => x"00000000",
         17156 => x"00000000",
         17157 => x"00000000",
         17158 => x"00000000",
         17159 => x"00000000",
         17160 => x"00000000",
         17161 => x"00000000",
         17162 => x"00000000",
         17163 => x"00000000",
         17164 => x"00000000",
         17165 => x"00000000",
         17166 => x"00000000",
         17167 => x"00000000",
         17168 => x"00000000",
         17169 => x"00000000",
         17170 => x"00000000",
         17171 => x"00000000",
         17172 => x"00000000",
         17173 => x"00000000",
         17174 => x"00000000",
         17175 => x"00000000",
         17176 => x"00000000",
         17177 => x"00000000",
         17178 => x"00000000",
         17179 => x"00000000",
         17180 => x"00000000",
         17181 => x"00000000",
         17182 => x"00000000",
         17183 => x"00000000",
         17184 => x"00000000",
         17185 => x"00000000",
         17186 => x"00000000",
         17187 => x"00000000",
         17188 => x"00000000",
         17189 => x"00000000",
         17190 => x"00000000",
         17191 => x"00000000",
         17192 => x"00000000",
         17193 => x"00000000",
         17194 => x"00000000",
         17195 => x"00000000",
         17196 => x"00000000",
         17197 => x"00000000",
         17198 => x"00000000",
         17199 => x"00000000",
         17200 => x"00000000",
         17201 => x"00000000",
         17202 => x"00000000",
         17203 => x"00000000",
         17204 => x"00000000",
         17205 => x"00000000",
         17206 => x"00000000",
         17207 => x"00000000",
         17208 => x"00000000",
         17209 => x"00000000",
         17210 => x"00000000",
         17211 => x"00000000",
         17212 => x"00000000",
         17213 => x"00000000",
         17214 => x"00000000",
         17215 => x"00000000",
         17216 => x"00000000",
         17217 => x"00000000",
         17218 => x"00000000",
         17219 => x"00000000",
         17220 => x"00000000",
         17221 => x"00000000",
         17222 => x"00000000",
         17223 => x"00000000",
         17224 => x"00000000",
         17225 => x"00000000",
         17226 => x"00000000",
         17227 => x"00000000",
         17228 => x"00000000",
         17229 => x"00000000",
         17230 => x"00000000",
         17231 => x"00000000",
         17232 => x"00000000",
         17233 => x"00000000",
         17234 => x"00000000",
         17235 => x"00000000",
         17236 => x"00000000",
         17237 => x"00000000",
         17238 => x"00000000",
         17239 => x"00000000",
         17240 => x"00000000",
         17241 => x"00000000",
         17242 => x"00000000",
         17243 => x"00000000",
         17244 => x"00000000",
         17245 => x"00000000",
         17246 => x"00000000",
         17247 => x"00000000",
         17248 => x"00000000",
         17249 => x"00000000",
         17250 => x"00000000",
         17251 => x"00000000",
         17252 => x"00000000",
         17253 => x"00000000",
         17254 => x"00000000",
         17255 => x"00000000",
         17256 => x"00000000",
         17257 => x"00000000",
         17258 => x"00000000",
         17259 => x"00000000",
         17260 => x"00000000",
         17261 => x"00000000",
         17262 => x"00000000",
         17263 => x"00000000",
         17264 => x"00000000",
         17265 => x"00000000",
         17266 => x"00000000",
         17267 => x"00000000",
         17268 => x"00000000",
         17269 => x"00000000",
         17270 => x"00000000",
         17271 => x"00000000",
         17272 => x"00000000",
         17273 => x"00000000",
         17274 => x"00000000",
         17275 => x"00000000",
         17276 => x"00000000",
         17277 => x"00000000",
         17278 => x"00000000",
         17279 => x"00000000",
         17280 => x"00000000",
         17281 => x"00000000",
         17282 => x"00000000",
         17283 => x"00000000",
         17284 => x"00000000",
         17285 => x"00000000",
         17286 => x"00000000",
         17287 => x"00000000",
         17288 => x"00000000",
         17289 => x"00000000",
         17290 => x"00000000",
         17291 => x"00000000",
         17292 => x"00000000",
         17293 => x"00000000",
         17294 => x"00000000",
         17295 => x"00000000",
         17296 => x"00000000",
         17297 => x"00000000",
         17298 => x"00000000",
         17299 => x"00000000",
         17300 => x"00000000",
         17301 => x"00000000",
         17302 => x"00000000",
         17303 => x"00000000",
         17304 => x"00000000",
         17305 => x"00000000",
         17306 => x"00000000",
         17307 => x"00000000",
         17308 => x"00000000",
         17309 => x"00000000",
         17310 => x"00000000",
         17311 => x"00000000",
         17312 => x"00000000",
         17313 => x"00000000",
         17314 => x"00000000",
         17315 => x"00000000",
         17316 => x"00000000",
         17317 => x"00000000",
         17318 => x"00000000",
         17319 => x"00000000",
         17320 => x"00000000",
         17321 => x"00000000",
         17322 => x"00000000",
         17323 => x"00000000",
         17324 => x"00000000",
         17325 => x"00000000",
         17326 => x"00000000",
         17327 => x"00000000",
         17328 => x"00000000",
         17329 => x"00000000",
         17330 => x"00000000",
         17331 => x"00000000",
         17332 => x"00000000",
         17333 => x"00000000",
         17334 => x"00000000",
         17335 => x"00000000",
         17336 => x"00000000",
         17337 => x"00000000",
         17338 => x"00000000",
         17339 => x"00000000",
         17340 => x"00000000",
         17341 => x"00000000",
         17342 => x"00000000",
         17343 => x"00000000",
         17344 => x"00000000",
         17345 => x"00000000",
         17346 => x"00000000",
         17347 => x"00000000",
         17348 => x"00000000",
         17349 => x"00000000",
         17350 => x"00000000",
         17351 => x"00000000",
         17352 => x"00000000",
         17353 => x"00000000",
         17354 => x"00000000",
         17355 => x"00000000",
         17356 => x"00000000",
         17357 => x"00000000",
         17358 => x"00000000",
         17359 => x"00000000",
         17360 => x"00000000",
         17361 => x"00000000",
         17362 => x"00000000",
         17363 => x"00000000",
         17364 => x"00000000",
         17365 => x"00000000",
         17366 => x"00000000",
         17367 => x"00000000",
         17368 => x"00000000",
         17369 => x"00000000",
         17370 => x"00000000",
         17371 => x"00000000",
         17372 => x"00000000",
         17373 => x"00000000",
         17374 => x"00000000",
         17375 => x"00000000",
         17376 => x"00000000",
         17377 => x"00000000",
         17378 => x"00000000",
         17379 => x"00000000",
         17380 => x"00000000",
         17381 => x"00000000",
         17382 => x"00000000",
         17383 => x"00000000",
         17384 => x"00000000",
         17385 => x"00000000",
         17386 => x"00000000",
         17387 => x"00000000",
         17388 => x"00000000",
         17389 => x"00000000",
         17390 => x"00000000",
         17391 => x"00000000",
         17392 => x"00000000",
         17393 => x"00000000",
         17394 => x"00000000",
         17395 => x"00000000",
         17396 => x"00000000",
         17397 => x"00000000",
         17398 => x"00000000",
         17399 => x"00000000",
         17400 => x"00000000",
         17401 => x"00000000",
         17402 => x"00000000",
         17403 => x"00000000",
         17404 => x"00000000",
         17405 => x"00000000",
         17406 => x"00000000",
         17407 => x"00000000",
         17408 => x"00000000",
         17409 => x"00000000",
         17410 => x"00000000",
         17411 => x"00000000",
         17412 => x"00000000",
         17413 => x"00000000",
         17414 => x"00000000",
         17415 => x"00000000",
         17416 => x"00000000",
         17417 => x"00000000",
         17418 => x"00000000",
         17419 => x"00000000",
         17420 => x"00000000",
         17421 => x"00000000",
         17422 => x"00000000",
         17423 => x"00000000",
         17424 => x"00000000",
         17425 => x"00000000",
         17426 => x"00000000",
         17427 => x"00000000",
         17428 => x"00000000",
         17429 => x"00000000",
         17430 => x"00000000",
         17431 => x"00000000",
         17432 => x"00000000",
         17433 => x"00000000",
         17434 => x"00000000",
         17435 => x"00000000",
         17436 => x"00000000",
         17437 => x"00000000",
         17438 => x"00000000",
         17439 => x"00000000",
         17440 => x"00000000",
         17441 => x"00000000",
         17442 => x"00000000",
         17443 => x"00000000",
         17444 => x"00000000",
         17445 => x"00000000",
         17446 => x"00000000",
         17447 => x"00000000",
         17448 => x"00000000",
         17449 => x"00000000",
         17450 => x"00000000",
         17451 => x"00000000",
         17452 => x"00000000",
         17453 => x"00000000",
         17454 => x"00000000",
         17455 => x"00000000",
         17456 => x"00000000",
         17457 => x"00000000",
         17458 => x"00000000",
         17459 => x"00000000",
         17460 => x"00000000",
         17461 => x"00000000",
         17462 => x"00000000",
         17463 => x"00000000",
         17464 => x"00000000",
         17465 => x"00000000",
         17466 => x"00000000",
         17467 => x"00000000",
         17468 => x"00000000",
         17469 => x"00000000",
         17470 => x"00000000",
         17471 => x"00000000",
         17472 => x"00000000",
         17473 => x"00000000",
         17474 => x"00000000",
         17475 => x"00000000",
         17476 => x"00000000",
         17477 => x"00000000",
         17478 => x"00000000",
         17479 => x"00000000",
         17480 => x"00000000",
         17481 => x"00000000",
         17482 => x"00000000",
         17483 => x"00000000",
         17484 => x"00000000",
         17485 => x"00000000",
         17486 => x"00000000",
         17487 => x"00000000",
         17488 => x"00000000",
         17489 => x"00000000",
         17490 => x"00000000",
         17491 => x"00000000",
         17492 => x"00000000",
         17493 => x"00000000",
         17494 => x"00000000",
         17495 => x"00000000",
         17496 => x"00000000",
         17497 => x"00000000",
         17498 => x"00000000",
         17499 => x"00000000",
         17500 => x"00000000",
         17501 => x"00000000",
         17502 => x"00000000",
         17503 => x"00000000",
         17504 => x"00000000",
         17505 => x"00000000",
         17506 => x"00000000",
         17507 => x"00000000",
         17508 => x"00000000",
         17509 => x"00000000",
         17510 => x"00000000",
         17511 => x"00000000",
         17512 => x"00000000",
         17513 => x"00000000",
         17514 => x"00000000",
         17515 => x"00000000",
         17516 => x"00000000",
         17517 => x"00000000",
         17518 => x"00000000",
         17519 => x"00000000",
         17520 => x"00000000",
         17521 => x"00000000",
         17522 => x"00000000",
         17523 => x"00000000",
         17524 => x"00000000",
         17525 => x"00000000",
         17526 => x"00000000",
         17527 => x"00000000",
         17528 => x"00000000",
         17529 => x"00000000",
         17530 => x"00000000",
         17531 => x"00000000",
         17532 => x"00000000",
         17533 => x"00000000",
         17534 => x"00000000",
         17535 => x"00000000",
         17536 => x"00000000",
         17537 => x"00000000",
         17538 => x"00000000",
         17539 => x"00000000",
         17540 => x"00000000",
         17541 => x"00000000",
         17542 => x"00000000",
         17543 => x"00000000",
         17544 => x"00000000",
         17545 => x"00000000",
         17546 => x"00000000",
         17547 => x"00000000",
         17548 => x"00000000",
         17549 => x"00000000",
         17550 => x"00000000",
         17551 => x"00000000",
         17552 => x"00000000",
         17553 => x"00000000",
         17554 => x"00000000",
         17555 => x"00000000",
         17556 => x"00000000",
         17557 => x"00000000",
         17558 => x"00000000",
         17559 => x"00000000",
         17560 => x"00000000",
         17561 => x"00000000",
         17562 => x"00000000",
         17563 => x"00000000",
         17564 => x"00000000",
         17565 => x"00000000",
         17566 => x"00000000",
         17567 => x"00000000",
         17568 => x"00000000",
         17569 => x"00000000",
         17570 => x"00000000",
         17571 => x"00000000",
         17572 => x"00000000",
         17573 => x"00000000",
         17574 => x"00000000",
         17575 => x"00000000",
         17576 => x"00000000",
         17577 => x"00000000",
         17578 => x"00000000",
         17579 => x"00000000",
         17580 => x"00000000",
         17581 => x"00000000",
         17582 => x"00000000",
         17583 => x"00000000",
         17584 => x"00000000",
         17585 => x"00000000",
         17586 => x"00000000",
         17587 => x"00000000",
         17588 => x"00000000",
         17589 => x"00000000",
         17590 => x"00000000",
         17591 => x"00000000",
         17592 => x"00000000",
         17593 => x"00000000",
         17594 => x"00000000",
         17595 => x"00000000",
         17596 => x"00000000",
         17597 => x"00000000",
         17598 => x"00000000",
         17599 => x"00000000",
         17600 => x"00000000",
         17601 => x"00000000",
         17602 => x"00000000",
         17603 => x"00000000",
         17604 => x"00000000",
         17605 => x"00000000",
         17606 => x"00000000",
         17607 => x"00000000",
         17608 => x"00000000",
         17609 => x"00000000",
         17610 => x"00000000",
         17611 => x"00000000",
         17612 => x"00000000",
         17613 => x"00000000",
         17614 => x"00000000",
         17615 => x"00000000",
         17616 => x"00000000",
         17617 => x"00000000",
         17618 => x"00000000",
         17619 => x"00000000",
         17620 => x"00000000",
         17621 => x"00000000",
         17622 => x"00000000",
         17623 => x"00000000",
         17624 => x"00000000",
         17625 => x"00000000",
         17626 => x"00000000",
         17627 => x"00000000",
         17628 => x"00000000",
         17629 => x"00000000",
         17630 => x"00000000",
         17631 => x"00000000",
         17632 => x"00000000",
         17633 => x"00000000",
         17634 => x"00000000",
         17635 => x"00000000",
         17636 => x"00000000",
         17637 => x"00000000",
         17638 => x"00000000",
         17639 => x"00000000",
         17640 => x"00000000",
         17641 => x"00000000",
         17642 => x"00000000",
         17643 => x"00000000",
         17644 => x"00000000",
         17645 => x"00000000",
         17646 => x"00000000",
         17647 => x"00000000",
         17648 => x"00000000",
         17649 => x"00000000",
         17650 => x"00000000",
         17651 => x"00000000",
         17652 => x"00000000",
         17653 => x"00000000",
         17654 => x"00000000",
         17655 => x"00000000",
         17656 => x"00000000",
         17657 => x"00000000",
         17658 => x"00000000",
         17659 => x"00000000",
         17660 => x"00000000",
         17661 => x"00000000",
         17662 => x"00000000",
         17663 => x"00000000",
         17664 => x"00000000",
         17665 => x"00000000",
         17666 => x"00000000",
         17667 => x"00000000",
         17668 => x"00000000",
         17669 => x"00000000",
         17670 => x"00000000",
         17671 => x"00000000",
         17672 => x"00000000",
         17673 => x"00000000",
         17674 => x"00000000",
         17675 => x"00000000",
         17676 => x"00000000",
         17677 => x"00000000",
         17678 => x"00000000",
         17679 => x"00000000",
         17680 => x"00000000",
         17681 => x"00000000",
         17682 => x"00000000",
         17683 => x"00000000",
         17684 => x"00000000",
         17685 => x"00000000",
         17686 => x"00000000",
         17687 => x"00000000",
         17688 => x"00000000",
         17689 => x"00000000",
         17690 => x"00000000",
         17691 => x"00000000",
         17692 => x"00000000",
         17693 => x"00000000",
         17694 => x"00000000",
         17695 => x"00000000",
         17696 => x"00000000",
         17697 => x"00000000",
         17698 => x"00000000",
         17699 => x"00000000",
         17700 => x"00000000",
         17701 => x"00000000",
         17702 => x"00000000",
         17703 => x"00000000",
         17704 => x"00000000",
         17705 => x"00000000",
         17706 => x"00000000",
         17707 => x"00000000",
         17708 => x"00000000",
         17709 => x"00000000",
         17710 => x"00000000",
         17711 => x"00000000",
         17712 => x"00000000",
         17713 => x"00000000",
         17714 => x"00000000",
         17715 => x"00000000",
         17716 => x"00000000",
         17717 => x"00000000",
         17718 => x"00000000",
         17719 => x"00000000",
         17720 => x"00000000",
         17721 => x"00000000",
         17722 => x"00000000",
         17723 => x"00000000",
         17724 => x"00000000",
         17725 => x"00000000",
         17726 => x"00000000",
         17727 => x"00000000",
         17728 => x"00000000",
         17729 => x"00000000",
         17730 => x"00000000",
         17731 => x"00000000",
         17732 => x"00000000",
         17733 => x"00000000",
         17734 => x"00000000",
         17735 => x"00000000",
         17736 => x"00000000",
         17737 => x"00000000",
         17738 => x"00000000",
         17739 => x"00000000",
         17740 => x"00000000",
         17741 => x"00000000",
         17742 => x"00000000",
         17743 => x"00000000",
         17744 => x"00000000",
         17745 => x"00000000",
         17746 => x"00000000",
         17747 => x"00000000",
         17748 => x"00000000",
         17749 => x"00000000",
         17750 => x"00000000",
         17751 => x"00000000",
         17752 => x"00000000",
         17753 => x"00000000",
         17754 => x"00000000",
         17755 => x"00000000",
         17756 => x"00000000",
         17757 => x"00000000",
         17758 => x"00000000",
         17759 => x"00000000",
         17760 => x"00000000",
         17761 => x"00000000",
         17762 => x"00000000",
         17763 => x"00000000",
         17764 => x"00000000",
         17765 => x"00000000",
         17766 => x"00000000",
         17767 => x"00000000",
         17768 => x"00000000",
         17769 => x"00000000",
         17770 => x"00000000",
         17771 => x"00000000",
         17772 => x"00000000",
         17773 => x"00000000",
         17774 => x"00000000",
         17775 => x"00000000",
         17776 => x"00000000",
         17777 => x"00000000",
         17778 => x"00000000",
         17779 => x"00000000",
         17780 => x"00000000",
         17781 => x"00000000",
         17782 => x"00000000",
         17783 => x"00000000",
         17784 => x"00000000",
         17785 => x"00000000",
         17786 => x"00000000",
         17787 => x"00000000",
         17788 => x"00000000",
         17789 => x"00000000",
         17790 => x"00000000",
         17791 => x"00000000",
         17792 => x"00000000",
         17793 => x"00000000",
         17794 => x"00000000",
         17795 => x"00000000",
         17796 => x"00000000",
         17797 => x"00000000",
         17798 => x"00000000",
         17799 => x"00000000",
         17800 => x"00000000",
         17801 => x"00000000",
         17802 => x"00000000",
         17803 => x"00000000",
         17804 => x"00000000",
         17805 => x"00000000",
         17806 => x"00000000",
         17807 => x"00000000",
         17808 => x"00000000",
         17809 => x"00000000",
         17810 => x"00000000",
         17811 => x"00000000",
         17812 => x"00000000",
         17813 => x"00000000",
         17814 => x"00000000",
         17815 => x"00000000",
         17816 => x"00000000",
         17817 => x"00000000",
         17818 => x"00000000",
         17819 => x"00000000",
         17820 => x"00000000",
         17821 => x"00000000",
         17822 => x"00000000",
         17823 => x"00000000",
         17824 => x"00000000",
         17825 => x"00000000",
         17826 => x"00000000",
         17827 => x"00000000",
         17828 => x"00000000",
         17829 => x"00000000",
         17830 => x"00000000",
         17831 => x"00000000",
         17832 => x"00000000",
         17833 => x"00000000",
         17834 => x"00000000",
         17835 => x"00000000",
         17836 => x"00000000",
         17837 => x"00000000",
         17838 => x"00000000",
         17839 => x"00000000",
         17840 => x"00000000",
         17841 => x"00000000",
         17842 => x"00000000",
         17843 => x"00000000",
         17844 => x"00000000",
         17845 => x"00000000",
         17846 => x"00000000",
         17847 => x"00000000",
         17848 => x"00000000",
         17849 => x"00000000",
         17850 => x"00000000",
         17851 => x"00000000",
         17852 => x"00000000",
         17853 => x"00000000",
         17854 => x"00000000",
         17855 => x"00000000",
         17856 => x"00000000",
         17857 => x"00000000",
         17858 => x"00000000",
         17859 => x"00000000",
         17860 => x"00000000",
         17861 => x"00000000",
         17862 => x"00000000",
         17863 => x"00000000",
         17864 => x"00000000",
         17865 => x"00000000",
         17866 => x"00000000",
         17867 => x"00000000",
         17868 => x"00000000",
         17869 => x"00000000",
         17870 => x"00000000",
         17871 => x"00000000",
         17872 => x"00000000",
         17873 => x"00000000",
         17874 => x"00000000",
         17875 => x"00000000",
         17876 => x"00000000",
         17877 => x"00000000",
         17878 => x"00000000",
         17879 => x"00000000",
         17880 => x"00000000",
         17881 => x"00000000",
         17882 => x"00000000",
         17883 => x"00000000",
         17884 => x"00000000",
         17885 => x"00000000",
         17886 => x"00000000",
         17887 => x"00000000",
         17888 => x"00000000",
         17889 => x"00000000",
         17890 => x"00000000",
         17891 => x"00000000",
         17892 => x"00000000",
         17893 => x"00000000",
         17894 => x"00000000",
         17895 => x"00000000",
         17896 => x"00000000",
         17897 => x"00000000",
         17898 => x"00000000",
         17899 => x"00000000",
         17900 => x"00000000",
         17901 => x"00000000",
         17902 => x"00000000",
         17903 => x"00000000",
         17904 => x"00000000",
         17905 => x"00000000",
         17906 => x"00000000",
         17907 => x"00000000",
         17908 => x"00000000",
         17909 => x"00000000",
         17910 => x"00000000",
         17911 => x"00000000",
         17912 => x"00000000",
         17913 => x"00000000",
         17914 => x"00000000",
         17915 => x"00000000",
         17916 => x"00000000",
         17917 => x"00000000",
         17918 => x"00000000",
         17919 => x"00000000",
         17920 => x"00000000",
         17921 => x"00000000",
         17922 => x"00000000",
         17923 => x"00000000",
         17924 => x"00000000",
         17925 => x"00000000",
         17926 => x"00000000",
         17927 => x"00000000",
         17928 => x"00000000",
         17929 => x"00000000",
         17930 => x"00000000",
         17931 => x"00000000",
         17932 => x"00000000",
         17933 => x"00000000",
         17934 => x"00000000",
         17935 => x"00000000",
         17936 => x"00000000",
         17937 => x"00000000",
         17938 => x"00000000",
         17939 => x"00000000",
         17940 => x"00000000",
         17941 => x"00000000",
         17942 => x"00000000",
         17943 => x"00000000",
         17944 => x"00000000",
         17945 => x"00000000",
         17946 => x"00000000",
         17947 => x"00000000",
         17948 => x"00000000",
         17949 => x"00000000",
         17950 => x"00000000",
         17951 => x"00000000",
         17952 => x"00000000",
         17953 => x"00000000",
         17954 => x"00000000",
         17955 => x"00000000",
         17956 => x"00000000",
         17957 => x"00000000",
         17958 => x"00000000",
         17959 => x"00000000",
         17960 => x"00000000",
         17961 => x"00000000",
         17962 => x"00000000",
         17963 => x"00000000",
         17964 => x"00000000",
         17965 => x"00000000",
         17966 => x"00000000",
         17967 => x"00000000",
         17968 => x"00000000",
         17969 => x"00000000",
         17970 => x"00000000",
         17971 => x"00000000",
         17972 => x"00000000",
         17973 => x"00000000",
         17974 => x"00000000",
         17975 => x"00000000",
         17976 => x"00000000",
         17977 => x"00000000",
         17978 => x"00000000",
         17979 => x"00000000",
         17980 => x"00000000",
         17981 => x"00000000",
         17982 => x"00000000",
         17983 => x"00000000",
         17984 => x"00000000",
         17985 => x"00000000",
         17986 => x"00000000",
         17987 => x"00000000",
         17988 => x"00000000",
         17989 => x"00000000",
         17990 => x"00000000",
         17991 => x"00000000",
         17992 => x"00000000",
         17993 => x"00000000",
         17994 => x"00000000",
         17995 => x"00000000",
         17996 => x"00000000",
         17997 => x"00000000",
         17998 => x"00000000",
         17999 => x"00000000",
         18000 => x"00000000",
         18001 => x"00000000",
         18002 => x"00000000",
         18003 => x"00000000",
         18004 => x"00000000",
         18005 => x"00000000",
         18006 => x"00000000",
         18007 => x"00000000",
         18008 => x"00000000",
         18009 => x"00000000",
         18010 => x"00000000",
         18011 => x"00000000",
         18012 => x"00000000",
         18013 => x"00000000",
         18014 => x"00000000",
         18015 => x"00000000",
         18016 => x"00000000",
         18017 => x"00000000",
         18018 => x"00000000",
         18019 => x"00000000",
         18020 => x"00000000",
         18021 => x"00000000",
         18022 => x"00000000",
         18023 => x"00000000",
         18024 => x"00000000",
         18025 => x"00000000",
         18026 => x"00000000",
         18027 => x"00000000",
         18028 => x"00000000",
         18029 => x"00000000",
         18030 => x"00000000",
         18031 => x"00000000",
         18032 => x"00000000",
         18033 => x"00000000",
         18034 => x"00000000",
         18035 => x"00000000",
         18036 => x"00000000",
         18037 => x"00000000",
         18038 => x"00000000",
         18039 => x"00000000",
         18040 => x"00000000",
         18041 => x"00000000",
         18042 => x"00000000",
         18043 => x"00000000",
         18044 => x"00000000",
         18045 => x"00000000",
         18046 => x"00000000",
         18047 => x"00000000",
         18048 => x"00000000",
         18049 => x"00000000",
         18050 => x"00000000",
         18051 => x"00000000",
         18052 => x"00000000",
         18053 => x"00000000",
         18054 => x"00000000",
         18055 => x"00000000",
         18056 => x"00000000",
         18057 => x"00000000",
         18058 => x"00000000",
         18059 => x"00000000",
         18060 => x"00000000",
         18061 => x"00000000",
         18062 => x"00000000",
         18063 => x"00000000",
         18064 => x"00000000",
         18065 => x"00000000",
         18066 => x"00000000",
         18067 => x"00000000",
         18068 => x"00000000",
         18069 => x"00000000",
         18070 => x"00000000",
         18071 => x"00000000",
         18072 => x"00000000",
         18073 => x"00000000",
         18074 => x"00000000",
         18075 => x"00000000",
         18076 => x"00000000",
         18077 => x"00000000",
         18078 => x"00000000",
         18079 => x"00000000",
         18080 => x"00000000",
         18081 => x"00000000",
         18082 => x"00000000",
         18083 => x"00000000",
         18084 => x"00000000",
         18085 => x"00000000",
         18086 => x"00000000",
         18087 => x"00000000",
         18088 => x"00000000",
         18089 => x"00000000",
         18090 => x"00000000",
         18091 => x"00000000",
         18092 => x"00000000",
         18093 => x"00000000",
         18094 => x"00000000",
         18095 => x"00000000",
         18096 => x"00000000",
         18097 => x"00000000",
         18098 => x"00000000",
         18099 => x"00000000",
         18100 => x"00000000",
         18101 => x"00000000",
         18102 => x"00000000",
         18103 => x"00000000",
         18104 => x"00000000",
         18105 => x"00000000",
         18106 => x"00000000",
         18107 => x"00000000",
         18108 => x"00000000",
         18109 => x"00000000",
         18110 => x"00000000",
         18111 => x"00000000",
         18112 => x"00000000",
         18113 => x"00000000",
         18114 => x"00000000",
         18115 => x"00000000",
         18116 => x"00000000",
         18117 => x"00000000",
         18118 => x"00000000",
         18119 => x"00000000",
         18120 => x"00000000",
         18121 => x"00000000",
         18122 => x"00000000",
         18123 => x"00000000",
         18124 => x"00000000",
         18125 => x"00000000",
         18126 => x"00000000",
         18127 => x"00000000",
         18128 => x"00000000",
         18129 => x"00000000",
         18130 => x"00000000",
         18131 => x"00000000",
         18132 => x"00000000",
         18133 => x"00000000",
         18134 => x"00000000",
         18135 => x"00000000",
         18136 => x"00000000",
         18137 => x"00000000",
         18138 => x"00000000",
         18139 => x"00000000",
         18140 => x"00000000",
         18141 => x"00000000",
         18142 => x"00000000",
         18143 => x"00000000",
         18144 => x"00000000",
         18145 => x"00000000",
         18146 => x"00000000",
         18147 => x"00000000",
         18148 => x"00000000",
         18149 => x"00000000",
         18150 => x"00000000",
         18151 => x"00000000",
         18152 => x"00000000",
         18153 => x"00000000",
         18154 => x"00000000",
         18155 => x"00000000",
         18156 => x"00000000",
         18157 => x"00000000",
         18158 => x"00003219",
         18159 => x"50000100",
         18160 => x"00000000",
         18161 => x"cce0f2f3",
         18162 => x"cecff6f7",
         18163 => x"f8f9fafb",
         18164 => x"fcfdfeff",
         18165 => x"e1c1c2c3",
         18166 => x"c4c5c6e2",
         18167 => x"e3e4e5e6",
         18168 => x"ebeeeff4",
         18169 => x"00616263",
         18170 => x"64656667",
         18171 => x"68696b6a",
         18172 => x"2f2a2e2d",
         18173 => x"20212223",
         18174 => x"24252627",
         18175 => x"28294f2c",
         18176 => x"512b5749",
         18177 => x"55010203",
         18178 => x"04050607",
         18179 => x"08090a0b",
         18180 => x"0c0d0e0f",
         18181 => x"10111213",
         18182 => x"14151617",
         18183 => x"18191a52",
         18184 => x"5954be3c",
         18185 => x"c7818283",
         18186 => x"84858687",
         18187 => x"88898a8b",
         18188 => x"8c8d8e8f",
         18189 => x"90919293",
         18190 => x"94959697",
         18191 => x"98999abc",
         18192 => x"8040a5c0",
         18193 => x"00000000",
         18194 => x"00000000",
         18195 => x"00000000",
         18196 => x"00000000",
         18197 => x"00000000",
         18198 => x"00000000",
         18199 => x"00000000",
         18200 => x"00000000",
         18201 => x"00000000",
         18202 => x"00000000",
         18203 => x"00000000",
         18204 => x"00000000",
         18205 => x"00000000",
         18206 => x"00000000",
         18207 => x"00000000",
         18208 => x"00000000",
         18209 => x"00000000",
         18210 => x"00000000",
         18211 => x"00000000",
         18212 => x"00000000",
         18213 => x"00000000",
         18214 => x"00000000",
         18215 => x"00000000",
         18216 => x"00000000",
         18217 => x"00000000",
         18218 => x"00000000",
         18219 => x"00000000",
         18220 => x"00000000",
         18221 => x"00000000",
         18222 => x"00000000",
         18223 => x"00020003",
         18224 => x"00040101",
         18225 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

