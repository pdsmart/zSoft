-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b83ff",
             1 => x"f80d0b0b",
             2 => x"0b93b904",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"9d040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b9380",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b829a",
           162 => x"8c738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93850400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b80c3",
           171 => x"f42d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b80c5",
           179 => x"e02d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"95040b0b",
           269 => x"0b8ca404",
           270 => x"0b0b0b8c",
           271 => x"b3040b0b",
           272 => x"0b8cc204",
           273 => x"0b0b0b8c",
           274 => x"d1040b0b",
           275 => x"0b8ce004",
           276 => x"0b0b0b8c",
           277 => x"f0040b0b",
           278 => x"0b8d8004",
           279 => x"0b0b0b8d",
           280 => x"8f040b0b",
           281 => x"0b8d9e04",
           282 => x"0b0b0b8d",
           283 => x"ad040b0b",
           284 => x"0b8dbd04",
           285 => x"0b0b0b8d",
           286 => x"cd040b0b",
           287 => x"0b8ddd04",
           288 => x"0b0b0b8d",
           289 => x"ed040b0b",
           290 => x"0b8dfd04",
           291 => x"0b0b0b8e",
           292 => x"8d040b0b",
           293 => x"0b8e9d04",
           294 => x"0b0b0b8e",
           295 => x"ad040b0b",
           296 => x"0b8ebd04",
           297 => x"0b0b0b8e",
           298 => x"cd040b0b",
           299 => x"0b8edd04",
           300 => x"0b0b0b8e",
           301 => x"ed040b0b",
           302 => x"0b8efd04",
           303 => x"0b0b0b8f",
           304 => x"8d040b0b",
           305 => x"0b8f9d04",
           306 => x"0b0b0b8f",
           307 => x"ad040b0b",
           308 => x"0b8fbd04",
           309 => x"0b0b0b8f",
           310 => x"cd040b0b",
           311 => x"0b8fdd04",
           312 => x"0b0b0b8f",
           313 => x"ed040b0b",
           314 => x"0b8ffd04",
           315 => x"0b0b0b90",
           316 => x"8d040b0b",
           317 => x"0b909d04",
           318 => x"0b0b0b90",
           319 => x"ad040b0b",
           320 => x"0b90bd04",
           321 => x"0b0b0b90",
           322 => x"cd040b0b",
           323 => x"0b90dd04",
           324 => x"0b0b0b90",
           325 => x"ed040b0b",
           326 => x"0b90fd04",
           327 => x"0b0b0b91",
           328 => x"8d040b0b",
           329 => x"0b919d04",
           330 => x"0b0b0b91",
           331 => x"ad040b0b",
           332 => x"0b91bd04",
           333 => x"0b0b0b91",
           334 => x"cd040b0b",
           335 => x"0b91dd04",
           336 => x"0b0b0b91",
           337 => x"ed040b0b",
           338 => x"0b91fd04",
           339 => x"0b0b0b92",
           340 => x"8d040b0b",
           341 => x"0b929d04",
           342 => x"0b0b0b92",
           343 => x"ad040b0b",
           344 => x"0b92bd04",
           345 => x"0b0b0b92",
           346 => x"cd04ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0482bbe8",
           386 => x"0c80f98d",
           387 => x"2d82bbe8",
           388 => x"0882d890",
           389 => x"0482bbe8",
           390 => x"0cb3b22d",
           391 => x"82bbe808",
           392 => x"82d89004",
           393 => x"82bbe80c",
           394 => x"afe32d82",
           395 => x"bbe80882",
           396 => x"d8900482",
           397 => x"bbe80caf",
           398 => x"ad2d82bb",
           399 => x"e80882d8",
           400 => x"900482bb",
           401 => x"e80c94ad",
           402 => x"2d82bbe8",
           403 => x"0882d890",
           404 => x"0482bbe8",
           405 => x"0cb1c22d",
           406 => x"82bbe808",
           407 => x"82d89004",
           408 => x"82bbe80c",
           409 => x"80cfcc2d",
           410 => x"82bbe808",
           411 => x"82d89004",
           412 => x"82bbe80c",
           413 => x"80c9fb2d",
           414 => x"82bbe808",
           415 => x"82d89004",
           416 => x"82bbe80c",
           417 => x"93d82d82",
           418 => x"bbe80882",
           419 => x"d8900482",
           420 => x"bbe80c96",
           421 => x"c02d82bb",
           422 => x"e80882d8",
           423 => x"900482bb",
           424 => x"e80c97cd",
           425 => x"2d82bbe8",
           426 => x"0882d890",
           427 => x"0482bbe8",
           428 => x"0c80fcb7",
           429 => x"2d82bbe8",
           430 => x"0882d890",
           431 => x"0482bbe8",
           432 => x"0c80fd95",
           433 => x"2d82bbe8",
           434 => x"0882d890",
           435 => x"0482bbe8",
           436 => x"0c80f4d2",
           437 => x"2d82bbe8",
           438 => x"0882d890",
           439 => x"0482bbe8",
           440 => x"0c80f6c9",
           441 => x"2d82bbe8",
           442 => x"0882d890",
           443 => x"0482bbe8",
           444 => x"0c80f7fc",
           445 => x"2d82bbe8",
           446 => x"0882d890",
           447 => x"0482bbe8",
           448 => x"0c81dcf0",
           449 => x"2d82bbe8",
           450 => x"0882d890",
           451 => x"0482bbe8",
           452 => x"0c81e9e1",
           453 => x"2d82bbe8",
           454 => x"0882d890",
           455 => x"0482bbe8",
           456 => x"0c81e1d5",
           457 => x"2d82bbe8",
           458 => x"0882d890",
           459 => x"0482bbe8",
           460 => x"0c81e4d2",
           461 => x"2d82bbe8",
           462 => x"0882d890",
           463 => x"0482bbe8",
           464 => x"0c81eef0",
           465 => x"2d82bbe8",
           466 => x"0882d890",
           467 => x"0482bbe8",
           468 => x"0c81f7d0",
           469 => x"2d82bbe8",
           470 => x"0882d890",
           471 => x"0482bbe8",
           472 => x"0c81e8c3",
           473 => x"2d82bbe8",
           474 => x"0882d890",
           475 => x"0482bbe8",
           476 => x"0c81f28f",
           477 => x"2d82bbe8",
           478 => x"0882d890",
           479 => x"0482bbe8",
           480 => x"0c81f3ae",
           481 => x"2d82bbe8",
           482 => x"0882d890",
           483 => x"0482bbe8",
           484 => x"0c81f3cd",
           485 => x"2d82bbe8",
           486 => x"0882d890",
           487 => x"0482bbe8",
           488 => x"0c81fbb7",
           489 => x"2d82bbe8",
           490 => x"0882d890",
           491 => x"0482bbe8",
           492 => x"0c81f99d",
           493 => x"2d82bbe8",
           494 => x"0882d890",
           495 => x"0482bbe8",
           496 => x"0c81fe8b",
           497 => x"2d82bbe8",
           498 => x"0882d890",
           499 => x"0482bbe8",
           500 => x"0c81f4d1",
           501 => x"2d82bbe8",
           502 => x"0882d890",
           503 => x"0482bbe8",
           504 => x"0c82818b",
           505 => x"2d82bbe8",
           506 => x"0882d890",
           507 => x"0482bbe8",
           508 => x"0c82828c",
           509 => x"2d82bbe8",
           510 => x"0882d890",
           511 => x"0482bbe8",
           512 => x"0c81eac1",
           513 => x"2d82bbe8",
           514 => x"0882d890",
           515 => x"0482bbe8",
           516 => x"0c81ea9a",
           517 => x"2d82bbe8",
           518 => x"0882d890",
           519 => x"0482bbe8",
           520 => x"0c81ebc5",
           521 => x"2d82bbe8",
           522 => x"0882d890",
           523 => x"0482bbe8",
           524 => x"0c81f5a8",
           525 => x"2d82bbe8",
           526 => x"0882d890",
           527 => x"0482bbe8",
           528 => x"0c8282fd",
           529 => x"2d82bbe8",
           530 => x"0882d890",
           531 => x"0482bbe8",
           532 => x"0c828587",
           533 => x"2d82bbe8",
           534 => x"0882d890",
           535 => x"0482bbe8",
           536 => x"0c8288c9",
           537 => x"2d82bbe8",
           538 => x"0882d890",
           539 => x"0482bbe8",
           540 => x"0c81dc8f",
           541 => x"2d82bbe8",
           542 => x"0882d890",
           543 => x"0482bbe8",
           544 => x"0c828bb5",
           545 => x"2d82bbe8",
           546 => x"0882d890",
           547 => x"0482bbe8",
           548 => x"0c8299ea",
           549 => x"2d82bbe8",
           550 => x"0882d890",
           551 => x"0482bbe8",
           552 => x"0c8297d6",
           553 => x"2d82bbe8",
           554 => x"0882d890",
           555 => x"0482bbe8",
           556 => x"0c81adca",
           557 => x"2d82bbe8",
           558 => x"0882d890",
           559 => x"0482bbe8",
           560 => x"0c81afb4",
           561 => x"2d82bbe8",
           562 => x"0882d890",
           563 => x"0482bbe8",
           564 => x"0c81b198",
           565 => x"2d82bbe8",
           566 => x"0882d890",
           567 => x"0482bbe8",
           568 => x"0c80f4fb",
           569 => x"2d82bbe8",
           570 => x"0882d890",
           571 => x"0482bbe8",
           572 => x"0c80f69f",
           573 => x"2d82bbe8",
           574 => x"0882d890",
           575 => x"0482bbe8",
           576 => x"0c80fa82",
           577 => x"2d82bbe8",
           578 => x"0882d890",
           579 => x"0482bbe8",
           580 => x"0c80d698",
           581 => x"2d82bbe8",
           582 => x"0882d890",
           583 => x"0482bbe8",
           584 => x"0c81a7de",
           585 => x"2d82bbe8",
           586 => x"0882d890",
           587 => x"0482bbe8",
           588 => x"0c81a886",
           589 => x"2d82bbe8",
           590 => x"0882d890",
           591 => x"0482bbe8",
           592 => x"0c81abfe",
           593 => x"2d82bbe8",
           594 => x"0882d890",
           595 => x"0482bbe8",
           596 => x"0c81a4c8",
           597 => x"2d82bbe8",
           598 => x"0882d890",
           599 => x"043c0400",
           600 => x"00101010",
           601 => x"10101010",
           602 => x"10101010",
           603 => x"10101010",
           604 => x"10101010",
           605 => x"10101010",
           606 => x"10101010",
           607 => x"10101010",
           608 => x"53510400",
           609 => x"007381ff",
           610 => x"06738306",
           611 => x"09810583",
           612 => x"05101010",
           613 => x"2b0772fc",
           614 => x"060c5151",
           615 => x"04727280",
           616 => x"728106ff",
           617 => x"05097206",
           618 => x"05711052",
           619 => x"720a100a",
           620 => x"5372ed38",
           621 => x"51515351",
           622 => x"0482bbdc",
           623 => x"7082d3b8",
           624 => x"278e3880",
           625 => x"71708405",
           626 => x"530c0b0b",
           627 => x"0b93bc04",
           628 => x"8c815180",
           629 => x"f3950400",
           630 => x"82bbe808",
           631 => x"0282bbe8",
           632 => x"0cfb3d0d",
           633 => x"82bbe808",
           634 => x"8c057082",
           635 => x"bbe808fc",
           636 => x"050c82bb",
           637 => x"e808fc05",
           638 => x"085482bb",
           639 => x"e8088805",
           640 => x"085382d3",
           641 => x"b0085254",
           642 => x"849a3f82",
           643 => x"bbdc0870",
           644 => x"82bbe808",
           645 => x"f8050c82",
           646 => x"bbe808f8",
           647 => x"05087082",
           648 => x"bbdc0c51",
           649 => x"54873d0d",
           650 => x"82bbe80c",
           651 => x"0482bbe8",
           652 => x"080282bb",
           653 => x"e80cfb3d",
           654 => x"0d82bbe8",
           655 => x"08900508",
           656 => x"85113370",
           657 => x"81327081",
           658 => x"06515151",
           659 => x"52718f38",
           660 => x"800b82bb",
           661 => x"e8088c05",
           662 => x"08258338",
           663 => x"8d39800b",
           664 => x"82bbe808",
           665 => x"f4050c81",
           666 => x"c43982bb",
           667 => x"e8088c05",
           668 => x"08ff0582",
           669 => x"bbe8088c",
           670 => x"050c800b",
           671 => x"82bbe808",
           672 => x"f8050c82",
           673 => x"bbe80888",
           674 => x"050882bb",
           675 => x"e808fc05",
           676 => x"0c82bbe8",
           677 => x"08f80508",
           678 => x"8a2e80f6",
           679 => x"38800b82",
           680 => x"bbe8088c",
           681 => x"05082580",
           682 => x"e93882bb",
           683 => x"e8089005",
           684 => x"0851a090",
           685 => x"3f82bbdc",
           686 => x"087082bb",
           687 => x"e808f805",
           688 => x"0c5282bb",
           689 => x"e808f805",
           690 => x"08ff2e09",
           691 => x"81068d38",
           692 => x"800b82bb",
           693 => x"e808f405",
           694 => x"0c80d239",
           695 => x"82bbe808",
           696 => x"fc050882",
           697 => x"bbe808f8",
           698 => x"05085353",
           699 => x"71733482",
           700 => x"bbe8088c",
           701 => x"0508ff05",
           702 => x"82bbe808",
           703 => x"8c050c82",
           704 => x"bbe808fc",
           705 => x"05088105",
           706 => x"82bbe808",
           707 => x"fc050cff",
           708 => x"803982bb",
           709 => x"e808fc05",
           710 => x"08528072",
           711 => x"3482bbe8",
           712 => x"08880508",
           713 => x"7082bbe8",
           714 => x"08f4050c",
           715 => x"5282bbe8",
           716 => x"08f40508",
           717 => x"82bbdc0c",
           718 => x"873d0d82",
           719 => x"bbe80c04",
           720 => x"82bbe808",
           721 => x"0282bbe8",
           722 => x"0cf43d0d",
           723 => x"860b82bb",
           724 => x"e808e505",
           725 => x"3482bbe8",
           726 => x"08880508",
           727 => x"82bbe808",
           728 => x"e0050cfe",
           729 => x"0a0b82bb",
           730 => x"e808e805",
           731 => x"0c82bbe8",
           732 => x"08900570",
           733 => x"82bbe808",
           734 => x"fc050c82",
           735 => x"bbe808fc",
           736 => x"05085482",
           737 => x"bbe8088c",
           738 => x"05085382",
           739 => x"bbe808e0",
           740 => x"05705351",
           741 => x"54818d3f",
           742 => x"82bbdc08",
           743 => x"7082bbe8",
           744 => x"08dc050c",
           745 => x"82bbe808",
           746 => x"ec050882",
           747 => x"bbe80888",
           748 => x"05080551",
           749 => x"54807434",
           750 => x"82bbe808",
           751 => x"dc050870",
           752 => x"82bbdc0c",
           753 => x"548e3d0d",
           754 => x"82bbe80c",
           755 => x"0482bbe8",
           756 => x"080282bb",
           757 => x"e80cfb3d",
           758 => x"0d82bbe8",
           759 => x"08900570",
           760 => x"82bbe808",
           761 => x"fc050c82",
           762 => x"bbe808fc",
           763 => x"05085482",
           764 => x"bbe8088c",
           765 => x"05085382",
           766 => x"bbe80888",
           767 => x"05085254",
           768 => x"a33f82bb",
           769 => x"dc087082",
           770 => x"bbe808f8",
           771 => x"050c82bb",
           772 => x"e808f805",
           773 => x"087082bb",
           774 => x"dc0c5154",
           775 => x"873d0d82",
           776 => x"bbe80c04",
           777 => x"82bbe808",
           778 => x"0282bbe8",
           779 => x"0ced3d0d",
           780 => x"800b82bb",
           781 => x"e808e405",
           782 => x"2382bbe8",
           783 => x"08880508",
           784 => x"53800b8c",
           785 => x"140c82bb",
           786 => x"e8088805",
           787 => x"08851133",
           788 => x"70812a70",
           789 => x"81327081",
           790 => x"06515151",
           791 => x"51537280",
           792 => x"2e8d38ff",
           793 => x"0b82bbe8",
           794 => x"08e0050c",
           795 => x"96ac3982",
           796 => x"bbe8088c",
           797 => x"05085372",
           798 => x"33537282",
           799 => x"bbe808f8",
           800 => x"05347281",
           801 => x"ff065372",
           802 => x"802e95fa",
           803 => x"3882bbe8",
           804 => x"088c0508",
           805 => x"810582bb",
           806 => x"e8088c05",
           807 => x"0c82bbe8",
           808 => x"08e40522",
           809 => x"70810651",
           810 => x"5372802e",
           811 => x"958b3882",
           812 => x"bbe808f8",
           813 => x"053353af",
           814 => x"732781fc",
           815 => x"3882bbe8",
           816 => x"08f80533",
           817 => x"5372b926",
           818 => x"81ee3882",
           819 => x"bbe808f8",
           820 => x"05335372",
           821 => x"b02e0981",
           822 => x"0680c538",
           823 => x"82bbe808",
           824 => x"e8053370",
           825 => x"982b7098",
           826 => x"2c515153",
           827 => x"72b23882",
           828 => x"bbe808e4",
           829 => x"05227083",
           830 => x"2a708132",
           831 => x"70810651",
           832 => x"51515372",
           833 => x"802e9938",
           834 => x"82bbe808",
           835 => x"e4052270",
           836 => x"82800751",
           837 => x"537282bb",
           838 => x"e808e405",
           839 => x"23fed039",
           840 => x"82bbe808",
           841 => x"e8053370",
           842 => x"982b7098",
           843 => x"2c707083",
           844 => x"2b721173",
           845 => x"11515151",
           846 => x"53515553",
           847 => x"7282bbe8",
           848 => x"08e80534",
           849 => x"82bbe808",
           850 => x"e8053354",
           851 => x"82bbe808",
           852 => x"f8053370",
           853 => x"15d01151",
           854 => x"51537282",
           855 => x"bbe808e8",
           856 => x"053482bb",
           857 => x"e808e805",
           858 => x"3370982b",
           859 => x"70982c51",
           860 => x"51537280",
           861 => x"258b3880",
           862 => x"ff0b82bb",
           863 => x"e808e805",
           864 => x"3482bbe8",
           865 => x"08e40522",
           866 => x"70832a70",
           867 => x"81065151",
           868 => x"5372fddb",
           869 => x"3882bbe8",
           870 => x"08e80533",
           871 => x"70882b70",
           872 => x"902b7090",
           873 => x"2c70882c",
           874 => x"51515151",
           875 => x"537282bb",
           876 => x"e808ec05",
           877 => x"23fdb839",
           878 => x"82bbe808",
           879 => x"e4052270",
           880 => x"832a7081",
           881 => x"06515153",
           882 => x"72802e9d",
           883 => x"3882bbe8",
           884 => x"08e80533",
           885 => x"70982b70",
           886 => x"982c5151",
           887 => x"53728a38",
           888 => x"810b82bb",
           889 => x"e808e805",
           890 => x"3482bbe8",
           891 => x"08f80533",
           892 => x"e01182bb",
           893 => x"e808c405",
           894 => x"0c5382bb",
           895 => x"e808c405",
           896 => x"0880d826",
           897 => x"92943882",
           898 => x"bbe808c4",
           899 => x"05087082",
           900 => x"2b829bd8",
           901 => x"11700851",
           902 => x"51515372",
           903 => x"0482bbe8",
           904 => x"08e40522",
           905 => x"70900751",
           906 => x"537282bb",
           907 => x"e808e405",
           908 => x"2382bbe8",
           909 => x"08e40522",
           910 => x"70a00751",
           911 => x"537282bb",
           912 => x"e808e405",
           913 => x"23fca839",
           914 => x"82bbe808",
           915 => x"e4052270",
           916 => x"81800751",
           917 => x"537282bb",
           918 => x"e808e405",
           919 => x"23fc9039",
           920 => x"82bbe808",
           921 => x"e4052270",
           922 => x"80c00751",
           923 => x"537282bb",
           924 => x"e808e405",
           925 => x"23fbf839",
           926 => x"82bbe808",
           927 => x"e4052270",
           928 => x"88075153",
           929 => x"7282bbe8",
           930 => x"08e40523",
           931 => x"800b82bb",
           932 => x"e808e805",
           933 => x"34fbd839",
           934 => x"82bbe808",
           935 => x"e4052270",
           936 => x"84075153",
           937 => x"7282bbe8",
           938 => x"08e40523",
           939 => x"fbc139bf",
           940 => x"0b82bbe8",
           941 => x"08fc0534",
           942 => x"82bbe808",
           943 => x"ec0522ff",
           944 => x"11515372",
           945 => x"82bbe808",
           946 => x"ec052380",
           947 => x"e30b82bb",
           948 => x"e808f805",
           949 => x"348da839",
           950 => x"82bbe808",
           951 => x"90050882",
           952 => x"bbe80890",
           953 => x"05088405",
           954 => x"82bbe808",
           955 => x"90050c70",
           956 => x"08515372",
           957 => x"82bbe808",
           958 => x"fc053482",
           959 => x"bbe808ec",
           960 => x"0522ff11",
           961 => x"51537282",
           962 => x"bbe808ec",
           963 => x"05238cef",
           964 => x"3982bbe8",
           965 => x"08900508",
           966 => x"82bbe808",
           967 => x"90050884",
           968 => x"0582bbe8",
           969 => x"0890050c",
           970 => x"700882bb",
           971 => x"e808fc05",
           972 => x"0c82bbe8",
           973 => x"08e40522",
           974 => x"70832a70",
           975 => x"81065151",
           976 => x"51537280",
           977 => x"2eab3882",
           978 => x"bbe808e8",
           979 => x"05337098",
           980 => x"2b537298",
           981 => x"2c5382bb",
           982 => x"e808fc05",
           983 => x"085253a2",
           984 => x"d83f82bb",
           985 => x"dc085372",
           986 => x"82bbe808",
           987 => x"f4052399",
           988 => x"3982bbe8",
           989 => x"08fc0508",
           990 => x"519d8a3f",
           991 => x"82bbdc08",
           992 => x"537282bb",
           993 => x"e808f405",
           994 => x"2382bbe8",
           995 => x"08ec0522",
           996 => x"5382bbe8",
           997 => x"08f40522",
           998 => x"73713154",
           999 => x"547282bb",
          1000 => x"e808ec05",
          1001 => x"238bd839",
          1002 => x"82bbe808",
          1003 => x"90050882",
          1004 => x"bbe80890",
          1005 => x"05088405",
          1006 => x"82bbe808",
          1007 => x"90050c70",
          1008 => x"0882bbe8",
          1009 => x"08fc050c",
          1010 => x"82bbe808",
          1011 => x"e4052270",
          1012 => x"832a7081",
          1013 => x"06515151",
          1014 => x"5372802e",
          1015 => x"ab3882bb",
          1016 => x"e808e805",
          1017 => x"3370982b",
          1018 => x"5372982c",
          1019 => x"5382bbe8",
          1020 => x"08fc0508",
          1021 => x"5253a1c1",
          1022 => x"3f82bbdc",
          1023 => x"08537282",
          1024 => x"bbe808f4",
          1025 => x"05239939",
          1026 => x"82bbe808",
          1027 => x"fc050851",
          1028 => x"9bf33f82",
          1029 => x"bbdc0853",
          1030 => x"7282bbe8",
          1031 => x"08f40523",
          1032 => x"82bbe808",
          1033 => x"ec052253",
          1034 => x"82bbe808",
          1035 => x"f4052273",
          1036 => x"71315454",
          1037 => x"7282bbe8",
          1038 => x"08ec0523",
          1039 => x"8ac13982",
          1040 => x"bbe808e4",
          1041 => x"05227082",
          1042 => x"2a708106",
          1043 => x"51515372",
          1044 => x"802ea438",
          1045 => x"82bbe808",
          1046 => x"90050882",
          1047 => x"bbe80890",
          1048 => x"05088405",
          1049 => x"82bbe808",
          1050 => x"90050c70",
          1051 => x"0882bbe8",
          1052 => x"08dc050c",
          1053 => x"53a23982",
          1054 => x"bbe80890",
          1055 => x"050882bb",
          1056 => x"e8089005",
          1057 => x"08840582",
          1058 => x"bbe80890",
          1059 => x"050c7008",
          1060 => x"82bbe808",
          1061 => x"dc050c53",
          1062 => x"82bbe808",
          1063 => x"dc050882",
          1064 => x"bbe808fc",
          1065 => x"050c82bb",
          1066 => x"e808fc05",
          1067 => x"088025a4",
          1068 => x"3882bbe8",
          1069 => x"08e40522",
          1070 => x"70820751",
          1071 => x"537282bb",
          1072 => x"e808e405",
          1073 => x"2382bbe8",
          1074 => x"08fc0508",
          1075 => x"3082bbe8",
          1076 => x"08fc050c",
          1077 => x"82bbe808",
          1078 => x"e4052270",
          1079 => x"ffbf0651",
          1080 => x"537282bb",
          1081 => x"e808e405",
          1082 => x"2381af39",
          1083 => x"880b82bb",
          1084 => x"e808f405",
          1085 => x"23a93982",
          1086 => x"bbe808e4",
          1087 => x"05227080",
          1088 => x"c0075153",
          1089 => x"7282bbe8",
          1090 => x"08e40523",
          1091 => x"80f80b82",
          1092 => x"bbe808f8",
          1093 => x"0534900b",
          1094 => x"82bbe808",
          1095 => x"f4052382",
          1096 => x"bbe808e4",
          1097 => x"05227082",
          1098 => x"2a708106",
          1099 => x"51515372",
          1100 => x"802ea438",
          1101 => x"82bbe808",
          1102 => x"90050882",
          1103 => x"bbe80890",
          1104 => x"05088405",
          1105 => x"82bbe808",
          1106 => x"90050c70",
          1107 => x"0882bbe8",
          1108 => x"08d8050c",
          1109 => x"53a23982",
          1110 => x"bbe80890",
          1111 => x"050882bb",
          1112 => x"e8089005",
          1113 => x"08840582",
          1114 => x"bbe80890",
          1115 => x"050c7008",
          1116 => x"82bbe808",
          1117 => x"d8050c53",
          1118 => x"82bbe808",
          1119 => x"d8050882",
          1120 => x"bbe808fc",
          1121 => x"050c82bb",
          1122 => x"e808e405",
          1123 => x"2270cf06",
          1124 => x"51537282",
          1125 => x"bbe808e4",
          1126 => x"052382bb",
          1127 => x"ec0b82bb",
          1128 => x"e808f005",
          1129 => x"0c82bbe8",
          1130 => x"08f00508",
          1131 => x"82bbe808",
          1132 => x"f4052282",
          1133 => x"bbe808fc",
          1134 => x"05087155",
          1135 => x"70545654",
          1136 => x"55a3f33f",
          1137 => x"82bbdc08",
          1138 => x"53727534",
          1139 => x"82bbe808",
          1140 => x"f0050882",
          1141 => x"bbe808d4",
          1142 => x"050c82bb",
          1143 => x"e808f005",
          1144 => x"08703351",
          1145 => x"53897327",
          1146 => x"a43882bb",
          1147 => x"e808f005",
          1148 => x"08537233",
          1149 => x"5482bbe8",
          1150 => x"08f80533",
          1151 => x"7015df11",
          1152 => x"51515372",
          1153 => x"82bbe808",
          1154 => x"d0053497",
          1155 => x"3982bbe8",
          1156 => x"08f00508",
          1157 => x"537233b0",
          1158 => x"11515372",
          1159 => x"82bbe808",
          1160 => x"d0053482",
          1161 => x"bbe808d4",
          1162 => x"05085382",
          1163 => x"bbe808d0",
          1164 => x"05337334",
          1165 => x"82bbe808",
          1166 => x"f0050881",
          1167 => x"0582bbe8",
          1168 => x"08f0050c",
          1169 => x"82bbe808",
          1170 => x"f4052270",
          1171 => x"5382bbe8",
          1172 => x"08fc0508",
          1173 => x"5253a2ab",
          1174 => x"3f82bbdc",
          1175 => x"087082bb",
          1176 => x"e808fc05",
          1177 => x"0c5382bb",
          1178 => x"e808fc05",
          1179 => x"08802e84",
          1180 => x"38feb239",
          1181 => x"82bbe808",
          1182 => x"f0050882",
          1183 => x"bbec5455",
          1184 => x"72547470",
          1185 => x"75315153",
          1186 => x"7282bbe8",
          1187 => x"08fc0534",
          1188 => x"82bbe808",
          1189 => x"e4052270",
          1190 => x"b2065153",
          1191 => x"72802e94",
          1192 => x"3882bbe8",
          1193 => x"08ec0522",
          1194 => x"ff115153",
          1195 => x"7282bbe8",
          1196 => x"08ec0523",
          1197 => x"82bbe808",
          1198 => x"e4052270",
          1199 => x"862a7081",
          1200 => x"06515153",
          1201 => x"72802e80",
          1202 => x"e73882bb",
          1203 => x"e808ec05",
          1204 => x"2270902b",
          1205 => x"82bbe808",
          1206 => x"cc050c82",
          1207 => x"bbe808cc",
          1208 => x"0508902c",
          1209 => x"82bbe808",
          1210 => x"cc050c82",
          1211 => x"bbe808f4",
          1212 => x"05225153",
          1213 => x"72902e09",
          1214 => x"81069538",
          1215 => x"82bbe808",
          1216 => x"cc0508fe",
          1217 => x"05537282",
          1218 => x"bbe808c8",
          1219 => x"05239339",
          1220 => x"82bbe808",
          1221 => x"cc0508ff",
          1222 => x"05537282",
          1223 => x"bbe808c8",
          1224 => x"052382bb",
          1225 => x"e808c805",
          1226 => x"2282bbe8",
          1227 => x"08ec0523",
          1228 => x"82bbe808",
          1229 => x"e4052270",
          1230 => x"832a7081",
          1231 => x"06515153",
          1232 => x"72802e80",
          1233 => x"d03882bb",
          1234 => x"e808e805",
          1235 => x"3370982b",
          1236 => x"70982c82",
          1237 => x"bbe808fc",
          1238 => x"05335751",
          1239 => x"51537274",
          1240 => x"24973882",
          1241 => x"bbe808e4",
          1242 => x"052270f7",
          1243 => x"06515372",
          1244 => x"82bbe808",
          1245 => x"e405239d",
          1246 => x"3982bbe8",
          1247 => x"08e80533",
          1248 => x"5382bbe8",
          1249 => x"08fc0533",
          1250 => x"73713154",
          1251 => x"547282bb",
          1252 => x"e808e805",
          1253 => x"3482bbe8",
          1254 => x"08e40522",
          1255 => x"70832a70",
          1256 => x"81065151",
          1257 => x"5372802e",
          1258 => x"b13882bb",
          1259 => x"e808e805",
          1260 => x"3370882b",
          1261 => x"70902b70",
          1262 => x"902c7088",
          1263 => x"2c515151",
          1264 => x"51537254",
          1265 => x"82bbe808",
          1266 => x"ec052270",
          1267 => x"75315153",
          1268 => x"7282bbe8",
          1269 => x"08ec0523",
          1270 => x"af3982bb",
          1271 => x"e808fc05",
          1272 => x"3370882b",
          1273 => x"70902b70",
          1274 => x"902c7088",
          1275 => x"2c515151",
          1276 => x"51537254",
          1277 => x"82bbe808",
          1278 => x"ec052270",
          1279 => x"75315153",
          1280 => x"7282bbe8",
          1281 => x"08ec0523",
          1282 => x"82bbe808",
          1283 => x"e4052270",
          1284 => x"83800651",
          1285 => x"5372b038",
          1286 => x"82bbe808",
          1287 => x"ec0522ff",
          1288 => x"11545472",
          1289 => x"82bbe808",
          1290 => x"ec052373",
          1291 => x"902b7090",
          1292 => x"2c515380",
          1293 => x"73259038",
          1294 => x"82bbe808",
          1295 => x"88050852",
          1296 => x"a0518aee",
          1297 => x"3fd23982",
          1298 => x"bbe808e4",
          1299 => x"05227081",
          1300 => x"2a708106",
          1301 => x"51515372",
          1302 => x"802e9138",
          1303 => x"82bbe808",
          1304 => x"88050852",
          1305 => x"ad518aca",
          1306 => x"3f80c739",
          1307 => x"82bbe808",
          1308 => x"e4052270",
          1309 => x"842a7081",
          1310 => x"06515153",
          1311 => x"72802e90",
          1312 => x"3882bbe8",
          1313 => x"08880508",
          1314 => x"52ab518a",
          1315 => x"a53fa339",
          1316 => x"82bbe808",
          1317 => x"e4052270",
          1318 => x"852a7081",
          1319 => x"06515153",
          1320 => x"72802e8e",
          1321 => x"3882bbe8",
          1322 => x"08880508",
          1323 => x"52a0518a",
          1324 => x"813f82bb",
          1325 => x"e808e405",
          1326 => x"2270862a",
          1327 => x"70810651",
          1328 => x"51537280",
          1329 => x"2eb13882",
          1330 => x"bbe80888",
          1331 => x"050852b0",
          1332 => x"5189df3f",
          1333 => x"82bbe808",
          1334 => x"f4052253",
          1335 => x"72902e09",
          1336 => x"81069438",
          1337 => x"82bbe808",
          1338 => x"88050852",
          1339 => x"82bbe808",
          1340 => x"f8053351",
          1341 => x"89bc3f82",
          1342 => x"bbe808e4",
          1343 => x"05227088",
          1344 => x"2a708106",
          1345 => x"51515372",
          1346 => x"802eb038",
          1347 => x"82bbe808",
          1348 => x"ec0522ff",
          1349 => x"11545472",
          1350 => x"82bbe808",
          1351 => x"ec052373",
          1352 => x"902b7090",
          1353 => x"2c515380",
          1354 => x"73259038",
          1355 => x"82bbe808",
          1356 => x"88050852",
          1357 => x"b05188fa",
          1358 => x"3fd23982",
          1359 => x"bbe808e4",
          1360 => x"05227083",
          1361 => x"2a708106",
          1362 => x"51515372",
          1363 => x"802eb038",
          1364 => x"82bbe808",
          1365 => x"e80533ff",
          1366 => x"11545472",
          1367 => x"82bbe808",
          1368 => x"e8053473",
          1369 => x"982b7098",
          1370 => x"2c515380",
          1371 => x"73259038",
          1372 => x"82bbe808",
          1373 => x"88050852",
          1374 => x"b05188b6",
          1375 => x"3fd23982",
          1376 => x"bbe808e4",
          1377 => x"05227087",
          1378 => x"2a708106",
          1379 => x"51515372",
          1380 => x"b03882bb",
          1381 => x"e808ec05",
          1382 => x"22ff1154",
          1383 => x"547282bb",
          1384 => x"e808ec05",
          1385 => x"2373902b",
          1386 => x"70902c51",
          1387 => x"53807325",
          1388 => x"903882bb",
          1389 => x"e8088805",
          1390 => x"0852a051",
          1391 => x"87f43fd2",
          1392 => x"3982bbe8",
          1393 => x"08f80533",
          1394 => x"537280e3",
          1395 => x"2e098106",
          1396 => x"973882bb",
          1397 => x"e8088805",
          1398 => x"085282bb",
          1399 => x"e808fc05",
          1400 => x"335187ce",
          1401 => x"3f81ee39",
          1402 => x"82bbe808",
          1403 => x"f8053353",
          1404 => x"7280f32e",
          1405 => x"09810680",
          1406 => x"cb3882bb",
          1407 => x"e808f405",
          1408 => x"22ff1151",
          1409 => x"537282bb",
          1410 => x"e808f405",
          1411 => x"237283ff",
          1412 => x"ff065372",
          1413 => x"83ffff2e",
          1414 => x"81bb3882",
          1415 => x"bbe80888",
          1416 => x"05085282",
          1417 => x"bbe808fc",
          1418 => x"05087033",
          1419 => x"5282bbe8",
          1420 => x"08fc0508",
          1421 => x"810582bb",
          1422 => x"e808fc05",
          1423 => x"0c5386f2",
          1424 => x"3fffb739",
          1425 => x"82bbe808",
          1426 => x"f8053353",
          1427 => x"7280d32e",
          1428 => x"09810680",
          1429 => x"cb3882bb",
          1430 => x"e808f405",
          1431 => x"22ff1151",
          1432 => x"537282bb",
          1433 => x"e808f405",
          1434 => x"237283ff",
          1435 => x"ff065372",
          1436 => x"83ffff2e",
          1437 => x"80df3882",
          1438 => x"bbe80888",
          1439 => x"05085282",
          1440 => x"bbe808fc",
          1441 => x"05087033",
          1442 => x"525386a6",
          1443 => x"3f82bbe8",
          1444 => x"08fc0508",
          1445 => x"810582bb",
          1446 => x"e808fc05",
          1447 => x"0cffb739",
          1448 => x"82bbe808",
          1449 => x"f0050882",
          1450 => x"bbec2ea9",
          1451 => x"3882bbe8",
          1452 => x"08880508",
          1453 => x"5282bbe8",
          1454 => x"08f00508",
          1455 => x"ff0582bb",
          1456 => x"e808f005",
          1457 => x"0c82bbe8",
          1458 => x"08f00508",
          1459 => x"70335253",
          1460 => x"85e03fcc",
          1461 => x"3982bbe8",
          1462 => x"08e40522",
          1463 => x"70872a70",
          1464 => x"81065151",
          1465 => x"5372802e",
          1466 => x"80c33882",
          1467 => x"bbe808ec",
          1468 => x"0522ff11",
          1469 => x"54547282",
          1470 => x"bbe808ec",
          1471 => x"05237390",
          1472 => x"2b70902c",
          1473 => x"51538073",
          1474 => x"25a33882",
          1475 => x"bbe80888",
          1476 => x"050852a0",
          1477 => x"51859b3f",
          1478 => x"d23982bb",
          1479 => x"e8088805",
          1480 => x"085282bb",
          1481 => x"e808f805",
          1482 => x"33518586",
          1483 => x"3f800b82",
          1484 => x"bbe808e4",
          1485 => x"0523eab7",
          1486 => x"3982bbe8",
          1487 => x"08f80533",
          1488 => x"5372a52e",
          1489 => x"098106a8",
          1490 => x"38810b82",
          1491 => x"bbe808e4",
          1492 => x"0523800b",
          1493 => x"82bbe808",
          1494 => x"ec052380",
          1495 => x"0b82bbe8",
          1496 => x"08e80534",
          1497 => x"8a0b82bb",
          1498 => x"e808f405",
          1499 => x"23ea8039",
          1500 => x"82bbe808",
          1501 => x"88050852",
          1502 => x"82bbe808",
          1503 => x"f8053351",
          1504 => x"84b03fe9",
          1505 => x"ea3982bb",
          1506 => x"e8088805",
          1507 => x"088c1108",
          1508 => x"7082bbe8",
          1509 => x"08e0050c",
          1510 => x"515382bb",
          1511 => x"e808e005",
          1512 => x"0882bbdc",
          1513 => x"0c953d0d",
          1514 => x"82bbe80c",
          1515 => x"0482bbe8",
          1516 => x"080282bb",
          1517 => x"e80cfd3d",
          1518 => x"0d82d3ac",
          1519 => x"085382bb",
          1520 => x"e8088c05",
          1521 => x"085282bb",
          1522 => x"e8088805",
          1523 => x"0851e4dd",
          1524 => x"3f82bbdc",
          1525 => x"087082bb",
          1526 => x"dc0c5485",
          1527 => x"3d0d82bb",
          1528 => x"e80c0482",
          1529 => x"bbe80802",
          1530 => x"82bbe80c",
          1531 => x"fb3d0d80",
          1532 => x"0b82bbe8",
          1533 => x"08f8050c",
          1534 => x"82d3b008",
          1535 => x"85113370",
          1536 => x"812a7081",
          1537 => x"32708106",
          1538 => x"51515151",
          1539 => x"5372802e",
          1540 => x"8d38ff0b",
          1541 => x"82bbe808",
          1542 => x"f4050c81",
          1543 => x"923982bb",
          1544 => x"e8088805",
          1545 => x"08537233",
          1546 => x"82bbe808",
          1547 => x"88050881",
          1548 => x"0582bbe8",
          1549 => x"0888050c",
          1550 => x"537282bb",
          1551 => x"e808fc05",
          1552 => x"347281ff",
          1553 => x"06537280",
          1554 => x"2eb03882",
          1555 => x"d3b00882",
          1556 => x"d3b00853",
          1557 => x"82bbe808",
          1558 => x"fc053352",
          1559 => x"90110851",
          1560 => x"53722d82",
          1561 => x"bbdc0853",
          1562 => x"72802eff",
          1563 => x"b138ff0b",
          1564 => x"82bbe808",
          1565 => x"f8050cff",
          1566 => x"a53982d3",
          1567 => x"b00882d3",
          1568 => x"b0085353",
          1569 => x"8a519013",
          1570 => x"0853722d",
          1571 => x"82bbdc08",
          1572 => x"5372802e",
          1573 => x"8a38ff0b",
          1574 => x"82bbe808",
          1575 => x"f8050c82",
          1576 => x"bbe808f8",
          1577 => x"05087082",
          1578 => x"bbe808f4",
          1579 => x"050c5382",
          1580 => x"bbe808f4",
          1581 => x"050882bb",
          1582 => x"dc0c873d",
          1583 => x"0d82bbe8",
          1584 => x"0c0482bb",
          1585 => x"e8080282",
          1586 => x"bbe80cfb",
          1587 => x"3d0d800b",
          1588 => x"82bbe808",
          1589 => x"f8050c82",
          1590 => x"bbe8088c",
          1591 => x"05088511",
          1592 => x"3370812a",
          1593 => x"70813270",
          1594 => x"81065151",
          1595 => x"51515372",
          1596 => x"802e8d38",
          1597 => x"ff0b82bb",
          1598 => x"e808f405",
          1599 => x"0c80f339",
          1600 => x"82bbe808",
          1601 => x"88050853",
          1602 => x"723382bb",
          1603 => x"e8088805",
          1604 => x"08810582",
          1605 => x"bbe80888",
          1606 => x"050c5372",
          1607 => x"82bbe808",
          1608 => x"fc053472",
          1609 => x"81ff0653",
          1610 => x"72802eb6",
          1611 => x"3882bbe8",
          1612 => x"088c0508",
          1613 => x"82bbe808",
          1614 => x"8c050853",
          1615 => x"82bbe808",
          1616 => x"fc053352",
          1617 => x"90110851",
          1618 => x"53722d82",
          1619 => x"bbdc0853",
          1620 => x"72802eff",
          1621 => x"ab38ff0b",
          1622 => x"82bbe808",
          1623 => x"f8050cff",
          1624 => x"9f3982bb",
          1625 => x"e808f805",
          1626 => x"087082bb",
          1627 => x"e808f405",
          1628 => x"0c5382bb",
          1629 => x"e808f405",
          1630 => x"0882bbdc",
          1631 => x"0c873d0d",
          1632 => x"82bbe80c",
          1633 => x"0482bbe8",
          1634 => x"080282bb",
          1635 => x"e80cfe3d",
          1636 => x"0d82d3b0",
          1637 => x"085282bb",
          1638 => x"e8088805",
          1639 => x"0851933f",
          1640 => x"82bbdc08",
          1641 => x"7082bbdc",
          1642 => x"0c53843d",
          1643 => x"0d82bbe8",
          1644 => x"0c0482bb",
          1645 => x"e8080282",
          1646 => x"bbe80cfb",
          1647 => x"3d0d82bb",
          1648 => x"e8088c05",
          1649 => x"08851133",
          1650 => x"70812a70",
          1651 => x"81327081",
          1652 => x"06515151",
          1653 => x"51537280",
          1654 => x"2e8d38ff",
          1655 => x"0b82bbe8",
          1656 => x"08fc050c",
          1657 => x"81cb3982",
          1658 => x"bbe8088c",
          1659 => x"05088511",
          1660 => x"3370822a",
          1661 => x"70810651",
          1662 => x"51515372",
          1663 => x"802e80db",
          1664 => x"3882bbe8",
          1665 => x"088c0508",
          1666 => x"82bbe808",
          1667 => x"8c050854",
          1668 => x"548c1408",
          1669 => x"88140825",
          1670 => x"9f3882bb",
          1671 => x"e8088c05",
          1672 => x"08700870",
          1673 => x"82bbe808",
          1674 => x"88050852",
          1675 => x"57545472",
          1676 => x"75347308",
          1677 => x"8105740c",
          1678 => x"82bbe808",
          1679 => x"8c05088c",
          1680 => x"11088105",
          1681 => x"8c120c82",
          1682 => x"bbe80888",
          1683 => x"05087082",
          1684 => x"bbe808fc",
          1685 => x"050c5153",
          1686 => x"80d73982",
          1687 => x"bbe8088c",
          1688 => x"050882bb",
          1689 => x"e8088c05",
          1690 => x"085382bb",
          1691 => x"e8088805",
          1692 => x"087081ff",
          1693 => x"06539012",
          1694 => x"08515454",
          1695 => x"722d82bb",
          1696 => x"dc085372",
          1697 => x"a33882bb",
          1698 => x"e8088c05",
          1699 => x"088c1108",
          1700 => x"81058c12",
          1701 => x"0c82bbe8",
          1702 => x"08880508",
          1703 => x"7082bbe8",
          1704 => x"08fc050c",
          1705 => x"51538a39",
          1706 => x"ff0b82bb",
          1707 => x"e808fc05",
          1708 => x"0c82bbe8",
          1709 => x"08fc0508",
          1710 => x"82bbdc0c",
          1711 => x"873d0d82",
          1712 => x"bbe80c04",
          1713 => x"82bbe808",
          1714 => x"0282bbe8",
          1715 => x"0cf93d0d",
          1716 => x"82bbe808",
          1717 => x"88050885",
          1718 => x"11337081",
          1719 => x"32708106",
          1720 => x"51515152",
          1721 => x"71802e8d",
          1722 => x"38ff0b82",
          1723 => x"bbe808f8",
          1724 => x"050c8394",
          1725 => x"3982bbe8",
          1726 => x"08880508",
          1727 => x"85113370",
          1728 => x"862a7081",
          1729 => x"06515151",
          1730 => x"5271802e",
          1731 => x"80c53882",
          1732 => x"bbe80888",
          1733 => x"050882bb",
          1734 => x"e8088805",
          1735 => x"08535385",
          1736 => x"123370ff",
          1737 => x"bf065152",
          1738 => x"71851434",
          1739 => x"82bbe808",
          1740 => x"8805088c",
          1741 => x"11088105",
          1742 => x"8c120c82",
          1743 => x"bbe80888",
          1744 => x"05088411",
          1745 => x"337082bb",
          1746 => x"e808f805",
          1747 => x"0c515152",
          1748 => x"82b63982",
          1749 => x"bbe80888",
          1750 => x"05088511",
          1751 => x"3370822a",
          1752 => x"70810651",
          1753 => x"51515271",
          1754 => x"802e80d7",
          1755 => x"3882bbe8",
          1756 => x"08880508",
          1757 => x"70087033",
          1758 => x"82bbe808",
          1759 => x"fc050c51",
          1760 => x"5282bbe8",
          1761 => x"08fc0508",
          1762 => x"a93882bb",
          1763 => x"e8088805",
          1764 => x"0882bbe8",
          1765 => x"08880508",
          1766 => x"53538512",
          1767 => x"3370a007",
          1768 => x"51527185",
          1769 => x"1434ff0b",
          1770 => x"82bbe808",
          1771 => x"f8050c81",
          1772 => x"d73982bb",
          1773 => x"e8088805",
          1774 => x"08700881",
          1775 => x"05710c52",
          1776 => x"81a13982",
          1777 => x"bbe80888",
          1778 => x"050882bb",
          1779 => x"e8088805",
          1780 => x"08529411",
          1781 => x"08515271",
          1782 => x"2d82bbdc",
          1783 => x"087082bb",
          1784 => x"e808fc05",
          1785 => x"0c5282bb",
          1786 => x"e808fc05",
          1787 => x"08802580",
          1788 => x"f23882bb",
          1789 => x"e8088805",
          1790 => x"0882bbe8",
          1791 => x"08f4050c",
          1792 => x"82bbe808",
          1793 => x"88050885",
          1794 => x"113382bb",
          1795 => x"e808f005",
          1796 => x"0c5282bb",
          1797 => x"e808fc05",
          1798 => x"08ff2e09",
          1799 => x"81069538",
          1800 => x"82bbe808",
          1801 => x"f0050890",
          1802 => x"07527182",
          1803 => x"bbe808ec",
          1804 => x"05349339",
          1805 => x"82bbe808",
          1806 => x"f00508a0",
          1807 => x"07527182",
          1808 => x"bbe808ec",
          1809 => x"053482bb",
          1810 => x"e808f405",
          1811 => x"085282bb",
          1812 => x"e808ec05",
          1813 => x"33851334",
          1814 => x"ff0b82bb",
          1815 => x"e808f805",
          1816 => x"0ca63982",
          1817 => x"bbe80888",
          1818 => x"05088c11",
          1819 => x"0881058c",
          1820 => x"120c82bb",
          1821 => x"e808fc05",
          1822 => x"087081ff",
          1823 => x"067082bb",
          1824 => x"e808f805",
          1825 => x"0c515152",
          1826 => x"82bbe808",
          1827 => x"f8050882",
          1828 => x"bbdc0c89",
          1829 => x"3d0d82bb",
          1830 => x"e80c0482",
          1831 => x"bbe80802",
          1832 => x"82bbe80c",
          1833 => x"fd3d0d82",
          1834 => x"bbe80888",
          1835 => x"050882bb",
          1836 => x"e808fc05",
          1837 => x"0c82bbe8",
          1838 => x"088c0508",
          1839 => x"82bbe808",
          1840 => x"f8050c82",
          1841 => x"bbe80890",
          1842 => x"0508802e",
          1843 => x"82a23882",
          1844 => x"bbe808f8",
          1845 => x"050882bb",
          1846 => x"e808fc05",
          1847 => x"082681ac",
          1848 => x"3882bbe8",
          1849 => x"08f80508",
          1850 => x"82bbe808",
          1851 => x"90050805",
          1852 => x"5182bbe8",
          1853 => x"08fc0508",
          1854 => x"71278190",
          1855 => x"3882bbe8",
          1856 => x"08fc0508",
          1857 => x"82bbe808",
          1858 => x"90050805",
          1859 => x"82bbe808",
          1860 => x"fc050c82",
          1861 => x"bbe808f8",
          1862 => x"050882bb",
          1863 => x"e8089005",
          1864 => x"080582bb",
          1865 => x"e808f805",
          1866 => x"0c82bbe8",
          1867 => x"08900508",
          1868 => x"810582bb",
          1869 => x"e8089005",
          1870 => x"0c82bbe8",
          1871 => x"08900508",
          1872 => x"ff0582bb",
          1873 => x"e8089005",
          1874 => x"0c82bbe8",
          1875 => x"08900508",
          1876 => x"802e819c",
          1877 => x"3882bbe8",
          1878 => x"08fc0508",
          1879 => x"ff0582bb",
          1880 => x"e808fc05",
          1881 => x"0c82bbe8",
          1882 => x"08f80508",
          1883 => x"ff0582bb",
          1884 => x"e808f805",
          1885 => x"0c82bbe8",
          1886 => x"08fc0508",
          1887 => x"82bbe808",
          1888 => x"f8050853",
          1889 => x"51713371",
          1890 => x"34ffae39",
          1891 => x"82bbe808",
          1892 => x"90050881",
          1893 => x"0582bbe8",
          1894 => x"0890050c",
          1895 => x"82bbe808",
          1896 => x"900508ff",
          1897 => x"0582bbe8",
          1898 => x"0890050c",
          1899 => x"82bbe808",
          1900 => x"90050880",
          1901 => x"2eba3882",
          1902 => x"bbe808f8",
          1903 => x"05085170",
          1904 => x"3382bbe8",
          1905 => x"08f80508",
          1906 => x"810582bb",
          1907 => x"e808f805",
          1908 => x"0c82bbe8",
          1909 => x"08fc0508",
          1910 => x"52527171",
          1911 => x"3482bbe8",
          1912 => x"08fc0508",
          1913 => x"810582bb",
          1914 => x"e808fc05",
          1915 => x"0cffad39",
          1916 => x"82bbe808",
          1917 => x"88050870",
          1918 => x"82bbdc0c",
          1919 => x"51853d0d",
          1920 => x"82bbe80c",
          1921 => x"0482bbe8",
          1922 => x"080282bb",
          1923 => x"e80cfe3d",
          1924 => x"0d82bbe8",
          1925 => x"08880508",
          1926 => x"82bbe808",
          1927 => x"fc050c82",
          1928 => x"bbe808fc",
          1929 => x"05085271",
          1930 => x"3382bbe8",
          1931 => x"08fc0508",
          1932 => x"810582bb",
          1933 => x"e808fc05",
          1934 => x"0c7081ff",
          1935 => x"06515170",
          1936 => x"802e8338",
          1937 => x"da3982bb",
          1938 => x"e808fc05",
          1939 => x"08ff0582",
          1940 => x"bbe808fc",
          1941 => x"050c82bb",
          1942 => x"e808fc05",
          1943 => x"0882bbe8",
          1944 => x"08880508",
          1945 => x"317082bb",
          1946 => x"dc0c5184",
          1947 => x"3d0d82bb",
          1948 => x"e80c0482",
          1949 => x"bbe80802",
          1950 => x"82bbe80c",
          1951 => x"fe3d0d82",
          1952 => x"bbe80888",
          1953 => x"050882bb",
          1954 => x"e808fc05",
          1955 => x"0c82bbe8",
          1956 => x"088c0508",
          1957 => x"52713382",
          1958 => x"bbe8088c",
          1959 => x"05088105",
          1960 => x"82bbe808",
          1961 => x"8c050c82",
          1962 => x"bbe808fc",
          1963 => x"05085351",
          1964 => x"70723482",
          1965 => x"bbe808fc",
          1966 => x"05088105",
          1967 => x"82bbe808",
          1968 => x"fc050c70",
          1969 => x"81ff0651",
          1970 => x"70802e84",
          1971 => x"38ffbe39",
          1972 => x"82bbe808",
          1973 => x"88050870",
          1974 => x"82bbdc0c",
          1975 => x"51843d0d",
          1976 => x"82bbe80c",
          1977 => x"0482bbe8",
          1978 => x"080282bb",
          1979 => x"e80cfd3d",
          1980 => x"0d82bbe8",
          1981 => x"08880508",
          1982 => x"82bbe808",
          1983 => x"fc050c82",
          1984 => x"bbe8088c",
          1985 => x"050882bb",
          1986 => x"e808f805",
          1987 => x"0c82bbe8",
          1988 => x"08900508",
          1989 => x"802e80e5",
          1990 => x"3882bbe8",
          1991 => x"08900508",
          1992 => x"810582bb",
          1993 => x"e8089005",
          1994 => x"0c82bbe8",
          1995 => x"08900508",
          1996 => x"ff0582bb",
          1997 => x"e8089005",
          1998 => x"0c82bbe8",
          1999 => x"08900508",
          2000 => x"802eba38",
          2001 => x"82bbe808",
          2002 => x"f8050851",
          2003 => x"703382bb",
          2004 => x"e808f805",
          2005 => x"08810582",
          2006 => x"bbe808f8",
          2007 => x"050c82bb",
          2008 => x"e808fc05",
          2009 => x"08525271",
          2010 => x"713482bb",
          2011 => x"e808fc05",
          2012 => x"08810582",
          2013 => x"bbe808fc",
          2014 => x"050cffad",
          2015 => x"3982bbe8",
          2016 => x"08880508",
          2017 => x"7082bbdc",
          2018 => x"0c51853d",
          2019 => x"0d82bbe8",
          2020 => x"0c0482bb",
          2021 => x"e8080282",
          2022 => x"bbe80cfd",
          2023 => x"3d0d82bb",
          2024 => x"e8089005",
          2025 => x"08802e81",
          2026 => x"f43882bb",
          2027 => x"e8088c05",
          2028 => x"08527133",
          2029 => x"82bbe808",
          2030 => x"8c050881",
          2031 => x"0582bbe8",
          2032 => x"088c050c",
          2033 => x"82bbe808",
          2034 => x"88050870",
          2035 => x"337281ff",
          2036 => x"06535454",
          2037 => x"5171712e",
          2038 => x"843880ce",
          2039 => x"3982bbe8",
          2040 => x"08880508",
          2041 => x"52713382",
          2042 => x"bbe80888",
          2043 => x"05088105",
          2044 => x"82bbe808",
          2045 => x"88050c70",
          2046 => x"81ff0651",
          2047 => x"51708d38",
          2048 => x"800b82bb",
          2049 => x"e808fc05",
          2050 => x"0c819b39",
          2051 => x"82bbe808",
          2052 => x"900508ff",
          2053 => x"0582bbe8",
          2054 => x"0890050c",
          2055 => x"82bbe808",
          2056 => x"90050880",
          2057 => x"2e8438ff",
          2058 => x"813982bb",
          2059 => x"e8089005",
          2060 => x"08802e80",
          2061 => x"e83882bb",
          2062 => x"e8088805",
          2063 => x"08703352",
          2064 => x"53708d38",
          2065 => x"ff0b82bb",
          2066 => x"e808fc05",
          2067 => x"0c80d739",
          2068 => x"82bbe808",
          2069 => x"8c0508ff",
          2070 => x"0582bbe8",
          2071 => x"088c050c",
          2072 => x"82bbe808",
          2073 => x"8c050870",
          2074 => x"33525270",
          2075 => x"8c38810b",
          2076 => x"82bbe808",
          2077 => x"fc050cae",
          2078 => x"3982bbe8",
          2079 => x"08880508",
          2080 => x"703382bb",
          2081 => x"e8088c05",
          2082 => x"08703372",
          2083 => x"71317082",
          2084 => x"bbe808fc",
          2085 => x"050c5355",
          2086 => x"5252538a",
          2087 => x"39800b82",
          2088 => x"bbe808fc",
          2089 => x"050c82bb",
          2090 => x"e808fc05",
          2091 => x"0882bbdc",
          2092 => x"0c853d0d",
          2093 => x"82bbe80c",
          2094 => x"0482bbe8",
          2095 => x"080282bb",
          2096 => x"e80cfd3d",
          2097 => x"0d82bbe8",
          2098 => x"08880508",
          2099 => x"82bbe808",
          2100 => x"f8050c82",
          2101 => x"bbe8088c",
          2102 => x"05088d38",
          2103 => x"800b82bb",
          2104 => x"e808fc05",
          2105 => x"0c80ec39",
          2106 => x"82bbe808",
          2107 => x"f8050852",
          2108 => x"713382bb",
          2109 => x"e808f805",
          2110 => x"08810582",
          2111 => x"bbe808f8",
          2112 => x"050c7081",
          2113 => x"ff065151",
          2114 => x"70802e9f",
          2115 => x"3882bbe8",
          2116 => x"088c0508",
          2117 => x"ff0582bb",
          2118 => x"e8088c05",
          2119 => x"0c82bbe8",
          2120 => x"088c0508",
          2121 => x"ff2e8438",
          2122 => x"ffbe3982",
          2123 => x"bbe808f8",
          2124 => x"0508ff05",
          2125 => x"82bbe808",
          2126 => x"f8050c82",
          2127 => x"bbe808f8",
          2128 => x"050882bb",
          2129 => x"e8088805",
          2130 => x"08317082",
          2131 => x"bbe808fc",
          2132 => x"050c5182",
          2133 => x"bbe808fc",
          2134 => x"050882bb",
          2135 => x"dc0c853d",
          2136 => x"0d82bbe8",
          2137 => x"0c0482bb",
          2138 => x"e8080282",
          2139 => x"bbe80cfe",
          2140 => x"3d0d82bb",
          2141 => x"e8088805",
          2142 => x"0882bbe8",
          2143 => x"08fc050c",
          2144 => x"82bbe808",
          2145 => x"90050880",
          2146 => x"2e80d438",
          2147 => x"82bbe808",
          2148 => x"90050881",
          2149 => x"0582bbe8",
          2150 => x"0890050c",
          2151 => x"82bbe808",
          2152 => x"900508ff",
          2153 => x"0582bbe8",
          2154 => x"0890050c",
          2155 => x"82bbe808",
          2156 => x"90050880",
          2157 => x"2ea93882",
          2158 => x"bbe8088c",
          2159 => x"05085170",
          2160 => x"82bbe808",
          2161 => x"fc050852",
          2162 => x"52717134",
          2163 => x"82bbe808",
          2164 => x"fc050881",
          2165 => x"0582bbe8",
          2166 => x"08fc050c",
          2167 => x"ffbe3982",
          2168 => x"bbe80888",
          2169 => x"05087082",
          2170 => x"bbdc0c51",
          2171 => x"843d0d82",
          2172 => x"bbe80c04",
          2173 => x"82bbe808",
          2174 => x"0282bbe8",
          2175 => x"0cf93d0d",
          2176 => x"800b82bb",
          2177 => x"e808fc05",
          2178 => x"0c82bbe8",
          2179 => x"08880508",
          2180 => x"8025b938",
          2181 => x"82bbe808",
          2182 => x"88050830",
          2183 => x"82bbe808",
          2184 => x"88050c80",
          2185 => x"0b82bbe8",
          2186 => x"08f4050c",
          2187 => x"82bbe808",
          2188 => x"fc05088a",
          2189 => x"38810b82",
          2190 => x"bbe808f4",
          2191 => x"050c82bb",
          2192 => x"e808f405",
          2193 => x"0882bbe8",
          2194 => x"08fc050c",
          2195 => x"82bbe808",
          2196 => x"8c050880",
          2197 => x"25b93882",
          2198 => x"bbe8088c",
          2199 => x"05083082",
          2200 => x"bbe8088c",
          2201 => x"050c800b",
          2202 => x"82bbe808",
          2203 => x"f0050c82",
          2204 => x"bbe808fc",
          2205 => x"05088a38",
          2206 => x"810b82bb",
          2207 => x"e808f005",
          2208 => x"0c82bbe8",
          2209 => x"08f00508",
          2210 => x"82bbe808",
          2211 => x"fc050c80",
          2212 => x"5382bbe8",
          2213 => x"088c0508",
          2214 => x"5282bbe8",
          2215 => x"08880508",
          2216 => x"5182c53f",
          2217 => x"82bbdc08",
          2218 => x"7082bbe8",
          2219 => x"08f8050c",
          2220 => x"5482bbe8",
          2221 => x"08fc0508",
          2222 => x"802e9038",
          2223 => x"82bbe808",
          2224 => x"f8050830",
          2225 => x"82bbe808",
          2226 => x"f8050c82",
          2227 => x"bbe808f8",
          2228 => x"05087082",
          2229 => x"bbdc0c54",
          2230 => x"893d0d82",
          2231 => x"bbe80c04",
          2232 => x"82bbe808",
          2233 => x"0282bbe8",
          2234 => x"0cfb3d0d",
          2235 => x"800b82bb",
          2236 => x"e808fc05",
          2237 => x"0c82bbe8",
          2238 => x"08880508",
          2239 => x"80259938",
          2240 => x"82bbe808",
          2241 => x"88050830",
          2242 => x"82bbe808",
          2243 => x"88050c81",
          2244 => x"0b82bbe8",
          2245 => x"08fc050c",
          2246 => x"82bbe808",
          2247 => x"8c050880",
          2248 => x"25903882",
          2249 => x"bbe8088c",
          2250 => x"05083082",
          2251 => x"bbe8088c",
          2252 => x"050c8153",
          2253 => x"82bbe808",
          2254 => x"8c050852",
          2255 => x"82bbe808",
          2256 => x"88050851",
          2257 => x"81a23f82",
          2258 => x"bbdc0870",
          2259 => x"82bbe808",
          2260 => x"f8050c54",
          2261 => x"82bbe808",
          2262 => x"fc050880",
          2263 => x"2e903882",
          2264 => x"bbe808f8",
          2265 => x"05083082",
          2266 => x"bbe808f8",
          2267 => x"050c82bb",
          2268 => x"e808f805",
          2269 => x"087082bb",
          2270 => x"dc0c5487",
          2271 => x"3d0d82bb",
          2272 => x"e80c0482",
          2273 => x"bbe80802",
          2274 => x"82bbe80c",
          2275 => x"fd3d0d80",
          2276 => x"5382bbe8",
          2277 => x"088c0508",
          2278 => x"5282bbe8",
          2279 => x"08880508",
          2280 => x"5180c53f",
          2281 => x"82bbdc08",
          2282 => x"7082bbdc",
          2283 => x"0c54853d",
          2284 => x"0d82bbe8",
          2285 => x"0c0482bb",
          2286 => x"e8080282",
          2287 => x"bbe80cfd",
          2288 => x"3d0d8153",
          2289 => x"82bbe808",
          2290 => x"8c050852",
          2291 => x"82bbe808",
          2292 => x"88050851",
          2293 => x"933f82bb",
          2294 => x"dc087082",
          2295 => x"bbdc0c54",
          2296 => x"853d0d82",
          2297 => x"bbe80c04",
          2298 => x"82bbe808",
          2299 => x"0282bbe8",
          2300 => x"0cfd3d0d",
          2301 => x"810b82bb",
          2302 => x"e808fc05",
          2303 => x"0c800b82",
          2304 => x"bbe808f8",
          2305 => x"050c82bb",
          2306 => x"e8088c05",
          2307 => x"0882bbe8",
          2308 => x"08880508",
          2309 => x"27b93882",
          2310 => x"bbe808fc",
          2311 => x"0508802e",
          2312 => x"ae38800b",
          2313 => x"82bbe808",
          2314 => x"8c050824",
          2315 => x"a23882bb",
          2316 => x"e8088c05",
          2317 => x"081082bb",
          2318 => x"e8088c05",
          2319 => x"0c82bbe8",
          2320 => x"08fc0508",
          2321 => x"1082bbe8",
          2322 => x"08fc050c",
          2323 => x"ffb83982",
          2324 => x"bbe808fc",
          2325 => x"0508802e",
          2326 => x"80e13882",
          2327 => x"bbe8088c",
          2328 => x"050882bb",
          2329 => x"e8088805",
          2330 => x"0826ad38",
          2331 => x"82bbe808",
          2332 => x"88050882",
          2333 => x"bbe8088c",
          2334 => x"05083182",
          2335 => x"bbe80888",
          2336 => x"050c82bb",
          2337 => x"e808f805",
          2338 => x"0882bbe8",
          2339 => x"08fc0508",
          2340 => x"0782bbe8",
          2341 => x"08f8050c",
          2342 => x"82bbe808",
          2343 => x"fc050881",
          2344 => x"2a82bbe8",
          2345 => x"08fc050c",
          2346 => x"82bbe808",
          2347 => x"8c050881",
          2348 => x"2a82bbe8",
          2349 => x"088c050c",
          2350 => x"ff953982",
          2351 => x"bbe80890",
          2352 => x"0508802e",
          2353 => x"933882bb",
          2354 => x"e8088805",
          2355 => x"087082bb",
          2356 => x"e808f405",
          2357 => x"0c519139",
          2358 => x"82bbe808",
          2359 => x"f8050870",
          2360 => x"82bbe808",
          2361 => x"f4050c51",
          2362 => x"82bbe808",
          2363 => x"f4050882",
          2364 => x"bbdc0c85",
          2365 => x"3d0d82bb",
          2366 => x"e80c0482",
          2367 => x"bbe80802",
          2368 => x"82bbe80c",
          2369 => x"f73d0d80",
          2370 => x"0b82bbe8",
          2371 => x"08f00534",
          2372 => x"82bbe808",
          2373 => x"8c050853",
          2374 => x"80730c82",
          2375 => x"bbe80888",
          2376 => x"05087008",
          2377 => x"51537233",
          2378 => x"537282bb",
          2379 => x"e808f805",
          2380 => x"347281ff",
          2381 => x"065372a0",
          2382 => x"2e098106",
          2383 => x"913882bb",
          2384 => x"e8088805",
          2385 => x"08700881",
          2386 => x"05710c53",
          2387 => x"ce3982bb",
          2388 => x"e808f805",
          2389 => x"335372ad",
          2390 => x"2e098106",
          2391 => x"a438810b",
          2392 => x"82bbe808",
          2393 => x"f0053482",
          2394 => x"bbe80888",
          2395 => x"05087008",
          2396 => x"8105710c",
          2397 => x"70085153",
          2398 => x"723382bb",
          2399 => x"e808f805",
          2400 => x"3482bbe8",
          2401 => x"08f80533",
          2402 => x"5372b02e",
          2403 => x"09810681",
          2404 => x"dc3882bb",
          2405 => x"e8088805",
          2406 => x"08700881",
          2407 => x"05710c70",
          2408 => x"08515372",
          2409 => x"3382bbe8",
          2410 => x"08f80534",
          2411 => x"82bbe808",
          2412 => x"f8053382",
          2413 => x"bbe808e8",
          2414 => x"050c82bb",
          2415 => x"e808e805",
          2416 => x"0880e22e",
          2417 => x"b63882bb",
          2418 => x"e808e805",
          2419 => x"0880f82e",
          2420 => x"843880cd",
          2421 => x"39900b82",
          2422 => x"bbe808f4",
          2423 => x"053482bb",
          2424 => x"e8088805",
          2425 => x"08700881",
          2426 => x"05710c70",
          2427 => x"08515372",
          2428 => x"3382bbe8",
          2429 => x"08f80534",
          2430 => x"81a43982",
          2431 => x"0b82bbe8",
          2432 => x"08f40534",
          2433 => x"82bbe808",
          2434 => x"88050870",
          2435 => x"08810571",
          2436 => x"0c700851",
          2437 => x"53723382",
          2438 => x"bbe808f8",
          2439 => x"053480fe",
          2440 => x"3982bbe8",
          2441 => x"08f80533",
          2442 => x"5372a026",
          2443 => x"8d38810b",
          2444 => x"82bbe808",
          2445 => x"ec050c83",
          2446 => x"803982bb",
          2447 => x"e808f805",
          2448 => x"3353af73",
          2449 => x"27903882",
          2450 => x"bbe808f8",
          2451 => x"05335372",
          2452 => x"b9268338",
          2453 => x"8d39800b",
          2454 => x"82bbe808",
          2455 => x"ec050c82",
          2456 => x"d839880b",
          2457 => x"82bbe808",
          2458 => x"f40534b2",
          2459 => x"3982bbe8",
          2460 => x"08f80533",
          2461 => x"53af7327",
          2462 => x"903882bb",
          2463 => x"e808f805",
          2464 => x"335372b9",
          2465 => x"2683388d",
          2466 => x"39800b82",
          2467 => x"bbe808ec",
          2468 => x"050c82a5",
          2469 => x"398a0b82",
          2470 => x"bbe808f4",
          2471 => x"0534800b",
          2472 => x"82bbe808",
          2473 => x"fc050c82",
          2474 => x"bbe808f8",
          2475 => x"053353a0",
          2476 => x"732781cf",
          2477 => x"3882bbe8",
          2478 => x"08f80533",
          2479 => x"5380e073",
          2480 => x"27943882",
          2481 => x"bbe808f8",
          2482 => x"0533e011",
          2483 => x"51537282",
          2484 => x"bbe808f8",
          2485 => x"053482bb",
          2486 => x"e808f805",
          2487 => x"33d01151",
          2488 => x"537282bb",
          2489 => x"e808f805",
          2490 => x"3482bbe8",
          2491 => x"08f80533",
          2492 => x"53907327",
          2493 => x"ad3882bb",
          2494 => x"e808f805",
          2495 => x"33f91151",
          2496 => x"537282bb",
          2497 => x"e808f805",
          2498 => x"3482bbe8",
          2499 => x"08f80533",
          2500 => x"53728926",
          2501 => x"8d38800b",
          2502 => x"82bbe808",
          2503 => x"ec050c81",
          2504 => x"983982bb",
          2505 => x"e808f805",
          2506 => x"3382bbe8",
          2507 => x"08f40533",
          2508 => x"54547274",
          2509 => x"268d3880",
          2510 => x"0b82bbe8",
          2511 => x"08ec050c",
          2512 => x"80f73982",
          2513 => x"bbe808f4",
          2514 => x"05337082",
          2515 => x"bbe808fc",
          2516 => x"05082982",
          2517 => x"bbe808f8",
          2518 => x"05337012",
          2519 => x"82bbe808",
          2520 => x"fc050c82",
          2521 => x"bbe80888",
          2522 => x"05087008",
          2523 => x"8105710c",
          2524 => x"70085151",
          2525 => x"52555372",
          2526 => x"3382bbe8",
          2527 => x"08f80534",
          2528 => x"fea53982",
          2529 => x"bbe808f0",
          2530 => x"05335372",
          2531 => x"802e9038",
          2532 => x"82bbe808",
          2533 => x"fc050830",
          2534 => x"82bbe808",
          2535 => x"fc050c82",
          2536 => x"bbe8088c",
          2537 => x"050882bb",
          2538 => x"e808fc05",
          2539 => x"08710c53",
          2540 => x"810b82bb",
          2541 => x"e808ec05",
          2542 => x"0c82bbe8",
          2543 => x"08ec0508",
          2544 => x"82bbdc0c",
          2545 => x"8b3d0d82",
          2546 => x"bbe80c04",
          2547 => x"82bbe808",
          2548 => x"0282bbe8",
          2549 => x"0cf73d0d",
          2550 => x"800b82bb",
          2551 => x"e808f005",
          2552 => x"3482bbe8",
          2553 => x"088c0508",
          2554 => x"5380730c",
          2555 => x"82bbe808",
          2556 => x"88050870",
          2557 => x"08515372",
          2558 => x"33537282",
          2559 => x"bbe808f8",
          2560 => x"05347281",
          2561 => x"ff065372",
          2562 => x"a02e0981",
          2563 => x"06913882",
          2564 => x"bbe80888",
          2565 => x"05087008",
          2566 => x"8105710c",
          2567 => x"53ce3982",
          2568 => x"bbe808f8",
          2569 => x"05335372",
          2570 => x"ad2e0981",
          2571 => x"06a43881",
          2572 => x"0b82bbe8",
          2573 => x"08f00534",
          2574 => x"82bbe808",
          2575 => x"88050870",
          2576 => x"08810571",
          2577 => x"0c700851",
          2578 => x"53723382",
          2579 => x"bbe808f8",
          2580 => x"053482bb",
          2581 => x"e808f805",
          2582 => x"335372b0",
          2583 => x"2e098106",
          2584 => x"81dc3882",
          2585 => x"bbe80888",
          2586 => x"05087008",
          2587 => x"8105710c",
          2588 => x"70085153",
          2589 => x"723382bb",
          2590 => x"e808f805",
          2591 => x"3482bbe8",
          2592 => x"08f80533",
          2593 => x"82bbe808",
          2594 => x"e8050c82",
          2595 => x"bbe808e8",
          2596 => x"050880e2",
          2597 => x"2eb63882",
          2598 => x"bbe808e8",
          2599 => x"050880f8",
          2600 => x"2e843880",
          2601 => x"cd39900b",
          2602 => x"82bbe808",
          2603 => x"f4053482",
          2604 => x"bbe80888",
          2605 => x"05087008",
          2606 => x"8105710c",
          2607 => x"70085153",
          2608 => x"723382bb",
          2609 => x"e808f805",
          2610 => x"3481a439",
          2611 => x"820b82bb",
          2612 => x"e808f405",
          2613 => x"3482bbe8",
          2614 => x"08880508",
          2615 => x"70088105",
          2616 => x"710c7008",
          2617 => x"51537233",
          2618 => x"82bbe808",
          2619 => x"f8053480",
          2620 => x"fe3982bb",
          2621 => x"e808f805",
          2622 => x"335372a0",
          2623 => x"268d3881",
          2624 => x"0b82bbe8",
          2625 => x"08ec050c",
          2626 => x"83803982",
          2627 => x"bbe808f8",
          2628 => x"053353af",
          2629 => x"73279038",
          2630 => x"82bbe808",
          2631 => x"f8053353",
          2632 => x"72b92683",
          2633 => x"388d3980",
          2634 => x"0b82bbe8",
          2635 => x"08ec050c",
          2636 => x"82d83988",
          2637 => x"0b82bbe8",
          2638 => x"08f40534",
          2639 => x"b23982bb",
          2640 => x"e808f805",
          2641 => x"3353af73",
          2642 => x"27903882",
          2643 => x"bbe808f8",
          2644 => x"05335372",
          2645 => x"b9268338",
          2646 => x"8d39800b",
          2647 => x"82bbe808",
          2648 => x"ec050c82",
          2649 => x"a5398a0b",
          2650 => x"82bbe808",
          2651 => x"f4053480",
          2652 => x"0b82bbe8",
          2653 => x"08fc050c",
          2654 => x"82bbe808",
          2655 => x"f8053353",
          2656 => x"a0732781",
          2657 => x"cf3882bb",
          2658 => x"e808f805",
          2659 => x"335380e0",
          2660 => x"73279438",
          2661 => x"82bbe808",
          2662 => x"f80533e0",
          2663 => x"11515372",
          2664 => x"82bbe808",
          2665 => x"f8053482",
          2666 => x"bbe808f8",
          2667 => x"0533d011",
          2668 => x"51537282",
          2669 => x"bbe808f8",
          2670 => x"053482bb",
          2671 => x"e808f805",
          2672 => x"33539073",
          2673 => x"27ad3882",
          2674 => x"bbe808f8",
          2675 => x"0533f911",
          2676 => x"51537282",
          2677 => x"bbe808f8",
          2678 => x"053482bb",
          2679 => x"e808f805",
          2680 => x"33537289",
          2681 => x"268d3880",
          2682 => x"0b82bbe8",
          2683 => x"08ec050c",
          2684 => x"81983982",
          2685 => x"bbe808f8",
          2686 => x"053382bb",
          2687 => x"e808f405",
          2688 => x"33545472",
          2689 => x"74268d38",
          2690 => x"800b82bb",
          2691 => x"e808ec05",
          2692 => x"0c80f739",
          2693 => x"82bbe808",
          2694 => x"f4053370",
          2695 => x"82bbe808",
          2696 => x"fc050829",
          2697 => x"82bbe808",
          2698 => x"f8053370",
          2699 => x"1282bbe8",
          2700 => x"08fc050c",
          2701 => x"82bbe808",
          2702 => x"88050870",
          2703 => x"08810571",
          2704 => x"0c700851",
          2705 => x"51525553",
          2706 => x"723382bb",
          2707 => x"e808f805",
          2708 => x"34fea539",
          2709 => x"82bbe808",
          2710 => x"f0053353",
          2711 => x"72802e90",
          2712 => x"3882bbe8",
          2713 => x"08fc0508",
          2714 => x"3082bbe8",
          2715 => x"08fc050c",
          2716 => x"82bbe808",
          2717 => x"8c050882",
          2718 => x"bbe808fc",
          2719 => x"0508710c",
          2720 => x"53810b82",
          2721 => x"bbe808ec",
          2722 => x"050c82bb",
          2723 => x"e808ec05",
          2724 => x"0882bbdc",
          2725 => x"0c8b3d0d",
          2726 => x"82bbe80c",
          2727 => x"04f93d0d",
          2728 => x"79700870",
          2729 => x"56565874",
          2730 => x"802e80e3",
          2731 => x"38953975",
          2732 => x"0851e6d1",
          2733 => x"3f82bbdc",
          2734 => x"0815780c",
          2735 => x"85163354",
          2736 => x"80cd3974",
          2737 => x"335473a0",
          2738 => x"2e098106",
          2739 => x"86388115",
          2740 => x"55f13980",
          2741 => x"57769029",
          2742 => x"82b6dc05",
          2743 => x"70085256",
          2744 => x"e6a33f82",
          2745 => x"bbdc0853",
          2746 => x"74527508",
          2747 => x"51e9a33f",
          2748 => x"82bbdc08",
          2749 => x"8b388416",
          2750 => x"33547381",
          2751 => x"2effb038",
          2752 => x"81177081",
          2753 => x"ff065854",
          2754 => x"997727c9",
          2755 => x"38ff5473",
          2756 => x"82bbdc0c",
          2757 => x"893d0d04",
          2758 => x"ff3d0d73",
          2759 => x"52719326",
          2760 => x"818e3871",
          2761 => x"8429829a",
          2762 => x"9c055271",
          2763 => x"0804829f",
          2764 => x"e8518180",
          2765 => x"39829ff4",
          2766 => x"5180f939",
          2767 => x"82a08451",
          2768 => x"80f23982",
          2769 => x"a0945180",
          2770 => x"eb3982a0",
          2771 => x"a45180e4",
          2772 => x"3982a0b4",
          2773 => x"5180dd39",
          2774 => x"82a0c851",
          2775 => x"80d63982",
          2776 => x"a0d85180",
          2777 => x"cf3982a0",
          2778 => x"f05180c8",
          2779 => x"3982a188",
          2780 => x"5180c139",
          2781 => x"82a1a051",
          2782 => x"bb3982a1",
          2783 => x"bc51b539",
          2784 => x"82a1d051",
          2785 => x"af3982a1",
          2786 => x"f851a939",
          2787 => x"82a28851",
          2788 => x"a33982a2",
          2789 => x"a8519d39",
          2790 => x"82a2b851",
          2791 => x"973982a2",
          2792 => x"d0519139",
          2793 => x"82a2e851",
          2794 => x"8b3982a3",
          2795 => x"80518539",
          2796 => x"82a38c51",
          2797 => x"d8ad3f83",
          2798 => x"3d0d04fb",
          2799 => x"3d0d7779",
          2800 => x"56567487",
          2801 => x"e7268a38",
          2802 => x"74527587",
          2803 => x"e8295190",
          2804 => x"3987e852",
          2805 => x"7451efab",
          2806 => x"3f82bbdc",
          2807 => x"08527551",
          2808 => x"efa13f82",
          2809 => x"bbdc0854",
          2810 => x"79537552",
          2811 => x"82a39c51",
          2812 => x"ffbbe53f",
          2813 => x"873d0d04",
          2814 => x"ec3d0d66",
          2815 => x"02840580",
          2816 => x"e305335b",
          2817 => x"57806878",
          2818 => x"30707a07",
          2819 => x"73255157",
          2820 => x"59597856",
          2821 => x"7787ff26",
          2822 => x"83388156",
          2823 => x"74760770",
          2824 => x"81ff0651",
          2825 => x"55935674",
          2826 => x"81823881",
          2827 => x"5376528c",
          2828 => x"3d705256",
          2829 => x"8184b93f",
          2830 => x"82bbdc08",
          2831 => x"5782bbdc",
          2832 => x"08b93882",
          2833 => x"bbdc0887",
          2834 => x"c098880c",
          2835 => x"82bbdc08",
          2836 => x"59963dd4",
          2837 => x"05548480",
          2838 => x"53775275",
          2839 => x"518188f5",
          2840 => x"3f82bbdc",
          2841 => x"085782bb",
          2842 => x"dc089038",
          2843 => x"7a557480",
          2844 => x"2e893874",
          2845 => x"19751959",
          2846 => x"59d73996",
          2847 => x"3dd80551",
          2848 => x"8190de3f",
          2849 => x"76307078",
          2850 => x"0780257b",
          2851 => x"30709f2a",
          2852 => x"72065157",
          2853 => x"51567480",
          2854 => x"2e903882",
          2855 => x"a3c05387",
          2856 => x"c0988808",
          2857 => x"527851fe",
          2858 => x"923f7656",
          2859 => x"7582bbdc",
          2860 => x"0c963d0d",
          2861 => x"04f83d0d",
          2862 => x"7c028405",
          2863 => x"b7053358",
          2864 => x"59ff5880",
          2865 => x"537b527a",
          2866 => x"51fead3f",
          2867 => x"82bbdc08",
          2868 => x"a8387680",
          2869 => x"2e883876",
          2870 => x"812e9c38",
          2871 => x"9c3982d3",
          2872 => x"ac566155",
          2873 => x"605482bb",
          2874 => x"dc537f52",
          2875 => x"7e51782d",
          2876 => x"82bbdc08",
          2877 => x"58833978",
          2878 => x"047782bb",
          2879 => x"dc0c8a3d",
          2880 => x"0d04f33d",
          2881 => x"0d7f6163",
          2882 => x"028c0580",
          2883 => x"cf053373",
          2884 => x"73156841",
          2885 => x"5f5c5c5e",
          2886 => x"5e5e7a52",
          2887 => x"82a3c851",
          2888 => x"ffb9b53f",
          2889 => x"82a3d051",
          2890 => x"ffb9ad3f",
          2891 => x"80557479",
          2892 => x"27818038",
          2893 => x"7b902e89",
          2894 => x"387ba02e",
          2895 => x"a73880c6",
          2896 => x"39741853",
          2897 => x"727a278e",
          2898 => x"38722252",
          2899 => x"82a3d451",
          2900 => x"ffb9853f",
          2901 => x"893982a3",
          2902 => x"e051ffb8",
          2903 => x"fb3f8215",
          2904 => x"5580c339",
          2905 => x"74185372",
          2906 => x"7a278e38",
          2907 => x"72085282",
          2908 => x"a3c851ff",
          2909 => x"b8e23f89",
          2910 => x"3982a3dc",
          2911 => x"51ffb8d8",
          2912 => x"3f841555",
          2913 => x"a1397418",
          2914 => x"53727a27",
          2915 => x"8e387233",
          2916 => x"5282a3e8",
          2917 => x"51ffb8c0",
          2918 => x"3f893982",
          2919 => x"a3f051ff",
          2920 => x"b8b63f81",
          2921 => x"155582d3",
          2922 => x"b00852a0",
          2923 => x"51d8833f",
          2924 => x"fefc3982",
          2925 => x"a3f451ff",
          2926 => x"b89e3f80",
          2927 => x"55747927",
          2928 => x"80c63874",
          2929 => x"18703355",
          2930 => x"53805672",
          2931 => x"7a278338",
          2932 => x"81568053",
          2933 => x"9f742783",
          2934 => x"38815375",
          2935 => x"73067081",
          2936 => x"ff065153",
          2937 => x"72802e90",
          2938 => x"387380fe",
          2939 => x"268a3882",
          2940 => x"d3b00852",
          2941 => x"73518839",
          2942 => x"82d3b008",
          2943 => x"52a051d7",
          2944 => x"b13f8115",
          2945 => x"55ffb639",
          2946 => x"82a3f851",
          2947 => x"d3d53f78",
          2948 => x"18791c5c",
          2949 => x"58a0fe3f",
          2950 => x"82bbdc08",
          2951 => x"982b7098",
          2952 => x"2c515776",
          2953 => x"a02e0981",
          2954 => x"06aa38a0",
          2955 => x"e83f82bb",
          2956 => x"dc08982b",
          2957 => x"70982c70",
          2958 => x"a0327030",
          2959 => x"729b3270",
          2960 => x"30707207",
          2961 => x"73750706",
          2962 => x"51585859",
          2963 => x"57515780",
          2964 => x"7324d838",
          2965 => x"769b2e09",
          2966 => x"81068538",
          2967 => x"80538c39",
          2968 => x"7c1e5372",
          2969 => x"7826fdb2",
          2970 => x"38ff5372",
          2971 => x"82bbdc0c",
          2972 => x"8f3d0d04",
          2973 => x"fc3d0d02",
          2974 => x"9b053382",
          2975 => x"a3fc5382",
          2976 => x"a4845255",
          2977 => x"ffb6d13f",
          2978 => x"82bab422",
          2979 => x"51a9d93f",
          2980 => x"82a49054",
          2981 => x"82a49c53",
          2982 => x"82bab533",
          2983 => x"5282a4a4",
          2984 => x"51ffb6b4",
          2985 => x"3f74802e",
          2986 => x"8438a58b",
          2987 => x"3f863d0d",
          2988 => x"04fe3d0d",
          2989 => x"87c09680",
          2990 => x"0853aab6",
          2991 => x"3f81519c",
          2992 => x"c13f82a4",
          2993 => x"c0519dd6",
          2994 => x"3f80519c",
          2995 => x"b53f7281",
          2996 => x"2a708106",
          2997 => x"51527180",
          2998 => x"2e923881",
          2999 => x"519ca33f",
          3000 => x"82a4d851",
          3001 => x"9db83f80",
          3002 => x"519c973f",
          3003 => x"72822a70",
          3004 => x"81065152",
          3005 => x"71802e92",
          3006 => x"3881519c",
          3007 => x"853f82a4",
          3008 => x"e8519d9a",
          3009 => x"3f80519b",
          3010 => x"f93f7283",
          3011 => x"2a708106",
          3012 => x"51527180",
          3013 => x"2e923881",
          3014 => x"519be73f",
          3015 => x"82a4f851",
          3016 => x"9cfc3f80",
          3017 => x"519bdb3f",
          3018 => x"72842a70",
          3019 => x"81065152",
          3020 => x"71802e92",
          3021 => x"3881519b",
          3022 => x"c93f82a5",
          3023 => x"8c519cde",
          3024 => x"3f80519b",
          3025 => x"bd3f7285",
          3026 => x"2a708106",
          3027 => x"51527180",
          3028 => x"2e923881",
          3029 => x"519bab3f",
          3030 => x"82a5a051",
          3031 => x"9cc03f80",
          3032 => x"519b9f3f",
          3033 => x"72862a70",
          3034 => x"81065152",
          3035 => x"71802e92",
          3036 => x"3881519b",
          3037 => x"8d3f82a5",
          3038 => x"b4519ca2",
          3039 => x"3f80519b",
          3040 => x"813f7287",
          3041 => x"2a708106",
          3042 => x"51527180",
          3043 => x"2e923881",
          3044 => x"519aef3f",
          3045 => x"82a5c851",
          3046 => x"9c843f80",
          3047 => x"519ae33f",
          3048 => x"72882a70",
          3049 => x"81065152",
          3050 => x"71802e92",
          3051 => x"3881519a",
          3052 => x"d13f82a5",
          3053 => x"dc519be6",
          3054 => x"3f80519a",
          3055 => x"c53fa8ba",
          3056 => x"3f843d0d",
          3057 => x"04fb3d0d",
          3058 => x"77028405",
          3059 => x"a3053370",
          3060 => x"55565680",
          3061 => x"527551e3",
          3062 => x"8d3f0b0b",
          3063 => x"82b6d833",
          3064 => x"5473a938",
          3065 => x"815382a6",
          3066 => x"985282d2",
          3067 => x"dc5180fc",
          3068 => x"ff3f82bb",
          3069 => x"dc083070",
          3070 => x"82bbdc08",
          3071 => x"07802582",
          3072 => x"71315151",
          3073 => x"54730b0b",
          3074 => x"82b6d834",
          3075 => x"0b0b82b6",
          3076 => x"d8335473",
          3077 => x"812e0981",
          3078 => x"06af3882",
          3079 => x"d2dc5374",
          3080 => x"52755181",
          3081 => x"b7b03f82",
          3082 => x"bbdc0880",
          3083 => x"2e8b3882",
          3084 => x"bbdc0851",
          3085 => x"cfad3f91",
          3086 => x"3982d2dc",
          3087 => x"518189a1",
          3088 => x"3f820b0b",
          3089 => x"0b82b6d8",
          3090 => x"340b0b82",
          3091 => x"b6d83354",
          3092 => x"73822e09",
          3093 => x"81068c38",
          3094 => x"82a6a853",
          3095 => x"74527551",
          3096 => x"aeb23f80",
          3097 => x"0b82bbdc",
          3098 => x"0c873d0d",
          3099 => x"04ce3d0d",
          3100 => x"80707182",
          3101 => x"d2d80c5f",
          3102 => x"5d81527c",
          3103 => x"5180cbcb",
          3104 => x"3f82bbdc",
          3105 => x"0881ff06",
          3106 => x"59787d2e",
          3107 => x"098106a3",
          3108 => x"38963d59",
          3109 => x"835382a6",
          3110 => x"b4527851",
          3111 => x"dcc73f7c",
          3112 => x"53785282",
          3113 => x"bd885180",
          3114 => x"fae53f82",
          3115 => x"bbdc087d",
          3116 => x"2e883882",
          3117 => x"a6b85191",
          3118 => x"d5398170",
          3119 => x"5f5d82a6",
          3120 => x"f051ffb2",
          3121 => x"933f963d",
          3122 => x"70465a80",
          3123 => x"f8527951",
          3124 => x"fdf33fb4",
          3125 => x"3dff8405",
          3126 => x"51f3c23f",
          3127 => x"82bbdc08",
          3128 => x"902b7090",
          3129 => x"2c515978",
          3130 => x"80c12e89",
          3131 => x"d4387880",
          3132 => x"c12480d9",
          3133 => x"3878ab2e",
          3134 => x"83b93878",
          3135 => x"ab24a438",
          3136 => x"78822e81",
          3137 => x"b3387882",
          3138 => x"248a3878",
          3139 => x"802effae",
          3140 => x"388f8039",
          3141 => x"78842e82",
          3142 => x"83387894",
          3143 => x"2e82ad38",
          3144 => x"8ef13978",
          3145 => x"bd2e84fc",
          3146 => x"3878bd24",
          3147 => x"903878b0",
          3148 => x"2e83a638",
          3149 => x"78bc2e84",
          3150 => x"84388ed7",
          3151 => x"3978bf2e",
          3152 => x"85c43878",
          3153 => x"80c02e86",
          3154 => x"bd388ec7",
          3155 => x"397880d5",
          3156 => x"2e8da038",
          3157 => x"7880d524",
          3158 => x"b0387880",
          3159 => x"d02e8cd9",
          3160 => x"387880d0",
          3161 => x"24923878",
          3162 => x"80c22e89",
          3163 => x"fc387880",
          3164 => x"c32e8ba5",
          3165 => x"388e9c39",
          3166 => x"7880d12e",
          3167 => x"8cca3878",
          3168 => x"80d42e8c",
          3169 => x"d2388e8b",
          3170 => x"39788182",
          3171 => x"2e8de238",
          3172 => x"78818224",
          3173 => x"92387880",
          3174 => x"f82e8cf4",
          3175 => x"387880f9",
          3176 => x"2e8d9138",
          3177 => x"8ded3978",
          3178 => x"81832e8d",
          3179 => x"d3387881",
          3180 => x"852e8dd9",
          3181 => x"388ddc39",
          3182 => x"b43dff80",
          3183 => x"1153ff84",
          3184 => x"0551ec88",
          3185 => x"3f82bbdc",
          3186 => x"08883882",
          3187 => x"a6f4518f",
          3188 => x"bd39b43d",
          3189 => x"fefc1153",
          3190 => x"ff840551",
          3191 => x"ebee3f82",
          3192 => x"bbdc0880",
          3193 => x"2e883881",
          3194 => x"63258338",
          3195 => x"80430280",
          3196 => x"cb053352",
          3197 => x"0280cf05",
          3198 => x"335180c8",
          3199 => x"ce3f82bb",
          3200 => x"dc0881ff",
          3201 => x"0659788d",
          3202 => x"3882a784",
          3203 => x"51cbd43f",
          3204 => x"815efdaa",
          3205 => x"3982a794",
          3206 => x"518ef339",
          3207 => x"b43dff80",
          3208 => x"1153ff84",
          3209 => x"0551eba4",
          3210 => x"3f82bbdc",
          3211 => x"08802efd",
          3212 => x"8d388053",
          3213 => x"80520280",
          3214 => x"cf053351",
          3215 => x"80ccd93f",
          3216 => x"82bbdc08",
          3217 => x"5282a7ac",
          3218 => x"518c9f39",
          3219 => x"b43dff80",
          3220 => x"1153ff84",
          3221 => x"0551eaf4",
          3222 => x"3f82bbdc",
          3223 => x"08802e87",
          3224 => x"38638926",
          3225 => x"fcd838b4",
          3226 => x"3dfefc11",
          3227 => x"53ff8405",
          3228 => x"51ead93f",
          3229 => x"82bbdc08",
          3230 => x"863882bb",
          3231 => x"dc084363",
          3232 => x"5382a7b4",
          3233 => x"527951ff",
          3234 => x"b1b63f02",
          3235 => x"80cb0533",
          3236 => x"53795263",
          3237 => x"84b42982",
          3238 => x"bd880551",
          3239 => x"80f6f03f",
          3240 => x"82bbdc08",
          3241 => x"818c3882",
          3242 => x"a78451ca",
          3243 => x"b63f815d",
          3244 => x"fc8c39b4",
          3245 => x"3dff8405",
          3246 => x"518fc03f",
          3247 => x"82bbdc08",
          3248 => x"b53dff84",
          3249 => x"05525b90",
          3250 => x"d63f8153",
          3251 => x"82bbdc08",
          3252 => x"527a51f2",
          3253 => x"a33f80d1",
          3254 => x"39b43dff",
          3255 => x"8405518f",
          3256 => x"9a3f82bb",
          3257 => x"dc08b53d",
          3258 => x"ff840552",
          3259 => x"5b90b03f",
          3260 => x"82bbdc08",
          3261 => x"b53dff84",
          3262 => x"05525a90",
          3263 => x"a23f82bb",
          3264 => x"dc08b53d",
          3265 => x"ff840552",
          3266 => x"5990943f",
          3267 => x"82ba8058",
          3268 => x"82bc8c57",
          3269 => x"80568055",
          3270 => x"82bbdc08",
          3271 => x"81ff0654",
          3272 => x"78537952",
          3273 => x"7a51f38d",
          3274 => x"3f82bbdc",
          3275 => x"08802efb",
          3276 => x"8d3882bb",
          3277 => x"dc0851ef",
          3278 => x"df3ffb82",
          3279 => x"39b43dff",
          3280 => x"801153ff",
          3281 => x"840551e9",
          3282 => x"833f82bb",
          3283 => x"dc08802e",
          3284 => x"faec38b4",
          3285 => x"3dfefc11",
          3286 => x"53ff8405",
          3287 => x"51e8ed3f",
          3288 => x"82bbdc08",
          3289 => x"802efad6",
          3290 => x"38b43dfe",
          3291 => x"f81153ff",
          3292 => x"840551e8",
          3293 => x"d73f82bb",
          3294 => x"dc088638",
          3295 => x"82bbdc08",
          3296 => x"4282a7b8",
          3297 => x"51ffacd0",
          3298 => x"3f63635c",
          3299 => x"5a797b27",
          3300 => x"81ec3861",
          3301 => x"59787a70",
          3302 => x"84055c0c",
          3303 => x"7a7a26f5",
          3304 => x"3881db39",
          3305 => x"b43dff80",
          3306 => x"1153ff84",
          3307 => x"0551e89c",
          3308 => x"3f82bbdc",
          3309 => x"08802efa",
          3310 => x"8538b43d",
          3311 => x"fefc1153",
          3312 => x"ff840551",
          3313 => x"e8863f82",
          3314 => x"bbdc0880",
          3315 => x"2ef9ef38",
          3316 => x"b43dfef8",
          3317 => x"1153ff84",
          3318 => x"0551e7f0",
          3319 => x"3f82bbdc",
          3320 => x"08802ef9",
          3321 => x"d93882a7",
          3322 => x"c851ffab",
          3323 => x"eb3f635a",
          3324 => x"79632781",
          3325 => x"89386159",
          3326 => x"79708105",
          3327 => x"5b337934",
          3328 => x"61810542",
          3329 => x"eb39b43d",
          3330 => x"ff801153",
          3331 => x"ff840551",
          3332 => x"e7ba3f82",
          3333 => x"bbdc0880",
          3334 => x"2ef9a338",
          3335 => x"b43dfefc",
          3336 => x"1153ff84",
          3337 => x"0551e7a4",
          3338 => x"3f82bbdc",
          3339 => x"08802ef9",
          3340 => x"8d38b43d",
          3341 => x"fef81153",
          3342 => x"ff840551",
          3343 => x"e78e3f82",
          3344 => x"bbdc0880",
          3345 => x"2ef8f738",
          3346 => x"82a7d451",
          3347 => x"ffab893f",
          3348 => x"635a7963",
          3349 => x"27a83861",
          3350 => x"70337b33",
          3351 => x"5e5a5b78",
          3352 => x"7c2e9238",
          3353 => x"78557a54",
          3354 => x"79335379",
          3355 => x"5282a7e4",
          3356 => x"51ffaae4",
          3357 => x"3f811a62",
          3358 => x"8105435a",
          3359 => x"d5398a51",
          3360 => x"ca833ff8",
          3361 => x"b939b43d",
          3362 => x"ff801153",
          3363 => x"ff840551",
          3364 => x"e6ba3f82",
          3365 => x"bbdc0880",
          3366 => x"df3882ba",
          3367 => x"c8335978",
          3368 => x"802e8938",
          3369 => x"82ba8008",
          3370 => x"4480cd39",
          3371 => x"82bac933",
          3372 => x"5978802e",
          3373 => x"883882ba",
          3374 => x"880844bc",
          3375 => x"3982baca",
          3376 => x"33597880",
          3377 => x"2e883882",
          3378 => x"ba900844",
          3379 => x"ab3982ba",
          3380 => x"cb335978",
          3381 => x"802e8838",
          3382 => x"82ba9808",
          3383 => x"449a3982",
          3384 => x"bac63359",
          3385 => x"78802e88",
          3386 => x"3882baa0",
          3387 => x"08448939",
          3388 => x"82bab008",
          3389 => x"fc800544",
          3390 => x"b43dfefc",
          3391 => x"1153ff84",
          3392 => x"0551e5c8",
          3393 => x"3f82bbdc",
          3394 => x"0880de38",
          3395 => x"82bac833",
          3396 => x"5978802e",
          3397 => x"893882ba",
          3398 => x"84084380",
          3399 => x"cc3982ba",
          3400 => x"c9335978",
          3401 => x"802e8838",
          3402 => x"82ba8c08",
          3403 => x"43bb3982",
          3404 => x"baca3359",
          3405 => x"78802e88",
          3406 => x"3882ba94",
          3407 => x"0843aa39",
          3408 => x"82bacb33",
          3409 => x"5978802e",
          3410 => x"883882ba",
          3411 => x"9c084399",
          3412 => x"3982bac6",
          3413 => x"33597880",
          3414 => x"2e883882",
          3415 => x"baa40843",
          3416 => x"883982ba",
          3417 => x"b0088805",
          3418 => x"43b43dfe",
          3419 => x"f81153ff",
          3420 => x"840551e4",
          3421 => x"d73f82bb",
          3422 => x"dc08802e",
          3423 => x"a7388062",
          3424 => x"5c5c7a88",
          3425 => x"2e833881",
          3426 => x"5c7a9032",
          3427 => x"70307072",
          3428 => x"079f2a70",
          3429 => x"7f065151",
          3430 => x"5a5a7880",
          3431 => x"2e88387a",
          3432 => x"a02e8338",
          3433 => x"884282a8",
          3434 => x"8051c4b7",
          3435 => x"3fa05563",
          3436 => x"54615362",
          3437 => x"526351ee",
          3438 => x"c93f82a8",
          3439 => x"8c5187ce",
          3440 => x"39b43dff",
          3441 => x"801153ff",
          3442 => x"840551e3",
          3443 => x"ff3f82bb",
          3444 => x"dc08802e",
          3445 => x"f5e838b4",
          3446 => x"3dfefc11",
          3447 => x"53ff8405",
          3448 => x"51e3e93f",
          3449 => x"82bbdc08",
          3450 => x"802ea438",
          3451 => x"63590280",
          3452 => x"cb053379",
          3453 => x"34638105",
          3454 => x"44b43dfe",
          3455 => x"fc1153ff",
          3456 => x"840551e3",
          3457 => x"c73f82bb",
          3458 => x"dc08e138",
          3459 => x"f5b03963",
          3460 => x"70335452",
          3461 => x"82a89851",
          3462 => x"ffa7bd3f",
          3463 => x"82d3ac08",
          3464 => x"5380f852",
          3465 => x"7951ffa8",
          3466 => x"843f7945",
          3467 => x"79335978",
          3468 => x"ae2ef58a",
          3469 => x"389f7927",
          3470 => x"9f38b43d",
          3471 => x"fefc1153",
          3472 => x"ff840551",
          3473 => x"e3863f82",
          3474 => x"bbdc0880",
          3475 => x"2e913863",
          3476 => x"590280cb",
          3477 => x"05337934",
          3478 => x"63810544",
          3479 => x"ffb13982",
          3480 => x"a8a451c2",
          3481 => x"fe3fffa7",
          3482 => x"39b43dfe",
          3483 => x"f41153ff",
          3484 => x"840551dd",
          3485 => x"863f82bb",
          3486 => x"dc08802e",
          3487 => x"f4c038b4",
          3488 => x"3dfef011",
          3489 => x"53ff8405",
          3490 => x"51dcf03f",
          3491 => x"82bbdc08",
          3492 => x"802ea538",
          3493 => x"605902be",
          3494 => x"05227970",
          3495 => x"82055b23",
          3496 => x"7841b43d",
          3497 => x"fef01153",
          3498 => x"ff840551",
          3499 => x"dccd3f82",
          3500 => x"bbdc08e0",
          3501 => x"38f48739",
          3502 => x"60702254",
          3503 => x"5282a8a8",
          3504 => x"51ffa694",
          3505 => x"3f82d3ac",
          3506 => x"085380f8",
          3507 => x"527951ff",
          3508 => x"a6db3f79",
          3509 => x"45793359",
          3510 => x"78ae2ef3",
          3511 => x"e138789f",
          3512 => x"26873860",
          3513 => x"820541d0",
          3514 => x"39b43dfe",
          3515 => x"f01153ff",
          3516 => x"840551dc",
          3517 => x"863f82bb",
          3518 => x"dc08802e",
          3519 => x"92386059",
          3520 => x"02be0522",
          3521 => x"79708205",
          3522 => x"5b237841",
          3523 => x"ffaa3982",
          3524 => x"a8a451c1",
          3525 => x"ce3fffa0",
          3526 => x"39b43dfe",
          3527 => x"f41153ff",
          3528 => x"840551db",
          3529 => x"d63f82bb",
          3530 => x"dc08802e",
          3531 => x"f39038b4",
          3532 => x"3dfef011",
          3533 => x"53ff8405",
          3534 => x"51dbc03f",
          3535 => x"82bbdc08",
          3536 => x"802ea038",
          3537 => x"6060710c",
          3538 => x"59608405",
          3539 => x"41b43dfe",
          3540 => x"f01153ff",
          3541 => x"840551db",
          3542 => x"a23f82bb",
          3543 => x"dc08e538",
          3544 => x"f2dc3960",
          3545 => x"70085452",
          3546 => x"82a8b451",
          3547 => x"ffa4e93f",
          3548 => x"82d3ac08",
          3549 => x"5380f852",
          3550 => x"7951ffa5",
          3551 => x"b03f7945",
          3552 => x"79335978",
          3553 => x"ae2ef2b6",
          3554 => x"389f7927",
          3555 => x"9b38b43d",
          3556 => x"fef01153",
          3557 => x"ff840551",
          3558 => x"dae13f82",
          3559 => x"bbdc0880",
          3560 => x"2e8d3860",
          3561 => x"60710c59",
          3562 => x"60840541",
          3563 => x"ffb53982",
          3564 => x"a8a451c0",
          3565 => x"ae3fffab",
          3566 => x"3982a8c4",
          3567 => x"51c0a43f",
          3568 => x"82519889",
          3569 => x"3ff1f739",
          3570 => x"82a8dc51",
          3571 => x"c0953fa2",
          3572 => x"5197de3f",
          3573 => x"f1e83982",
          3574 => x"a8f051c0",
          3575 => x"863f8480",
          3576 => x"810b87c0",
          3577 => x"94840c84",
          3578 => x"80810b87",
          3579 => x"c094940c",
          3580 => x"f1cc3982",
          3581 => x"a98451ff",
          3582 => x"bfe93f8c",
          3583 => x"80830b87",
          3584 => x"c094840c",
          3585 => x"8c80830b",
          3586 => x"87c09494",
          3587 => x"0cf1af39",
          3588 => x"b43dff80",
          3589 => x"1153ff84",
          3590 => x"0551dfb0",
          3591 => x"3f82bbdc",
          3592 => x"08802ef1",
          3593 => x"99386352",
          3594 => x"82a99851",
          3595 => x"ffa3a93f",
          3596 => x"63597804",
          3597 => x"b43dff80",
          3598 => x"1153ff84",
          3599 => x"0551df8c",
          3600 => x"3f82bbdc",
          3601 => x"08802ef0",
          3602 => x"f5386352",
          3603 => x"82a9b451",
          3604 => x"ffa3853f",
          3605 => x"6359782d",
          3606 => x"82bbdc08",
          3607 => x"802ef0de",
          3608 => x"3882bbdc",
          3609 => x"085282a9",
          3610 => x"d051ffa2",
          3611 => x"eb3ff0ce",
          3612 => x"3982a9ec",
          3613 => x"51ffbeeb",
          3614 => x"3fffa2bd",
          3615 => x"3ff0bf39",
          3616 => x"82aa8851",
          3617 => x"ffbedc3f",
          3618 => x"8059ffa6",
          3619 => x"3991a83f",
          3620 => x"f0ac3979",
          3621 => x"45793359",
          3622 => x"78802ef0",
          3623 => x"a1387d7d",
          3624 => x"06597880",
          3625 => x"2e81cf38",
          3626 => x"b43dff84",
          3627 => x"055183cb",
          3628 => x"3f82bbdc",
          3629 => x"085b815c",
          3630 => x"7b822eb2",
          3631 => x"387b8224",
          3632 => x"89387b81",
          3633 => x"2e8c3880",
          3634 => x"ca397b83",
          3635 => x"2ead3880",
          3636 => x"c23982aa",
          3637 => x"9c567a55",
          3638 => x"82aaa054",
          3639 => x"805382aa",
          3640 => x"a452b43d",
          3641 => x"ffb00551",
          3642 => x"ffa4d53f",
          3643 => x"b8397a52",
          3644 => x"b43dffb0",
          3645 => x"0551cafb",
          3646 => x"3fab397a",
          3647 => x"5582aaa0",
          3648 => x"54805382",
          3649 => x"aab452b4",
          3650 => x"3dffb005",
          3651 => x"51ffa4b0",
          3652 => x"3f93397a",
          3653 => x"54805382",
          3654 => x"aac052b4",
          3655 => x"3dffb005",
          3656 => x"51ffa49c",
          3657 => x"3f82ba80",
          3658 => x"5882bc8c",
          3659 => x"57805664",
          3660 => x"55805482",
          3661 => x"d8805382",
          3662 => x"d88052b4",
          3663 => x"3dffb005",
          3664 => x"51e6f23f",
          3665 => x"82bbdc08",
          3666 => x"82bbdc08",
          3667 => x"09703070",
          3668 => x"72078025",
          3669 => x"515b5b5f",
          3670 => x"805a7b83",
          3671 => x"26833881",
          3672 => x"5a787a06",
          3673 => x"5978802e",
          3674 => x"8d38811c",
          3675 => x"7081ff06",
          3676 => x"5d597bfe",
          3677 => x"c3387d81",
          3678 => x"327d8132",
          3679 => x"0759788a",
          3680 => x"387eff2e",
          3681 => x"098106ee",
          3682 => x"b53882aa",
          3683 => x"c851ffbc",
          3684 => x"d23feeaa",
          3685 => x"39f53d0d",
          3686 => x"800b82bc",
          3687 => x"8c3487c0",
          3688 => x"948c7008",
          3689 => x"54558784",
          3690 => x"80527251",
          3691 => x"d3d53f82",
          3692 => x"bbdc0890",
          3693 => x"2b750855",
          3694 => x"53878480",
          3695 => x"527351d3",
          3696 => x"c23f7282",
          3697 => x"bbdc0807",
          3698 => x"750c87c0",
          3699 => x"949c7008",
          3700 => x"54558784",
          3701 => x"80527251",
          3702 => x"d3a93f82",
          3703 => x"bbdc0890",
          3704 => x"2b750855",
          3705 => x"53878480",
          3706 => x"527351d3",
          3707 => x"963f7282",
          3708 => x"bbdc0807",
          3709 => x"750c8c80",
          3710 => x"830b87c0",
          3711 => x"94840c8c",
          3712 => x"80830b87",
          3713 => x"c094940c",
          3714 => x"80fa9a5a",
          3715 => x"80fd865b",
          3716 => x"83028405",
          3717 => x"99053480",
          3718 => x"5c82d3ac",
          3719 => x"0b873d70",
          3720 => x"88130c70",
          3721 => x"720c82d3",
          3722 => x"b00c5489",
          3723 => x"be3f93c2",
          3724 => x"3f82aad8",
          3725 => x"51ffbbab",
          3726 => x"3f82aae4",
          3727 => x"51ffbba3",
          3728 => x"3f80ddb1",
          3729 => x"5192e53f",
          3730 => x"8151e8a8",
          3731 => x"3fec9e3f",
          3732 => x"8004fe3d",
          3733 => x"0d805283",
          3734 => x"5371882b",
          3735 => x"5287d83f",
          3736 => x"82bbdc08",
          3737 => x"81ff0672",
          3738 => x"07ff1454",
          3739 => x"52728025",
          3740 => x"e8387182",
          3741 => x"bbdc0c84",
          3742 => x"3d0d04fc",
          3743 => x"3d0d7670",
          3744 => x"08545580",
          3745 => x"73525472",
          3746 => x"742e818a",
          3747 => x"38723351",
          3748 => x"70a02e09",
          3749 => x"81068638",
          3750 => x"811353f1",
          3751 => x"39723351",
          3752 => x"70a22e09",
          3753 => x"81068638",
          3754 => x"81135381",
          3755 => x"54725273",
          3756 => x"812e0981",
          3757 => x"069f3884",
          3758 => x"39811252",
          3759 => x"80723352",
          3760 => x"5470a22e",
          3761 => x"83388154",
          3762 => x"70802e9d",
          3763 => x"3873ea38",
          3764 => x"98398112",
          3765 => x"52807233",
          3766 => x"525470a0",
          3767 => x"2e833881",
          3768 => x"5470802e",
          3769 => x"843873ea",
          3770 => x"38807233",
          3771 => x"525470a0",
          3772 => x"2e098106",
          3773 => x"83388154",
          3774 => x"70a23270",
          3775 => x"30708025",
          3776 => x"76075151",
          3777 => x"5170802e",
          3778 => x"88388072",
          3779 => x"70810554",
          3780 => x"3471750c",
          3781 => x"72517082",
          3782 => x"bbdc0c86",
          3783 => x"3d0d04fc",
          3784 => x"3d0d7653",
          3785 => x"7208802e",
          3786 => x"9138863d",
          3787 => x"fc055272",
          3788 => x"51d3c83f",
          3789 => x"82bbdc08",
          3790 => x"85388053",
          3791 => x"83397453",
          3792 => x"7282bbdc",
          3793 => x"0c863d0d",
          3794 => x"04fc3d0d",
          3795 => x"76821133",
          3796 => x"ff055253",
          3797 => x"8152708b",
          3798 => x"26819838",
          3799 => x"831333ff",
          3800 => x"05518252",
          3801 => x"709e2681",
          3802 => x"8a388413",
          3803 => x"33518352",
          3804 => x"70972680",
          3805 => x"fe388513",
          3806 => x"33518452",
          3807 => x"70bb2680",
          3808 => x"f2388613",
          3809 => x"33518552",
          3810 => x"70bb2680",
          3811 => x"e6388813",
          3812 => x"22558652",
          3813 => x"7487e726",
          3814 => x"80d9388a",
          3815 => x"13225487",
          3816 => x"527387e7",
          3817 => x"2680cc38",
          3818 => x"810b87c0",
          3819 => x"989c0c72",
          3820 => x"2287c098",
          3821 => x"bc0c8213",
          3822 => x"3387c098",
          3823 => x"b80c8313",
          3824 => x"3387c098",
          3825 => x"b40c8413",
          3826 => x"3387c098",
          3827 => x"b00c8513",
          3828 => x"3387c098",
          3829 => x"ac0c8613",
          3830 => x"3387c098",
          3831 => x"a80c7487",
          3832 => x"c098a40c",
          3833 => x"7387c098",
          3834 => x"a00c800b",
          3835 => x"87c0989c",
          3836 => x"0c805271",
          3837 => x"82bbdc0c",
          3838 => x"863d0d04",
          3839 => x"f33d0d7f",
          3840 => x"5b87c098",
          3841 => x"9c5d817d",
          3842 => x"0c87c098",
          3843 => x"bc085e7d",
          3844 => x"7b2387c0",
          3845 => x"98b8085a",
          3846 => x"79821c34",
          3847 => x"87c098b4",
          3848 => x"085a7983",
          3849 => x"1c3487c0",
          3850 => x"98b0085a",
          3851 => x"79841c34",
          3852 => x"87c098ac",
          3853 => x"085a7985",
          3854 => x"1c3487c0",
          3855 => x"98a8085a",
          3856 => x"79861c34",
          3857 => x"87c098a4",
          3858 => x"085c7b88",
          3859 => x"1c2387c0",
          3860 => x"98a0085a",
          3861 => x"798a1c23",
          3862 => x"807d0c79",
          3863 => x"83ffff06",
          3864 => x"597b83ff",
          3865 => x"ff065886",
          3866 => x"1b335785",
          3867 => x"1b335684",
          3868 => x"1b335583",
          3869 => x"1b335482",
          3870 => x"1b33537d",
          3871 => x"83ffff06",
          3872 => x"5282aafc",
          3873 => x"51ff9ad0",
          3874 => x"3f8f3d0d",
          3875 => x"04fb3d0d",
          3876 => x"029f0533",
          3877 => x"82b9fc33",
          3878 => x"7081ff06",
          3879 => x"58555587",
          3880 => x"c0948451",
          3881 => x"75802e86",
          3882 => x"3887c094",
          3883 => x"94517008",
          3884 => x"70962a70",
          3885 => x"81065354",
          3886 => x"5270802e",
          3887 => x"8c387191",
          3888 => x"2a708106",
          3889 => x"515170d7",
          3890 => x"38728132",
          3891 => x"70810651",
          3892 => x"5170802e",
          3893 => x"8d387193",
          3894 => x"2a708106",
          3895 => x"515170ff",
          3896 => x"be387381",
          3897 => x"ff065187",
          3898 => x"c0948052",
          3899 => x"70802e86",
          3900 => x"3887c094",
          3901 => x"90527472",
          3902 => x"0c7482bb",
          3903 => x"dc0c873d",
          3904 => x"0d04ff3d",
          3905 => x"0d028f05",
          3906 => x"33703070",
          3907 => x"9f2a5152",
          3908 => x"527082b9",
          3909 => x"fc34833d",
          3910 => x"0d04f93d",
          3911 => x"0d02a705",
          3912 => x"3358778a",
          3913 => x"2e098106",
          3914 => x"87387a52",
          3915 => x"8d51eb3f",
          3916 => x"82b9fc33",
          3917 => x"7081ff06",
          3918 => x"585687c0",
          3919 => x"94845376",
          3920 => x"802e8638",
          3921 => x"87c09494",
          3922 => x"53720870",
          3923 => x"962a7081",
          3924 => x"06555654",
          3925 => x"72802e8c",
          3926 => x"3873912a",
          3927 => x"70810651",
          3928 => x"5372d738",
          3929 => x"74813270",
          3930 => x"81065153",
          3931 => x"72802e8d",
          3932 => x"3873932a",
          3933 => x"70810651",
          3934 => x"5372ffbe",
          3935 => x"387581ff",
          3936 => x"065387c0",
          3937 => x"94805472",
          3938 => x"802e8638",
          3939 => x"87c09490",
          3940 => x"5477740c",
          3941 => x"800b82bb",
          3942 => x"dc0c893d",
          3943 => x"0d04f93d",
          3944 => x"0d795480",
          3945 => x"74337081",
          3946 => x"ff065353",
          3947 => x"5770772e",
          3948 => x"80fc3871",
          3949 => x"81ff0681",
          3950 => x"1582b9fc",
          3951 => x"337081ff",
          3952 => x"06595755",
          3953 => x"5887c094",
          3954 => x"84517580",
          3955 => x"2e863887",
          3956 => x"c0949451",
          3957 => x"70087096",
          3958 => x"2a708106",
          3959 => x"53545270",
          3960 => x"802e8c38",
          3961 => x"71912a70",
          3962 => x"81065151",
          3963 => x"70d73872",
          3964 => x"81327081",
          3965 => x"06515170",
          3966 => x"802e8d38",
          3967 => x"71932a70",
          3968 => x"81065151",
          3969 => x"70ffbe38",
          3970 => x"7481ff06",
          3971 => x"5187c094",
          3972 => x"80527080",
          3973 => x"2e863887",
          3974 => x"c0949052",
          3975 => x"77720c81",
          3976 => x"17743370",
          3977 => x"81ff0653",
          3978 => x"535770ff",
          3979 => x"86387682",
          3980 => x"bbdc0c89",
          3981 => x"3d0d04fe",
          3982 => x"3d0d82b9",
          3983 => x"fc337081",
          3984 => x"ff065452",
          3985 => x"87c09484",
          3986 => x"5172802e",
          3987 => x"863887c0",
          3988 => x"94945170",
          3989 => x"0870822a",
          3990 => x"70810651",
          3991 => x"51517080",
          3992 => x"2ee23871",
          3993 => x"81ff0651",
          3994 => x"87c09480",
          3995 => x"5270802e",
          3996 => x"863887c0",
          3997 => x"94905271",
          3998 => x"087081ff",
          3999 => x"0682bbdc",
          4000 => x"0c51843d",
          4001 => x"0d04ffaf",
          4002 => x"3f82bbdc",
          4003 => x"0881ff06",
          4004 => x"82bbdc0c",
          4005 => x"04fe3d0d",
          4006 => x"82b9fc33",
          4007 => x"7081ff06",
          4008 => x"525387c0",
          4009 => x"94845270",
          4010 => x"802e8638",
          4011 => x"87c09494",
          4012 => x"52710870",
          4013 => x"822a7081",
          4014 => x"06515151",
          4015 => x"ff527080",
          4016 => x"2ea03872",
          4017 => x"81ff0651",
          4018 => x"87c09480",
          4019 => x"5270802e",
          4020 => x"863887c0",
          4021 => x"94905271",
          4022 => x"0870982b",
          4023 => x"70982c51",
          4024 => x"53517182",
          4025 => x"bbdc0c84",
          4026 => x"3d0d04ff",
          4027 => x"3d0d87c0",
          4028 => x"9e800870",
          4029 => x"9c2a8a06",
          4030 => x"51517080",
          4031 => x"2e84b438",
          4032 => x"87c09ea4",
          4033 => x"0882ba80",
          4034 => x"0c87c09e",
          4035 => x"a80882ba",
          4036 => x"840c87c0",
          4037 => x"9e940882",
          4038 => x"ba880c87",
          4039 => x"c09e9808",
          4040 => x"82ba8c0c",
          4041 => x"87c09e9c",
          4042 => x"0882ba90",
          4043 => x"0c87c09e",
          4044 => x"a00882ba",
          4045 => x"940c87c0",
          4046 => x"9eac0882",
          4047 => x"ba980c87",
          4048 => x"c09eb008",
          4049 => x"82ba9c0c",
          4050 => x"87c09eb4",
          4051 => x"0882baa0",
          4052 => x"0c87c09e",
          4053 => x"b80882ba",
          4054 => x"a40c87c0",
          4055 => x"9ebc0882",
          4056 => x"baa80c87",
          4057 => x"c09ec008",
          4058 => x"82baac0c",
          4059 => x"87c09ec4",
          4060 => x"0882bab0",
          4061 => x"0c87c09e",
          4062 => x"80085170",
          4063 => x"82bab423",
          4064 => x"87c09e84",
          4065 => x"0882bab8",
          4066 => x"0c87c09e",
          4067 => x"880882ba",
          4068 => x"bc0c87c0",
          4069 => x"9e8c0882",
          4070 => x"bac00c81",
          4071 => x"0b82bac4",
          4072 => x"34800b87",
          4073 => x"c09e9008",
          4074 => x"7084800a",
          4075 => x"06515252",
          4076 => x"70802e83",
          4077 => x"38815271",
          4078 => x"82bac534",
          4079 => x"800b87c0",
          4080 => x"9e900870",
          4081 => x"88800a06",
          4082 => x"51525270",
          4083 => x"802e8338",
          4084 => x"81527182",
          4085 => x"bac63480",
          4086 => x"0b87c09e",
          4087 => x"90087090",
          4088 => x"800a0651",
          4089 => x"52527080",
          4090 => x"2e833881",
          4091 => x"527182ba",
          4092 => x"c734800b",
          4093 => x"87c09e90",
          4094 => x"08708880",
          4095 => x"80065152",
          4096 => x"5270802e",
          4097 => x"83388152",
          4098 => x"7182bac8",
          4099 => x"34800b87",
          4100 => x"c09e9008",
          4101 => x"70a08080",
          4102 => x"06515252",
          4103 => x"70802e83",
          4104 => x"38815271",
          4105 => x"82bac934",
          4106 => x"800b87c0",
          4107 => x"9e900870",
          4108 => x"90808006",
          4109 => x"51525270",
          4110 => x"802e8338",
          4111 => x"81527182",
          4112 => x"baca3480",
          4113 => x"0b87c09e",
          4114 => x"90087084",
          4115 => x"80800651",
          4116 => x"52527080",
          4117 => x"2e833881",
          4118 => x"527182ba",
          4119 => x"cb34800b",
          4120 => x"87c09e90",
          4121 => x"08708280",
          4122 => x"80065152",
          4123 => x"5270802e",
          4124 => x"83388152",
          4125 => x"7182bacc",
          4126 => x"34800b87",
          4127 => x"c09e9008",
          4128 => x"70818080",
          4129 => x"06515252",
          4130 => x"70802e83",
          4131 => x"38815271",
          4132 => x"82bacd34",
          4133 => x"800b87c0",
          4134 => x"9e900870",
          4135 => x"80c08006",
          4136 => x"51525270",
          4137 => x"802e8338",
          4138 => x"81527182",
          4139 => x"bace3480",
          4140 => x"0b87c09e",
          4141 => x"900870a0",
          4142 => x"80065152",
          4143 => x"5270802e",
          4144 => x"83388152",
          4145 => x"7182bacf",
          4146 => x"3487c09e",
          4147 => x"90087098",
          4148 => x"8006708a",
          4149 => x"2a515151",
          4150 => x"7082bad0",
          4151 => x"34800b87",
          4152 => x"c09e9008",
          4153 => x"70848006",
          4154 => x"51525270",
          4155 => x"802e8338",
          4156 => x"81527182",
          4157 => x"bad13487",
          4158 => x"c09e9008",
          4159 => x"7083f006",
          4160 => x"70842a51",
          4161 => x"51517082",
          4162 => x"bad23480",
          4163 => x"0b87c09e",
          4164 => x"90087088",
          4165 => x"06515252",
          4166 => x"70802e83",
          4167 => x"38815271",
          4168 => x"82bad334",
          4169 => x"87c09e90",
          4170 => x"08708706",
          4171 => x"51517082",
          4172 => x"bad43483",
          4173 => x"3d0d04fb",
          4174 => x"3d0d82ab",
          4175 => x"9451ffad",
          4176 => x"a23f82ba",
          4177 => x"c4335473",
          4178 => x"802e8938",
          4179 => x"82aba851",
          4180 => x"ffad903f",
          4181 => x"82abbc51",
          4182 => x"ffad883f",
          4183 => x"82bac633",
          4184 => x"5473802e",
          4185 => x"943882ba",
          4186 => x"a00882ba",
          4187 => x"a4081154",
          4188 => x"5282abd4",
          4189 => x"51ff90e0",
          4190 => x"3f82bacb",
          4191 => x"33547380",
          4192 => x"2e943882",
          4193 => x"ba980882",
          4194 => x"ba9c0811",
          4195 => x"545282ab",
          4196 => x"f051ff90",
          4197 => x"c33f82ba",
          4198 => x"c8335473",
          4199 => x"802e9438",
          4200 => x"82ba8008",
          4201 => x"82ba8408",
          4202 => x"11545282",
          4203 => x"ac8c51ff",
          4204 => x"90a63f82",
          4205 => x"bac93354",
          4206 => x"73802e94",
          4207 => x"3882ba88",
          4208 => x"0882ba8c",
          4209 => x"08115452",
          4210 => x"82aca851",
          4211 => x"ff90893f",
          4212 => x"82baca33",
          4213 => x"5473802e",
          4214 => x"943882ba",
          4215 => x"900882ba",
          4216 => x"94081154",
          4217 => x"5282acc4",
          4218 => x"51ff8fec",
          4219 => x"3f82bacf",
          4220 => x"33547380",
          4221 => x"2e8e3882",
          4222 => x"bad03352",
          4223 => x"82ace051",
          4224 => x"ff8fd53f",
          4225 => x"82bad333",
          4226 => x"5473802e",
          4227 => x"8e3882ba",
          4228 => x"d4335282",
          4229 => x"ad8051ff",
          4230 => x"8fbe3f82",
          4231 => x"bad13354",
          4232 => x"73802e8e",
          4233 => x"3882bad2",
          4234 => x"335282ad",
          4235 => x"a051ff8f",
          4236 => x"a73f82ba",
          4237 => x"c5335473",
          4238 => x"802e8938",
          4239 => x"82adc051",
          4240 => x"ffaba03f",
          4241 => x"82bac733",
          4242 => x"5473802e",
          4243 => x"893882ad",
          4244 => x"d451ffab",
          4245 => x"8e3f82ba",
          4246 => x"cc335473",
          4247 => x"802e8938",
          4248 => x"82ade051",
          4249 => x"ffaafc3f",
          4250 => x"82bacd33",
          4251 => x"5473802e",
          4252 => x"893882ad",
          4253 => x"ec51ffaa",
          4254 => x"ea3f82ba",
          4255 => x"ce335473",
          4256 => x"802e8938",
          4257 => x"82adf851",
          4258 => x"ffaad83f",
          4259 => x"82ae8451",
          4260 => x"ffaad03f",
          4261 => x"82baa808",
          4262 => x"5282ae90",
          4263 => x"51ff8eb8",
          4264 => x"3f82baac",
          4265 => x"085282ae",
          4266 => x"b851ff8e",
          4267 => x"ab3f82ba",
          4268 => x"b0085282",
          4269 => x"aee051ff",
          4270 => x"8e9e3f82",
          4271 => x"af8851ff",
          4272 => x"aaa13f82",
          4273 => x"bab42252",
          4274 => x"82af9051",
          4275 => x"ff8e893f",
          4276 => x"82bab808",
          4277 => x"56bd84c0",
          4278 => x"527551c1",
          4279 => x"a63f82bb",
          4280 => x"dc08bd84",
          4281 => x"c0297671",
          4282 => x"31545482",
          4283 => x"bbdc0852",
          4284 => x"82afb851",
          4285 => x"ff8de13f",
          4286 => x"82bacb33",
          4287 => x"5473802e",
          4288 => x"a93882ba",
          4289 => x"bc0856bd",
          4290 => x"84c05275",
          4291 => x"51c0f43f",
          4292 => x"82bbdc08",
          4293 => x"bd84c029",
          4294 => x"76713154",
          4295 => x"5482bbdc",
          4296 => x"085282af",
          4297 => x"e451ff8d",
          4298 => x"af3f82ba",
          4299 => x"c6335473",
          4300 => x"802ea938",
          4301 => x"82bac008",
          4302 => x"56bd84c0",
          4303 => x"527551c0",
          4304 => x"c23f82bb",
          4305 => x"dc08bd84",
          4306 => x"c0297671",
          4307 => x"31545482",
          4308 => x"bbdc0852",
          4309 => x"82b09051",
          4310 => x"ff8cfd3f",
          4311 => x"82a7fc51",
          4312 => x"ffa9803f",
          4313 => x"873d0d04",
          4314 => x"fe3d0d02",
          4315 => x"920533ff",
          4316 => x"05527184",
          4317 => x"26aa3871",
          4318 => x"8429829a",
          4319 => x"ec055271",
          4320 => x"080482b0",
          4321 => x"bc519d39",
          4322 => x"82b0c451",
          4323 => x"973982b0",
          4324 => x"cc519139",
          4325 => x"82b0d451",
          4326 => x"8b3982b0",
          4327 => x"d8518539",
          4328 => x"82b0e051",
          4329 => x"ffa8bc3f",
          4330 => x"843d0d04",
          4331 => x"7188800c",
          4332 => x"04ff3d0d",
          4333 => x"87c09684",
          4334 => x"70085252",
          4335 => x"80720c70",
          4336 => x"74077082",
          4337 => x"bad80c72",
          4338 => x"0c833d0d",
          4339 => x"04ff3d0d",
          4340 => x"87c09684",
          4341 => x"700882ba",
          4342 => x"d80c5280",
          4343 => x"720c7309",
          4344 => x"7082bad8",
          4345 => x"08067082",
          4346 => x"bad80c73",
          4347 => x"0c51833d",
          4348 => x"0d04800b",
          4349 => x"87c09684",
          4350 => x"0c0482ba",
          4351 => x"d80887c0",
          4352 => x"96840c04",
          4353 => x"fd3d0d76",
          4354 => x"982b7098",
          4355 => x"2c79982b",
          4356 => x"70982c72",
          4357 => x"10137082",
          4358 => x"2b515351",
          4359 => x"54515180",
          4360 => x"0b82b0ec",
          4361 => x"12335553",
          4362 => x"7174259c",
          4363 => x"3882b0e8",
          4364 => x"11081202",
          4365 => x"84059705",
          4366 => x"33713352",
          4367 => x"52527072",
          4368 => x"2e098106",
          4369 => x"83388153",
          4370 => x"7282bbdc",
          4371 => x"0c853d0d",
          4372 => x"04fb3d0d",
          4373 => x"79028405",
          4374 => x"a3053371",
          4375 => x"33555654",
          4376 => x"72802eb1",
          4377 => x"3882d3b0",
          4378 => x"08528851",
          4379 => x"ffaac33f",
          4380 => x"82d3b008",
          4381 => x"52a051ff",
          4382 => x"aab83f82",
          4383 => x"d3b00852",
          4384 => x"8851ffaa",
          4385 => x"ad3f7333",
          4386 => x"ff055372",
          4387 => x"74347281",
          4388 => x"ff0653cc",
          4389 => x"397751ff",
          4390 => x"8abe3f74",
          4391 => x"7434873d",
          4392 => x"0d04f63d",
          4393 => x"0d7c0284",
          4394 => x"05b70533",
          4395 => x"028805bb",
          4396 => x"053382bb",
          4397 => x"b4337084",
          4398 => x"2982badc",
          4399 => x"05700851",
          4400 => x"59595a58",
          4401 => x"5974802e",
          4402 => x"86387451",
          4403 => x"9afa3f82",
          4404 => x"bbb43370",
          4405 => x"842982ba",
          4406 => x"dc058119",
          4407 => x"70545856",
          4408 => x"5a9dfb3f",
          4409 => x"82bbdc08",
          4410 => x"750c82bb",
          4411 => x"b4337084",
          4412 => x"2982badc",
          4413 => x"05700851",
          4414 => x"565a7480",
          4415 => x"2ea73875",
          4416 => x"53785274",
          4417 => x"51ffb3dd",
          4418 => x"3f82bbb4",
          4419 => x"33810555",
          4420 => x"7482bbb4",
          4421 => x"347481ff",
          4422 => x"06559375",
          4423 => x"27873880",
          4424 => x"0b82bbb4",
          4425 => x"3477802e",
          4426 => x"b63882bb",
          4427 => x"b0085675",
          4428 => x"802eac38",
          4429 => x"82bbac33",
          4430 => x"5574a438",
          4431 => x"8c3dfc05",
          4432 => x"54765378",
          4433 => x"52755180",
          4434 => x"da883f82",
          4435 => x"bbb00852",
          4436 => x"8a51818f",
          4437 => x"953f82bb",
          4438 => x"b0085180",
          4439 => x"dde53f8c",
          4440 => x"3d0d04fd",
          4441 => x"3d0d82ba",
          4442 => x"dc539354",
          4443 => x"72085271",
          4444 => x"802e8938",
          4445 => x"715199d0",
          4446 => x"3f80730c",
          4447 => x"ff148414",
          4448 => x"54547380",
          4449 => x"25e63880",
          4450 => x"0b82bbb4",
          4451 => x"3482bbb0",
          4452 => x"08527180",
          4453 => x"2e953871",
          4454 => x"5180dec5",
          4455 => x"3f82bbb0",
          4456 => x"085199a4",
          4457 => x"3f800b82",
          4458 => x"bbb00c85",
          4459 => x"3d0d04dc",
          4460 => x"3d0d8157",
          4461 => x"805282bb",
          4462 => x"b0085180",
          4463 => x"e3b23f82",
          4464 => x"bbdc0880",
          4465 => x"d33882bb",
          4466 => x"b0085380",
          4467 => x"f852883d",
          4468 => x"70525681",
          4469 => x"8c803f82",
          4470 => x"bbdc0880",
          4471 => x"2eba3875",
          4472 => x"51ffb0a1",
          4473 => x"3f82bbdc",
          4474 => x"0855800b",
          4475 => x"82bbdc08",
          4476 => x"259d3882",
          4477 => x"bbdc08ff",
          4478 => x"05701755",
          4479 => x"55807434",
          4480 => x"75537652",
          4481 => x"811782b3",
          4482 => x"dc5257ff",
          4483 => x"87ca3f74",
          4484 => x"ff2e0981",
          4485 => x"06ffaf38",
          4486 => x"a63d0d04",
          4487 => x"d93d0daa",
          4488 => x"3d08ad3d",
          4489 => x"085a5a81",
          4490 => x"70585880",
          4491 => x"5282bbb0",
          4492 => x"085180e2",
          4493 => x"bb3f82bb",
          4494 => x"dc088195",
          4495 => x"38ff0b82",
          4496 => x"bbb00854",
          4497 => x"5580f852",
          4498 => x"8b3d7052",
          4499 => x"56818b86",
          4500 => x"3f82bbdc",
          4501 => x"08802ea5",
          4502 => x"387551ff",
          4503 => x"afa73f82",
          4504 => x"bbdc0881",
          4505 => x"18585580",
          4506 => x"0b82bbdc",
          4507 => x"08258e38",
          4508 => x"82bbdc08",
          4509 => x"ff057017",
          4510 => x"55558074",
          4511 => x"34740970",
          4512 => x"30707207",
          4513 => x"9f2a5155",
          4514 => x"5578772e",
          4515 => x"853873ff",
          4516 => x"ac3882bb",
          4517 => x"b0088c11",
          4518 => x"08535180",
          4519 => x"e1d23f82",
          4520 => x"bbdc0880",
          4521 => x"2e893882",
          4522 => x"b3e851ff",
          4523 => x"86aa3f78",
          4524 => x"772e0981",
          4525 => x"069b3875",
          4526 => x"527951ff",
          4527 => x"afb53f79",
          4528 => x"51ffaec1",
          4529 => x"3fab3d08",
          4530 => x"5482bbdc",
          4531 => x"08743480",
          4532 => x"587782bb",
          4533 => x"dc0ca93d",
          4534 => x"0d04f63d",
          4535 => x"0d7c7e71",
          4536 => x"5c717233",
          4537 => x"57595a58",
          4538 => x"73a02e09",
          4539 => x"8106a238",
          4540 => x"78337805",
          4541 => x"56777627",
          4542 => x"98388117",
          4543 => x"705b7071",
          4544 => x"33565855",
          4545 => x"73a02e09",
          4546 => x"81068638",
          4547 => x"757526ea",
          4548 => x"38805473",
          4549 => x"882982bb",
          4550 => x"b8057008",
          4551 => x"5255ffad",
          4552 => x"e43f82bb",
          4553 => x"dc085379",
          4554 => x"52740851",
          4555 => x"ffb0e33f",
          4556 => x"82bbdc08",
          4557 => x"80c53884",
          4558 => x"15335574",
          4559 => x"812e8838",
          4560 => x"74822e88",
          4561 => x"38b539fc",
          4562 => x"e63fac39",
          4563 => x"811a5a8c",
          4564 => x"3dfc1153",
          4565 => x"f80551c0",
          4566 => x"f33f82bb",
          4567 => x"dc08802e",
          4568 => x"9a38ff1b",
          4569 => x"53785277",
          4570 => x"51fdb13f",
          4571 => x"82bbdc08",
          4572 => x"81ff0655",
          4573 => x"74853874",
          4574 => x"54913981",
          4575 => x"147081ff",
          4576 => x"06515482",
          4577 => x"7427ff8b",
          4578 => x"38805473",
          4579 => x"82bbdc0c",
          4580 => x"8c3d0d04",
          4581 => x"d33d0db0",
          4582 => x"3d08b23d",
          4583 => x"08b43d08",
          4584 => x"595f5a80",
          4585 => x"0baf3d34",
          4586 => x"82bbb433",
          4587 => x"82bbb008",
          4588 => x"555b7381",
          4589 => x"cb387382",
          4590 => x"bbac3355",
          4591 => x"55738338",
          4592 => x"81557680",
          4593 => x"2e81bc38",
          4594 => x"81707606",
          4595 => x"55567380",
          4596 => x"2e81ad38",
          4597 => x"a8519886",
          4598 => x"3f82bbdc",
          4599 => x"0882bbb0",
          4600 => x"0c82bbdc",
          4601 => x"08802e81",
          4602 => x"92389353",
          4603 => x"765282bb",
          4604 => x"dc085180",
          4605 => x"ccfa3f82",
          4606 => x"bbdc0880",
          4607 => x"2e8c3882",
          4608 => x"b49451ff",
          4609 => x"9fdd3f80",
          4610 => x"f73982bb",
          4611 => x"dc085b82",
          4612 => x"bbb00853",
          4613 => x"80f85290",
          4614 => x"3d705254",
          4615 => x"8187b73f",
          4616 => x"82bbdc08",
          4617 => x"5682bbdc",
          4618 => x"08742e09",
          4619 => x"810680d0",
          4620 => x"3882bbdc",
          4621 => x"0851ffab",
          4622 => x"cc3f82bb",
          4623 => x"dc085580",
          4624 => x"0b82bbdc",
          4625 => x"0825a938",
          4626 => x"82bbdc08",
          4627 => x"ff057017",
          4628 => x"55558074",
          4629 => x"34805374",
          4630 => x"81ff0652",
          4631 => x"7551f8c2",
          4632 => x"3f811b70",
          4633 => x"81ff065c",
          4634 => x"54937b27",
          4635 => x"8338805b",
          4636 => x"74ff2e09",
          4637 => x"8106ff97",
          4638 => x"38863975",
          4639 => x"82bbac34",
          4640 => x"768c3882",
          4641 => x"bbb00880",
          4642 => x"2e8438f9",
          4643 => x"d63f8f3d",
          4644 => x"5dec823f",
          4645 => x"82bbdc08",
          4646 => x"982b7098",
          4647 => x"2c515978",
          4648 => x"ff2eee38",
          4649 => x"7881ff06",
          4650 => x"82d38833",
          4651 => x"70982b70",
          4652 => x"982c82d3",
          4653 => x"84337098",
          4654 => x"2b70972c",
          4655 => x"71982c05",
          4656 => x"70842982",
          4657 => x"b0e80570",
          4658 => x"08157033",
          4659 => x"51515151",
          4660 => x"59595159",
          4661 => x"5d588156",
          4662 => x"73782e80",
          4663 => x"e9387774",
          4664 => x"27b43874",
          4665 => x"81800a29",
          4666 => x"81ff0a05",
          4667 => x"70982c51",
          4668 => x"55807524",
          4669 => x"80ce3876",
          4670 => x"53745277",
          4671 => x"51f6853f",
          4672 => x"82bbdc08",
          4673 => x"81ff0654",
          4674 => x"73802ed7",
          4675 => x"387482d3",
          4676 => x"84348156",
          4677 => x"b1397481",
          4678 => x"800a2981",
          4679 => x"800a0570",
          4680 => x"982c7081",
          4681 => x"ff065651",
          4682 => x"55739526",
          4683 => x"97387653",
          4684 => x"74527751",
          4685 => x"f5ce3f82",
          4686 => x"bbdc0881",
          4687 => x"ff065473",
          4688 => x"cc38d339",
          4689 => x"80567580",
          4690 => x"2e80ca38",
          4691 => x"811c5574",
          4692 => x"82d38834",
          4693 => x"74982b70",
          4694 => x"982c82d3",
          4695 => x"84337098",
          4696 => x"2b70982c",
          4697 => x"70101170",
          4698 => x"822b82b0",
          4699 => x"ec11335e",
          4700 => x"51515157",
          4701 => x"58515574",
          4702 => x"772e0981",
          4703 => x"06fe9238",
          4704 => x"82b0f014",
          4705 => x"087d0c80",
          4706 => x"0b82d388",
          4707 => x"34800b82",
          4708 => x"d3843492",
          4709 => x"397582d3",
          4710 => x"88347582",
          4711 => x"d3843478",
          4712 => x"af3d3475",
          4713 => x"7d0c7e54",
          4714 => x"739526fd",
          4715 => x"e1387384",
          4716 => x"29829b80",
          4717 => x"05547308",
          4718 => x"0482d390",
          4719 => x"3354737e",
          4720 => x"2efdcb38",
          4721 => x"82d38c33",
          4722 => x"55737527",
          4723 => x"ab387498",
          4724 => x"2b70982c",
          4725 => x"51557375",
          4726 => x"249e3874",
          4727 => x"1a547333",
          4728 => x"81153474",
          4729 => x"81800a29",
          4730 => x"81ff0a05",
          4731 => x"70982c82",
          4732 => x"d3903356",
          4733 => x"5155df39",
          4734 => x"82d39033",
          4735 => x"81115654",
          4736 => x"7482d390",
          4737 => x"34731a54",
          4738 => x"ae3d3374",
          4739 => x"3482d38c",
          4740 => x"3354737e",
          4741 => x"25893881",
          4742 => x"14547382",
          4743 => x"d38c3482",
          4744 => x"d3903370",
          4745 => x"81800a29",
          4746 => x"81ff0a05",
          4747 => x"70982c82",
          4748 => x"d38c335a",
          4749 => x"51565674",
          4750 => x"7725a838",
          4751 => x"82d3b008",
          4752 => x"52741a70",
          4753 => x"335254ff",
          4754 => x"9ee83f74",
          4755 => x"81800a29",
          4756 => x"81800a05",
          4757 => x"70982c82",
          4758 => x"d38c3356",
          4759 => x"51557375",
          4760 => x"24da3882",
          4761 => x"d3903370",
          4762 => x"982b7098",
          4763 => x"2c82d38c",
          4764 => x"335a5156",
          4765 => x"56747725",
          4766 => x"fc943882",
          4767 => x"d3b00852",
          4768 => x"8851ff9e",
          4769 => x"ad3f7481",
          4770 => x"800a2981",
          4771 => x"800a0570",
          4772 => x"982c82d3",
          4773 => x"8c335651",
          4774 => x"55737524",
          4775 => x"de38fbee",
          4776 => x"39837a34",
          4777 => x"800b811b",
          4778 => x"3482d390",
          4779 => x"53805282",
          4780 => x"a3bc51f3",
          4781 => x"9c3f81fd",
          4782 => x"3982d390",
          4783 => x"337081ff",
          4784 => x"06555573",
          4785 => x"802efbc6",
          4786 => x"3882d38c",
          4787 => x"33ff0554",
          4788 => x"7382d38c",
          4789 => x"34ff1554",
          4790 => x"7382d390",
          4791 => x"3482d3b0",
          4792 => x"08528851",
          4793 => x"ff9dcb3f",
          4794 => x"82d39033",
          4795 => x"70982b70",
          4796 => x"982c82d3",
          4797 => x"8c335751",
          4798 => x"56577474",
          4799 => x"25ad3874",
          4800 => x"1a548114",
          4801 => x"33743482",
          4802 => x"d3b00852",
          4803 => x"733351ff",
          4804 => x"9da03f74",
          4805 => x"81800a29",
          4806 => x"81800a05",
          4807 => x"70982c82",
          4808 => x"d38c3358",
          4809 => x"51557575",
          4810 => x"24d53882",
          4811 => x"d3b00852",
          4812 => x"a051ff9c",
          4813 => x"fd3f82d3",
          4814 => x"90337098",
          4815 => x"2b70982c",
          4816 => x"82d38c33",
          4817 => x"57515657",
          4818 => x"747424fa",
          4819 => x"c13882d3",
          4820 => x"b0085288",
          4821 => x"51ff9cda",
          4822 => x"3f748180",
          4823 => x"0a298180",
          4824 => x"0a057098",
          4825 => x"2c82d38c",
          4826 => x"33585155",
          4827 => x"757525de",
          4828 => x"38fa9b39",
          4829 => x"82d38c33",
          4830 => x"7a055480",
          4831 => x"743482d3",
          4832 => x"b008528a",
          4833 => x"51ff9caa",
          4834 => x"3f82d38c",
          4835 => x"527951f6",
          4836 => x"c93f82bb",
          4837 => x"dc0881ff",
          4838 => x"06547396",
          4839 => x"3882d38c",
          4840 => x"33547380",
          4841 => x"2e8f3881",
          4842 => x"53735279",
          4843 => x"51f1f33f",
          4844 => x"8439807a",
          4845 => x"34800b82",
          4846 => x"d3903480",
          4847 => x"0b82d38c",
          4848 => x"347982bb",
          4849 => x"dc0caf3d",
          4850 => x"0d0482d3",
          4851 => x"90335473",
          4852 => x"802ef9ba",
          4853 => x"3882d3b0",
          4854 => x"08528851",
          4855 => x"ff9bd33f",
          4856 => x"82d39033",
          4857 => x"ff055473",
          4858 => x"82d39034",
          4859 => x"7381ff06",
          4860 => x"54dd3982",
          4861 => x"d3903382",
          4862 => x"d38c3355",
          4863 => x"5573752e",
          4864 => x"f98c38ff",
          4865 => x"14547382",
          4866 => x"d38c3474",
          4867 => x"982b7098",
          4868 => x"2c7581ff",
          4869 => x"06565155",
          4870 => x"747425ad",
          4871 => x"38741a54",
          4872 => x"81143374",
          4873 => x"3482d3b0",
          4874 => x"08527333",
          4875 => x"51ff9b82",
          4876 => x"3f748180",
          4877 => x"0a298180",
          4878 => x"0a057098",
          4879 => x"2c82d38c",
          4880 => x"33585155",
          4881 => x"757524d5",
          4882 => x"3882d3b0",
          4883 => x"0852a051",
          4884 => x"ff9adf3f",
          4885 => x"82d39033",
          4886 => x"70982b70",
          4887 => x"982c82d3",
          4888 => x"8c335751",
          4889 => x"56577474",
          4890 => x"24f8a338",
          4891 => x"82d3b008",
          4892 => x"528851ff",
          4893 => x"9abc3f74",
          4894 => x"81800a29",
          4895 => x"81800a05",
          4896 => x"70982c82",
          4897 => x"d38c3358",
          4898 => x"51557575",
          4899 => x"25de38f7",
          4900 => x"fd3982d3",
          4901 => x"90337081",
          4902 => x"ff0682d3",
          4903 => x"8c335956",
          4904 => x"54747727",
          4905 => x"f7e83882",
          4906 => x"d3b00852",
          4907 => x"81145473",
          4908 => x"82d39034",
          4909 => x"741a7033",
          4910 => x"5254ff99",
          4911 => x"f53f82d3",
          4912 => x"90337081",
          4913 => x"ff0682d3",
          4914 => x"8c335856",
          4915 => x"54757526",
          4916 => x"d638f7ba",
          4917 => x"3982d390",
          4918 => x"53805282",
          4919 => x"a3bc51ee",
          4920 => x"f03f800b",
          4921 => x"82d39034",
          4922 => x"800b82d3",
          4923 => x"8c34f79e",
          4924 => x"397ab038",
          4925 => x"82bba808",
          4926 => x"5574802e",
          4927 => x"a6387451",
          4928 => x"ffa2823f",
          4929 => x"82bbdc08",
          4930 => x"82d38c34",
          4931 => x"82bbdc08",
          4932 => x"81ff0681",
          4933 => x"05537452",
          4934 => x"7951ffa3",
          4935 => x"c83f935b",
          4936 => x"81c0397a",
          4937 => x"842982ba",
          4938 => x"dc05fc11",
          4939 => x"08565474",
          4940 => x"802ea738",
          4941 => x"7451ffa1",
          4942 => x"cc3f82bb",
          4943 => x"dc0882d3",
          4944 => x"8c3482bb",
          4945 => x"dc0881ff",
          4946 => x"06810553",
          4947 => x"74527951",
          4948 => x"ffa3923f",
          4949 => x"ff1b5480",
          4950 => x"fa397308",
          4951 => x"5574802e",
          4952 => x"f6ac3874",
          4953 => x"51ffa19d",
          4954 => x"3f99397a",
          4955 => x"932e0981",
          4956 => x"06ae3882",
          4957 => x"badc0855",
          4958 => x"74802ea4",
          4959 => x"387451ff",
          4960 => x"a1833f82",
          4961 => x"bbdc0882",
          4962 => x"d38c3482",
          4963 => x"bbdc0881",
          4964 => x"ff068105",
          4965 => x"53745279",
          4966 => x"51ffa2c9",
          4967 => x"3f80c339",
          4968 => x"7a842982",
          4969 => x"bae00570",
          4970 => x"08565474",
          4971 => x"802eab38",
          4972 => x"7451ffa0",
          4973 => x"d03f82bb",
          4974 => x"dc0882d3",
          4975 => x"8c3482bb",
          4976 => x"dc0881ff",
          4977 => x"06810553",
          4978 => x"74527951",
          4979 => x"ffa2963f",
          4980 => x"811b5473",
          4981 => x"81ff065b",
          4982 => x"89397482",
          4983 => x"d38c3474",
          4984 => x"7a3482d3",
          4985 => x"905382d3",
          4986 => x"8c335279",
          4987 => x"51ece23f",
          4988 => x"f59c3982",
          4989 => x"d3903370",
          4990 => x"81ff0682",
          4991 => x"d38c3359",
          4992 => x"56547477",
          4993 => x"27f58738",
          4994 => x"82d3b008",
          4995 => x"52811454",
          4996 => x"7382d390",
          4997 => x"34741a70",
          4998 => x"335254ff",
          4999 => x"97943ff4",
          5000 => x"ed3982d3",
          5001 => x"90335473",
          5002 => x"802ef4e2",
          5003 => x"3882d3b0",
          5004 => x"08528851",
          5005 => x"ff96fb3f",
          5006 => x"82d39033",
          5007 => x"ff055473",
          5008 => x"82d39034",
          5009 => x"f4c839f9",
          5010 => x"3d0d83c0",
          5011 => x"800b82bb",
          5012 => x"d40c8480",
          5013 => x"0b82bbd0",
          5014 => x"23a08053",
          5015 => x"805283c0",
          5016 => x"8051ffa6",
          5017 => x"813f82bb",
          5018 => x"d4085480",
          5019 => x"58777434",
          5020 => x"81577681",
          5021 => x"153482bb",
          5022 => x"d4085477",
          5023 => x"84153476",
          5024 => x"85153482",
          5025 => x"bbd40854",
          5026 => x"77861534",
          5027 => x"76871534",
          5028 => x"82bbd408",
          5029 => x"82bbd022",
          5030 => x"ff05fe80",
          5031 => x"80077083",
          5032 => x"ffff0670",
          5033 => x"882a5851",
          5034 => x"55567488",
          5035 => x"17347389",
          5036 => x"173482bb",
          5037 => x"d0227088",
          5038 => x"2982bbd4",
          5039 => x"0805f811",
          5040 => x"51555577",
          5041 => x"82153476",
          5042 => x"83153489",
          5043 => x"3d0d04ff",
          5044 => x"3d0d7352",
          5045 => x"81518472",
          5046 => x"278f38fb",
          5047 => x"12832a82",
          5048 => x"117083ff",
          5049 => x"ff065151",
          5050 => x"517082bb",
          5051 => x"dc0c833d",
          5052 => x"0d04f93d",
          5053 => x"0d02a605",
          5054 => x"22028405",
          5055 => x"aa052271",
          5056 => x"0582bbd4",
          5057 => x"0871832b",
          5058 => x"71117483",
          5059 => x"2b731170",
          5060 => x"33811233",
          5061 => x"71882b07",
          5062 => x"02a405ae",
          5063 => x"05227181",
          5064 => x"ffff0607",
          5065 => x"70882a53",
          5066 => x"51525954",
          5067 => x"5b5b5753",
          5068 => x"54557177",
          5069 => x"34708118",
          5070 => x"3482bbd4",
          5071 => x"08147588",
          5072 => x"2a525470",
          5073 => x"82153474",
          5074 => x"83153482",
          5075 => x"bbd40870",
          5076 => x"17703381",
          5077 => x"12337188",
          5078 => x"2b077083",
          5079 => x"2b8ffff8",
          5080 => x"06515256",
          5081 => x"52710573",
          5082 => x"83ffff06",
          5083 => x"70882a54",
          5084 => x"54517182",
          5085 => x"12347281",
          5086 => x"ff065372",
          5087 => x"83123482",
          5088 => x"bbd40816",
          5089 => x"56717634",
          5090 => x"72811734",
          5091 => x"893d0d04",
          5092 => x"fb3d0d82",
          5093 => x"bbd40802",
          5094 => x"84059e05",
          5095 => x"2270832b",
          5096 => x"72118611",
          5097 => x"33871233",
          5098 => x"718b2b71",
          5099 => x"832b0758",
          5100 => x"5b595255",
          5101 => x"52720584",
          5102 => x"12338513",
          5103 => x"3371882b",
          5104 => x"0770882a",
          5105 => x"54565652",
          5106 => x"70841334",
          5107 => x"73851334",
          5108 => x"82bbd408",
          5109 => x"70148411",
          5110 => x"33851233",
          5111 => x"718b2b71",
          5112 => x"832b0756",
          5113 => x"59575272",
          5114 => x"05861233",
          5115 => x"87133371",
          5116 => x"882b0770",
          5117 => x"882a5456",
          5118 => x"56527086",
          5119 => x"13347387",
          5120 => x"133482bb",
          5121 => x"d4081370",
          5122 => x"33811233",
          5123 => x"71882b07",
          5124 => x"7081ffff",
          5125 => x"0670882a",
          5126 => x"53515353",
          5127 => x"53717334",
          5128 => x"70811434",
          5129 => x"873d0d04",
          5130 => x"fa3d0d02",
          5131 => x"a2052282",
          5132 => x"bbd40871",
          5133 => x"832b7111",
          5134 => x"70338112",
          5135 => x"3371882b",
          5136 => x"07708829",
          5137 => x"15703381",
          5138 => x"12337198",
          5139 => x"2b71902b",
          5140 => x"07535f53",
          5141 => x"55525a56",
          5142 => x"57535471",
          5143 => x"802580f6",
          5144 => x"387251fe",
          5145 => x"ab3f82bb",
          5146 => x"d4087016",
          5147 => x"70338112",
          5148 => x"33718b2b",
          5149 => x"71832b07",
          5150 => x"74117033",
          5151 => x"81123371",
          5152 => x"882b0770",
          5153 => x"832b8fff",
          5154 => x"f8065152",
          5155 => x"5451535a",
          5156 => x"58537205",
          5157 => x"74882a54",
          5158 => x"52728213",
          5159 => x"34738313",
          5160 => x"3482bbd4",
          5161 => x"08701670",
          5162 => x"33811233",
          5163 => x"718b2b71",
          5164 => x"832b0756",
          5165 => x"59575572",
          5166 => x"05703381",
          5167 => x"12337188",
          5168 => x"2b077081",
          5169 => x"ffff0670",
          5170 => x"882a5751",
          5171 => x"52585272",
          5172 => x"74347181",
          5173 => x"1534883d",
          5174 => x"0d04fb3d",
          5175 => x"0d82bbd4",
          5176 => x"08028405",
          5177 => x"9e052270",
          5178 => x"832b7211",
          5179 => x"82113383",
          5180 => x"1233718b",
          5181 => x"2b71832b",
          5182 => x"07595b59",
          5183 => x"52565273",
          5184 => x"05713381",
          5185 => x"13337188",
          5186 => x"2b07028c",
          5187 => x"05a20522",
          5188 => x"71077088",
          5189 => x"2a535153",
          5190 => x"53537173",
          5191 => x"34708114",
          5192 => x"3482bbd4",
          5193 => x"08701570",
          5194 => x"33811233",
          5195 => x"718b2b71",
          5196 => x"832b0756",
          5197 => x"59575272",
          5198 => x"05821233",
          5199 => x"83133371",
          5200 => x"882b0770",
          5201 => x"882a5455",
          5202 => x"56527082",
          5203 => x"13347283",
          5204 => x"133482bb",
          5205 => x"d4081482",
          5206 => x"11338312",
          5207 => x"3371882b",
          5208 => x"0782bbdc",
          5209 => x"0c525487",
          5210 => x"3d0d04f7",
          5211 => x"3d0d7b82",
          5212 => x"bbd40831",
          5213 => x"832a7083",
          5214 => x"ffff0670",
          5215 => x"535753fd",
          5216 => x"a73f82bb",
          5217 => x"d4087683",
          5218 => x"2b711182",
          5219 => x"11338312",
          5220 => x"33718b2b",
          5221 => x"71832b07",
          5222 => x"75117033",
          5223 => x"81123371",
          5224 => x"982b7190",
          5225 => x"2b075342",
          5226 => x"4051535b",
          5227 => x"58555954",
          5228 => x"7280258d",
          5229 => x"38828080",
          5230 => x"527551fe",
          5231 => x"9d3f8184",
          5232 => x"39841433",
          5233 => x"85153371",
          5234 => x"8b2b7183",
          5235 => x"2b077611",
          5236 => x"79882a53",
          5237 => x"51555855",
          5238 => x"76861434",
          5239 => x"7581ff06",
          5240 => x"56758714",
          5241 => x"3482bbd4",
          5242 => x"08701984",
          5243 => x"12338513",
          5244 => x"3371882b",
          5245 => x"0770882a",
          5246 => x"54575b56",
          5247 => x"53728416",
          5248 => x"34738516",
          5249 => x"3482bbd4",
          5250 => x"08185380",
          5251 => x"0b861434",
          5252 => x"800b8714",
          5253 => x"3482bbd4",
          5254 => x"08537684",
          5255 => x"14347585",
          5256 => x"143482bb",
          5257 => x"d4081870",
          5258 => x"33811233",
          5259 => x"71882b07",
          5260 => x"70828080",
          5261 => x"0770882a",
          5262 => x"53515556",
          5263 => x"54747434",
          5264 => x"72811534",
          5265 => x"8b3d0d04",
          5266 => x"ff3d0d73",
          5267 => x"5282bbd4",
          5268 => x"088438f7",
          5269 => x"f23f7180",
          5270 => x"2e863871",
          5271 => x"51fe8c3f",
          5272 => x"833d0d04",
          5273 => x"f53d0d80",
          5274 => x"7e5258f8",
          5275 => x"e23f82bb",
          5276 => x"dc0883ff",
          5277 => x"ff0682bb",
          5278 => x"d4088411",
          5279 => x"33851233",
          5280 => x"71882b07",
          5281 => x"705f5956",
          5282 => x"585a81ff",
          5283 => x"ff597578",
          5284 => x"2e80cb38",
          5285 => x"75882917",
          5286 => x"70338112",
          5287 => x"3371882b",
          5288 => x"077081ff",
          5289 => x"ff067931",
          5290 => x"7083ffff",
          5291 => x"06707f27",
          5292 => x"52535156",
          5293 => x"59557779",
          5294 => x"278a3873",
          5295 => x"802e8538",
          5296 => x"75785a5b",
          5297 => x"84153385",
          5298 => x"16337188",
          5299 => x"2b075754",
          5300 => x"75c23878",
          5301 => x"81ffff2e",
          5302 => x"85387a79",
          5303 => x"59568076",
          5304 => x"832b82bb",
          5305 => x"d4081170",
          5306 => x"33811233",
          5307 => x"71882b07",
          5308 => x"7081ffff",
          5309 => x"0651525a",
          5310 => x"565c5573",
          5311 => x"752e8338",
          5312 => x"81558054",
          5313 => x"79782681",
          5314 => x"cc387454",
          5315 => x"74802e81",
          5316 => x"c438777a",
          5317 => x"2e098106",
          5318 => x"89387551",
          5319 => x"f8f23f81",
          5320 => x"ac398280",
          5321 => x"80537952",
          5322 => x"7551f7c6",
          5323 => x"3f82bbd4",
          5324 => x"08701c86",
          5325 => x"11338712",
          5326 => x"33718b2b",
          5327 => x"71832b07",
          5328 => x"535a5e55",
          5329 => x"74057a17",
          5330 => x"7083ffff",
          5331 => x"0670882a",
          5332 => x"5c595654",
          5333 => x"78841534",
          5334 => x"7681ff06",
          5335 => x"57768515",
          5336 => x"3482bbd4",
          5337 => x"0875832b",
          5338 => x"7111721e",
          5339 => x"86113387",
          5340 => x"12337188",
          5341 => x"2b077088",
          5342 => x"2a535b5e",
          5343 => x"535a5654",
          5344 => x"73861934",
          5345 => x"75871934",
          5346 => x"82bbd408",
          5347 => x"701c8411",
          5348 => x"33851233",
          5349 => x"718b2b71",
          5350 => x"832b0753",
          5351 => x"5d5a5574",
          5352 => x"05547886",
          5353 => x"15347687",
          5354 => x"153482bb",
          5355 => x"d4087016",
          5356 => x"711d8411",
          5357 => x"33851233",
          5358 => x"71882b07",
          5359 => x"70882a53",
          5360 => x"5a5f5256",
          5361 => x"54738416",
          5362 => x"34758516",
          5363 => x"3482bbd4",
          5364 => x"081b8405",
          5365 => x"547382bb",
          5366 => x"dc0c8d3d",
          5367 => x"0d04fe3d",
          5368 => x"0d745282",
          5369 => x"bbd40884",
          5370 => x"38f4dc3f",
          5371 => x"71537180",
          5372 => x"2e8b3871",
          5373 => x"51fced3f",
          5374 => x"82bbdc08",
          5375 => x"537282bb",
          5376 => x"dc0c843d",
          5377 => x"0d04ee3d",
          5378 => x"0d646640",
          5379 => x"5c807042",
          5380 => x"4082bbd4",
          5381 => x"08602e09",
          5382 => x"81068438",
          5383 => x"f4a93f7b",
          5384 => x"8e387e51",
          5385 => x"ffb83f82",
          5386 => x"bbdc0854",
          5387 => x"83c7397e",
          5388 => x"8b387b51",
          5389 => x"fc923f7e",
          5390 => x"5483ba39",
          5391 => x"7e51f58f",
          5392 => x"3f82bbdc",
          5393 => x"0883ffff",
          5394 => x"0682bbd4",
          5395 => x"087d7131",
          5396 => x"832a7083",
          5397 => x"ffff0670",
          5398 => x"832b7311",
          5399 => x"70338112",
          5400 => x"3371882b",
          5401 => x"07707531",
          5402 => x"7083ffff",
          5403 => x"06708829",
          5404 => x"fc057388",
          5405 => x"291a7033",
          5406 => x"81123371",
          5407 => x"882b0770",
          5408 => x"902b5344",
          5409 => x"4e534841",
          5410 => x"525c545b",
          5411 => x"415c565b",
          5412 => x"5b738025",
          5413 => x"8f387681",
          5414 => x"ffff0675",
          5415 => x"317083ff",
          5416 => x"ff064254",
          5417 => x"82163383",
          5418 => x"17337188",
          5419 => x"2b077088",
          5420 => x"291c7033",
          5421 => x"81123371",
          5422 => x"982b7190",
          5423 => x"2b075347",
          5424 => x"45525654",
          5425 => x"7380258b",
          5426 => x"38787531",
          5427 => x"7083ffff",
          5428 => x"06415477",
          5429 => x"7b2781fe",
          5430 => x"38601854",
          5431 => x"737b2e09",
          5432 => x"81068f38",
          5433 => x"7851f6c0",
          5434 => x"3f7a83ff",
          5435 => x"ff065881",
          5436 => x"e5397f8e",
          5437 => x"387a7424",
          5438 => x"89387851",
          5439 => x"f6aa3f81",
          5440 => x"a5397f18",
          5441 => x"557a7524",
          5442 => x"80c83879",
          5443 => x"1d821133",
          5444 => x"83123371",
          5445 => x"882b0753",
          5446 => x"5754f4f4",
          5447 => x"3f805278",
          5448 => x"51f7b73f",
          5449 => x"82bbdc08",
          5450 => x"83ffff06",
          5451 => x"7e547c53",
          5452 => x"70832b82",
          5453 => x"bbd40811",
          5454 => x"84055355",
          5455 => x"59ff8edb",
          5456 => x"3f82bbd4",
          5457 => x"08148405",
          5458 => x"7583ffff",
          5459 => x"06595c81",
          5460 => x"85396015",
          5461 => x"547a7424",
          5462 => x"80d43878",
          5463 => x"51f5c93f",
          5464 => x"82bbd408",
          5465 => x"1d821133",
          5466 => x"83123371",
          5467 => x"882b0753",
          5468 => x"4354f49c",
          5469 => x"3f805278",
          5470 => x"51f6df3f",
          5471 => x"82bbdc08",
          5472 => x"83ffff06",
          5473 => x"7e547c53",
          5474 => x"70832b82",
          5475 => x"bbd40811",
          5476 => x"84055355",
          5477 => x"59ff8e83",
          5478 => x"3f82bbd4",
          5479 => x"08148405",
          5480 => x"60620519",
          5481 => x"555c7383",
          5482 => x"ffff0658",
          5483 => x"a9397b7f",
          5484 => x"5254f9b0",
          5485 => x"3f82bbdc",
          5486 => x"085c82bb",
          5487 => x"dc08802e",
          5488 => x"93387d53",
          5489 => x"735282bb",
          5490 => x"dc0851ff",
          5491 => x"92973f73",
          5492 => x"51f7983f",
          5493 => x"7a587a78",
          5494 => x"27993880",
          5495 => x"537a5278",
          5496 => x"51f28f3f",
          5497 => x"7a19832b",
          5498 => x"82bbd408",
          5499 => x"05840551",
          5500 => x"f6f93f7b",
          5501 => x"547382bb",
          5502 => x"dc0c943d",
          5503 => x"0d04fc3d",
          5504 => x"0d777729",
          5505 => x"705254fb",
          5506 => x"d53f82bb",
          5507 => x"dc085582",
          5508 => x"bbdc0880",
          5509 => x"2e8e3873",
          5510 => x"53805282",
          5511 => x"bbdc0851",
          5512 => x"ff96c33f",
          5513 => x"7482bbdc",
          5514 => x"0c863d0d",
          5515 => x"04ff3d0d",
          5516 => x"028f0533",
          5517 => x"51815270",
          5518 => x"72268738",
          5519 => x"82bbd811",
          5520 => x"33527182",
          5521 => x"bbdc0c83",
          5522 => x"3d0d04fc",
          5523 => x"3d0d029b",
          5524 => x"05330284",
          5525 => x"059f0533",
          5526 => x"56538351",
          5527 => x"72812680",
          5528 => x"e0387284",
          5529 => x"2b87c092",
          5530 => x"8c115351",
          5531 => x"88547480",
          5532 => x"2e843881",
          5533 => x"88547372",
          5534 => x"0c87c092",
          5535 => x"8c115181",
          5536 => x"710c850b",
          5537 => x"87c0988c",
          5538 => x"0c705271",
          5539 => x"08708206",
          5540 => x"51517080",
          5541 => x"2e8a3887",
          5542 => x"c0988c08",
          5543 => x"5170ec38",
          5544 => x"7108fc80",
          5545 => x"80065271",
          5546 => x"923887c0",
          5547 => x"988c0851",
          5548 => x"70802e87",
          5549 => x"387182bb",
          5550 => x"d8143482",
          5551 => x"bbd81333",
          5552 => x"517082bb",
          5553 => x"dc0c863d",
          5554 => x"0d04f33d",
          5555 => x"0d606264",
          5556 => x"028c05bf",
          5557 => x"05335740",
          5558 => x"585b8374",
          5559 => x"525afecd",
          5560 => x"3f82bbdc",
          5561 => x"0881067a",
          5562 => x"54527181",
          5563 => x"be387172",
          5564 => x"75842b87",
          5565 => x"c0928011",
          5566 => x"87c0928c",
          5567 => x"1287c092",
          5568 => x"8413415a",
          5569 => x"40575a58",
          5570 => x"850b87c0",
          5571 => x"988c0c76",
          5572 => x"7d0c8476",
          5573 => x"0c750870",
          5574 => x"852a7081",
          5575 => x"06515354",
          5576 => x"71802e8e",
          5577 => x"387b0852",
          5578 => x"717b7081",
          5579 => x"055d3481",
          5580 => x"19598074",
          5581 => x"a2065353",
          5582 => x"71732e83",
          5583 => x"38815378",
          5584 => x"83ff268f",
          5585 => x"3872802e",
          5586 => x"8a3887c0",
          5587 => x"988c0852",
          5588 => x"71c33887",
          5589 => x"c0988c08",
          5590 => x"5271802e",
          5591 => x"87387884",
          5592 => x"802e9938",
          5593 => x"81760c87",
          5594 => x"c0928c15",
          5595 => x"53720870",
          5596 => x"82065152",
          5597 => x"71f738ff",
          5598 => x"1a5a8d39",
          5599 => x"84801781",
          5600 => x"197081ff",
          5601 => x"065a5357",
          5602 => x"79802e90",
          5603 => x"3873fc80",
          5604 => x"80065271",
          5605 => x"87387d78",
          5606 => x"26feed38",
          5607 => x"73fc8080",
          5608 => x"06527180",
          5609 => x"2e833881",
          5610 => x"52715372",
          5611 => x"82bbdc0c",
          5612 => x"8f3d0d04",
          5613 => x"f33d0d60",
          5614 => x"6264028c",
          5615 => x"05bf0533",
          5616 => x"5740585b",
          5617 => x"83598074",
          5618 => x"5258fce1",
          5619 => x"3f82bbdc",
          5620 => x"08810679",
          5621 => x"54527178",
          5622 => x"2e098106",
          5623 => x"81b13877",
          5624 => x"74842b87",
          5625 => x"c0928011",
          5626 => x"87c0928c",
          5627 => x"1287c092",
          5628 => x"84134059",
          5629 => x"5f565a85",
          5630 => x"0b87c098",
          5631 => x"8c0c767d",
          5632 => x"0c82760c",
          5633 => x"80587508",
          5634 => x"70842a70",
          5635 => x"81065153",
          5636 => x"5471802e",
          5637 => x"8c387a70",
          5638 => x"81055c33",
          5639 => x"7c0c8118",
          5640 => x"5873812a",
          5641 => x"70810651",
          5642 => x"5271802e",
          5643 => x"8a3887c0",
          5644 => x"988c0852",
          5645 => x"71d03887",
          5646 => x"c0988c08",
          5647 => x"5271802e",
          5648 => x"87387784",
          5649 => x"802e9938",
          5650 => x"81760c87",
          5651 => x"c0928c15",
          5652 => x"53720870",
          5653 => x"82065152",
          5654 => x"71f738ff",
          5655 => x"19598d39",
          5656 => x"811a7081",
          5657 => x"ff068480",
          5658 => x"19595b52",
          5659 => x"78802e90",
          5660 => x"3873fc80",
          5661 => x"80065271",
          5662 => x"87387d7a",
          5663 => x"26fef838",
          5664 => x"73fc8080",
          5665 => x"06527180",
          5666 => x"2e833881",
          5667 => x"52715372",
          5668 => x"82bbdc0c",
          5669 => x"8f3d0d04",
          5670 => x"fa3d0d7a",
          5671 => x"028405a3",
          5672 => x"05330288",
          5673 => x"05a70533",
          5674 => x"71545456",
          5675 => x"57fafe3f",
          5676 => x"82bbdc08",
          5677 => x"81065383",
          5678 => x"547280fe",
          5679 => x"38850b87",
          5680 => x"c0988c0c",
          5681 => x"81567176",
          5682 => x"2e80dc38",
          5683 => x"71762493",
          5684 => x"3874842b",
          5685 => x"87c0928c",
          5686 => x"11545471",
          5687 => x"802e8d38",
          5688 => x"80d43971",
          5689 => x"832e80c6",
          5690 => x"3880cb39",
          5691 => x"72087081",
          5692 => x"2a708106",
          5693 => x"51515271",
          5694 => x"802e8a38",
          5695 => x"87c0988c",
          5696 => x"085271e8",
          5697 => x"3887c098",
          5698 => x"8c085271",
          5699 => x"96388173",
          5700 => x"0c87c092",
          5701 => x"8c145372",
          5702 => x"08708206",
          5703 => x"515271f7",
          5704 => x"38963980",
          5705 => x"56923988",
          5706 => x"800a770c",
          5707 => x"85398180",
          5708 => x"770c7256",
          5709 => x"83398456",
          5710 => x"75547382",
          5711 => x"bbdc0c88",
          5712 => x"3d0d04fe",
          5713 => x"3d0d7481",
          5714 => x"11337133",
          5715 => x"71882b07",
          5716 => x"82bbdc0c",
          5717 => x"5351843d",
          5718 => x"0d04fd3d",
          5719 => x"0d758311",
          5720 => x"33821233",
          5721 => x"71902b71",
          5722 => x"882b0781",
          5723 => x"14337072",
          5724 => x"07882b75",
          5725 => x"33710782",
          5726 => x"bbdc0c52",
          5727 => x"53545654",
          5728 => x"52853d0d",
          5729 => x"04ff3d0d",
          5730 => x"73028405",
          5731 => x"92052252",
          5732 => x"52707270",
          5733 => x"81055434",
          5734 => x"70882a51",
          5735 => x"70723483",
          5736 => x"3d0d04ff",
          5737 => x"3d0d7375",
          5738 => x"52527072",
          5739 => x"70810554",
          5740 => x"3470882a",
          5741 => x"51707270",
          5742 => x"81055434",
          5743 => x"70882a51",
          5744 => x"70727081",
          5745 => x"05543470",
          5746 => x"882a5170",
          5747 => x"7234833d",
          5748 => x"0d04fe3d",
          5749 => x"0d767577",
          5750 => x"54545170",
          5751 => x"802e9238",
          5752 => x"71708105",
          5753 => x"53337370",
          5754 => x"81055534",
          5755 => x"ff1151eb",
          5756 => x"39843d0d",
          5757 => x"04fe3d0d",
          5758 => x"75777654",
          5759 => x"52537272",
          5760 => x"70810554",
          5761 => x"34ff1151",
          5762 => x"70f43884",
          5763 => x"3d0d04fc",
          5764 => x"3d0d7877",
          5765 => x"79565653",
          5766 => x"74708105",
          5767 => x"56337470",
          5768 => x"81055633",
          5769 => x"717131ff",
          5770 => x"16565252",
          5771 => x"5272802e",
          5772 => x"86387180",
          5773 => x"2ee23871",
          5774 => x"82bbdc0c",
          5775 => x"863d0d04",
          5776 => x"fe3d0d74",
          5777 => x"76545189",
          5778 => x"3971732e",
          5779 => x"8a388111",
          5780 => x"51703352",
          5781 => x"71f33870",
          5782 => x"3382bbdc",
          5783 => x"0c843d0d",
          5784 => x"04800b82",
          5785 => x"bbdc0c04",
          5786 => x"800b82bb",
          5787 => x"dc0c04f7",
          5788 => x"3d0d7b56",
          5789 => x"800b8317",
          5790 => x"33565a74",
          5791 => x"7a2e80d6",
          5792 => x"388154b0",
          5793 => x"160853b4",
          5794 => x"16705381",
          5795 => x"17335259",
          5796 => x"faa23f82",
          5797 => x"bbdc087a",
          5798 => x"2e098106",
          5799 => x"b73882bb",
          5800 => x"dc088317",
          5801 => x"34b01608",
          5802 => x"70a41808",
          5803 => x"319c1808",
          5804 => x"59565874",
          5805 => x"77279f38",
          5806 => x"82163355",
          5807 => x"74822e09",
          5808 => x"81069338",
          5809 => x"81547618",
          5810 => x"53785281",
          5811 => x"163351f9",
          5812 => x"e33f8339",
          5813 => x"815a7982",
          5814 => x"bbdc0c8b",
          5815 => x"3d0d04fa",
          5816 => x"3d0d787a",
          5817 => x"56568057",
          5818 => x"74b01708",
          5819 => x"2eaf3875",
          5820 => x"51fefc3f",
          5821 => x"82bbdc08",
          5822 => x"5782bbdc",
          5823 => x"089f3881",
          5824 => x"547453b4",
          5825 => x"16528116",
          5826 => x"3351f7be",
          5827 => x"3f82bbdc",
          5828 => x"08802e85",
          5829 => x"38ff5581",
          5830 => x"5774b017",
          5831 => x"0c7682bb",
          5832 => x"dc0c883d",
          5833 => x"0d04f83d",
          5834 => x"0d7a7052",
          5835 => x"57fec03f",
          5836 => x"82bbdc08",
          5837 => x"5882bbdc",
          5838 => x"08819138",
          5839 => x"76335574",
          5840 => x"832e0981",
          5841 => x"0680f038",
          5842 => x"84173359",
          5843 => x"78812e09",
          5844 => x"810680e3",
          5845 => x"38848053",
          5846 => x"82bbdc08",
          5847 => x"52b41770",
          5848 => x"5256fd91",
          5849 => x"3f82d4d5",
          5850 => x"5284b217",
          5851 => x"51fc963f",
          5852 => x"848b85a4",
          5853 => x"d2527551",
          5854 => x"fca93f86",
          5855 => x"8a85e4f2",
          5856 => x"52849817",
          5857 => x"51fc9c3f",
          5858 => x"90170852",
          5859 => x"849c1751",
          5860 => x"fc913f8c",
          5861 => x"17085284",
          5862 => x"a01751fc",
          5863 => x"863fa017",
          5864 => x"08810570",
          5865 => x"b0190c79",
          5866 => x"55537552",
          5867 => x"81173351",
          5868 => x"f8823f77",
          5869 => x"84183480",
          5870 => x"53805281",
          5871 => x"173351f9",
          5872 => x"d73f82bb",
          5873 => x"dc08802e",
          5874 => x"83388158",
          5875 => x"7782bbdc",
          5876 => x"0c8a3d0d",
          5877 => x"04fb3d0d",
          5878 => x"77fe1a98",
          5879 => x"1208fe05",
          5880 => x"55565480",
          5881 => x"56747327",
          5882 => x"8d388a14",
          5883 => x"22757129",
          5884 => x"ac160805",
          5885 => x"57537582",
          5886 => x"bbdc0c87",
          5887 => x"3d0d04f9",
          5888 => x"3d0d7a7a",
          5889 => x"70085654",
          5890 => x"57817727",
          5891 => x"81df3876",
          5892 => x"98150827",
          5893 => x"81d738ff",
          5894 => x"74335458",
          5895 => x"72822e80",
          5896 => x"f5387282",
          5897 => x"24893872",
          5898 => x"812e8d38",
          5899 => x"81bf3972",
          5900 => x"832e818e",
          5901 => x"3881b639",
          5902 => x"76812a17",
          5903 => x"70892aa4",
          5904 => x"16080553",
          5905 => x"745255fd",
          5906 => x"963f82bb",
          5907 => x"dc08819f",
          5908 => x"387483ff",
          5909 => x"0614b411",
          5910 => x"33811770",
          5911 => x"892aa418",
          5912 => x"08055576",
          5913 => x"54575753",
          5914 => x"fcf53f82",
          5915 => x"bbdc0880",
          5916 => x"fe387483",
          5917 => x"ff0614b4",
          5918 => x"11337088",
          5919 => x"2b780779",
          5920 => x"81067184",
          5921 => x"2a5c5258",
          5922 => x"51537280",
          5923 => x"e238759f",
          5924 => x"ff065880",
          5925 => x"da397688",
          5926 => x"2aa41508",
          5927 => x"05527351",
          5928 => x"fcbd3f82",
          5929 => x"bbdc0880",
          5930 => x"c6387610",
          5931 => x"83fe0674",
          5932 => x"05b40551",
          5933 => x"f98d3f82",
          5934 => x"bbdc0883",
          5935 => x"ffff0658",
          5936 => x"ae397687",
          5937 => x"2aa41508",
          5938 => x"05527351",
          5939 => x"fc913f82",
          5940 => x"bbdc089b",
          5941 => x"3876822b",
          5942 => x"83fc0674",
          5943 => x"05b40551",
          5944 => x"f8f83f82",
          5945 => x"bbdc08f0",
          5946 => x"0a065883",
          5947 => x"39815877",
          5948 => x"82bbdc0c",
          5949 => x"893d0d04",
          5950 => x"f83d0d7a",
          5951 => x"7c7e5a58",
          5952 => x"56825981",
          5953 => x"7727829e",
          5954 => x"38769817",
          5955 => x"08278296",
          5956 => x"38753353",
          5957 => x"72792e81",
          5958 => x"9d387279",
          5959 => x"24893872",
          5960 => x"812e8d38",
          5961 => x"82803972",
          5962 => x"832e81b8",
          5963 => x"3881f739",
          5964 => x"76812a17",
          5965 => x"70892aa4",
          5966 => x"18080553",
          5967 => x"765255fb",
          5968 => x"9e3f82bb",
          5969 => x"dc085982",
          5970 => x"bbdc0881",
          5971 => x"d9387483",
          5972 => x"ff0616b4",
          5973 => x"05811678",
          5974 => x"81065956",
          5975 => x"54775376",
          5976 => x"802e8f38",
          5977 => x"77842b9f",
          5978 => x"f0067433",
          5979 => x"8f067107",
          5980 => x"51537274",
          5981 => x"34810b83",
          5982 => x"17347489",
          5983 => x"2aa41708",
          5984 => x"05527551",
          5985 => x"fad93f82",
          5986 => x"bbdc0859",
          5987 => x"82bbdc08",
          5988 => x"81943874",
          5989 => x"83ff0616",
          5990 => x"b4057884",
          5991 => x"2a545476",
          5992 => x"8f387788",
          5993 => x"2a743381",
          5994 => x"f006718f",
          5995 => x"06075153",
          5996 => x"72743480",
          5997 => x"ec397688",
          5998 => x"2aa41708",
          5999 => x"05527551",
          6000 => x"fa9d3f82",
          6001 => x"bbdc0859",
          6002 => x"82bbdc08",
          6003 => x"80d83877",
          6004 => x"83ffff06",
          6005 => x"52761083",
          6006 => x"fe067605",
          6007 => x"b40551f7",
          6008 => x"a43fbe39",
          6009 => x"76872aa4",
          6010 => x"17080552",
          6011 => x"7551f9ef",
          6012 => x"3f82bbdc",
          6013 => x"085982bb",
          6014 => x"dc08ab38",
          6015 => x"77f00a06",
          6016 => x"77822b83",
          6017 => x"fc067018",
          6018 => x"b4057054",
          6019 => x"515454f6",
          6020 => x"c93f82bb",
          6021 => x"dc088f0a",
          6022 => x"06740752",
          6023 => x"7251f783",
          6024 => x"3f810b83",
          6025 => x"17347882",
          6026 => x"bbdc0c8a",
          6027 => x"3d0d04f8",
          6028 => x"3d0d7a7c",
          6029 => x"7e720859",
          6030 => x"56565981",
          6031 => x"7527a438",
          6032 => x"74981708",
          6033 => x"279d3873",
          6034 => x"802eaa38",
          6035 => x"ff537352",
          6036 => x"7551fda4",
          6037 => x"3f82bbdc",
          6038 => x"085482bb",
          6039 => x"dc0880f2",
          6040 => x"38933982",
          6041 => x"5480eb39",
          6042 => x"815480e6",
          6043 => x"3982bbdc",
          6044 => x"085480de",
          6045 => x"39745278",
          6046 => x"51fb843f",
          6047 => x"82bbdc08",
          6048 => x"5882bbdc",
          6049 => x"08802e80",
          6050 => x"c73882bb",
          6051 => x"dc08812e",
          6052 => x"d23882bb",
          6053 => x"dc08ff2e",
          6054 => x"cf388053",
          6055 => x"74527551",
          6056 => x"fcd63f82",
          6057 => x"bbdc08c5",
          6058 => x"38981608",
          6059 => x"fe119018",
          6060 => x"08575557",
          6061 => x"74742790",
          6062 => x"38811590",
          6063 => x"170c8416",
          6064 => x"33810754",
          6065 => x"73841734",
          6066 => x"77557678",
          6067 => x"26ffa638",
          6068 => x"80547382",
          6069 => x"bbdc0c8a",
          6070 => x"3d0d04f6",
          6071 => x"3d0d7c7e",
          6072 => x"7108595b",
          6073 => x"5b799538",
          6074 => x"8c170858",
          6075 => x"77802e88",
          6076 => x"38981708",
          6077 => x"7826b238",
          6078 => x"8158ae39",
          6079 => x"79527a51",
          6080 => x"f9fd3f81",
          6081 => x"557482bb",
          6082 => x"dc082782",
          6083 => x"e03882bb",
          6084 => x"dc085582",
          6085 => x"bbdc08ff",
          6086 => x"2e82d238",
          6087 => x"98170882",
          6088 => x"bbdc0826",
          6089 => x"82c73879",
          6090 => x"58901708",
          6091 => x"70565473",
          6092 => x"802e82b9",
          6093 => x"38777a2e",
          6094 => x"09810680",
          6095 => x"e238811a",
          6096 => x"56981708",
          6097 => x"76268338",
          6098 => x"82567552",
          6099 => x"7a51f9af",
          6100 => x"3f805982",
          6101 => x"bbdc0881",
          6102 => x"2e098106",
          6103 => x"863882bb",
          6104 => x"dc085982",
          6105 => x"bbdc0809",
          6106 => x"70307072",
          6107 => x"07802570",
          6108 => x"7c0782bb",
          6109 => x"dc085451",
          6110 => x"51555573",
          6111 => x"81ef3882",
          6112 => x"bbdc0880",
          6113 => x"2e95388c",
          6114 => x"17085481",
          6115 => x"74279038",
          6116 => x"73981808",
          6117 => x"27893873",
          6118 => x"58853975",
          6119 => x"80db3877",
          6120 => x"56811656",
          6121 => x"98170876",
          6122 => x"26893882",
          6123 => x"56757826",
          6124 => x"81ac3875",
          6125 => x"527a51f8",
          6126 => x"c63f82bb",
          6127 => x"dc08802e",
          6128 => x"b8388059",
          6129 => x"82bbdc08",
          6130 => x"812e0981",
          6131 => x"06863882",
          6132 => x"bbdc0859",
          6133 => x"82bbdc08",
          6134 => x"09703070",
          6135 => x"72078025",
          6136 => x"707c0751",
          6137 => x"51555573",
          6138 => x"80f83875",
          6139 => x"782e0981",
          6140 => x"06ffae38",
          6141 => x"735580f5",
          6142 => x"39ff5375",
          6143 => x"527651f9",
          6144 => x"f73f82bb",
          6145 => x"dc0882bb",
          6146 => x"dc083070",
          6147 => x"82bbdc08",
          6148 => x"07802551",
          6149 => x"55557980",
          6150 => x"2e943873",
          6151 => x"802e8f38",
          6152 => x"75537952",
          6153 => x"7651f9d0",
          6154 => x"3f82bbdc",
          6155 => x"085574a5",
          6156 => x"38758c18",
          6157 => x"0c981708",
          6158 => x"fe059018",
          6159 => x"08565474",
          6160 => x"74268638",
          6161 => x"ff159018",
          6162 => x"0c841733",
          6163 => x"81075473",
          6164 => x"84183497",
          6165 => x"39ff5674",
          6166 => x"812e9038",
          6167 => x"8c398055",
          6168 => x"8c3982bb",
          6169 => x"dc085585",
          6170 => x"39815675",
          6171 => x"557482bb",
          6172 => x"dc0c8c3d",
          6173 => x"0d04f83d",
          6174 => x"0d7a7052",
          6175 => x"55f3f03f",
          6176 => x"82bbdc08",
          6177 => x"58815682",
          6178 => x"bbdc0880",
          6179 => x"d8387b52",
          6180 => x"7451f6c1",
          6181 => x"3f82bbdc",
          6182 => x"0882bbdc",
          6183 => x"08b0170c",
          6184 => x"59848053",
          6185 => x"7752b415",
          6186 => x"705257f2",
          6187 => x"c83f7756",
          6188 => x"84398116",
          6189 => x"568a1522",
          6190 => x"58757827",
          6191 => x"97388154",
          6192 => x"75195376",
          6193 => x"52811533",
          6194 => x"51ede93f",
          6195 => x"82bbdc08",
          6196 => x"802edf38",
          6197 => x"8a152276",
          6198 => x"32703070",
          6199 => x"7207709f",
          6200 => x"2a535156",
          6201 => x"567582bb",
          6202 => x"dc0c8a3d",
          6203 => x"0d04f83d",
          6204 => x"0d7a7c71",
          6205 => x"08585657",
          6206 => x"74f0800a",
          6207 => x"2680f138",
          6208 => x"749f0653",
          6209 => x"7280e938",
          6210 => x"7490180c",
          6211 => x"88170854",
          6212 => x"73aa3875",
          6213 => x"33538273",
          6214 => x"278838a8",
          6215 => x"16085473",
          6216 => x"9b387485",
          6217 => x"2a53820b",
          6218 => x"8817225a",
          6219 => x"58727927",
          6220 => x"80fe38a8",
          6221 => x"16089818",
          6222 => x"0c80cd39",
          6223 => x"8a162270",
          6224 => x"892b5458",
          6225 => x"727526b2",
          6226 => x"38735276",
          6227 => x"51f5b03f",
          6228 => x"82bbdc08",
          6229 => x"5482bbdc",
          6230 => x"08ff2ebd",
          6231 => x"38810b82",
          6232 => x"bbdc0827",
          6233 => x"8b389816",
          6234 => x"0882bbdc",
          6235 => x"08268538",
          6236 => x"8258bd39",
          6237 => x"74733155",
          6238 => x"cb397352",
          6239 => x"7551f4d5",
          6240 => x"3f82bbdc",
          6241 => x"0898180c",
          6242 => x"7394180c",
          6243 => x"98170853",
          6244 => x"82587280",
          6245 => x"2e9a3885",
          6246 => x"39815894",
          6247 => x"3974892a",
          6248 => x"1398180c",
          6249 => x"7483ff06",
          6250 => x"16b4059c",
          6251 => x"180c8058",
          6252 => x"7782bbdc",
          6253 => x"0c8a3d0d",
          6254 => x"04f83d0d",
          6255 => x"7a700890",
          6256 => x"1208a005",
          6257 => x"595754f0",
          6258 => x"800a7727",
          6259 => x"8638800b",
          6260 => x"98150c98",
          6261 => x"14085384",
          6262 => x"5572802e",
          6263 => x"81cb3876",
          6264 => x"83ff0658",
          6265 => x"7781b538",
          6266 => x"81139815",
          6267 => x"0c941408",
          6268 => x"55749238",
          6269 => x"76852a88",
          6270 => x"17225653",
          6271 => x"74732681",
          6272 => x"9b3880c0",
          6273 => x"398a1622",
          6274 => x"ff057789",
          6275 => x"2a065372",
          6276 => x"818a3874",
          6277 => x"527351f3",
          6278 => x"e63f82bb",
          6279 => x"dc085382",
          6280 => x"55810b82",
          6281 => x"bbdc0827",
          6282 => x"80ff3881",
          6283 => x"5582bbdc",
          6284 => x"08ff2e80",
          6285 => x"f4389816",
          6286 => x"0882bbdc",
          6287 => x"082680ca",
          6288 => x"387b8a38",
          6289 => x"7798150c",
          6290 => x"845580dd",
          6291 => x"39941408",
          6292 => x"527351f9",
          6293 => x"863f82bb",
          6294 => x"dc085387",
          6295 => x"5582bbdc",
          6296 => x"08802e80",
          6297 => x"c4388255",
          6298 => x"82bbdc08",
          6299 => x"812eba38",
          6300 => x"815582bb",
          6301 => x"dc08ff2e",
          6302 => x"b03882bb",
          6303 => x"dc085275",
          6304 => x"51fbf33f",
          6305 => x"82bbdc08",
          6306 => x"a0387294",
          6307 => x"150c7252",
          6308 => x"7551f2c1",
          6309 => x"3f82bbdc",
          6310 => x"0898150c",
          6311 => x"7690150c",
          6312 => x"7716b405",
          6313 => x"9c150c80",
          6314 => x"557482bb",
          6315 => x"dc0c8a3d",
          6316 => x"0d04f73d",
          6317 => x"0d7b7d71",
          6318 => x"085b5b57",
          6319 => x"80527651",
          6320 => x"fcac3f82",
          6321 => x"bbdc0854",
          6322 => x"82bbdc08",
          6323 => x"80ec3882",
          6324 => x"bbdc0856",
          6325 => x"98170852",
          6326 => x"7851f083",
          6327 => x"3f82bbdc",
          6328 => x"085482bb",
          6329 => x"dc0880d2",
          6330 => x"3882bbdc",
          6331 => x"089c1808",
          6332 => x"70335154",
          6333 => x"587281e5",
          6334 => x"2e098106",
          6335 => x"83388158",
          6336 => x"82bbdc08",
          6337 => x"55728338",
          6338 => x"81557775",
          6339 => x"07537280",
          6340 => x"2e8e3881",
          6341 => x"1656757a",
          6342 => x"2e098106",
          6343 => x"8838a539",
          6344 => x"82bbdc08",
          6345 => x"56815276",
          6346 => x"51fd8e3f",
          6347 => x"82bbdc08",
          6348 => x"5482bbdc",
          6349 => x"08802eff",
          6350 => x"9b387384",
          6351 => x"2e098106",
          6352 => x"83388754",
          6353 => x"7382bbdc",
          6354 => x"0c8b3d0d",
          6355 => x"04fd3d0d",
          6356 => x"769a1152",
          6357 => x"54ebec3f",
          6358 => x"82bbdc08",
          6359 => x"83ffff06",
          6360 => x"76703351",
          6361 => x"53537183",
          6362 => x"2e098106",
          6363 => x"90389414",
          6364 => x"51ebd03f",
          6365 => x"82bbdc08",
          6366 => x"902b7307",
          6367 => x"537282bb",
          6368 => x"dc0c853d",
          6369 => x"0d04fc3d",
          6370 => x"0d777970",
          6371 => x"83ffff06",
          6372 => x"549a1253",
          6373 => x"5555ebed",
          6374 => x"3f767033",
          6375 => x"51537283",
          6376 => x"2e098106",
          6377 => x"8b387390",
          6378 => x"2a529415",
          6379 => x"51ebd63f",
          6380 => x"863d0d04",
          6381 => x"f73d0d7b",
          6382 => x"7d5b5584",
          6383 => x"75085a58",
          6384 => x"98150880",
          6385 => x"2e818a38",
          6386 => x"98150852",
          6387 => x"7851ee8f",
          6388 => x"3f82bbdc",
          6389 => x"085882bb",
          6390 => x"dc0880f5",
          6391 => x"389c1508",
          6392 => x"70335553",
          6393 => x"73863884",
          6394 => x"5880e639",
          6395 => x"8b133370",
          6396 => x"bf067081",
          6397 => x"ff065851",
          6398 => x"53728616",
          6399 => x"3482bbdc",
          6400 => x"08537381",
          6401 => x"e52e8338",
          6402 => x"815373ae",
          6403 => x"2ea93881",
          6404 => x"70740654",
          6405 => x"5772802e",
          6406 => x"9e38758f",
          6407 => x"2e993882",
          6408 => x"bbdc0876",
          6409 => x"df065454",
          6410 => x"72882e09",
          6411 => x"81068338",
          6412 => x"7654737a",
          6413 => x"2ea03880",
          6414 => x"527451fa",
          6415 => x"fc3f82bb",
          6416 => x"dc085882",
          6417 => x"bbdc0889",
          6418 => x"38981508",
          6419 => x"fefa3886",
          6420 => x"39800b98",
          6421 => x"160c7782",
          6422 => x"bbdc0c8b",
          6423 => x"3d0d04fb",
          6424 => x"3d0d7770",
          6425 => x"08575481",
          6426 => x"527351fc",
          6427 => x"c53f82bb",
          6428 => x"dc085582",
          6429 => x"bbdc08b4",
          6430 => x"38981408",
          6431 => x"527551ec",
          6432 => x"de3f82bb",
          6433 => x"dc085582",
          6434 => x"bbdc08a0",
          6435 => x"38a05382",
          6436 => x"bbdc0852",
          6437 => x"9c140851",
          6438 => x"eadb3f8b",
          6439 => x"53a01452",
          6440 => x"9c140851",
          6441 => x"eaac3f81",
          6442 => x"0b831734",
          6443 => x"7482bbdc",
          6444 => x"0c873d0d",
          6445 => x"04fd3d0d",
          6446 => x"75700898",
          6447 => x"12085470",
          6448 => x"535553ec",
          6449 => x"9a3f82bb",
          6450 => x"dc088d38",
          6451 => x"9c130853",
          6452 => x"e5733481",
          6453 => x"0b831534",
          6454 => x"853d0d04",
          6455 => x"fa3d0d78",
          6456 => x"7a575780",
          6457 => x"0b891734",
          6458 => x"98170880",
          6459 => x"2e818238",
          6460 => x"80708918",
          6461 => x"5555559c",
          6462 => x"17081470",
          6463 => x"33811656",
          6464 => x"515271a0",
          6465 => x"2ea83871",
          6466 => x"852e0981",
          6467 => x"06843881",
          6468 => x"e5527389",
          6469 => x"2e098106",
          6470 => x"8b38ae73",
          6471 => x"70810555",
          6472 => x"34811555",
          6473 => x"71737081",
          6474 => x"05553481",
          6475 => x"15558a74",
          6476 => x"27c53875",
          6477 => x"15880552",
          6478 => x"800b8113",
          6479 => x"349c1708",
          6480 => x"528b1233",
          6481 => x"8817349c",
          6482 => x"17089c11",
          6483 => x"5252e88a",
          6484 => x"3f82bbdc",
          6485 => x"08760c96",
          6486 => x"1251e7e7",
          6487 => x"3f82bbdc",
          6488 => x"08861723",
          6489 => x"981251e7",
          6490 => x"da3f82bb",
          6491 => x"dc088417",
          6492 => x"23883d0d",
          6493 => x"04f33d0d",
          6494 => x"7f70085e",
          6495 => x"5b806170",
          6496 => x"33515555",
          6497 => x"73af2e83",
          6498 => x"38815573",
          6499 => x"80dc2e91",
          6500 => x"3874802e",
          6501 => x"8c38941d",
          6502 => x"08881c0c",
          6503 => x"aa398115",
          6504 => x"41806170",
          6505 => x"33565656",
          6506 => x"73af2e09",
          6507 => x"81068338",
          6508 => x"81567380",
          6509 => x"dc327030",
          6510 => x"70802578",
          6511 => x"07515154",
          6512 => x"73dc3873",
          6513 => x"881c0c60",
          6514 => x"70335154",
          6515 => x"739f2696",
          6516 => x"38ff800b",
          6517 => x"ab1c3480",
          6518 => x"527a51f6",
          6519 => x"913f82bb",
          6520 => x"dc085585",
          6521 => x"9839913d",
          6522 => x"61a01d5c",
          6523 => x"5a5e8b53",
          6524 => x"a0527951",
          6525 => x"e7ff3f80",
          6526 => x"70595788",
          6527 => x"7933555c",
          6528 => x"73ae2e09",
          6529 => x"810680d4",
          6530 => x"38781870",
          6531 => x"33811a71",
          6532 => x"ae327030",
          6533 => x"709f2a73",
          6534 => x"82260751",
          6535 => x"51535a57",
          6536 => x"54738c38",
          6537 => x"79175475",
          6538 => x"74348117",
          6539 => x"57db3975",
          6540 => x"af327030",
          6541 => x"709f2a51",
          6542 => x"51547580",
          6543 => x"dc2e8c38",
          6544 => x"73802e87",
          6545 => x"3875a026",
          6546 => x"82bd3877",
          6547 => x"197e0ca4",
          6548 => x"54a07627",
          6549 => x"82bd38a0",
          6550 => x"5482b839",
          6551 => x"78187033",
          6552 => x"811a5a57",
          6553 => x"54a07627",
          6554 => x"81fc3875",
          6555 => x"af327030",
          6556 => x"7780dc32",
          6557 => x"70307280",
          6558 => x"25718025",
          6559 => x"07515156",
          6560 => x"51557380",
          6561 => x"2eac3884",
          6562 => x"39811858",
          6563 => x"80781a70",
          6564 => x"33515555",
          6565 => x"73af2e09",
          6566 => x"81068338",
          6567 => x"81557380",
          6568 => x"dc327030",
          6569 => x"70802577",
          6570 => x"07515154",
          6571 => x"73db3881",
          6572 => x"b53975ae",
          6573 => x"2e098106",
          6574 => x"83388154",
          6575 => x"767c2774",
          6576 => x"07547380",
          6577 => x"2ea2387b",
          6578 => x"8b327030",
          6579 => x"77ae3270",
          6580 => x"30728025",
          6581 => x"719f2a07",
          6582 => x"53515651",
          6583 => x"557481a7",
          6584 => x"3888578b",
          6585 => x"5cfef539",
          6586 => x"75982b54",
          6587 => x"7380258c",
          6588 => x"387580ff",
          6589 => x"0682b5a4",
          6590 => x"11335754",
          6591 => x"7551e6e1",
          6592 => x"3f82bbdc",
          6593 => x"08802eb2",
          6594 => x"38781870",
          6595 => x"33811a71",
          6596 => x"545a5654",
          6597 => x"e6d23f82",
          6598 => x"bbdc0880",
          6599 => x"2e80e838",
          6600 => x"ff1c5476",
          6601 => x"742780df",
          6602 => x"38791754",
          6603 => x"75743481",
          6604 => x"177a1155",
          6605 => x"57747434",
          6606 => x"a7397552",
          6607 => x"82b4c451",
          6608 => x"e5fe3f82",
          6609 => x"bbdc08bf",
          6610 => x"38ff9f16",
          6611 => x"54739926",
          6612 => x"8938e016",
          6613 => x"7081ff06",
          6614 => x"57547917",
          6615 => x"54757434",
          6616 => x"811757fd",
          6617 => x"f7397719",
          6618 => x"7e0c7680",
          6619 => x"2e993879",
          6620 => x"33547381",
          6621 => x"e52e0981",
          6622 => x"06843885",
          6623 => x"7a348454",
          6624 => x"a076278f",
          6625 => x"388b3986",
          6626 => x"5581f239",
          6627 => x"845680f3",
          6628 => x"39805473",
          6629 => x"8b1b3480",
          6630 => x"7b085852",
          6631 => x"7a51f2ce",
          6632 => x"3f82bbdc",
          6633 => x"085682bb",
          6634 => x"dc0880d7",
          6635 => x"38981b08",
          6636 => x"527651e6",
          6637 => x"aa3f82bb",
          6638 => x"dc085682",
          6639 => x"bbdc0880",
          6640 => x"c2389c1b",
          6641 => x"08703355",
          6642 => x"5573802e",
          6643 => x"ffbe388b",
          6644 => x"1533bf06",
          6645 => x"5473861c",
          6646 => x"348b1533",
          6647 => x"70832a70",
          6648 => x"81065155",
          6649 => x"58739238",
          6650 => x"8b537952",
          6651 => x"7451e49f",
          6652 => x"3f82bbdc",
          6653 => x"08802e8b",
          6654 => x"3875527a",
          6655 => x"51f3ba3f",
          6656 => x"ff9f3975",
          6657 => x"ab1c3357",
          6658 => x"5574802e",
          6659 => x"bb387484",
          6660 => x"2e098106",
          6661 => x"80e73875",
          6662 => x"852a7081",
          6663 => x"0677822a",
          6664 => x"58515473",
          6665 => x"802e9638",
          6666 => x"75810654",
          6667 => x"73802efb",
          6668 => x"b538ff80",
          6669 => x"0bab1c34",
          6670 => x"805580c1",
          6671 => x"39758106",
          6672 => x"5473ba38",
          6673 => x"8555b639",
          6674 => x"75822a70",
          6675 => x"81065154",
          6676 => x"73ab3886",
          6677 => x"1b337084",
          6678 => x"2a708106",
          6679 => x"51555573",
          6680 => x"802ee138",
          6681 => x"901b0883",
          6682 => x"ff061db4",
          6683 => x"05527c51",
          6684 => x"f5db3f82",
          6685 => x"bbdc0888",
          6686 => x"1c0cfaea",
          6687 => x"397482bb",
          6688 => x"dc0c8f3d",
          6689 => x"0d04f63d",
          6690 => x"0d7c5bff",
          6691 => x"7b087071",
          6692 => x"7355595c",
          6693 => x"55597380",
          6694 => x"2e81c638",
          6695 => x"75708105",
          6696 => x"573370a0",
          6697 => x"26525271",
          6698 => x"ba2e8d38",
          6699 => x"70ee3871",
          6700 => x"ba2e0981",
          6701 => x"0681a538",
          6702 => x"7333d011",
          6703 => x"7081ff06",
          6704 => x"51525370",
          6705 => x"89269138",
          6706 => x"82147381",
          6707 => x"ff06d005",
          6708 => x"56527176",
          6709 => x"2e80f738",
          6710 => x"800b82b5",
          6711 => x"94595577",
          6712 => x"087a5557",
          6713 => x"76708105",
          6714 => x"58337470",
          6715 => x"81055633",
          6716 => x"ff9f1253",
          6717 => x"53537099",
          6718 => x"268938e0",
          6719 => x"137081ff",
          6720 => x"065451ff",
          6721 => x"9f125170",
          6722 => x"99268938",
          6723 => x"e0127081",
          6724 => x"ff065351",
          6725 => x"7230709f",
          6726 => x"2a515172",
          6727 => x"722e0981",
          6728 => x"06853870",
          6729 => x"ffbe3872",
          6730 => x"30747732",
          6731 => x"70307072",
          6732 => x"079f2a73",
          6733 => x"9f2a0753",
          6734 => x"54545170",
          6735 => x"802e8f38",
          6736 => x"81158419",
          6737 => x"59558375",
          6738 => x"25ff9438",
          6739 => x"8b397483",
          6740 => x"24863874",
          6741 => x"767c0c59",
          6742 => x"78518639",
          6743 => x"82d3a833",
          6744 => x"517082bb",
          6745 => x"dc0c8c3d",
          6746 => x"0d04fa3d",
          6747 => x"0d785680",
          6748 => x"0b831734",
          6749 => x"ff0bb017",
          6750 => x"0c795275",
          6751 => x"51e2e03f",
          6752 => x"845582bb",
          6753 => x"dc088180",
          6754 => x"3884b216",
          6755 => x"51dfb43f",
          6756 => x"82bbdc08",
          6757 => x"83ffff06",
          6758 => x"54835573",
          6759 => x"82d4d52e",
          6760 => x"09810680",
          6761 => x"e338800b",
          6762 => x"b4173356",
          6763 => x"577481e9",
          6764 => x"2e098106",
          6765 => x"83388157",
          6766 => x"7481eb32",
          6767 => x"70307080",
          6768 => x"25790751",
          6769 => x"5154738a",
          6770 => x"387481e8",
          6771 => x"2e098106",
          6772 => x"b5388353",
          6773 => x"82b4d452",
          6774 => x"80ea1651",
          6775 => x"e0b13f82",
          6776 => x"bbdc0855",
          6777 => x"82bbdc08",
          6778 => x"802e9d38",
          6779 => x"855382b4",
          6780 => x"d8528186",
          6781 => x"1651e097",
          6782 => x"3f82bbdc",
          6783 => x"085582bb",
          6784 => x"dc08802e",
          6785 => x"83388255",
          6786 => x"7482bbdc",
          6787 => x"0c883d0d",
          6788 => x"04f23d0d",
          6789 => x"61028405",
          6790 => x"80cb0533",
          6791 => x"58558075",
          6792 => x"0c6051fc",
          6793 => x"e13f82bb",
          6794 => x"dc08588b",
          6795 => x"56800b82",
          6796 => x"bbdc0824",
          6797 => x"86fc3882",
          6798 => x"bbdc0884",
          6799 => x"2982d394",
          6800 => x"05700855",
          6801 => x"538c5673",
          6802 => x"802e86e6",
          6803 => x"3873750c",
          6804 => x"7681fe06",
          6805 => x"74335457",
          6806 => x"72802eae",
          6807 => x"38811433",
          6808 => x"51d7ca3f",
          6809 => x"82bbdc08",
          6810 => x"81ff0670",
          6811 => x"81065455",
          6812 => x"72983876",
          6813 => x"802e86b8",
          6814 => x"3874822a",
          6815 => x"70810651",
          6816 => x"538a5672",
          6817 => x"86ac3886",
          6818 => x"a7398074",
          6819 => x"34778115",
          6820 => x"34815281",
          6821 => x"143351d7",
          6822 => x"b23f82bb",
          6823 => x"dc0881ff",
          6824 => x"06708106",
          6825 => x"54558356",
          6826 => x"72868738",
          6827 => x"76802e8f",
          6828 => x"3874822a",
          6829 => x"70810651",
          6830 => x"538a5672",
          6831 => x"85f43880",
          6832 => x"70537452",
          6833 => x"5bfda33f",
          6834 => x"82bbdc08",
          6835 => x"81ff0657",
          6836 => x"76822e09",
          6837 => x"810680e2",
          6838 => x"388c3d74",
          6839 => x"56588356",
          6840 => x"83f61533",
          6841 => x"70585372",
          6842 => x"802e8d38",
          6843 => x"83fa1551",
          6844 => x"dce83f82",
          6845 => x"bbdc0857",
          6846 => x"76787084",
          6847 => x"055a0cff",
          6848 => x"16901656",
          6849 => x"56758025",
          6850 => x"d738800b",
          6851 => x"8d3d5456",
          6852 => x"72708405",
          6853 => x"54085b83",
          6854 => x"577a802e",
          6855 => x"95387a52",
          6856 => x"7351fcc6",
          6857 => x"3f82bbdc",
          6858 => x"0881ff06",
          6859 => x"57817727",
          6860 => x"89388116",
          6861 => x"56837627",
          6862 => x"d7388156",
          6863 => x"76842e84",
          6864 => x"f1388d56",
          6865 => x"76812684",
          6866 => x"e938bf14",
          6867 => x"51dbf43f",
          6868 => x"82bbdc08",
          6869 => x"83ffff06",
          6870 => x"53728480",
          6871 => x"2e098106",
          6872 => x"84d03880",
          6873 => x"ca1451db",
          6874 => x"da3f82bb",
          6875 => x"dc0883ff",
          6876 => x"ff065877",
          6877 => x"8d3880d8",
          6878 => x"1451dbde",
          6879 => x"3f82bbdc",
          6880 => x"0858779c",
          6881 => x"150c80c4",
          6882 => x"14338215",
          6883 => x"3480c414",
          6884 => x"33ff1170",
          6885 => x"81ff0651",
          6886 => x"54558d56",
          6887 => x"72812684",
          6888 => x"91387481",
          6889 => x"ff067871",
          6890 => x"2980c116",
          6891 => x"33525953",
          6892 => x"728a1523",
          6893 => x"72802e8b",
          6894 => x"38ff1373",
          6895 => x"06537280",
          6896 => x"2e86388d",
          6897 => x"5683eb39",
          6898 => x"80c51451",
          6899 => x"daf53f82",
          6900 => x"bbdc0853",
          6901 => x"82bbdc08",
          6902 => x"88152372",
          6903 => x"8f06578d",
          6904 => x"567683ce",
          6905 => x"3880c714",
          6906 => x"51dad83f",
          6907 => x"82bbdc08",
          6908 => x"83ffff06",
          6909 => x"55748d38",
          6910 => x"80d41451",
          6911 => x"dadc3f82",
          6912 => x"bbdc0855",
          6913 => x"80c21451",
          6914 => x"dab93f82",
          6915 => x"bbdc0883",
          6916 => x"ffff0653",
          6917 => x"8d567280",
          6918 => x"2e839738",
          6919 => x"88142278",
          6920 => x"1471842a",
          6921 => x"055a5a78",
          6922 => x"75268386",
          6923 => x"388a1422",
          6924 => x"52747931",
          6925 => x"51feeecb",
          6926 => x"3f82bbdc",
          6927 => x"085582bb",
          6928 => x"dc08802e",
          6929 => x"82ec3882",
          6930 => x"bbdc0880",
          6931 => x"fffffff5",
          6932 => x"26833883",
          6933 => x"577483ff",
          6934 => x"f5268338",
          6935 => x"8257749f",
          6936 => x"f5268538",
          6937 => x"81578939",
          6938 => x"8d567680",
          6939 => x"2e82c338",
          6940 => x"82157098",
          6941 => x"160c7ba0",
          6942 => x"160c731c",
          6943 => x"70a4170c",
          6944 => x"7a1dac17",
          6945 => x"0c545576",
          6946 => x"832e0981",
          6947 => x"06af3880",
          6948 => x"de1451d9",
          6949 => x"ae3f82bb",
          6950 => x"dc0883ff",
          6951 => x"ff06538d",
          6952 => x"5672828e",
          6953 => x"3879828a",
          6954 => x"3880e014",
          6955 => x"51d9ab3f",
          6956 => x"82bbdc08",
          6957 => x"a8150c74",
          6958 => x"822b53a2",
          6959 => x"398d5679",
          6960 => x"802e81ee",
          6961 => x"387713a8",
          6962 => x"150c7415",
          6963 => x"5376822e",
          6964 => x"8d387410",
          6965 => x"1570812a",
          6966 => x"76810605",
          6967 => x"515383ff",
          6968 => x"13892a53",
          6969 => x"8d56729c",
          6970 => x"15082681",
          6971 => x"c538ff0b",
          6972 => x"90150cff",
          6973 => x"0b8c150c",
          6974 => x"ff800b84",
          6975 => x"15347683",
          6976 => x"2e098106",
          6977 => x"81923880",
          6978 => x"e41451d8",
          6979 => x"b63f82bb",
          6980 => x"dc0883ff",
          6981 => x"ff065372",
          6982 => x"812e0981",
          6983 => x"0680f938",
          6984 => x"811b5273",
          6985 => x"51dbb83f",
          6986 => x"82bbdc08",
          6987 => x"80ea3882",
          6988 => x"bbdc0884",
          6989 => x"153484b2",
          6990 => x"1451d887",
          6991 => x"3f82bbdc",
          6992 => x"0883ffff",
          6993 => x"06537282",
          6994 => x"d4d52e09",
          6995 => x"810680c8",
          6996 => x"38b41451",
          6997 => x"d8843f82",
          6998 => x"bbdc0884",
          6999 => x"8b85a4d2",
          7000 => x"2e098106",
          7001 => x"b3388498",
          7002 => x"1451d7ee",
          7003 => x"3f82bbdc",
          7004 => x"08868a85",
          7005 => x"e4f22e09",
          7006 => x"81069d38",
          7007 => x"849c1451",
          7008 => x"d7d83f82",
          7009 => x"bbdc0890",
          7010 => x"150c84a0",
          7011 => x"1451d7ca",
          7012 => x"3f82bbdc",
          7013 => x"088c150c",
          7014 => x"76743482",
          7015 => x"d3a42281",
          7016 => x"05537282",
          7017 => x"d3a42372",
          7018 => x"86152380",
          7019 => x"0b94150c",
          7020 => x"80567582",
          7021 => x"bbdc0c90",
          7022 => x"3d0d04fb",
          7023 => x"3d0d7754",
          7024 => x"89557380",
          7025 => x"2eb93873",
          7026 => x"08537280",
          7027 => x"2eb13872",
          7028 => x"33527180",
          7029 => x"2ea93886",
          7030 => x"13228415",
          7031 => x"22575271",
          7032 => x"762e0981",
          7033 => x"06993881",
          7034 => x"133351d0",
          7035 => x"c03f82bb",
          7036 => x"dc088106",
          7037 => x"52718838",
          7038 => x"71740854",
          7039 => x"55833980",
          7040 => x"53787371",
          7041 => x"0c527482",
          7042 => x"bbdc0c87",
          7043 => x"3d0d04fa",
          7044 => x"3d0d02ab",
          7045 => x"05337a58",
          7046 => x"893dfc05",
          7047 => x"5256f4e6",
          7048 => x"3f8b5480",
          7049 => x"0b82bbdc",
          7050 => x"0824bc38",
          7051 => x"82bbdc08",
          7052 => x"842982d3",
          7053 => x"94057008",
          7054 => x"55557380",
          7055 => x"2e843880",
          7056 => x"74347854",
          7057 => x"73802e84",
          7058 => x"38807434",
          7059 => x"78750c75",
          7060 => x"5475802e",
          7061 => x"92388053",
          7062 => x"893d7053",
          7063 => x"840551f7",
          7064 => x"b03f82bb",
          7065 => x"dc085473",
          7066 => x"82bbdc0c",
          7067 => x"883d0d04",
          7068 => x"eb3d0d67",
          7069 => x"02840580",
          7070 => x"e7053359",
          7071 => x"59895478",
          7072 => x"802e84c8",
          7073 => x"3877bf06",
          7074 => x"7054983d",
          7075 => x"d0055399",
          7076 => x"3d840552",
          7077 => x"58f6fa3f",
          7078 => x"82bbdc08",
          7079 => x"5582bbdc",
          7080 => x"0884a438",
          7081 => x"7a5c6852",
          7082 => x"8c3d7052",
          7083 => x"56edc63f",
          7084 => x"82bbdc08",
          7085 => x"5582bbdc",
          7086 => x"08923802",
          7087 => x"80d70533",
          7088 => x"70982b55",
          7089 => x"57738025",
          7090 => x"83388655",
          7091 => x"779c0654",
          7092 => x"73802e81",
          7093 => x"ab387480",
          7094 => x"2e953874",
          7095 => x"842e0981",
          7096 => x"06aa3875",
          7097 => x"51eaf83f",
          7098 => x"82bbdc08",
          7099 => x"559e3902",
          7100 => x"b2053391",
          7101 => x"06547381",
          7102 => x"b8387782",
          7103 => x"2a708106",
          7104 => x"51547380",
          7105 => x"2e8e3888",
          7106 => x"5583bc39",
          7107 => x"77880758",
          7108 => x"7483b438",
          7109 => x"77832a70",
          7110 => x"81065154",
          7111 => x"73802e81",
          7112 => x"af386252",
          7113 => x"7a51e8a5",
          7114 => x"3f82bbdc",
          7115 => x"08568288",
          7116 => x"b20a5262",
          7117 => x"8e0551d4",
          7118 => x"ea3f6254",
          7119 => x"a00b8b15",
          7120 => x"34805362",
          7121 => x"527a51e8",
          7122 => x"bd3f8052",
          7123 => x"629c0551",
          7124 => x"d4d13f7a",
          7125 => x"54810b83",
          7126 => x"15347580",
          7127 => x"2e80f138",
          7128 => x"7ab01108",
          7129 => x"51548053",
          7130 => x"7552973d",
          7131 => x"d40551dd",
          7132 => x"be3f82bb",
          7133 => x"dc085582",
          7134 => x"bbdc0882",
          7135 => x"ca38b739",
          7136 => x"7482c438",
          7137 => x"02b20533",
          7138 => x"70842a70",
          7139 => x"81065155",
          7140 => x"5673802e",
          7141 => x"86388455",
          7142 => x"82ad3977",
          7143 => x"812a7081",
          7144 => x"06515473",
          7145 => x"802ea938",
          7146 => x"75810654",
          7147 => x"73802ea0",
          7148 => x"38875582",
          7149 => x"92397352",
          7150 => x"7a51d6a3",
          7151 => x"3f82bbdc",
          7152 => x"087bff18",
          7153 => x"8c120c55",
          7154 => x"5582bbdc",
          7155 => x"0881f838",
          7156 => x"77832a70",
          7157 => x"81065154",
          7158 => x"73802e86",
          7159 => x"387780c0",
          7160 => x"07587ab0",
          7161 => x"1108a01b",
          7162 => x"0c63a41b",
          7163 => x"0c635370",
          7164 => x"5257e6d9",
          7165 => x"3f82bbdc",
          7166 => x"0882bbdc",
          7167 => x"08881b0c",
          7168 => x"639c0552",
          7169 => x"5ad2d33f",
          7170 => x"82bbdc08",
          7171 => x"82bbdc08",
          7172 => x"8c1b0c77",
          7173 => x"7a0c5686",
          7174 => x"1722841a",
          7175 => x"2377901a",
          7176 => x"34800b91",
          7177 => x"1a34800b",
          7178 => x"9c1a0c80",
          7179 => x"0b941a0c",
          7180 => x"77852a70",
          7181 => x"81065154",
          7182 => x"73802e81",
          7183 => x"8d3882bb",
          7184 => x"dc08802e",
          7185 => x"81843882",
          7186 => x"bbdc0894",
          7187 => x"1a0c8a17",
          7188 => x"2270892b",
          7189 => x"7b525957",
          7190 => x"a8397652",
          7191 => x"7851d79f",
          7192 => x"3f82bbdc",
          7193 => x"085782bb",
          7194 => x"dc088126",
          7195 => x"83388255",
          7196 => x"82bbdc08",
          7197 => x"ff2e0981",
          7198 => x"06833879",
          7199 => x"55757831",
          7200 => x"56743070",
          7201 => x"76078025",
          7202 => x"51547776",
          7203 => x"278a3881",
          7204 => x"70750655",
          7205 => x"5a73c338",
          7206 => x"76981a0c",
          7207 => x"74a93875",
          7208 => x"83ff0654",
          7209 => x"73802ea2",
          7210 => x"3876527a",
          7211 => x"51d6a63f",
          7212 => x"82bbdc08",
          7213 => x"85388255",
          7214 => x"8e397589",
          7215 => x"2a82bbdc",
          7216 => x"08059c1a",
          7217 => x"0c843980",
          7218 => x"790c7454",
          7219 => x"7382bbdc",
          7220 => x"0c973d0d",
          7221 => x"04f23d0d",
          7222 => x"60636564",
          7223 => x"40405d59",
          7224 => x"807e0c90",
          7225 => x"3dfc0552",
          7226 => x"7851f9cf",
          7227 => x"3f82bbdc",
          7228 => x"085582bb",
          7229 => x"dc088a38",
          7230 => x"91193355",
          7231 => x"74802e86",
          7232 => x"38745682",
          7233 => x"c4399019",
          7234 => x"33810655",
          7235 => x"87567480",
          7236 => x"2e82b638",
          7237 => x"9539820b",
          7238 => x"911a3482",
          7239 => x"5682aa39",
          7240 => x"810b911a",
          7241 => x"34815682",
          7242 => x"a0398c19",
          7243 => x"08941a08",
          7244 => x"3155747c",
          7245 => x"27833874",
          7246 => x"5c7b802e",
          7247 => x"82893894",
          7248 => x"19087083",
          7249 => x"ff065656",
          7250 => x"7481b238",
          7251 => x"7e8a1122",
          7252 => x"ff057789",
          7253 => x"2a065b55",
          7254 => x"79a83875",
          7255 => x"87388819",
          7256 => x"08558f39",
          7257 => x"98190852",
          7258 => x"7851d593",
          7259 => x"3f82bbdc",
          7260 => x"08558175",
          7261 => x"27ff9f38",
          7262 => x"74ff2eff",
          7263 => x"a3387498",
          7264 => x"1a0c9819",
          7265 => x"08527e51",
          7266 => x"d4cb3f82",
          7267 => x"bbdc0880",
          7268 => x"2eff8338",
          7269 => x"82bbdc08",
          7270 => x"1a7c892a",
          7271 => x"59577780",
          7272 => x"2e80d638",
          7273 => x"771a7f8a",
          7274 => x"1122585c",
          7275 => x"55757527",
          7276 => x"8538757a",
          7277 => x"31587754",
          7278 => x"76537c52",
          7279 => x"811b3351",
          7280 => x"ca883f82",
          7281 => x"bbdc08fe",
          7282 => x"d7387e83",
          7283 => x"11335656",
          7284 => x"74802e9f",
          7285 => x"38b01608",
          7286 => x"77315574",
          7287 => x"78279438",
          7288 => x"848053b4",
          7289 => x"1652b016",
          7290 => x"08773189",
          7291 => x"2b7d0551",
          7292 => x"cfe03f77",
          7293 => x"892b56b9",
          7294 => x"39769c1a",
          7295 => x"0c941908",
          7296 => x"83ff0684",
          7297 => x"80713157",
          7298 => x"557b7627",
          7299 => x"83387b56",
          7300 => x"9c190852",
          7301 => x"7e51d1c7",
          7302 => x"3f82bbdc",
          7303 => x"08fe8138",
          7304 => x"75539419",
          7305 => x"0883ff06",
          7306 => x"1fb40552",
          7307 => x"7c51cfa2",
          7308 => x"3f7b7631",
          7309 => x"7e08177f",
          7310 => x"0c761e94",
          7311 => x"1b081894",
          7312 => x"1c0c5e5c",
          7313 => x"fdf33980",
          7314 => x"567582bb",
          7315 => x"dc0c903d",
          7316 => x"0d04f23d",
          7317 => x"0d606365",
          7318 => x"6440405d",
          7319 => x"58807e0c",
          7320 => x"903dfc05",
          7321 => x"527751f6",
          7322 => x"d23f82bb",
          7323 => x"dc085582",
          7324 => x"bbdc088a",
          7325 => x"38911833",
          7326 => x"5574802e",
          7327 => x"86387456",
          7328 => x"83b83990",
          7329 => x"18337081",
          7330 => x"2a708106",
          7331 => x"51565687",
          7332 => x"5674802e",
          7333 => x"83a43895",
          7334 => x"39820b91",
          7335 => x"19348256",
          7336 => x"83983981",
          7337 => x"0b911934",
          7338 => x"8156838e",
          7339 => x"39941808",
          7340 => x"7c115656",
          7341 => x"74762784",
          7342 => x"3875095c",
          7343 => x"7b802e82",
          7344 => x"ec389418",
          7345 => x"087083ff",
          7346 => x"06565674",
          7347 => x"81fd387e",
          7348 => x"8a1122ff",
          7349 => x"0577892a",
          7350 => x"065c557a",
          7351 => x"bf38758c",
          7352 => x"38881808",
          7353 => x"55749c38",
          7354 => x"7a528539",
          7355 => x"98180852",
          7356 => x"7751d7e7",
          7357 => x"3f82bbdc",
          7358 => x"085582bb",
          7359 => x"dc08802e",
          7360 => x"82ab3874",
          7361 => x"812eff91",
          7362 => x"3874ff2e",
          7363 => x"ff953874",
          7364 => x"98190c88",
          7365 => x"18088538",
          7366 => x"7488190c",
          7367 => x"7e55b015",
          7368 => x"089c1908",
          7369 => x"2e098106",
          7370 => x"8d387451",
          7371 => x"cec13f82",
          7372 => x"bbdc08fe",
          7373 => x"ee389818",
          7374 => x"08527e51",
          7375 => x"d1973f82",
          7376 => x"bbdc0880",
          7377 => x"2efed238",
          7378 => x"82bbdc08",
          7379 => x"1b7c892a",
          7380 => x"5a577880",
          7381 => x"2e80d538",
          7382 => x"781b7f8a",
          7383 => x"1122585b",
          7384 => x"55757527",
          7385 => x"8538757b",
          7386 => x"31597854",
          7387 => x"76537c52",
          7388 => x"811a3351",
          7389 => x"c8be3f82",
          7390 => x"bbdc08fe",
          7391 => x"a6387eb0",
          7392 => x"11087831",
          7393 => x"56567479",
          7394 => x"279b3884",
          7395 => x"8053b016",
          7396 => x"08773189",
          7397 => x"2b7d0552",
          7398 => x"b41651cc",
          7399 => x"b53f7e55",
          7400 => x"800b8316",
          7401 => x"3478892b",
          7402 => x"5680db39",
          7403 => x"8c180894",
          7404 => x"19082693",
          7405 => x"387e51cd",
          7406 => x"b63f82bb",
          7407 => x"dc08fde3",
          7408 => x"387e77b0",
          7409 => x"120c5576",
          7410 => x"9c190c94",
          7411 => x"180883ff",
          7412 => x"06848071",
          7413 => x"3157557b",
          7414 => x"76278338",
          7415 => x"7b569c18",
          7416 => x"08527e51",
          7417 => x"cdf93f82",
          7418 => x"bbdc08fd",
          7419 => x"b6387553",
          7420 => x"7c529418",
          7421 => x"0883ff06",
          7422 => x"1fb40551",
          7423 => x"cbd43f7e",
          7424 => x"55810b83",
          7425 => x"16347b76",
          7426 => x"317e0817",
          7427 => x"7f0c761e",
          7428 => x"941a0818",
          7429 => x"70941c0c",
          7430 => x"8c1b0858",
          7431 => x"585e5c74",
          7432 => x"76278338",
          7433 => x"7555748c",
          7434 => x"190cfd90",
          7435 => x"39901833",
          7436 => x"80c00755",
          7437 => x"74901934",
          7438 => x"80567582",
          7439 => x"bbdc0c90",
          7440 => x"3d0d04f8",
          7441 => x"3d0d7a8b",
          7442 => x"3dfc0553",
          7443 => x"705256f2",
          7444 => x"ea3f82bb",
          7445 => x"dc085782",
          7446 => x"bbdc0880",
          7447 => x"fb389016",
          7448 => x"3370862a",
          7449 => x"70810651",
          7450 => x"55557380",
          7451 => x"2e80e938",
          7452 => x"a0160852",
          7453 => x"7851cce7",
          7454 => x"3f82bbdc",
          7455 => x"085782bb",
          7456 => x"dc0880d4",
          7457 => x"38a41608",
          7458 => x"8b1133a0",
          7459 => x"07555573",
          7460 => x"8b163488",
          7461 => x"16085374",
          7462 => x"52750851",
          7463 => x"dde83f8c",
          7464 => x"1608529c",
          7465 => x"1551c9fb",
          7466 => x"3f8288b2",
          7467 => x"0a529615",
          7468 => x"51c9f03f",
          7469 => x"76529215",
          7470 => x"51c9ca3f",
          7471 => x"7854810b",
          7472 => x"83153478",
          7473 => x"51ccdf3f",
          7474 => x"82bbdc08",
          7475 => x"90173381",
          7476 => x"bf065557",
          7477 => x"73901734",
          7478 => x"7682bbdc",
          7479 => x"0c8a3d0d",
          7480 => x"04fc3d0d",
          7481 => x"76705254",
          7482 => x"fed93f82",
          7483 => x"bbdc0853",
          7484 => x"82bbdc08",
          7485 => x"9c38863d",
          7486 => x"fc055273",
          7487 => x"51f1bc3f",
          7488 => x"82bbdc08",
          7489 => x"5382bbdc",
          7490 => x"08873882",
          7491 => x"bbdc0874",
          7492 => x"0c7282bb",
          7493 => x"dc0c863d",
          7494 => x"0d04ff3d",
          7495 => x"0d843d51",
          7496 => x"e6e43f8b",
          7497 => x"52800b82",
          7498 => x"bbdc0824",
          7499 => x"8b3882bb",
          7500 => x"dc0882d3",
          7501 => x"a8348052",
          7502 => x"7182bbdc",
          7503 => x"0c833d0d",
          7504 => x"04ef3d0d",
          7505 => x"8053933d",
          7506 => x"d0055294",
          7507 => x"3d51e9c1",
          7508 => x"3f82bbdc",
          7509 => x"085582bb",
          7510 => x"dc0880e0",
          7511 => x"38765863",
          7512 => x"52933dd4",
          7513 => x"0551e08d",
          7514 => x"3f82bbdc",
          7515 => x"085582bb",
          7516 => x"dc08bc38",
          7517 => x"0280c705",
          7518 => x"3370982b",
          7519 => x"55567380",
          7520 => x"25893876",
          7521 => x"7a94120c",
          7522 => x"54b23902",
          7523 => x"a2053370",
          7524 => x"842a7081",
          7525 => x"06515556",
          7526 => x"73802e9e",
          7527 => x"38767f53",
          7528 => x"705254db",
          7529 => x"a83f82bb",
          7530 => x"dc089415",
          7531 => x"0c8e3982",
          7532 => x"bbdc0884",
          7533 => x"2e098106",
          7534 => x"83388555",
          7535 => x"7482bbdc",
          7536 => x"0c933d0d",
          7537 => x"04e43d0d",
          7538 => x"6f6f5b5b",
          7539 => x"807a3480",
          7540 => x"539e3dff",
          7541 => x"b805529f",
          7542 => x"3d51e8b5",
          7543 => x"3f82bbdc",
          7544 => x"085782bb",
          7545 => x"dc0882fc",
          7546 => x"387b437a",
          7547 => x"7c941108",
          7548 => x"47555864",
          7549 => x"5473802e",
          7550 => x"81ed38a0",
          7551 => x"52933d70",
          7552 => x"5255d5ea",
          7553 => x"3f82bbdc",
          7554 => x"085782bb",
          7555 => x"dc0882d4",
          7556 => x"3868527b",
          7557 => x"51c9c83f",
          7558 => x"82bbdc08",
          7559 => x"5782bbdc",
          7560 => x"0882c138",
          7561 => x"69527b51",
          7562 => x"daa33f82",
          7563 => x"bbdc0845",
          7564 => x"76527451",
          7565 => x"d5b83f82",
          7566 => x"bbdc0857",
          7567 => x"82bbdc08",
          7568 => x"82a23880",
          7569 => x"527451da",
          7570 => x"eb3f82bb",
          7571 => x"dc085782",
          7572 => x"bbdc08a4",
          7573 => x"3869527b",
          7574 => x"51d9f23f",
          7575 => x"7382bbdc",
          7576 => x"082ea638",
          7577 => x"76527451",
          7578 => x"d6cf3f82",
          7579 => x"bbdc0857",
          7580 => x"82bbdc08",
          7581 => x"802ecc38",
          7582 => x"76842e09",
          7583 => x"81068638",
          7584 => x"825781e0",
          7585 => x"397681dc",
          7586 => x"389e3dff",
          7587 => x"bc055274",
          7588 => x"51dcc93f",
          7589 => x"76903d78",
          7590 => x"11811133",
          7591 => x"51565a56",
          7592 => x"73802e91",
          7593 => x"3802b905",
          7594 => x"55811681",
          7595 => x"16703356",
          7596 => x"565673f5",
          7597 => x"38811654",
          7598 => x"73782681",
          7599 => x"90387580",
          7600 => x"2e993878",
          7601 => x"16810555",
          7602 => x"ff186f11",
          7603 => x"ff18ff18",
          7604 => x"58585558",
          7605 => x"74337434",
          7606 => x"75ee38ff",
          7607 => x"186f1155",
          7608 => x"58af7434",
          7609 => x"fe8d3977",
          7610 => x"7b2e0981",
          7611 => x"068a38ff",
          7612 => x"186f1155",
          7613 => x"58af7434",
          7614 => x"800b82d3",
          7615 => x"a8337084",
          7616 => x"2982b594",
          7617 => x"05700870",
          7618 => x"33525c56",
          7619 => x"56567376",
          7620 => x"2e8d3881",
          7621 => x"16701a70",
          7622 => x"33515556",
          7623 => x"73f53882",
          7624 => x"16547378",
          7625 => x"26a73880",
          7626 => x"55747627",
          7627 => x"91387419",
          7628 => x"5473337a",
          7629 => x"7081055c",
          7630 => x"34811555",
          7631 => x"ec39ba7a",
          7632 => x"7081055c",
          7633 => x"3474ff2e",
          7634 => x"09810685",
          7635 => x"38915794",
          7636 => x"396e1881",
          7637 => x"19595473",
          7638 => x"337a7081",
          7639 => x"055c347a",
          7640 => x"7826ee38",
          7641 => x"807a3476",
          7642 => x"82bbdc0c",
          7643 => x"9e3d0d04",
          7644 => x"f73d0d7b",
          7645 => x"7d8d3dfc",
          7646 => x"05547153",
          7647 => x"5755ecbb",
          7648 => x"3f82bbdc",
          7649 => x"085382bb",
          7650 => x"dc0882fa",
          7651 => x"38911533",
          7652 => x"537282f2",
          7653 => x"388c1508",
          7654 => x"54737627",
          7655 => x"92389015",
          7656 => x"3370812a",
          7657 => x"70810651",
          7658 => x"54577283",
          7659 => x"38735694",
          7660 => x"15085480",
          7661 => x"7094170c",
          7662 => x"5875782e",
          7663 => x"82973879",
          7664 => x"8a112270",
          7665 => x"892b5951",
          7666 => x"5373782e",
          7667 => x"b7387652",
          7668 => x"ff1651fe",
          7669 => x"d7ad3f82",
          7670 => x"bbdc08ff",
          7671 => x"15785470",
          7672 => x"535553fe",
          7673 => x"d79d3f82",
          7674 => x"bbdc0873",
          7675 => x"26963876",
          7676 => x"30707506",
          7677 => x"7094180c",
          7678 => x"77713198",
          7679 => x"18085758",
          7680 => x"5153b139",
          7681 => x"88150854",
          7682 => x"73a63873",
          7683 => x"527451cd",
          7684 => x"ca3f82bb",
          7685 => x"dc085482",
          7686 => x"bbdc0881",
          7687 => x"2e819a38",
          7688 => x"82bbdc08",
          7689 => x"ff2e819b",
          7690 => x"3882bbdc",
          7691 => x"0888160c",
          7692 => x"7398160c",
          7693 => x"73802e81",
          7694 => x"9c387676",
          7695 => x"2780dc38",
          7696 => x"75773194",
          7697 => x"16081894",
          7698 => x"170c9016",
          7699 => x"3370812a",
          7700 => x"70810651",
          7701 => x"555a5672",
          7702 => x"802e9a38",
          7703 => x"73527451",
          7704 => x"ccf93f82",
          7705 => x"bbdc0854",
          7706 => x"82bbdc08",
          7707 => x"943882bb",
          7708 => x"dc0856a7",
          7709 => x"39735274",
          7710 => x"51c7843f",
          7711 => x"82bbdc08",
          7712 => x"5473ff2e",
          7713 => x"be388174",
          7714 => x"27af3879",
          7715 => x"53739814",
          7716 => x"0827a638",
          7717 => x"7398160c",
          7718 => x"ffa03994",
          7719 => x"15081694",
          7720 => x"160c7583",
          7721 => x"ff065372",
          7722 => x"802eaa38",
          7723 => x"73527951",
          7724 => x"c6a33f82",
          7725 => x"bbdc0894",
          7726 => x"38820b91",
          7727 => x"16348253",
          7728 => x"80c43981",
          7729 => x"0b911634",
          7730 => x"8153bb39",
          7731 => x"75892a82",
          7732 => x"bbdc0805",
          7733 => x"58941508",
          7734 => x"548c1508",
          7735 => x"74279038",
          7736 => x"738c160c",
          7737 => x"90153380",
          7738 => x"c0075372",
          7739 => x"90163473",
          7740 => x"83ff0653",
          7741 => x"72802e8c",
          7742 => x"38779c16",
          7743 => x"082e8538",
          7744 => x"779c160c",
          7745 => x"80537282",
          7746 => x"bbdc0c8b",
          7747 => x"3d0d04f9",
          7748 => x"3d0d7956",
          7749 => x"89547580",
          7750 => x"2e818a38",
          7751 => x"8053893d",
          7752 => x"fc05528a",
          7753 => x"3d840551",
          7754 => x"e1e73f82",
          7755 => x"bbdc0855",
          7756 => x"82bbdc08",
          7757 => x"80ea3877",
          7758 => x"760c7a52",
          7759 => x"7551d8b5",
          7760 => x"3f82bbdc",
          7761 => x"085582bb",
          7762 => x"dc0880c3",
          7763 => x"38ab1633",
          7764 => x"70982b55",
          7765 => x"57807424",
          7766 => x"a2388616",
          7767 => x"3370842a",
          7768 => x"70810651",
          7769 => x"55577380",
          7770 => x"2ead389c",
          7771 => x"16085277",
          7772 => x"51d3da3f",
          7773 => x"82bbdc08",
          7774 => x"88170c77",
          7775 => x"54861422",
          7776 => x"84172374",
          7777 => x"527551ce",
          7778 => x"e53f82bb",
          7779 => x"dc085574",
          7780 => x"842e0981",
          7781 => x"06853885",
          7782 => x"55863974",
          7783 => x"802e8438",
          7784 => x"80760c74",
          7785 => x"547382bb",
          7786 => x"dc0c893d",
          7787 => x"0d04fc3d",
          7788 => x"0d76873d",
          7789 => x"fc055370",
          7790 => x"5253e7ff",
          7791 => x"3f82bbdc",
          7792 => x"08873882",
          7793 => x"bbdc0873",
          7794 => x"0c863d0d",
          7795 => x"04fb3d0d",
          7796 => x"7779893d",
          7797 => x"fc055471",
          7798 => x"535654e7",
          7799 => x"de3f82bb",
          7800 => x"dc085382",
          7801 => x"bbdc0880",
          7802 => x"df387493",
          7803 => x"3882bbdc",
          7804 => x"08527351",
          7805 => x"cdf83f82",
          7806 => x"bbdc0853",
          7807 => x"80ca3982",
          7808 => x"bbdc0852",
          7809 => x"7351d3ac",
          7810 => x"3f82bbdc",
          7811 => x"085382bb",
          7812 => x"dc08842e",
          7813 => x"09810685",
          7814 => x"38805387",
          7815 => x"3982bbdc",
          7816 => x"08a63874",
          7817 => x"527351d5",
          7818 => x"b33f7252",
          7819 => x"7351cf89",
          7820 => x"3f82bbdc",
          7821 => x"08843270",
          7822 => x"30707207",
          7823 => x"9f2c7082",
          7824 => x"bbdc0806",
          7825 => x"51515454",
          7826 => x"7282bbdc",
          7827 => x"0c873d0d",
          7828 => x"04ee3d0d",
          7829 => x"65578053",
          7830 => x"893d7053",
          7831 => x"963d5256",
          7832 => x"dfaf3f82",
          7833 => x"bbdc0855",
          7834 => x"82bbdc08",
          7835 => x"b2386452",
          7836 => x"7551d681",
          7837 => x"3f82bbdc",
          7838 => x"085582bb",
          7839 => x"dc08a038",
          7840 => x"0280cb05",
          7841 => x"3370982b",
          7842 => x"55587380",
          7843 => x"25853886",
          7844 => x"558d3976",
          7845 => x"802e8838",
          7846 => x"76527551",
          7847 => x"d4be3f74",
          7848 => x"82bbdc0c",
          7849 => x"943d0d04",
          7850 => x"f03d0d63",
          7851 => x"65555c80",
          7852 => x"53923dec",
          7853 => x"0552933d",
          7854 => x"51ded63f",
          7855 => x"82bbdc08",
          7856 => x"5b82bbdc",
          7857 => x"08828038",
          7858 => x"7c740c73",
          7859 => x"08981108",
          7860 => x"fe119013",
          7861 => x"08595658",
          7862 => x"55757426",
          7863 => x"9138757c",
          7864 => x"0c81e439",
          7865 => x"815b81cc",
          7866 => x"39825b81",
          7867 => x"c73982bb",
          7868 => x"dc087533",
          7869 => x"55597381",
          7870 => x"2e098106",
          7871 => x"bf388275",
          7872 => x"5f577652",
          7873 => x"923df005",
          7874 => x"51c1f43f",
          7875 => x"82bbdc08",
          7876 => x"ff2ed138",
          7877 => x"82bbdc08",
          7878 => x"812ece38",
          7879 => x"82bbdc08",
          7880 => x"307082bb",
          7881 => x"dc080780",
          7882 => x"257a0581",
          7883 => x"197f5359",
          7884 => x"5a549814",
          7885 => x"087726ca",
          7886 => x"3880f939",
          7887 => x"a4150882",
          7888 => x"bbdc0857",
          7889 => x"58759838",
          7890 => x"77528118",
          7891 => x"7d5258ff",
          7892 => x"bf8d3f82",
          7893 => x"bbdc085b",
          7894 => x"82bbdc08",
          7895 => x"80d6387c",
          7896 => x"70337712",
          7897 => x"ff1a5d52",
          7898 => x"56547482",
          7899 => x"2e098106",
          7900 => x"9e38b414",
          7901 => x"51ffbbcb",
          7902 => x"3f82bbdc",
          7903 => x"0883ffff",
          7904 => x"06703070",
          7905 => x"80251b82",
          7906 => x"19595b51",
          7907 => x"549b39b4",
          7908 => x"1451ffbb",
          7909 => x"c53f82bb",
          7910 => x"dc08f00a",
          7911 => x"06703070",
          7912 => x"80251b84",
          7913 => x"19595b51",
          7914 => x"547583ff",
          7915 => x"067a5856",
          7916 => x"79ff9238",
          7917 => x"787c0c7c",
          7918 => x"7990120c",
          7919 => x"84113381",
          7920 => x"07565474",
          7921 => x"8415347a",
          7922 => x"82bbdc0c",
          7923 => x"923d0d04",
          7924 => x"f93d0d79",
          7925 => x"8a3dfc05",
          7926 => x"53705257",
          7927 => x"e3dd3f82",
          7928 => x"bbdc0856",
          7929 => x"82bbdc08",
          7930 => x"81a83891",
          7931 => x"17335675",
          7932 => x"81a03890",
          7933 => x"17337081",
          7934 => x"2a708106",
          7935 => x"51555587",
          7936 => x"5573802e",
          7937 => x"818e3894",
          7938 => x"17085473",
          7939 => x"8c180827",
          7940 => x"81803873",
          7941 => x"9b3882bb",
          7942 => x"dc085388",
          7943 => x"17085276",
          7944 => x"51c48c3f",
          7945 => x"82bbdc08",
          7946 => x"7488190c",
          7947 => x"5680c939",
          7948 => x"98170852",
          7949 => x"7651ffbf",
          7950 => x"c63f82bb",
          7951 => x"dc08ff2e",
          7952 => x"09810683",
          7953 => x"38815682",
          7954 => x"bbdc0881",
          7955 => x"2e098106",
          7956 => x"85388256",
          7957 => x"a33975a0",
          7958 => x"38775482",
          7959 => x"bbdc0898",
          7960 => x"15082794",
          7961 => x"38981708",
          7962 => x"5382bbdc",
          7963 => x"08527651",
          7964 => x"c3bd3f82",
          7965 => x"bbdc0856",
          7966 => x"9417088c",
          7967 => x"180c9017",
          7968 => x"3380c007",
          7969 => x"54739018",
          7970 => x"3475802e",
          7971 => x"85387591",
          7972 => x"18347555",
          7973 => x"7482bbdc",
          7974 => x"0c893d0d",
          7975 => x"04e23d0d",
          7976 => x"8253a03d",
          7977 => x"ffa40552",
          7978 => x"a13d51da",
          7979 => x"e43f82bb",
          7980 => x"dc085582",
          7981 => x"bbdc0881",
          7982 => x"f5387845",
          7983 => x"a13d0852",
          7984 => x"953d7052",
          7985 => x"58d1ae3f",
          7986 => x"82bbdc08",
          7987 => x"5582bbdc",
          7988 => x"0881db38",
          7989 => x"0280fb05",
          7990 => x"3370852a",
          7991 => x"70810651",
          7992 => x"55568655",
          7993 => x"7381c738",
          7994 => x"75982b54",
          7995 => x"80742481",
          7996 => x"bd380280",
          7997 => x"d6053370",
          7998 => x"81065854",
          7999 => x"87557681",
          8000 => x"ad386b52",
          8001 => x"7851ccc5",
          8002 => x"3f82bbdc",
          8003 => x"0874842a",
          8004 => x"70810651",
          8005 => x"55567380",
          8006 => x"2e80d438",
          8007 => x"785482bb",
          8008 => x"dc089415",
          8009 => x"082e8186",
          8010 => x"38735a82",
          8011 => x"bbdc085c",
          8012 => x"76528a3d",
          8013 => x"705254c7",
          8014 => x"b53f82bb",
          8015 => x"dc085582",
          8016 => x"bbdc0880",
          8017 => x"e93882bb",
          8018 => x"dc085273",
          8019 => x"51cce53f",
          8020 => x"82bbdc08",
          8021 => x"5582bbdc",
          8022 => x"08863887",
          8023 => x"5580cf39",
          8024 => x"82bbdc08",
          8025 => x"842e8838",
          8026 => x"82bbdc08",
          8027 => x"80c03877",
          8028 => x"51cec23f",
          8029 => x"82bbdc08",
          8030 => x"82bbdc08",
          8031 => x"307082bb",
          8032 => x"dc080780",
          8033 => x"25515555",
          8034 => x"75802e94",
          8035 => x"3873802e",
          8036 => x"8f388053",
          8037 => x"75527751",
          8038 => x"c1953f82",
          8039 => x"bbdc0855",
          8040 => x"748c3878",
          8041 => x"51ffbafe",
          8042 => x"3f82bbdc",
          8043 => x"08557482",
          8044 => x"bbdc0ca0",
          8045 => x"3d0d04e9",
          8046 => x"3d0d8253",
          8047 => x"993dc005",
          8048 => x"529a3d51",
          8049 => x"d8cb3f82",
          8050 => x"bbdc0854",
          8051 => x"82bbdc08",
          8052 => x"82b03878",
          8053 => x"5e69528e",
          8054 => x"3d705258",
          8055 => x"cf973f82",
          8056 => x"bbdc0854",
          8057 => x"82bbdc08",
          8058 => x"86388854",
          8059 => x"82943982",
          8060 => x"bbdc0884",
          8061 => x"2e098106",
          8062 => x"82883802",
          8063 => x"80df0533",
          8064 => x"70852a81",
          8065 => x"06515586",
          8066 => x"547481f6",
          8067 => x"38785a74",
          8068 => x"528a3d70",
          8069 => x"5257c1c3",
          8070 => x"3f82bbdc",
          8071 => x"08755556",
          8072 => x"82bbdc08",
          8073 => x"83388754",
          8074 => x"82bbdc08",
          8075 => x"812e0981",
          8076 => x"06833882",
          8077 => x"5482bbdc",
          8078 => x"08ff2e09",
          8079 => x"81068638",
          8080 => x"815481b4",
          8081 => x"397381b0",
          8082 => x"3882bbdc",
          8083 => x"08527851",
          8084 => x"c4a43f82",
          8085 => x"bbdc0854",
          8086 => x"82bbdc08",
          8087 => x"819a388b",
          8088 => x"53a052b4",
          8089 => x"1951ffb7",
          8090 => x"8c3f7854",
          8091 => x"ae0bb415",
          8092 => x"34785490",
          8093 => x"0bbf1534",
          8094 => x"8288b20a",
          8095 => x"5280ca19",
          8096 => x"51ffb69f",
          8097 => x"3f755378",
          8098 => x"b4115351",
          8099 => x"c9f83fa0",
          8100 => x"5378b411",
          8101 => x"5380d405",
          8102 => x"51ffb6b6",
          8103 => x"3f7854ae",
          8104 => x"0b80d515",
          8105 => x"347f5378",
          8106 => x"80d41153",
          8107 => x"51c9d73f",
          8108 => x"7854810b",
          8109 => x"83153477",
          8110 => x"51cba43f",
          8111 => x"82bbdc08",
          8112 => x"5482bbdc",
          8113 => x"08b23882",
          8114 => x"88b20a52",
          8115 => x"64960551",
          8116 => x"ffb5d03f",
          8117 => x"75536452",
          8118 => x"7851c9aa",
          8119 => x"3f645490",
          8120 => x"0b8b1534",
          8121 => x"7854810b",
          8122 => x"83153478",
          8123 => x"51ffb8b6",
          8124 => x"3f82bbdc",
          8125 => x"08548b39",
          8126 => x"80537552",
          8127 => x"7651ffbe",
          8128 => x"ae3f7382",
          8129 => x"bbdc0c99",
          8130 => x"3d0d04da",
          8131 => x"3d0da93d",
          8132 => x"840551d2",
          8133 => x"f13f8253",
          8134 => x"a83dff84",
          8135 => x"0552a93d",
          8136 => x"51d5ee3f",
          8137 => x"82bbdc08",
          8138 => x"5582bbdc",
          8139 => x"0882d338",
          8140 => x"784da93d",
          8141 => x"08529d3d",
          8142 => x"705258cc",
          8143 => x"b83f82bb",
          8144 => x"dc085582",
          8145 => x"bbdc0882",
          8146 => x"b9380281",
          8147 => x"9b053381",
          8148 => x"a0065486",
          8149 => x"557382aa",
          8150 => x"38a053a4",
          8151 => x"3d0852a8",
          8152 => x"3dff8805",
          8153 => x"51ffb4ea",
          8154 => x"3fac5377",
          8155 => x"52923d70",
          8156 => x"5254ffb4",
          8157 => x"dd3faa3d",
          8158 => x"08527351",
          8159 => x"cbf73f82",
          8160 => x"bbdc0855",
          8161 => x"82bbdc08",
          8162 => x"9538636f",
          8163 => x"2e098106",
          8164 => x"883865a2",
          8165 => x"3d082e92",
          8166 => x"38885581",
          8167 => x"e53982bb",
          8168 => x"dc08842e",
          8169 => x"09810681",
          8170 => x"b8387351",
          8171 => x"c9b13f82",
          8172 => x"bbdc0855",
          8173 => x"82bbdc08",
          8174 => x"81c83868",
          8175 => x"569353a8",
          8176 => x"3dff9505",
          8177 => x"528d1651",
          8178 => x"ffb4873f",
          8179 => x"02af0533",
          8180 => x"8b17348b",
          8181 => x"16337084",
          8182 => x"2a708106",
          8183 => x"51555573",
          8184 => x"893874a0",
          8185 => x"0754738b",
          8186 => x"17347854",
          8187 => x"810b8315",
          8188 => x"348b1633",
          8189 => x"70842a70",
          8190 => x"81065155",
          8191 => x"5573802e",
          8192 => x"80e5386e",
          8193 => x"642e80df",
          8194 => x"38755278",
          8195 => x"51c6be3f",
          8196 => x"82bbdc08",
          8197 => x"527851ff",
          8198 => x"b7bb3f82",
          8199 => x"5582bbdc",
          8200 => x"08802e80",
          8201 => x"dd3882bb",
          8202 => x"dc085278",
          8203 => x"51ffb5af",
          8204 => x"3f82bbdc",
          8205 => x"087980d4",
          8206 => x"11585855",
          8207 => x"82bbdc08",
          8208 => x"80c03881",
          8209 => x"16335473",
          8210 => x"ae2e0981",
          8211 => x"06993863",
          8212 => x"53755276",
          8213 => x"51c6af3f",
          8214 => x"7854810b",
          8215 => x"83153487",
          8216 => x"3982bbdc",
          8217 => x"089c3877",
          8218 => x"51c8ca3f",
          8219 => x"82bbdc08",
          8220 => x"5582bbdc",
          8221 => x"088c3878",
          8222 => x"51ffb5aa",
          8223 => x"3f82bbdc",
          8224 => x"08557482",
          8225 => x"bbdc0ca8",
          8226 => x"3d0d04ed",
          8227 => x"3d0d0280",
          8228 => x"db053302",
          8229 => x"840580df",
          8230 => x"05335757",
          8231 => x"8253953d",
          8232 => x"d0055296",
          8233 => x"3d51d2e9",
          8234 => x"3f82bbdc",
          8235 => x"085582bb",
          8236 => x"dc0880cf",
          8237 => x"38785a65",
          8238 => x"52953dd4",
          8239 => x"0551c9b5",
          8240 => x"3f82bbdc",
          8241 => x"085582bb",
          8242 => x"dc08b838",
          8243 => x"0280cf05",
          8244 => x"3381a006",
          8245 => x"54865573",
          8246 => x"aa3875a7",
          8247 => x"06617109",
          8248 => x"8b123371",
          8249 => x"067a7406",
          8250 => x"07515755",
          8251 => x"56748b15",
          8252 => x"34785481",
          8253 => x"0b831534",
          8254 => x"7851ffb4",
          8255 => x"a93f82bb",
          8256 => x"dc085574",
          8257 => x"82bbdc0c",
          8258 => x"953d0d04",
          8259 => x"ef3d0d64",
          8260 => x"56825393",
          8261 => x"3dd00552",
          8262 => x"943d51d1",
          8263 => x"f43f82bb",
          8264 => x"dc085582",
          8265 => x"bbdc0880",
          8266 => x"cb387658",
          8267 => x"6352933d",
          8268 => x"d40551c8",
          8269 => x"c03f82bb",
          8270 => x"dc085582",
          8271 => x"bbdc08b4",
          8272 => x"380280c7",
          8273 => x"053381a0",
          8274 => x"06548655",
          8275 => x"73a63884",
          8276 => x"16228617",
          8277 => x"2271902b",
          8278 => x"07535496",
          8279 => x"1f51ffb0",
          8280 => x"c23f7654",
          8281 => x"810b8315",
          8282 => x"347651ff",
          8283 => x"b3b83f82",
          8284 => x"bbdc0855",
          8285 => x"7482bbdc",
          8286 => x"0c933d0d",
          8287 => x"04ea3d0d",
          8288 => x"696b5c5a",
          8289 => x"8053983d",
          8290 => x"d0055299",
          8291 => x"3d51d181",
          8292 => x"3f82bbdc",
          8293 => x"0882bbdc",
          8294 => x"08307082",
          8295 => x"bbdc0807",
          8296 => x"80255155",
          8297 => x"5779802e",
          8298 => x"81853881",
          8299 => x"70750655",
          8300 => x"5573802e",
          8301 => x"80f9387b",
          8302 => x"5d805f80",
          8303 => x"528d3d70",
          8304 => x"5254ffbe",
          8305 => x"a93f82bb",
          8306 => x"dc085782",
          8307 => x"bbdc0880",
          8308 => x"d1387452",
          8309 => x"7351c3dc",
          8310 => x"3f82bbdc",
          8311 => x"085782bb",
          8312 => x"dc08bf38",
          8313 => x"82bbdc08",
          8314 => x"82bbdc08",
          8315 => x"655b5956",
          8316 => x"78188119",
          8317 => x"7b185659",
          8318 => x"55743374",
          8319 => x"34811656",
          8320 => x"8a7827ec",
          8321 => x"388b5675",
          8322 => x"1a548074",
          8323 => x"3475802e",
          8324 => x"9e38ff16",
          8325 => x"701b7033",
          8326 => x"51555673",
          8327 => x"a02ee838",
          8328 => x"8e397684",
          8329 => x"2e098106",
          8330 => x"8638807a",
          8331 => x"34805776",
          8332 => x"30707807",
          8333 => x"80255154",
          8334 => x"7a802e80",
          8335 => x"c1387380",
          8336 => x"2ebc387b",
          8337 => x"a0110853",
          8338 => x"51ffb193",
          8339 => x"3f82bbdc",
          8340 => x"085782bb",
          8341 => x"dc08a738",
          8342 => x"7b703355",
          8343 => x"5580c356",
          8344 => x"73832e8b",
          8345 => x"3880e456",
          8346 => x"73842e83",
          8347 => x"38a75675",
          8348 => x"15b40551",
          8349 => x"ffade33f",
          8350 => x"82bbdc08",
          8351 => x"7b0c7682",
          8352 => x"bbdc0c98",
          8353 => x"3d0d04e6",
          8354 => x"3d0d8253",
          8355 => x"9c3dffb8",
          8356 => x"05529d3d",
          8357 => x"51cefa3f",
          8358 => x"82bbdc08",
          8359 => x"82bbdc08",
          8360 => x"565482bb",
          8361 => x"dc088398",
          8362 => x"388b53a0",
          8363 => x"528b3d70",
          8364 => x"5259ffae",
          8365 => x"c03f736d",
          8366 => x"70337081",
          8367 => x"ff065257",
          8368 => x"55579f74",
          8369 => x"2781bc38",
          8370 => x"78587481",
          8371 => x"ff066d81",
          8372 => x"054e7052",
          8373 => x"55ffaf89",
          8374 => x"3f82bbdc",
          8375 => x"08802ea5",
          8376 => x"386c7033",
          8377 => x"70535754",
          8378 => x"ffaefd3f",
          8379 => x"82bbdc08",
          8380 => x"802e8d38",
          8381 => x"74882b76",
          8382 => x"076d8105",
          8383 => x"4e558639",
          8384 => x"82bbdc08",
          8385 => x"55ff9f15",
          8386 => x"7083ffff",
          8387 => x"06515473",
          8388 => x"99268a38",
          8389 => x"e0157083",
          8390 => x"ffff0656",
          8391 => x"5480ff75",
          8392 => x"27873882",
          8393 => x"b4a41533",
          8394 => x"5574802e",
          8395 => x"a3387452",
          8396 => x"82b6a451",
          8397 => x"ffae893f",
          8398 => x"82bbdc08",
          8399 => x"933881ff",
          8400 => x"75278838",
          8401 => x"76892688",
          8402 => x"388b398a",
          8403 => x"77278638",
          8404 => x"865581ec",
          8405 => x"3981ff75",
          8406 => x"278f3874",
          8407 => x"882a5473",
          8408 => x"78708105",
          8409 => x"5a348117",
          8410 => x"57747870",
          8411 => x"81055a34",
          8412 => x"81176d70",
          8413 => x"337081ff",
          8414 => x"06525755",
          8415 => x"57739f26",
          8416 => x"fec8388b",
          8417 => x"3d335486",
          8418 => x"557381e5",
          8419 => x"2e81b138",
          8420 => x"76802e99",
          8421 => x"3802a705",
          8422 => x"55761570",
          8423 => x"33515473",
          8424 => x"a02e0981",
          8425 => x"068738ff",
          8426 => x"175776ed",
          8427 => x"38794180",
          8428 => x"43805291",
          8429 => x"3d705255",
          8430 => x"ffbab33f",
          8431 => x"82bbdc08",
          8432 => x"5482bbdc",
          8433 => x"0880f738",
          8434 => x"81527451",
          8435 => x"ffbfe53f",
          8436 => x"82bbdc08",
          8437 => x"5482bbdc",
          8438 => x"088d3876",
          8439 => x"80c43867",
          8440 => x"54e57434",
          8441 => x"80c63982",
          8442 => x"bbdc0884",
          8443 => x"2e098106",
          8444 => x"80cc3880",
          8445 => x"5476742e",
          8446 => x"80c43881",
          8447 => x"527451ff",
          8448 => x"bdb03f82",
          8449 => x"bbdc0854",
          8450 => x"82bbdc08",
          8451 => x"b138a053",
          8452 => x"82bbdc08",
          8453 => x"526751ff",
          8454 => x"abdb3f67",
          8455 => x"54880b8b",
          8456 => x"15348b53",
          8457 => x"78526751",
          8458 => x"ffaba73f",
          8459 => x"7954810b",
          8460 => x"83153479",
          8461 => x"51ffadee",
          8462 => x"3f82bbdc",
          8463 => x"08547355",
          8464 => x"7482bbdc",
          8465 => x"0c9c3d0d",
          8466 => x"04f23d0d",
          8467 => x"60620288",
          8468 => x"0580cb05",
          8469 => x"33933dfc",
          8470 => x"05557254",
          8471 => x"405e5ad2",
          8472 => x"da3f82bb",
          8473 => x"dc085882",
          8474 => x"bbdc0882",
          8475 => x"bd38911a",
          8476 => x"33587782",
          8477 => x"b5387c80",
          8478 => x"2e97388c",
          8479 => x"1a085978",
          8480 => x"9038901a",
          8481 => x"3370812a",
          8482 => x"70810651",
          8483 => x"55557390",
          8484 => x"38875482",
          8485 => x"97398258",
          8486 => x"82903981",
          8487 => x"58828b39",
          8488 => x"7e8a1122",
          8489 => x"70892b70",
          8490 => x"557f5456",
          8491 => x"5656febd",
          8492 => x"d23fff14",
          8493 => x"7d067030",
          8494 => x"7072079f",
          8495 => x"2a82bbdc",
          8496 => x"08058c19",
          8497 => x"087c405a",
          8498 => x"5d555581",
          8499 => x"77278838",
          8500 => x"98160877",
          8501 => x"26833882",
          8502 => x"57767756",
          8503 => x"59805674",
          8504 => x"527951ff",
          8505 => x"ae993f81",
          8506 => x"157f5555",
          8507 => x"98140875",
          8508 => x"26833882",
          8509 => x"5582bbdc",
          8510 => x"08812eff",
          8511 => x"993882bb",
          8512 => x"dc08ff2e",
          8513 => x"ff953882",
          8514 => x"bbdc088e",
          8515 => x"38811656",
          8516 => x"757b2e09",
          8517 => x"81068738",
          8518 => x"93397459",
          8519 => x"80567477",
          8520 => x"2e098106",
          8521 => x"ffb93887",
          8522 => x"5880ff39",
          8523 => x"7d802eba",
          8524 => x"38787b55",
          8525 => x"557a802e",
          8526 => x"b4388115",
          8527 => x"5673812e",
          8528 => x"09810683",
          8529 => x"38ff5675",
          8530 => x"5374527e",
          8531 => x"51ffafa8",
          8532 => x"3f82bbdc",
          8533 => x"085882bb",
          8534 => x"dc0880ce",
          8535 => x"38748116",
          8536 => x"ff165656",
          8537 => x"5c73d338",
          8538 => x"8439ff19",
          8539 => x"5c7e7c8c",
          8540 => x"120c557d",
          8541 => x"802eb338",
          8542 => x"78881b0c",
          8543 => x"7c8c1b0c",
          8544 => x"901a3380",
          8545 => x"c0075473",
          8546 => x"901b3498",
          8547 => x"1508fe05",
          8548 => x"90160857",
          8549 => x"54757426",
          8550 => x"9138757b",
          8551 => x"3190160c",
          8552 => x"84153381",
          8553 => x"07547384",
          8554 => x"16347754",
          8555 => x"7382bbdc",
          8556 => x"0c903d0d",
          8557 => x"04e93d0d",
          8558 => x"6b6d0288",
          8559 => x"0580eb05",
          8560 => x"339d3d54",
          8561 => x"5a5c59c5",
          8562 => x"bd3f8b56",
          8563 => x"800b82bb",
          8564 => x"dc08248b",
          8565 => x"f83882bb",
          8566 => x"dc088429",
          8567 => x"82d39405",
          8568 => x"70085155",
          8569 => x"74802e84",
          8570 => x"38807534",
          8571 => x"82bbdc08",
          8572 => x"81ff065f",
          8573 => x"81527e51",
          8574 => x"ffa0d03f",
          8575 => x"82bbdc08",
          8576 => x"81ff0670",
          8577 => x"81065657",
          8578 => x"8356748b",
          8579 => x"c0387682",
          8580 => x"2a708106",
          8581 => x"51558a56",
          8582 => x"748bb238",
          8583 => x"993dfc05",
          8584 => x"5383527e",
          8585 => x"51ffa4f0",
          8586 => x"3f82bbdc",
          8587 => x"08993867",
          8588 => x"5574802e",
          8589 => x"92387482",
          8590 => x"8080268b",
          8591 => x"38ff1575",
          8592 => x"06557480",
          8593 => x"2e833881",
          8594 => x"4878802e",
          8595 => x"87388480",
          8596 => x"79269238",
          8597 => x"7881800a",
          8598 => x"268b38ff",
          8599 => x"19790655",
          8600 => x"74802e86",
          8601 => x"3893568a",
          8602 => x"e4397889",
          8603 => x"2a6e892a",
          8604 => x"70892b77",
          8605 => x"59484359",
          8606 => x"7a833881",
          8607 => x"56613070",
          8608 => x"80257707",
          8609 => x"51559156",
          8610 => x"748ac238",
          8611 => x"993df805",
          8612 => x"5381527e",
          8613 => x"51ffa480",
          8614 => x"3f815682",
          8615 => x"bbdc088a",
          8616 => x"ac387783",
          8617 => x"2a707706",
          8618 => x"82bbdc08",
          8619 => x"43564574",
          8620 => x"8338bf41",
          8621 => x"66558e56",
          8622 => x"6075268a",
          8623 => x"90387461",
          8624 => x"31704855",
          8625 => x"80ff7527",
          8626 => x"8a833893",
          8627 => x"56788180",
          8628 => x"2689fa38",
          8629 => x"77812a70",
          8630 => x"81065643",
          8631 => x"74802e95",
          8632 => x"38778706",
          8633 => x"5574822e",
          8634 => x"838d3877",
          8635 => x"81065574",
          8636 => x"802e8383",
          8637 => x"38778106",
          8638 => x"55935682",
          8639 => x"5e74802e",
          8640 => x"89cb3878",
          8641 => x"5a7d832e",
          8642 => x"09810680",
          8643 => x"e13878ae",
          8644 => x"3866912a",
          8645 => x"57810b82",
          8646 => x"b6c82256",
          8647 => x"5a74802e",
          8648 => x"9d387477",
          8649 => x"26983882",
          8650 => x"b6c85679",
          8651 => x"10821770",
          8652 => x"2257575a",
          8653 => x"74802e86",
          8654 => x"38767527",
          8655 => x"ee387952",
          8656 => x"6651feb8",
          8657 => x"be3f82bb",
          8658 => x"dc088429",
          8659 => x"84870570",
          8660 => x"892a5e55",
          8661 => x"a05c800b",
          8662 => x"82bbdc08",
          8663 => x"fc808a05",
          8664 => x"5644fdff",
          8665 => x"f00a7527",
          8666 => x"80ec3888",
          8667 => x"d33978ae",
          8668 => x"38668c2a",
          8669 => x"57810b82",
          8670 => x"b6b82256",
          8671 => x"5a74802e",
          8672 => x"9d387477",
          8673 => x"26983882",
          8674 => x"b6b85679",
          8675 => x"10821770",
          8676 => x"2257575a",
          8677 => x"74802e86",
          8678 => x"38767527",
          8679 => x"ee387952",
          8680 => x"6651feb7",
          8681 => x"de3f82bb",
          8682 => x"dc081084",
          8683 => x"055782bb",
          8684 => x"dc089ff5",
          8685 => x"26963881",
          8686 => x"0b82bbdc",
          8687 => x"081082bb",
          8688 => x"dc080571",
          8689 => x"11722a83",
          8690 => x"0559565e",
          8691 => x"83ff1789",
          8692 => x"2a5d815c",
          8693 => x"a044601c",
          8694 => x"7d116505",
          8695 => x"697012ff",
          8696 => x"05713070",
          8697 => x"72067431",
          8698 => x"5c525957",
          8699 => x"59407d83",
          8700 => x"2e098106",
          8701 => x"8938761c",
          8702 => x"6018415c",
          8703 => x"8439761d",
          8704 => x"5d799029",
          8705 => x"18706231",
          8706 => x"68585155",
          8707 => x"74762687",
          8708 => x"af38757c",
          8709 => x"317d317a",
          8710 => x"53706531",
          8711 => x"5255feb6",
          8712 => x"e23f82bb",
          8713 => x"dc08587d",
          8714 => x"832e0981",
          8715 => x"069b3882",
          8716 => x"bbdc0883",
          8717 => x"fff52680",
          8718 => x"dd387887",
          8719 => x"83387981",
          8720 => x"2a5978fd",
          8721 => x"be3886f8",
          8722 => x"397d822e",
          8723 => x"09810680",
          8724 => x"c53883ff",
          8725 => x"f50b82bb",
          8726 => x"dc0827a0",
          8727 => x"38788f38",
          8728 => x"791a5574",
          8729 => x"80c02686",
          8730 => x"387459fd",
          8731 => x"96396281",
          8732 => x"06557480",
          8733 => x"2e8f3883",
          8734 => x"5efd8839",
          8735 => x"82bbdc08",
          8736 => x"9ff52692",
          8737 => x"387886b8",
          8738 => x"38791a59",
          8739 => x"81807927",
          8740 => x"fcf13886",
          8741 => x"ab398055",
          8742 => x"7d812e09",
          8743 => x"81068338",
          8744 => x"7d559ff5",
          8745 => x"78278b38",
          8746 => x"74810655",
          8747 => x"8e567486",
          8748 => x"9c388480",
          8749 => x"5380527a",
          8750 => x"51ffa2b9",
          8751 => x"3f8b5382",
          8752 => x"b4e0527a",
          8753 => x"51ffa28a",
          8754 => x"3f848052",
          8755 => x"8b1b51ff",
          8756 => x"a1b33f79",
          8757 => x"8d1c347b",
          8758 => x"83ffff06",
          8759 => x"528e1b51",
          8760 => x"ffa1a23f",
          8761 => x"810b901c",
          8762 => x"347d8332",
          8763 => x"70307096",
          8764 => x"2a848006",
          8765 => x"54515591",
          8766 => x"1b51ffa1",
          8767 => x"883f6655",
          8768 => x"7483ffff",
          8769 => x"26903874",
          8770 => x"83ffff06",
          8771 => x"52931b51",
          8772 => x"ffa0f23f",
          8773 => x"8a397452",
          8774 => x"a01b51ff",
          8775 => x"a1853ff8",
          8776 => x"0b951c34",
          8777 => x"bf52981b",
          8778 => x"51ffa0d9",
          8779 => x"3f81ff52",
          8780 => x"9a1b51ff",
          8781 => x"a0cf3f60",
          8782 => x"529c1b51",
          8783 => x"ffa0e43f",
          8784 => x"7d832e09",
          8785 => x"810680cb",
          8786 => x"388288b2",
          8787 => x"0a5280c3",
          8788 => x"1b51ffa0",
          8789 => x"ce3f7c52",
          8790 => x"a41b51ff",
          8791 => x"a0c53f82",
          8792 => x"52ac1b51",
          8793 => x"ffa0bc3f",
          8794 => x"8152b01b",
          8795 => x"51ffa095",
          8796 => x"3f8652b2",
          8797 => x"1b51ffa0",
          8798 => x"8c3fff80",
          8799 => x"0b80c01c",
          8800 => x"34a90b80",
          8801 => x"c21c3493",
          8802 => x"5382b4ec",
          8803 => x"5280c71b",
          8804 => x"51ae3982",
          8805 => x"88b20a52",
          8806 => x"a71b51ff",
          8807 => x"a0853f7c",
          8808 => x"83ffff06",
          8809 => x"52961b51",
          8810 => x"ff9fda3f",
          8811 => x"ff800ba4",
          8812 => x"1c34a90b",
          8813 => x"a61c3493",
          8814 => x"5382b580",
          8815 => x"52ab1b51",
          8816 => x"ffa08f3f",
          8817 => x"82d4d552",
          8818 => x"83fe1b70",
          8819 => x"5259ff9f",
          8820 => x"b43f8154",
          8821 => x"60537a52",
          8822 => x"7e51ff9b",
          8823 => x"d73f8156",
          8824 => x"82bbdc08",
          8825 => x"83e7387d",
          8826 => x"832e0981",
          8827 => x"0680ee38",
          8828 => x"75546086",
          8829 => x"05537a52",
          8830 => x"7e51ff9b",
          8831 => x"b73f8480",
          8832 => x"5380527a",
          8833 => x"51ff9fed",
          8834 => x"3f848b85",
          8835 => x"a4d2527a",
          8836 => x"51ff9f8f",
          8837 => x"3f868a85",
          8838 => x"e4f25283",
          8839 => x"e41b51ff",
          8840 => x"9f813fff",
          8841 => x"185283e8",
          8842 => x"1b51ff9e",
          8843 => x"f63f8252",
          8844 => x"83ec1b51",
          8845 => x"ff9eec3f",
          8846 => x"82d4d552",
          8847 => x"7851ff9e",
          8848 => x"c43f7554",
          8849 => x"60870553",
          8850 => x"7a527e51",
          8851 => x"ff9ae53f",
          8852 => x"75546016",
          8853 => x"537a527e",
          8854 => x"51ff9ad8",
          8855 => x"3f655380",
          8856 => x"527a51ff",
          8857 => x"9f8f3f7f",
          8858 => x"5680587d",
          8859 => x"832e0981",
          8860 => x"069a38f8",
          8861 => x"527a51ff",
          8862 => x"9ea93fff",
          8863 => x"52841b51",
          8864 => x"ff9ea03f",
          8865 => x"f00a5288",
          8866 => x"1b519139",
          8867 => x"87fffff8",
          8868 => x"557d812e",
          8869 => x"8338f855",
          8870 => x"74527a51",
          8871 => x"ff9e843f",
          8872 => x"7c556157",
          8873 => x"74622683",
          8874 => x"38745776",
          8875 => x"5475537a",
          8876 => x"527e51ff",
          8877 => x"99fe3f82",
          8878 => x"bbdc0882",
          8879 => x"87388480",
          8880 => x"5382bbdc",
          8881 => x"08527a51",
          8882 => x"ff9eaa3f",
          8883 => x"76167578",
          8884 => x"31565674",
          8885 => x"cd388118",
          8886 => x"5877802e",
          8887 => x"ff8d3879",
          8888 => x"557d832e",
          8889 => x"83386355",
          8890 => x"61577462",
          8891 => x"26833874",
          8892 => x"57765475",
          8893 => x"537a527e",
          8894 => x"51ff99b8",
          8895 => x"3f82bbdc",
          8896 => x"0881c138",
          8897 => x"76167578",
          8898 => x"31565674",
          8899 => x"db388c56",
          8900 => x"7d832e93",
          8901 => x"38865666",
          8902 => x"83ffff26",
          8903 => x"8a388456",
          8904 => x"7d822e83",
          8905 => x"38815664",
          8906 => x"81065877",
          8907 => x"80fe3884",
          8908 => x"80537752",
          8909 => x"7a51ff9d",
          8910 => x"bc3f82d4",
          8911 => x"d5527851",
          8912 => x"ff9cc23f",
          8913 => x"83be1b55",
          8914 => x"77753481",
          8915 => x"0b811634",
          8916 => x"810b8216",
          8917 => x"34778316",
          8918 => x"34758416",
          8919 => x"34606705",
          8920 => x"5680fdc1",
          8921 => x"527551fe",
          8922 => x"b0993ffe",
          8923 => x"0b851634",
          8924 => x"82bbdc08",
          8925 => x"822abf07",
          8926 => x"56758616",
          8927 => x"3482bbdc",
          8928 => x"08871634",
          8929 => x"605283c6",
          8930 => x"1b51ff9c",
          8931 => x"963f6652",
          8932 => x"83ca1b51",
          8933 => x"ff9c8c3f",
          8934 => x"81547753",
          8935 => x"7a527e51",
          8936 => x"ff98913f",
          8937 => x"815682bb",
          8938 => x"dc08a238",
          8939 => x"80538052",
          8940 => x"7e51ff99",
          8941 => x"e33f8156",
          8942 => x"82bbdc08",
          8943 => x"90388939",
          8944 => x"8e568a39",
          8945 => x"81568639",
          8946 => x"82bbdc08",
          8947 => x"567582bb",
          8948 => x"dc0c993d",
          8949 => x"0d04f53d",
          8950 => x"0d7d605b",
          8951 => x"59807960",
          8952 => x"ff055a57",
          8953 => x"57767825",
          8954 => x"b4388d3d",
          8955 => x"f8115555",
          8956 => x"8153fc15",
          8957 => x"527951c9",
          8958 => x"dc3f7a81",
          8959 => x"2e098106",
          8960 => x"9c388c3d",
          8961 => x"3355748d",
          8962 => x"2edb3874",
          8963 => x"76708105",
          8964 => x"58348117",
          8965 => x"57748a2e",
          8966 => x"098106c9",
          8967 => x"38807634",
          8968 => x"78557683",
          8969 => x"38765574",
          8970 => x"82bbdc0c",
          8971 => x"8d3d0d04",
          8972 => x"f73d0d7b",
          8973 => x"028405b3",
          8974 => x"05335957",
          8975 => x"778a2e09",
          8976 => x"81068738",
          8977 => x"8d527651",
          8978 => x"e73f8417",
          8979 => x"08568076",
          8980 => x"24be3888",
          8981 => x"17087717",
          8982 => x"8c055659",
          8983 => x"77753481",
          8984 => x"1656bb76",
          8985 => x"25a1388b",
          8986 => x"3dfc0554",
          8987 => x"75538c17",
          8988 => x"52760851",
          8989 => x"cbdc3f79",
          8990 => x"76327030",
          8991 => x"7072079f",
          8992 => x"2a703053",
          8993 => x"51565675",
          8994 => x"84180c81",
          8995 => x"1988180c",
          8996 => x"8b3d0d04",
          8997 => x"f93d0d79",
          8998 => x"84110856",
          8999 => x"56807524",
          9000 => x"a738893d",
          9001 => x"fc055474",
          9002 => x"538c1652",
          9003 => x"750851cb",
          9004 => x"a13f82bb",
          9005 => x"dc089138",
          9006 => x"84160878",
          9007 => x"2e098106",
          9008 => x"87388816",
          9009 => x"08558339",
          9010 => x"ff557482",
          9011 => x"bbdc0c89",
          9012 => x"3d0d04fd",
          9013 => x"3d0d7554",
          9014 => x"80cc5380",
          9015 => x"527351ff",
          9016 => x"9a933f76",
          9017 => x"740c853d",
          9018 => x"0d04ea3d",
          9019 => x"0d0280e3",
          9020 => x"05336a53",
          9021 => x"863d7053",
          9022 => x"5454d83f",
          9023 => x"73527251",
          9024 => x"feae3f72",
          9025 => x"51ff8d3f",
          9026 => x"983d0d04",
          9027 => x"00ffffff",
          9028 => x"ff00ffff",
          9029 => x"ffff00ff",
          9030 => x"ffffff00",
          9031 => x"00002baa",
          9032 => x"00002b2e",
          9033 => x"00002b35",
          9034 => x"00002b3c",
          9035 => x"00002b43",
          9036 => x"00002b4a",
          9037 => x"00002b51",
          9038 => x"00002b58",
          9039 => x"00002b5f",
          9040 => x"00002b66",
          9041 => x"00002b6d",
          9042 => x"00002b74",
          9043 => x"00002b7a",
          9044 => x"00002b80",
          9045 => x"00002b86",
          9046 => x"00002b8c",
          9047 => x"00002b92",
          9048 => x"00002b98",
          9049 => x"00002b9e",
          9050 => x"00002ba4",
          9051 => x"00004382",
          9052 => x"00004388",
          9053 => x"0000438e",
          9054 => x"00004394",
          9055 => x"0000439a",
          9056 => x"000049b9",
          9057 => x"00004ab9",
          9058 => x"00004bca",
          9059 => x"00004e22",
          9060 => x"00004aa1",
          9061 => x"0000488e",
          9062 => x"00004c92",
          9063 => x"00004df3",
          9064 => x"00004cd5",
          9065 => x"00004d6b",
          9066 => x"00004cf1",
          9067 => x"00004b74",
          9068 => x"0000488e",
          9069 => x"00004bca",
          9070 => x"00004bf3",
          9071 => x"00004c92",
          9072 => x"0000488e",
          9073 => x"0000488e",
          9074 => x"00004cf1",
          9075 => x"00004d6b",
          9076 => x"00004df3",
          9077 => x"00004e22",
          9078 => x"00000e31",
          9079 => x"0000171a",
          9080 => x"0000171a",
          9081 => x"00000e60",
          9082 => x"0000171a",
          9083 => x"0000171a",
          9084 => x"0000171a",
          9085 => x"0000171a",
          9086 => x"0000171a",
          9087 => x"0000171a",
          9088 => x"0000171a",
          9089 => x"00000e1d",
          9090 => x"0000171a",
          9091 => x"00000e48",
          9092 => x"00000e78",
          9093 => x"0000171a",
          9094 => x"0000171a",
          9095 => x"0000171a",
          9096 => x"0000171a",
          9097 => x"0000171a",
          9098 => x"0000171a",
          9099 => x"0000171a",
          9100 => x"0000171a",
          9101 => x"0000171a",
          9102 => x"0000171a",
          9103 => x"0000171a",
          9104 => x"0000171a",
          9105 => x"0000171a",
          9106 => x"0000171a",
          9107 => x"0000171a",
          9108 => x"0000171a",
          9109 => x"0000171a",
          9110 => x"0000171a",
          9111 => x"0000171a",
          9112 => x"0000171a",
          9113 => x"0000171a",
          9114 => x"0000171a",
          9115 => x"0000171a",
          9116 => x"0000171a",
          9117 => x"0000171a",
          9118 => x"0000171a",
          9119 => x"0000171a",
          9120 => x"0000171a",
          9121 => x"0000171a",
          9122 => x"0000171a",
          9123 => x"0000171a",
          9124 => x"0000171a",
          9125 => x"0000171a",
          9126 => x"0000171a",
          9127 => x"0000171a",
          9128 => x"0000171a",
          9129 => x"00000fa8",
          9130 => x"0000171a",
          9131 => x"0000171a",
          9132 => x"0000171a",
          9133 => x"0000171a",
          9134 => x"00001116",
          9135 => x"0000171a",
          9136 => x"0000171a",
          9137 => x"0000171a",
          9138 => x"0000171a",
          9139 => x"0000171a",
          9140 => x"0000171a",
          9141 => x"0000171a",
          9142 => x"0000171a",
          9143 => x"0000171a",
          9144 => x"0000171a",
          9145 => x"00000ed8",
          9146 => x"0000103f",
          9147 => x"00000eaf",
          9148 => x"00000eaf",
          9149 => x"00000eaf",
          9150 => x"0000171a",
          9151 => x"0000103f",
          9152 => x"0000171a",
          9153 => x"0000171a",
          9154 => x"00000e98",
          9155 => x"0000171a",
          9156 => x"0000171a",
          9157 => x"000010ec",
          9158 => x"000010f7",
          9159 => x"0000171a",
          9160 => x"0000171a",
          9161 => x"00000f11",
          9162 => x"0000171a",
          9163 => x"0000111f",
          9164 => x"0000171a",
          9165 => x"0000171a",
          9166 => x"00001116",
          9167 => x"64696e69",
          9168 => x"74000000",
          9169 => x"64696f63",
          9170 => x"746c0000",
          9171 => x"66696e69",
          9172 => x"74000000",
          9173 => x"666c6f61",
          9174 => x"64000000",
          9175 => x"66657865",
          9176 => x"63000000",
          9177 => x"6d636c65",
          9178 => x"61720000",
          9179 => x"6d636f70",
          9180 => x"79000000",
          9181 => x"6d646966",
          9182 => x"66000000",
          9183 => x"6d64756d",
          9184 => x"70000000",
          9185 => x"6d656200",
          9186 => x"6d656800",
          9187 => x"6d657700",
          9188 => x"68696400",
          9189 => x"68696500",
          9190 => x"68666400",
          9191 => x"68666500",
          9192 => x"63616c6c",
          9193 => x"00000000",
          9194 => x"6a6d7000",
          9195 => x"72657374",
          9196 => x"61727400",
          9197 => x"72657365",
          9198 => x"74000000",
          9199 => x"696e666f",
          9200 => x"00000000",
          9201 => x"74657374",
          9202 => x"00000000",
          9203 => x"74626173",
          9204 => x"69630000",
          9205 => x"6d626173",
          9206 => x"69630000",
          9207 => x"6b696c6f",
          9208 => x"00000000",
          9209 => x"65640000",
          9210 => x"4469736b",
          9211 => x"20457272",
          9212 => x"6f720000",
          9213 => x"496e7465",
          9214 => x"726e616c",
          9215 => x"20657272",
          9216 => x"6f722e00",
          9217 => x"4469736b",
          9218 => x"206e6f74",
          9219 => x"20726561",
          9220 => x"64792e00",
          9221 => x"4e6f2066",
          9222 => x"696c6520",
          9223 => x"666f756e",
          9224 => x"642e0000",
          9225 => x"4e6f2070",
          9226 => x"61746820",
          9227 => x"666f756e",
          9228 => x"642e0000",
          9229 => x"496e7661",
          9230 => x"6c696420",
          9231 => x"66696c65",
          9232 => x"6e616d65",
          9233 => x"2e000000",
          9234 => x"41636365",
          9235 => x"73732064",
          9236 => x"656e6965",
          9237 => x"642e0000",
          9238 => x"46696c65",
          9239 => x"20616c72",
          9240 => x"65616479",
          9241 => x"20657869",
          9242 => x"7374732e",
          9243 => x"00000000",
          9244 => x"46696c65",
          9245 => x"2068616e",
          9246 => x"646c6520",
          9247 => x"696e7661",
          9248 => x"6c69642e",
          9249 => x"00000000",
          9250 => x"53442069",
          9251 => x"73207772",
          9252 => x"69746520",
          9253 => x"70726f74",
          9254 => x"65637465",
          9255 => x"642e0000",
          9256 => x"44726976",
          9257 => x"65206e75",
          9258 => x"6d626572",
          9259 => x"20697320",
          9260 => x"696e7661",
          9261 => x"6c69642e",
          9262 => x"00000000",
          9263 => x"4469736b",
          9264 => x"206e6f74",
          9265 => x"20656e61",
          9266 => x"626c6564",
          9267 => x"2e000000",
          9268 => x"4e6f2063",
          9269 => x"6f6d7061",
          9270 => x"7469626c",
          9271 => x"65206669",
          9272 => x"6c657379",
          9273 => x"7374656d",
          9274 => x"20666f75",
          9275 => x"6e64206f",
          9276 => x"6e206469",
          9277 => x"736b2e00",
          9278 => x"466f726d",
          9279 => x"61742061",
          9280 => x"626f7274",
          9281 => x"65642e00",
          9282 => x"54696d65",
          9283 => x"6f75742c",
          9284 => x"206f7065",
          9285 => x"72617469",
          9286 => x"6f6e2063",
          9287 => x"616e6365",
          9288 => x"6c6c6564",
          9289 => x"2e000000",
          9290 => x"46696c65",
          9291 => x"20697320",
          9292 => x"6c6f636b",
          9293 => x"65642e00",
          9294 => x"496e7375",
          9295 => x"66666963",
          9296 => x"69656e74",
          9297 => x"206d656d",
          9298 => x"6f72792e",
          9299 => x"00000000",
          9300 => x"546f6f20",
          9301 => x"6d616e79",
          9302 => x"206f7065",
          9303 => x"6e206669",
          9304 => x"6c65732e",
          9305 => x"00000000",
          9306 => x"50617261",
          9307 => x"6d657465",
          9308 => x"72732069",
          9309 => x"6e636f72",
          9310 => x"72656374",
          9311 => x"2e000000",
          9312 => x"53756363",
          9313 => x"6573732e",
          9314 => x"00000000",
          9315 => x"556e6b6e",
          9316 => x"6f776e20",
          9317 => x"6572726f",
          9318 => x"722e0000",
          9319 => x"0a256c75",
          9320 => x"20627974",
          9321 => x"65732025",
          9322 => x"73206174",
          9323 => x"20256c75",
          9324 => x"20627974",
          9325 => x"65732f73",
          9326 => x"65632e0a",
          9327 => x"00000000",
          9328 => x"72656164",
          9329 => x"00000000",
          9330 => x"2530386c",
          9331 => x"58000000",
          9332 => x"3a202000",
          9333 => x"25303458",
          9334 => x"00000000",
          9335 => x"20202020",
          9336 => x"20202020",
          9337 => x"00000000",
          9338 => x"25303258",
          9339 => x"00000000",
          9340 => x"20200000",
          9341 => x"207c0000",
          9342 => x"7c000000",
          9343 => x"5a505554",
          9344 => x"41000000",
          9345 => x"0a2a2a20",
          9346 => x"25732028",
          9347 => x"00000000",
          9348 => x"30322f30",
          9349 => x"352f3230",
          9350 => x"32300000",
          9351 => x"76312e35",
          9352 => x"32000000",
          9353 => x"205a5055",
          9354 => x"2c207265",
          9355 => x"76202530",
          9356 => x"32782920",
          9357 => x"25732025",
          9358 => x"73202a2a",
          9359 => x"0a0a0000",
          9360 => x"5a505554",
          9361 => x"4120496e",
          9362 => x"74657272",
          9363 => x"75707420",
          9364 => x"48616e64",
          9365 => x"6c657200",
          9366 => x"54696d65",
          9367 => x"7220696e",
          9368 => x"74657272",
          9369 => x"75707400",
          9370 => x"50533220",
          9371 => x"696e7465",
          9372 => x"72727570",
          9373 => x"74000000",
          9374 => x"494f4354",
          9375 => x"4c205244",
          9376 => x"20696e74",
          9377 => x"65727275",
          9378 => x"70740000",
          9379 => x"494f4354",
          9380 => x"4c205752",
          9381 => x"20696e74",
          9382 => x"65727275",
          9383 => x"70740000",
          9384 => x"55415254",
          9385 => x"30205258",
          9386 => x"20696e74",
          9387 => x"65727275",
          9388 => x"70740000",
          9389 => x"55415254",
          9390 => x"30205458",
          9391 => x"20696e74",
          9392 => x"65727275",
          9393 => x"70740000",
          9394 => x"55415254",
          9395 => x"31205258",
          9396 => x"20696e74",
          9397 => x"65727275",
          9398 => x"70740000",
          9399 => x"55415254",
          9400 => x"31205458",
          9401 => x"20696e74",
          9402 => x"65727275",
          9403 => x"70740000",
          9404 => x"53657474",
          9405 => x"696e6720",
          9406 => x"75702074",
          9407 => x"696d6572",
          9408 => x"2e2e2e00",
          9409 => x"456e6162",
          9410 => x"6c696e67",
          9411 => x"2074696d",
          9412 => x"65722e2e",
          9413 => x"2e000000",
          9414 => x"6175746f",
          9415 => x"65786563",
          9416 => x"2e626174",
          9417 => x"00000000",
          9418 => x"7a707574",
          9419 => x"612e6873",
          9420 => x"74000000",
          9421 => x"303a0000",
          9422 => x"4661696c",
          9423 => x"65642074",
          9424 => x"6f20696e",
          9425 => x"69746961",
          9426 => x"6c697365",
          9427 => x"20736420",
          9428 => x"63617264",
          9429 => x"20302c20",
          9430 => x"706c6561",
          9431 => x"73652069",
          9432 => x"6e697420",
          9433 => x"6d616e75",
          9434 => x"616c6c79",
          9435 => x"2e000000",
          9436 => x"2a200000",
          9437 => x"42616420",
          9438 => x"6469736b",
          9439 => x"20696421",
          9440 => x"00000000",
          9441 => x"496e6974",
          9442 => x"69616c69",
          9443 => x"7365642e",
          9444 => x"00000000",
          9445 => x"4661696c",
          9446 => x"65642074",
          9447 => x"6f20696e",
          9448 => x"69746961",
          9449 => x"6c697365",
          9450 => x"2e000000",
          9451 => x"72633d25",
          9452 => x"640a0000",
          9453 => x"25753a00",
          9454 => x"436c6561",
          9455 => x"72696e67",
          9456 => x"2e2e2e2e",
          9457 => x"00000000",
          9458 => x"436f7079",
          9459 => x"696e672e",
          9460 => x"2e2e0000",
          9461 => x"436f6d70",
          9462 => x"6172696e",
          9463 => x"672e2e2e",
          9464 => x"00000000",
          9465 => x"2530386c",
          9466 => x"78282530",
          9467 => x"3878292d",
          9468 => x"3e253038",
          9469 => x"6c782825",
          9470 => x"30387829",
          9471 => x"0a000000",
          9472 => x"44756d70",
          9473 => x"204d656d",
          9474 => x"6f727900",
          9475 => x"0a436f6d",
          9476 => x"706c6574",
          9477 => x"652e0000",
          9478 => x"2530386c",
          9479 => x"58202530",
          9480 => x"32582d00",
          9481 => x"3f3f3f00",
          9482 => x"2530386c",
          9483 => x"58202530",
          9484 => x"34582d00",
          9485 => x"2530386c",
          9486 => x"58202530",
          9487 => x"386c582d",
          9488 => x"00000000",
          9489 => x"44697361",
          9490 => x"626c696e",
          9491 => x"6720696e",
          9492 => x"74657272",
          9493 => x"75707473",
          9494 => x"00000000",
          9495 => x"456e6162",
          9496 => x"6c696e67",
          9497 => x"20696e74",
          9498 => x"65727275",
          9499 => x"70747300",
          9500 => x"44697361",
          9501 => x"626c6564",
          9502 => x"20756172",
          9503 => x"74206669",
          9504 => x"666f0000",
          9505 => x"456e6162",
          9506 => x"6c696e67",
          9507 => x"20756172",
          9508 => x"74206669",
          9509 => x"666f0000",
          9510 => x"45786563",
          9511 => x"7574696e",
          9512 => x"6720636f",
          9513 => x"64652040",
          9514 => x"20253038",
          9515 => x"6c78202e",
          9516 => x"2e2e0a00",
          9517 => x"43616c6c",
          9518 => x"696e6720",
          9519 => x"636f6465",
          9520 => x"20402025",
          9521 => x"30386c78",
          9522 => x"202e2e2e",
          9523 => x"0a000000",
          9524 => x"43616c6c",
          9525 => x"20726574",
          9526 => x"75726e65",
          9527 => x"6420636f",
          9528 => x"64652028",
          9529 => x"2564292e",
          9530 => x"0a000000",
          9531 => x"52657374",
          9532 => x"61727469",
          9533 => x"6e672061",
          9534 => x"70706c69",
          9535 => x"63617469",
          9536 => x"6f6e2e2e",
          9537 => x"2e000000",
          9538 => x"436f6c64",
          9539 => x"20726562",
          9540 => x"6f6f7469",
          9541 => x"6e672e2e",
          9542 => x"2e000000",
          9543 => x"5a505500",
          9544 => x"62696e00",
          9545 => x"25643a5c",
          9546 => x"25735c25",
          9547 => x"732e2573",
          9548 => x"00000000",
          9549 => x"25643a5c",
          9550 => x"25735c25",
          9551 => x"73000000",
          9552 => x"25643a5c",
          9553 => x"25730000",
          9554 => x"42616420",
          9555 => x"636f6d6d",
          9556 => x"616e642e",
          9557 => x"00000000",
          9558 => x"52756e6e",
          9559 => x"696e672e",
          9560 => x"2e2e0000",
          9561 => x"456e6162",
          9562 => x"6c696e67",
          9563 => x"20696e74",
          9564 => x"65727275",
          9565 => x"7074732e",
          9566 => x"2e2e0000",
          9567 => x"25642f25",
          9568 => x"642f2564",
          9569 => x"2025643a",
          9570 => x"25643a25",
          9571 => x"642e2564",
          9572 => x"25640a00",
          9573 => x"536f4320",
          9574 => x"436f6e66",
          9575 => x"69677572",
          9576 => x"6174696f",
          9577 => x"6e000000",
          9578 => x"20286672",
          9579 => x"6f6d2053",
          9580 => x"6f432063",
          9581 => x"6f6e6669",
          9582 => x"67290000",
          9583 => x"3a0a4465",
          9584 => x"76696365",
          9585 => x"7320696d",
          9586 => x"706c656d",
          9587 => x"656e7465",
          9588 => x"643a0a00",
          9589 => x"20202020",
          9590 => x"57422053",
          9591 => x"4452414d",
          9592 => x"20202825",
          9593 => x"3038583a",
          9594 => x"25303858",
          9595 => x"292e0a00",
          9596 => x"20202020",
          9597 => x"53445241",
          9598 => x"4d202020",
          9599 => x"20202825",
          9600 => x"3038583a",
          9601 => x"25303858",
          9602 => x"292e0a00",
          9603 => x"20202020",
          9604 => x"494e534e",
          9605 => x"20425241",
          9606 => x"4d202825",
          9607 => x"3038583a",
          9608 => x"25303858",
          9609 => x"292e0a00",
          9610 => x"20202020",
          9611 => x"4252414d",
          9612 => x"20202020",
          9613 => x"20202825",
          9614 => x"3038583a",
          9615 => x"25303858",
          9616 => x"292e0a00",
          9617 => x"20202020",
          9618 => x"52414d20",
          9619 => x"20202020",
          9620 => x"20202825",
          9621 => x"3038583a",
          9622 => x"25303858",
          9623 => x"292e0a00",
          9624 => x"20202020",
          9625 => x"53442043",
          9626 => x"41524420",
          9627 => x"20202844",
          9628 => x"65766963",
          9629 => x"6573203d",
          9630 => x"25303264",
          9631 => x"292e0a00",
          9632 => x"20202020",
          9633 => x"54494d45",
          9634 => x"52312020",
          9635 => x"20202854",
          9636 => x"696d6572",
          9637 => x"7320203d",
          9638 => x"25303264",
          9639 => x"292e0a00",
          9640 => x"20202020",
          9641 => x"494e5452",
          9642 => x"20435452",
          9643 => x"4c202843",
          9644 => x"68616e6e",
          9645 => x"656c733d",
          9646 => x"25303264",
          9647 => x"292e0a00",
          9648 => x"20202020",
          9649 => x"57495348",
          9650 => x"424f4e45",
          9651 => x"20425553",
          9652 => x"0a000000",
          9653 => x"20202020",
          9654 => x"57422049",
          9655 => x"32430a00",
          9656 => x"20202020",
          9657 => x"494f4354",
          9658 => x"4c0a0000",
          9659 => x"20202020",
          9660 => x"5053320a",
          9661 => x"00000000",
          9662 => x"20202020",
          9663 => x"5350490a",
          9664 => x"00000000",
          9665 => x"41646472",
          9666 => x"65737365",
          9667 => x"733a0a00",
          9668 => x"20202020",
          9669 => x"43505520",
          9670 => x"52657365",
          9671 => x"74205665",
          9672 => x"63746f72",
          9673 => x"20416464",
          9674 => x"72657373",
          9675 => x"203d2025",
          9676 => x"3038580a",
          9677 => x"00000000",
          9678 => x"20202020",
          9679 => x"43505520",
          9680 => x"4d656d6f",
          9681 => x"72792053",
          9682 => x"74617274",
          9683 => x"20416464",
          9684 => x"72657373",
          9685 => x"203d2025",
          9686 => x"3038580a",
          9687 => x"00000000",
          9688 => x"20202020",
          9689 => x"53746163",
          9690 => x"6b205374",
          9691 => x"61727420",
          9692 => x"41646472",
          9693 => x"65737320",
          9694 => x"20202020",
          9695 => x"203d2025",
          9696 => x"3038580a",
          9697 => x"00000000",
          9698 => x"4d697363",
          9699 => x"3a0a0000",
          9700 => x"20202020",
          9701 => x"5a505520",
          9702 => x"49642020",
          9703 => x"20202020",
          9704 => x"20202020",
          9705 => x"20202020",
          9706 => x"20202020",
          9707 => x"203d2025",
          9708 => x"3034580a",
          9709 => x"00000000",
          9710 => x"20202020",
          9711 => x"53797374",
          9712 => x"656d2043",
          9713 => x"6c6f636b",
          9714 => x"20467265",
          9715 => x"71202020",
          9716 => x"20202020",
          9717 => x"203d2025",
          9718 => x"642e2530",
          9719 => x"34644d48",
          9720 => x"7a0a0000",
          9721 => x"20202020",
          9722 => x"53445241",
          9723 => x"4d20436c",
          9724 => x"6f636b20",
          9725 => x"46726571",
          9726 => x"20202020",
          9727 => x"20202020",
          9728 => x"203d2025",
          9729 => x"642e2530",
          9730 => x"34644d48",
          9731 => x"7a0a0000",
          9732 => x"20202020",
          9733 => x"57697368",
          9734 => x"626f6e65",
          9735 => x"20534452",
          9736 => x"414d2043",
          9737 => x"6c6f636b",
          9738 => x"20467265",
          9739 => x"713d2025",
          9740 => x"642e2530",
          9741 => x"34644d48",
          9742 => x"7a0a0000",
          9743 => x"536d616c",
          9744 => x"6c000000",
          9745 => x"4d656469",
          9746 => x"756d0000",
          9747 => x"466c6578",
          9748 => x"00000000",
          9749 => x"45564f00",
          9750 => x"45564f6d",
          9751 => x"696e0000",
          9752 => x"556e6b6e",
          9753 => x"6f776e00",
          9754 => x"000099c4",
          9755 => x"01000000",
          9756 => x"00000002",
          9757 => x"000099c0",
          9758 => x"01000000",
          9759 => x"00000003",
          9760 => x"000099bc",
          9761 => x"01000000",
          9762 => x"00000004",
          9763 => x"000099b8",
          9764 => x"01000000",
          9765 => x"00000005",
          9766 => x"000099b4",
          9767 => x"01000000",
          9768 => x"00000006",
          9769 => x"000099b0",
          9770 => x"01000000",
          9771 => x"00000007",
          9772 => x"000099ac",
          9773 => x"01000000",
          9774 => x"00000001",
          9775 => x"000099a8",
          9776 => x"01000000",
          9777 => x"00000008",
          9778 => x"000099a4",
          9779 => x"01000000",
          9780 => x"0000000b",
          9781 => x"000099a0",
          9782 => x"01000000",
          9783 => x"00000009",
          9784 => x"0000999c",
          9785 => x"01000000",
          9786 => x"0000000a",
          9787 => x"00009998",
          9788 => x"04000000",
          9789 => x"0000000d",
          9790 => x"00009994",
          9791 => x"04000000",
          9792 => x"0000000c",
          9793 => x"00009990",
          9794 => x"04000000",
          9795 => x"0000000e",
          9796 => x"0000998c",
          9797 => x"03000000",
          9798 => x"0000000f",
          9799 => x"00009988",
          9800 => x"04000000",
          9801 => x"0000000f",
          9802 => x"00009984",
          9803 => x"04000000",
          9804 => x"00000010",
          9805 => x"00009980",
          9806 => x"04000000",
          9807 => x"00000011",
          9808 => x"0000997c",
          9809 => x"03000000",
          9810 => x"00000012",
          9811 => x"00009978",
          9812 => x"03000000",
          9813 => x"00000013",
          9814 => x"00009974",
          9815 => x"03000000",
          9816 => x"00000014",
          9817 => x"00009970",
          9818 => x"03000000",
          9819 => x"00000015",
          9820 => x"1b5b4400",
          9821 => x"1b5b4300",
          9822 => x"1b5b4200",
          9823 => x"1b5b4100",
          9824 => x"1b5b367e",
          9825 => x"1b5b357e",
          9826 => x"1b5b347e",
          9827 => x"1b304600",
          9828 => x"1b5b337e",
          9829 => x"1b5b327e",
          9830 => x"1b5b317e",
          9831 => x"10000000",
          9832 => x"0e000000",
          9833 => x"0d000000",
          9834 => x"0b000000",
          9835 => x"08000000",
          9836 => x"06000000",
          9837 => x"05000000",
          9838 => x"04000000",
          9839 => x"03000000",
          9840 => x"02000000",
          9841 => x"01000000",
          9842 => x"68697374",
          9843 => x"6f727900",
          9844 => x"68697374",
          9845 => x"00000000",
          9846 => x"21000000",
          9847 => x"2530346c",
          9848 => x"75202025",
          9849 => x"730a0000",
          9850 => x"4661696c",
          9851 => x"65642074",
          9852 => x"6f207265",
          9853 => x"73657420",
          9854 => x"74686520",
          9855 => x"68697374",
          9856 => x"6f727920",
          9857 => x"66696c65",
          9858 => x"20746f20",
          9859 => x"454f462e",
          9860 => x"00000000",
          9861 => x"43616e6e",
          9862 => x"6f74206f",
          9863 => x"70656e2f",
          9864 => x"63726561",
          9865 => x"74652068",
          9866 => x"6973746f",
          9867 => x"72792066",
          9868 => x"696c652c",
          9869 => x"20646973",
          9870 => x"61626c69",
          9871 => x"6e672e00",
          9872 => x"53440000",
          9873 => x"222a2b2c",
          9874 => x"3a3b3c3d",
          9875 => x"3e3f5b5d",
          9876 => x"7c7f0000",
          9877 => x"46415400",
          9878 => x"46415433",
          9879 => x"32000000",
          9880 => x"ebfe904d",
          9881 => x"53444f53",
          9882 => x"352e3000",
          9883 => x"4e4f204e",
          9884 => x"414d4520",
          9885 => x"20202046",
          9886 => x"41543332",
          9887 => x"20202000",
          9888 => x"4e4f204e",
          9889 => x"414d4520",
          9890 => x"20202046",
          9891 => x"41542020",
          9892 => x"20202000",
          9893 => x"00009a40",
          9894 => x"00000000",
          9895 => x"00000000",
          9896 => x"00000000",
          9897 => x"809a4541",
          9898 => x"8e418f80",
          9899 => x"45454549",
          9900 => x"49498e8f",
          9901 => x"9092924f",
          9902 => x"994f5555",
          9903 => x"59999a9b",
          9904 => x"9c9d9e9f",
          9905 => x"41494f55",
          9906 => x"a5a5a6a7",
          9907 => x"a8a9aaab",
          9908 => x"acadaeaf",
          9909 => x"b0b1b2b3",
          9910 => x"b4b5b6b7",
          9911 => x"b8b9babb",
          9912 => x"bcbdbebf",
          9913 => x"c0c1c2c3",
          9914 => x"c4c5c6c7",
          9915 => x"c8c9cacb",
          9916 => x"cccdcecf",
          9917 => x"d0d1d2d3",
          9918 => x"d4d5d6d7",
          9919 => x"d8d9dadb",
          9920 => x"dcdddedf",
          9921 => x"e0e1e2e3",
          9922 => x"e4e5e6e7",
          9923 => x"e8e9eaeb",
          9924 => x"ecedeeef",
          9925 => x"f0f1f2f3",
          9926 => x"f4f5f6f7",
          9927 => x"f8f9fafb",
          9928 => x"fcfdfeff",
          9929 => x"2b2e2c3b",
          9930 => x"3d5b5d2f",
          9931 => x"5c222a3a",
          9932 => x"3c3e3f7c",
          9933 => x"7f000000",
          9934 => x"00010004",
          9935 => x"00100040",
          9936 => x"01000200",
          9937 => x"00000000",
          9938 => x"00010002",
          9939 => x"00040008",
          9940 => x"00100020",
          9941 => x"00000000",
          9942 => x"00000000",
          9943 => x"00008f3c",
          9944 => x"01020100",
          9945 => x"00000000",
          9946 => x"00000000",
          9947 => x"00008f44",
          9948 => x"01040100",
          9949 => x"00000000",
          9950 => x"00000000",
          9951 => x"00008f4c",
          9952 => x"01140300",
          9953 => x"00000000",
          9954 => x"00000000",
          9955 => x"00008f54",
          9956 => x"012b0300",
          9957 => x"00000000",
          9958 => x"00000000",
          9959 => x"00008f5c",
          9960 => x"01300300",
          9961 => x"00000000",
          9962 => x"00000000",
          9963 => x"00008f64",
          9964 => x"013c0400",
          9965 => x"00000000",
          9966 => x"00000000",
          9967 => x"00008f6c",
          9968 => x"013d0400",
          9969 => x"00000000",
          9970 => x"00000000",
          9971 => x"00008f74",
          9972 => x"013f0400",
          9973 => x"00000000",
          9974 => x"00000000",
          9975 => x"00008f7c",
          9976 => x"01400400",
          9977 => x"00000000",
          9978 => x"00000000",
          9979 => x"00008f84",
          9980 => x"01410400",
          9981 => x"00000000",
          9982 => x"00000000",
          9983 => x"00008f88",
          9984 => x"01420400",
          9985 => x"00000000",
          9986 => x"00000000",
          9987 => x"00008f8c",
          9988 => x"01430400",
          9989 => x"00000000",
          9990 => x"00000000",
          9991 => x"00008f90",
          9992 => x"01500500",
          9993 => x"00000000",
          9994 => x"00000000",
          9995 => x"00008f94",
          9996 => x"01510500",
          9997 => x"00000000",
          9998 => x"00000000",
          9999 => x"00008f98",
         10000 => x"01540500",
         10001 => x"00000000",
         10002 => x"00000000",
         10003 => x"00008f9c",
         10004 => x"01550500",
         10005 => x"00000000",
         10006 => x"00000000",
         10007 => x"00008fa0",
         10008 => x"01790700",
         10009 => x"00000000",
         10010 => x"00000000",
         10011 => x"00008fa8",
         10012 => x"01780700",
         10013 => x"00000000",
         10014 => x"00000000",
         10015 => x"00008fac",
         10016 => x"01820800",
         10017 => x"00000000",
         10018 => x"00000000",
         10019 => x"00008fb4",
         10020 => x"01830800",
         10021 => x"00000000",
         10022 => x"00000000",
         10023 => x"00008fbc",
         10024 => x"01850800",
         10025 => x"00000000",
         10026 => x"00000000",
         10027 => x"00008fc4",
         10028 => x"01870800",
         10029 => x"00000000",
         10030 => x"00000000",
         10031 => x"00008fcc",
         10032 => x"018c0900",
         10033 => x"00000000",
         10034 => x"00000000",
         10035 => x"00008fd4",
         10036 => x"018d0900",
         10037 => x"00000000",
         10038 => x"00000000",
         10039 => x"00008fdc",
         10040 => x"018e0900",
         10041 => x"00000000",
         10042 => x"00000000",
         10043 => x"00008fe4",
         10044 => x"018f0900",
         10045 => x"00000000",
         10046 => x"00000000",
         10047 => x"00000000",
         10048 => x"00000000",
         10049 => x"00007fff",
         10050 => x"00000000",
         10051 => x"00007fff",
         10052 => x"00010000",
         10053 => x"00007fff",
         10054 => x"00010000",
         10055 => x"00810000",
         10056 => x"01000000",
         10057 => x"017fffff",
         10058 => x"00000000",
         10059 => x"00000000",
         10060 => x"00007800",
         10061 => x"00000000",
         10062 => x"05f5e100",
         10063 => x"05f5e100",
         10064 => x"05f5e100",
         10065 => x"00000000",
         10066 => x"01010101",
         10067 => x"01010101",
         10068 => x"01011001",
         10069 => x"01000000",
         10070 => x"00000000",
         10071 => x"00000000",
         10072 => x"00000000",
         10073 => x"00000000",
         10074 => x"00000000",
         10075 => x"00000000",
         10076 => x"00000000",
         10077 => x"00000000",
         10078 => x"00000000",
         10079 => x"00000000",
         10080 => x"00000000",
         10081 => x"00000000",
         10082 => x"00000000",
         10083 => x"00000000",
         10084 => x"00000000",
         10085 => x"00000000",
         10086 => x"00000000",
         10087 => x"00000000",
         10088 => x"00000000",
         10089 => x"00000000",
         10090 => x"00000000",
         10091 => x"00000000",
         10092 => x"00000000",
         10093 => x"00000000",
         10094 => x"000099c8",
         10095 => x"01000000",
         10096 => x"000099d0",
         10097 => x"01000000",
         10098 => x"000099d8",
         10099 => x"02000000",
         10100 => x"00000000",
         10101 => x"00000000",
         10102 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

