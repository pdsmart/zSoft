-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b0b93",
          2049 => x"8c040000",
          2050 => x"00000000",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b92",
          2121 => x"f0040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b92d3",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b81e1",
          2210 => x"b0738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"92d80400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b0b94",
          2219 => x"912d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b0b95",
          2227 => x"fd2d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"94040b0b",
          2317 => x"0b8ca304",
          2318 => x"0b0b0b8c",
          2319 => x"b2040b0b",
          2320 => x"0b8cc104",
          2321 => x"0b0b0b8c",
          2322 => x"d0040b0b",
          2323 => x"0b8cdf04",
          2324 => x"0b0b0b8c",
          2325 => x"ee040b0b",
          2326 => x"0b8cfd04",
          2327 => x"0b0b0b8d",
          2328 => x"8c040b0b",
          2329 => x"0b8d9b04",
          2330 => x"0b0b0b8d",
          2331 => x"aa040b0b",
          2332 => x"0b8db904",
          2333 => x"0b0b0b8d",
          2334 => x"c8040b0b",
          2335 => x"0b8dd704",
          2336 => x"0b0b0b8d",
          2337 => x"e6040b0b",
          2338 => x"0b8df504",
          2339 => x"0b0b0b8e",
          2340 => x"84040b0b",
          2341 => x"0b8e9304",
          2342 => x"0b0b0b8e",
          2343 => x"a3040b0b",
          2344 => x"0b8eb304",
          2345 => x"0b0b0b8e",
          2346 => x"c3040b0b",
          2347 => x"0b8ed304",
          2348 => x"0b0b0b8e",
          2349 => x"e3040b0b",
          2350 => x"0b8ef304",
          2351 => x"0b0b0b8f",
          2352 => x"83040b0b",
          2353 => x"0b8f9304",
          2354 => x"0b0b0b8f",
          2355 => x"a3040b0b",
          2356 => x"0b8fb304",
          2357 => x"0b0b0b8f",
          2358 => x"c3040b0b",
          2359 => x"0b8fd304",
          2360 => x"0b0b0b8f",
          2361 => x"e3040b0b",
          2362 => x"0b8ff304",
          2363 => x"0b0b0b90",
          2364 => x"83040b0b",
          2365 => x"0b909304",
          2366 => x"0b0b0b90",
          2367 => x"a3040b0b",
          2368 => x"0b90b304",
          2369 => x"0b0b0b90",
          2370 => x"c3040b0b",
          2371 => x"0b90d304",
          2372 => x"0b0b0b90",
          2373 => x"e3040b0b",
          2374 => x"0b90f304",
          2375 => x"0b0b0b91",
          2376 => x"83040b0b",
          2377 => x"0b919304",
          2378 => x"0b0b0b91",
          2379 => x"a3040b0b",
          2380 => x"0b91b304",
          2381 => x"0b0b0b91",
          2382 => x"c3040b0b",
          2383 => x"0b91d304",
          2384 => x"0b0b0b91",
          2385 => x"e3040b0b",
          2386 => x"0b91f304",
          2387 => x"0b0b0b92",
          2388 => x"82040b0b",
          2389 => x"0b929104",
          2390 => x"0b0b0b92",
          2391 => x"a004ffff",
          2392 => x"ffffffff",
          2393 => x"ffffffff",
          2394 => x"ffffffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0481fefc",
          2434 => x"0ca3ff2d",
          2435 => x"81fefc08",
          2436 => x"83809004",
          2437 => x"81fefc0c",
          2438 => x"b5c82d81",
          2439 => x"fefc0883",
          2440 => x"80900481",
          2441 => x"fefc0cb6",
          2442 => x"872d81fe",
          2443 => x"fc088380",
          2444 => x"900481fe",
          2445 => x"fc0cb6a5",
          2446 => x"2d81fefc",
          2447 => x"08838090",
          2448 => x"0481fefc",
          2449 => x"0cbce32d",
          2450 => x"81fefc08",
          2451 => x"83809004",
          2452 => x"81fefc0c",
          2453 => x"bde12d81",
          2454 => x"fefc0883",
          2455 => x"80900481",
          2456 => x"fefc0cb6",
          2457 => x"c82d81fe",
          2458 => x"fc088380",
          2459 => x"900481fe",
          2460 => x"fc0cbdfe",
          2461 => x"2d81fefc",
          2462 => x"08838090",
          2463 => x"0481fefc",
          2464 => x"0cbff02d",
          2465 => x"81fefc08",
          2466 => x"83809004",
          2467 => x"81fefc0c",
          2468 => x"bc892d81",
          2469 => x"fefc0883",
          2470 => x"80900481",
          2471 => x"fefc0cb6",
          2472 => x"fa2d81fe",
          2473 => x"fc088380",
          2474 => x"900481fe",
          2475 => x"fc0cbc9f",
          2476 => x"2d81fefc",
          2477 => x"08838090",
          2478 => x"0481fefc",
          2479 => x"0cbcc32d",
          2480 => x"81fefc08",
          2481 => x"83809004",
          2482 => x"81fefc0c",
          2483 => x"a68c2d81",
          2484 => x"fefc0883",
          2485 => x"80900481",
          2486 => x"fefc0ca6",
          2487 => x"dd2d81fe",
          2488 => x"fc088380",
          2489 => x"900481fe",
          2490 => x"fc0c9ef9",
          2491 => x"2d81fefc",
          2492 => x"08838090",
          2493 => x"0481fefc",
          2494 => x"0ca0ae2d",
          2495 => x"81fefc08",
          2496 => x"83809004",
          2497 => x"81fefc0c",
          2498 => x"a1e12d81",
          2499 => x"fefc0883",
          2500 => x"80900481",
          2501 => x"fefc0c81",
          2502 => x"84c32d81",
          2503 => x"fefc0883",
          2504 => x"80900481",
          2505 => x"fefc0c81",
          2506 => x"91b42d81",
          2507 => x"fefc0883",
          2508 => x"80900481",
          2509 => x"fefc0c81",
          2510 => x"89a82d81",
          2511 => x"fefc0883",
          2512 => x"80900481",
          2513 => x"fefc0c81",
          2514 => x"8ca52d81",
          2515 => x"fefc0883",
          2516 => x"80900481",
          2517 => x"fefc0c81",
          2518 => x"96c32d81",
          2519 => x"fefc0883",
          2520 => x"80900481",
          2521 => x"fefc0c81",
          2522 => x"9fa32d81",
          2523 => x"fefc0883",
          2524 => x"80900481",
          2525 => x"fefc0c81",
          2526 => x"90962d81",
          2527 => x"fefc0883",
          2528 => x"80900481",
          2529 => x"fefc0c81",
          2530 => x"99e22d81",
          2531 => x"fefc0883",
          2532 => x"80900481",
          2533 => x"fefc0c81",
          2534 => x"9b812d81",
          2535 => x"fefc0883",
          2536 => x"80900481",
          2537 => x"fefc0c81",
          2538 => x"9ba02d81",
          2539 => x"fefc0883",
          2540 => x"80900481",
          2541 => x"fefc0c81",
          2542 => x"a38a2d81",
          2543 => x"fefc0883",
          2544 => x"80900481",
          2545 => x"fefc0c81",
          2546 => x"a0f02d81",
          2547 => x"fefc0883",
          2548 => x"80900481",
          2549 => x"fefc0c81",
          2550 => x"a5de2d81",
          2551 => x"fefc0883",
          2552 => x"80900481",
          2553 => x"fefc0c81",
          2554 => x"9ca42d81",
          2555 => x"fefc0883",
          2556 => x"80900481",
          2557 => x"fefc0c81",
          2558 => x"a8de2d81",
          2559 => x"fefc0883",
          2560 => x"80900481",
          2561 => x"fefc0c81",
          2562 => x"a9df2d81",
          2563 => x"fefc0883",
          2564 => x"80900481",
          2565 => x"fefc0c81",
          2566 => x"92942d81",
          2567 => x"fefc0883",
          2568 => x"80900481",
          2569 => x"fefc0c81",
          2570 => x"91ed2d81",
          2571 => x"fefc0883",
          2572 => x"80900481",
          2573 => x"fefc0c81",
          2574 => x"93982d81",
          2575 => x"fefc0883",
          2576 => x"80900481",
          2577 => x"fefc0c81",
          2578 => x"9cfb2d81",
          2579 => x"fefc0883",
          2580 => x"80900481",
          2581 => x"fefc0c81",
          2582 => x"aad02d81",
          2583 => x"fefc0883",
          2584 => x"80900481",
          2585 => x"fefc0c81",
          2586 => x"acda2d81",
          2587 => x"fefc0883",
          2588 => x"80900481",
          2589 => x"fefc0c81",
          2590 => x"b09c2d81",
          2591 => x"fefc0883",
          2592 => x"80900481",
          2593 => x"fefc0c81",
          2594 => x"83e22d81",
          2595 => x"fefc0883",
          2596 => x"80900481",
          2597 => x"fefc0c81",
          2598 => x"b3882d81",
          2599 => x"fefc0883",
          2600 => x"80900481",
          2601 => x"fefc0c81",
          2602 => x"c1bd2d81",
          2603 => x"fefc0883",
          2604 => x"80900481",
          2605 => x"fefc0c81",
          2606 => x"bfa92d81",
          2607 => x"fefc0883",
          2608 => x"80900481",
          2609 => x"fefc0c80",
          2610 => x"d59d2d81",
          2611 => x"fefc0883",
          2612 => x"80900481",
          2613 => x"fefc0c80",
          2614 => x"d7872d81",
          2615 => x"fefc0883",
          2616 => x"80900481",
          2617 => x"fefc0c80",
          2618 => x"d8eb2d81",
          2619 => x"fefc0883",
          2620 => x"80900481",
          2621 => x"fefc0c9f",
          2622 => x"a22d81fe",
          2623 => x"fc088380",
          2624 => x"900481fe",
          2625 => x"fc0ca084",
          2626 => x"2d81fefc",
          2627 => x"08838090",
          2628 => x"0481fefc",
          2629 => x"0ca2f12d",
          2630 => x"81fefc08",
          2631 => x"83809004",
          2632 => x"81fefc0c",
          2633 => x"81c2d82d",
          2634 => x"81fefc08",
          2635 => x"83809004",
          2636 => x"3c040000",
          2637 => x"10101010",
          2638 => x"10101010",
          2639 => x"10101010",
          2640 => x"10101010",
          2641 => x"10101010",
          2642 => x"10101010",
          2643 => x"10101010",
          2644 => x"10101053",
          2645 => x"51040000",
          2646 => x"7381ff06",
          2647 => x"73830609",
          2648 => x"81058305",
          2649 => x"1010102b",
          2650 => x"0772fc06",
          2651 => x"0c515104",
          2652 => x"72728072",
          2653 => x"8106ff05",
          2654 => x"09720605",
          2655 => x"71105272",
          2656 => x"0a100a53",
          2657 => x"72ed3851",
          2658 => x"51535104",
          2659 => x"81fef070",
          2660 => x"8296b027",
          2661 => x"8e388071",
          2662 => x"70840553",
          2663 => x"0c0b0b0b",
          2664 => x"938f048c",
          2665 => x"815181e0",
          2666 => x"80040081",
          2667 => x"fefc0802",
          2668 => x"81fefc0c",
          2669 => x"fd3d0d80",
          2670 => x"5381fefc",
          2671 => x"088c0508",
          2672 => x"5281fefc",
          2673 => x"08880508",
          2674 => x"5183d43f",
          2675 => x"81fef008",
          2676 => x"7081fef0",
          2677 => x"0c54853d",
          2678 => x"0d81fefc",
          2679 => x"0c0481fe",
          2680 => x"fc080281",
          2681 => x"fefc0cfd",
          2682 => x"3d0d8153",
          2683 => x"81fefc08",
          2684 => x"8c050852",
          2685 => x"81fefc08",
          2686 => x"88050851",
          2687 => x"83a13f81",
          2688 => x"fef00870",
          2689 => x"81fef00c",
          2690 => x"54853d0d",
          2691 => x"81fefc0c",
          2692 => x"0481fefc",
          2693 => x"080281fe",
          2694 => x"fc0cf93d",
          2695 => x"0d800b81",
          2696 => x"fefc08fc",
          2697 => x"050c81fe",
          2698 => x"fc088805",
          2699 => x"088025b9",
          2700 => x"3881fefc",
          2701 => x"08880508",
          2702 => x"3081fefc",
          2703 => x"0888050c",
          2704 => x"800b81fe",
          2705 => x"fc08f405",
          2706 => x"0c81fefc",
          2707 => x"08fc0508",
          2708 => x"8a38810b",
          2709 => x"81fefc08",
          2710 => x"f4050c81",
          2711 => x"fefc08f4",
          2712 => x"050881fe",
          2713 => x"fc08fc05",
          2714 => x"0c81fefc",
          2715 => x"088c0508",
          2716 => x"8025b938",
          2717 => x"81fefc08",
          2718 => x"8c050830",
          2719 => x"81fefc08",
          2720 => x"8c050c80",
          2721 => x"0b81fefc",
          2722 => x"08f0050c",
          2723 => x"81fefc08",
          2724 => x"fc05088a",
          2725 => x"38810b81",
          2726 => x"fefc08f0",
          2727 => x"050c81fe",
          2728 => x"fc08f005",
          2729 => x"0881fefc",
          2730 => x"08fc050c",
          2731 => x"805381fe",
          2732 => x"fc088c05",
          2733 => x"085281fe",
          2734 => x"fc088805",
          2735 => x"085181df",
          2736 => x"3f81fef0",
          2737 => x"087081fe",
          2738 => x"fc08f805",
          2739 => x"0c5481fe",
          2740 => x"fc08fc05",
          2741 => x"08802e90",
          2742 => x"3881fefc",
          2743 => x"08f80508",
          2744 => x"3081fefc",
          2745 => x"08f8050c",
          2746 => x"81fefc08",
          2747 => x"f8050870",
          2748 => x"81fef00c",
          2749 => x"54893d0d",
          2750 => x"81fefc0c",
          2751 => x"0481fefc",
          2752 => x"080281fe",
          2753 => x"fc0cfb3d",
          2754 => x"0d800b81",
          2755 => x"fefc08fc",
          2756 => x"050c81fe",
          2757 => x"fc088805",
          2758 => x"08802599",
          2759 => x"3881fefc",
          2760 => x"08880508",
          2761 => x"3081fefc",
          2762 => x"0888050c",
          2763 => x"810b81fe",
          2764 => x"fc08fc05",
          2765 => x"0c81fefc",
          2766 => x"088c0508",
          2767 => x"80259038",
          2768 => x"81fefc08",
          2769 => x"8c050830",
          2770 => x"81fefc08",
          2771 => x"8c050c81",
          2772 => x"5381fefc",
          2773 => x"088c0508",
          2774 => x"5281fefc",
          2775 => x"08880508",
          2776 => x"51bd3f81",
          2777 => x"fef00870",
          2778 => x"81fefc08",
          2779 => x"f8050c54",
          2780 => x"81fefc08",
          2781 => x"fc050880",
          2782 => x"2e903881",
          2783 => x"fefc08f8",
          2784 => x"05083081",
          2785 => x"fefc08f8",
          2786 => x"050c81fe",
          2787 => x"fc08f805",
          2788 => x"087081fe",
          2789 => x"f00c5487",
          2790 => x"3d0d81fe",
          2791 => x"fc0c0481",
          2792 => x"fefc0802",
          2793 => x"81fefc0c",
          2794 => x"fd3d0d81",
          2795 => x"0b81fefc",
          2796 => x"08fc050c",
          2797 => x"800b81fe",
          2798 => x"fc08f805",
          2799 => x"0c81fefc",
          2800 => x"088c0508",
          2801 => x"81fefc08",
          2802 => x"88050827",
          2803 => x"b93881fe",
          2804 => x"fc08fc05",
          2805 => x"08802eae",
          2806 => x"38800b81",
          2807 => x"fefc088c",
          2808 => x"050824a2",
          2809 => x"3881fefc",
          2810 => x"088c0508",
          2811 => x"1081fefc",
          2812 => x"088c050c",
          2813 => x"81fefc08",
          2814 => x"fc050810",
          2815 => x"81fefc08",
          2816 => x"fc050cff",
          2817 => x"b83981fe",
          2818 => x"fc08fc05",
          2819 => x"08802e80",
          2820 => x"e13881fe",
          2821 => x"fc088c05",
          2822 => x"0881fefc",
          2823 => x"08880508",
          2824 => x"26ad3881",
          2825 => x"fefc0888",
          2826 => x"050881fe",
          2827 => x"fc088c05",
          2828 => x"083181fe",
          2829 => x"fc088805",
          2830 => x"0c81fefc",
          2831 => x"08f80508",
          2832 => x"81fefc08",
          2833 => x"fc050807",
          2834 => x"81fefc08",
          2835 => x"f8050c81",
          2836 => x"fefc08fc",
          2837 => x"0508812a",
          2838 => x"81fefc08",
          2839 => x"fc050c81",
          2840 => x"fefc088c",
          2841 => x"0508812a",
          2842 => x"81fefc08",
          2843 => x"8c050cff",
          2844 => x"953981fe",
          2845 => x"fc089005",
          2846 => x"08802e93",
          2847 => x"3881fefc",
          2848 => x"08880508",
          2849 => x"7081fefc",
          2850 => x"08f4050c",
          2851 => x"51913981",
          2852 => x"fefc08f8",
          2853 => x"05087081",
          2854 => x"fefc08f4",
          2855 => x"050c5181",
          2856 => x"fefc08f4",
          2857 => x"050881fe",
          2858 => x"f00c853d",
          2859 => x"0d81fefc",
          2860 => x"0c04fc3d",
          2861 => x"0d767079",
          2862 => x"7b555555",
          2863 => x"558f7227",
          2864 => x"8c387275",
          2865 => x"07830651",
          2866 => x"70802ea9",
          2867 => x"38ff1252",
          2868 => x"71ff2e98",
          2869 => x"38727081",
          2870 => x"05543374",
          2871 => x"70810556",
          2872 => x"34ff1252",
          2873 => x"71ff2e09",
          2874 => x"8106ea38",
          2875 => x"7481fef0",
          2876 => x"0c863d0d",
          2877 => x"04745172",
          2878 => x"70840554",
          2879 => x"08717084",
          2880 => x"05530c72",
          2881 => x"70840554",
          2882 => x"08717084",
          2883 => x"05530c72",
          2884 => x"70840554",
          2885 => x"08717084",
          2886 => x"05530c72",
          2887 => x"70840554",
          2888 => x"08717084",
          2889 => x"05530cf0",
          2890 => x"1252718f",
          2891 => x"26c93883",
          2892 => x"72279538",
          2893 => x"72708405",
          2894 => x"54087170",
          2895 => x"8405530c",
          2896 => x"fc125271",
          2897 => x"8326ed38",
          2898 => x"7054ff81",
          2899 => x"39fc3d0d",
          2900 => x"76797102",
          2901 => x"8c059f05",
          2902 => x"33575553",
          2903 => x"55837227",
          2904 => x"8a387483",
          2905 => x"06517080",
          2906 => x"2ea438ff",
          2907 => x"125271ff",
          2908 => x"2e933873",
          2909 => x"73708105",
          2910 => x"5534ff12",
          2911 => x"5271ff2e",
          2912 => x"098106ef",
          2913 => x"387481fe",
          2914 => x"f00c863d",
          2915 => x"0d047474",
          2916 => x"882b7507",
          2917 => x"7071902b",
          2918 => x"07515451",
          2919 => x"8f7227a5",
          2920 => x"38727170",
          2921 => x"8405530c",
          2922 => x"72717084",
          2923 => x"05530c72",
          2924 => x"71708405",
          2925 => x"530c7271",
          2926 => x"70840553",
          2927 => x"0cf01252",
          2928 => x"718f26dd",
          2929 => x"38837227",
          2930 => x"90387271",
          2931 => x"70840553",
          2932 => x"0cfc1252",
          2933 => x"718326f2",
          2934 => x"387053ff",
          2935 => x"8e39fc3d",
          2936 => x"0d767079",
          2937 => x"70730783",
          2938 => x"06545454",
          2939 => x"557080c3",
          2940 => x"38717008",
          2941 => x"700970f7",
          2942 => x"fbfdff13",
          2943 => x"0670f884",
          2944 => x"82818006",
          2945 => x"51515353",
          2946 => x"5470a638",
          2947 => x"84147274",
          2948 => x"70840556",
          2949 => x"0c700870",
          2950 => x"0970f7fb",
          2951 => x"fdff1306",
          2952 => x"70f88482",
          2953 => x"81800651",
          2954 => x"51535354",
          2955 => x"70802edc",
          2956 => x"38735271",
          2957 => x"70810553",
          2958 => x"33517073",
          2959 => x"70810555",
          2960 => x"3470f038",
          2961 => x"7481fef0",
          2962 => x"0c863d0d",
          2963 => x"04fd3d0d",
          2964 => x"75707183",
          2965 => x"06535552",
          2966 => x"70b83871",
          2967 => x"70087009",
          2968 => x"f7fbfdff",
          2969 => x"120670f8",
          2970 => x"84828180",
          2971 => x"06515152",
          2972 => x"53709d38",
          2973 => x"84137008",
          2974 => x"7009f7fb",
          2975 => x"fdff1206",
          2976 => x"70f88482",
          2977 => x"81800651",
          2978 => x"51525370",
          2979 => x"802ee538",
          2980 => x"72527133",
          2981 => x"5170802e",
          2982 => x"8a388112",
          2983 => x"70335252",
          2984 => x"70f83871",
          2985 => x"743181fe",
          2986 => x"f00c853d",
          2987 => x"0d04fa3d",
          2988 => x"0d787a7c",
          2989 => x"70545555",
          2990 => x"5272802e",
          2991 => x"80d93871",
          2992 => x"74078306",
          2993 => x"5170802e",
          2994 => x"80d638ff",
          2995 => x"135372ff",
          2996 => x"2eb13871",
          2997 => x"33743356",
          2998 => x"5174712e",
          2999 => x"098106a9",
          3000 => x"3872802e",
          3001 => x"81893870",
          3002 => x"81ff0651",
          3003 => x"70802e80",
          3004 => x"fe388112",
          3005 => x"8115ff15",
          3006 => x"55555272",
          3007 => x"ff2e0981",
          3008 => x"06d13871",
          3009 => x"33743356",
          3010 => x"517081ff",
          3011 => x"067581ff",
          3012 => x"06717131",
          3013 => x"51525270",
          3014 => x"81fef00c",
          3015 => x"883d0d04",
          3016 => x"71745755",
          3017 => x"83732788",
          3018 => x"38710874",
          3019 => x"082e8838",
          3020 => x"74765552",
          3021 => x"ff9539fc",
          3022 => x"13537280",
          3023 => x"2eb13874",
          3024 => x"087009f7",
          3025 => x"fbfdff12",
          3026 => x"0670f884",
          3027 => x"82818006",
          3028 => x"51515170",
          3029 => x"9a388415",
          3030 => x"84175755",
          3031 => x"837327d0",
          3032 => x"38740876",
          3033 => x"082ed038",
          3034 => x"74765552",
          3035 => x"fedd3980",
          3036 => x"0b81fef0",
          3037 => x"0c883d0d",
          3038 => x"04fe3d0d",
          3039 => x"80528353",
          3040 => x"71882b52",
          3041 => x"87863f81",
          3042 => x"fef00881",
          3043 => x"ff067207",
          3044 => x"ff145452",
          3045 => x"728025e8",
          3046 => x"387181fe",
          3047 => x"f00c843d",
          3048 => x"0d04fb3d",
          3049 => x"0d777008",
          3050 => x"70535356",
          3051 => x"71802e80",
          3052 => x"ca387133",
          3053 => x"5170a02e",
          3054 => x"09810686",
          3055 => x"38811252",
          3056 => x"f1397153",
          3057 => x"84398113",
          3058 => x"53807333",
          3059 => x"7081ff06",
          3060 => x"53555570",
          3061 => x"a02e8338",
          3062 => x"81557080",
          3063 => x"2e843874",
          3064 => x"e5387381",
          3065 => x"ff065170",
          3066 => x"a02e0981",
          3067 => x"06883880",
          3068 => x"73708105",
          3069 => x"55347276",
          3070 => x"0c715170",
          3071 => x"81fef00c",
          3072 => x"873d0d04",
          3073 => x"fc3d0d76",
          3074 => x"53720880",
          3075 => x"2e913886",
          3076 => x"3dfc0552",
          3077 => x"72519fd8",
          3078 => x"3f81fef0",
          3079 => x"08853880",
          3080 => x"53833974",
          3081 => x"537281fe",
          3082 => x"f00c863d",
          3083 => x"0d04fc3d",
          3084 => x"0d768211",
          3085 => x"33ff0552",
          3086 => x"53815270",
          3087 => x"8b268198",
          3088 => x"38831333",
          3089 => x"ff055182",
          3090 => x"52709e26",
          3091 => x"818a3884",
          3092 => x"13335183",
          3093 => x"52709726",
          3094 => x"80fe3885",
          3095 => x"13335184",
          3096 => x"5270bb26",
          3097 => x"80f23886",
          3098 => x"13335185",
          3099 => x"5270bb26",
          3100 => x"80e63888",
          3101 => x"13225586",
          3102 => x"527487e7",
          3103 => x"2680d938",
          3104 => x"8a132254",
          3105 => x"87527387",
          3106 => x"e72680cc",
          3107 => x"38810b87",
          3108 => x"c0989c0c",
          3109 => x"722287c0",
          3110 => x"98bc0c82",
          3111 => x"133387c0",
          3112 => x"98b80c83",
          3113 => x"133387c0",
          3114 => x"98b40c84",
          3115 => x"133387c0",
          3116 => x"98b00c85",
          3117 => x"133387c0",
          3118 => x"98ac0c86",
          3119 => x"133387c0",
          3120 => x"98a80c74",
          3121 => x"87c098a4",
          3122 => x"0c7387c0",
          3123 => x"98a00c80",
          3124 => x"0b87c098",
          3125 => x"9c0c8052",
          3126 => x"7181fef0",
          3127 => x"0c863d0d",
          3128 => x"04f33d0d",
          3129 => x"7f5b87c0",
          3130 => x"989c5d81",
          3131 => x"7d0c87c0",
          3132 => x"98bc085e",
          3133 => x"7d7b2387",
          3134 => x"c098b808",
          3135 => x"5a79821c",
          3136 => x"3487c098",
          3137 => x"b4085a79",
          3138 => x"831c3487",
          3139 => x"c098b008",
          3140 => x"5a79841c",
          3141 => x"3487c098",
          3142 => x"ac085a79",
          3143 => x"851c3487",
          3144 => x"c098a808",
          3145 => x"5a79861c",
          3146 => x"3487c098",
          3147 => x"a4085c7b",
          3148 => x"881c2387",
          3149 => x"c098a008",
          3150 => x"5a798a1c",
          3151 => x"23807d0c",
          3152 => x"7983ffff",
          3153 => x"06597b83",
          3154 => x"ffff0658",
          3155 => x"861b3357",
          3156 => x"851b3356",
          3157 => x"841b3355",
          3158 => x"831b3354",
          3159 => x"821b3353",
          3160 => x"7d83ffff",
          3161 => x"065281e2",
          3162 => x"d451999d",
          3163 => x"3f8f3d0d",
          3164 => x"04ff3d0d",
          3165 => x"028f0533",
          3166 => x"7030709f",
          3167 => x"2a515252",
          3168 => x"700b0b81",
          3169 => x"f9e83483",
          3170 => x"3d0d04fb",
          3171 => x"3d0d770b",
          3172 => x"0b81f9e8",
          3173 => x"337081ff",
          3174 => x"06575556",
          3175 => x"87c09484",
          3176 => x"5174802e",
          3177 => x"863887c0",
          3178 => x"94945170",
          3179 => x"0870962a",
          3180 => x"70810653",
          3181 => x"54527080",
          3182 => x"2e8c3871",
          3183 => x"912a7081",
          3184 => x"06515170",
          3185 => x"d7387281",
          3186 => x"32708106",
          3187 => x"51517080",
          3188 => x"2e8d3871",
          3189 => x"932a7081",
          3190 => x"06515170",
          3191 => x"ffbe3873",
          3192 => x"81ff0651",
          3193 => x"87c09480",
          3194 => x"5270802e",
          3195 => x"863887c0",
          3196 => x"94905275",
          3197 => x"720c7581",
          3198 => x"fef00c87",
          3199 => x"3d0d04fb",
          3200 => x"3d0d029f",
          3201 => x"05330b0b",
          3202 => x"81f9e833",
          3203 => x"7081ff06",
          3204 => x"57555687",
          3205 => x"c0948451",
          3206 => x"74802e86",
          3207 => x"3887c094",
          3208 => x"94517008",
          3209 => x"70962a70",
          3210 => x"81065354",
          3211 => x"5270802e",
          3212 => x"8c387191",
          3213 => x"2a708106",
          3214 => x"515170d7",
          3215 => x"38728132",
          3216 => x"70810651",
          3217 => x"5170802e",
          3218 => x"8d387193",
          3219 => x"2a708106",
          3220 => x"515170ff",
          3221 => x"be387381",
          3222 => x"ff065187",
          3223 => x"c0948052",
          3224 => x"70802e86",
          3225 => x"3887c094",
          3226 => x"90527572",
          3227 => x"0c873d0d",
          3228 => x"04f93d0d",
          3229 => x"79548074",
          3230 => x"337081ff",
          3231 => x"06535357",
          3232 => x"70772e80",
          3233 => x"fe387181",
          3234 => x"ff068115",
          3235 => x"0b0b81f9",
          3236 => x"e8337081",
          3237 => x"ff065957",
          3238 => x"555887c0",
          3239 => x"94845175",
          3240 => x"802e8638",
          3241 => x"87c09494",
          3242 => x"51700870",
          3243 => x"962a7081",
          3244 => x"06535452",
          3245 => x"70802e8c",
          3246 => x"3871912a",
          3247 => x"70810651",
          3248 => x"5170d738",
          3249 => x"72813270",
          3250 => x"81065151",
          3251 => x"70802e8d",
          3252 => x"3871932a",
          3253 => x"70810651",
          3254 => x"5170ffbe",
          3255 => x"387481ff",
          3256 => x"065187c0",
          3257 => x"94805270",
          3258 => x"802e8638",
          3259 => x"87c09490",
          3260 => x"5277720c",
          3261 => x"81177433",
          3262 => x"7081ff06",
          3263 => x"53535770",
          3264 => x"ff843876",
          3265 => x"81fef00c",
          3266 => x"893d0d04",
          3267 => x"fe3d0d0b",
          3268 => x"0b81f9e8",
          3269 => x"337081ff",
          3270 => x"06545287",
          3271 => x"c0948451",
          3272 => x"72802e86",
          3273 => x"3887c094",
          3274 => x"94517008",
          3275 => x"70822a70",
          3276 => x"81065151",
          3277 => x"5170802e",
          3278 => x"e2387181",
          3279 => x"ff065187",
          3280 => x"c0948052",
          3281 => x"70802e86",
          3282 => x"3887c094",
          3283 => x"90527108",
          3284 => x"7081ff06",
          3285 => x"81fef00c",
          3286 => x"51843d0d",
          3287 => x"04fe3d0d",
          3288 => x"0b0b81f9",
          3289 => x"e8337081",
          3290 => x"ff065253",
          3291 => x"87c09484",
          3292 => x"5270802e",
          3293 => x"863887c0",
          3294 => x"94945271",
          3295 => x"0870822a",
          3296 => x"70810651",
          3297 => x"5151ff52",
          3298 => x"70802ea0",
          3299 => x"387281ff",
          3300 => x"065187c0",
          3301 => x"94805270",
          3302 => x"802e8638",
          3303 => x"87c09490",
          3304 => x"52710870",
          3305 => x"982b7098",
          3306 => x"2c515351",
          3307 => x"7181fef0",
          3308 => x"0c843d0d",
          3309 => x"04ff3d0d",
          3310 => x"87c09e80",
          3311 => x"08709c2a",
          3312 => x"8a065151",
          3313 => x"70802e84",
          3314 => x"b43887c0",
          3315 => x"9ea40881",
          3316 => x"f9ec0c87",
          3317 => x"c09ea808",
          3318 => x"81f9f00c",
          3319 => x"87c09e94",
          3320 => x"0881f9f4",
          3321 => x"0c87c09e",
          3322 => x"980881f9",
          3323 => x"f80c87c0",
          3324 => x"9e9c0881",
          3325 => x"f9fc0c87",
          3326 => x"c09ea008",
          3327 => x"81fa800c",
          3328 => x"87c09eac",
          3329 => x"0881fa84",
          3330 => x"0c87c09e",
          3331 => x"b00881fa",
          3332 => x"880c87c0",
          3333 => x"9eb40881",
          3334 => x"fa8c0c87",
          3335 => x"c09eb808",
          3336 => x"81fa900c",
          3337 => x"87c09ebc",
          3338 => x"0881fa94",
          3339 => x"0c87c09e",
          3340 => x"c00881fa",
          3341 => x"980c87c0",
          3342 => x"9ec40881",
          3343 => x"fa9c0c87",
          3344 => x"c09e8008",
          3345 => x"517081fa",
          3346 => x"a02387c0",
          3347 => x"9e840881",
          3348 => x"faa40c87",
          3349 => x"c09e8808",
          3350 => x"81faa80c",
          3351 => x"87c09e8c",
          3352 => x"0881faac",
          3353 => x"0c810b81",
          3354 => x"fab03480",
          3355 => x"0b87c09e",
          3356 => x"90087084",
          3357 => x"800a0651",
          3358 => x"52527080",
          3359 => x"2e833881",
          3360 => x"527181fa",
          3361 => x"b134800b",
          3362 => x"87c09e90",
          3363 => x"08708880",
          3364 => x"0a065152",
          3365 => x"5270802e",
          3366 => x"83388152",
          3367 => x"7181fab2",
          3368 => x"34800b87",
          3369 => x"c09e9008",
          3370 => x"7090800a",
          3371 => x"06515252",
          3372 => x"70802e83",
          3373 => x"38815271",
          3374 => x"81fab334",
          3375 => x"800b87c0",
          3376 => x"9e900870",
          3377 => x"88808006",
          3378 => x"51525270",
          3379 => x"802e8338",
          3380 => x"81527181",
          3381 => x"fab43480",
          3382 => x"0b87c09e",
          3383 => x"900870a0",
          3384 => x"80800651",
          3385 => x"52527080",
          3386 => x"2e833881",
          3387 => x"527181fa",
          3388 => x"b534800b",
          3389 => x"87c09e90",
          3390 => x"08709080",
          3391 => x"80065152",
          3392 => x"5270802e",
          3393 => x"83388152",
          3394 => x"7181fab6",
          3395 => x"34800b87",
          3396 => x"c09e9008",
          3397 => x"70848080",
          3398 => x"06515252",
          3399 => x"70802e83",
          3400 => x"38815271",
          3401 => x"81fab734",
          3402 => x"800b87c0",
          3403 => x"9e900870",
          3404 => x"82808006",
          3405 => x"51525270",
          3406 => x"802e8338",
          3407 => x"81527181",
          3408 => x"fab83480",
          3409 => x"0b87c09e",
          3410 => x"90087081",
          3411 => x"80800651",
          3412 => x"52527080",
          3413 => x"2e833881",
          3414 => x"527181fa",
          3415 => x"b934800b",
          3416 => x"87c09e90",
          3417 => x"087080c0",
          3418 => x"80065152",
          3419 => x"5270802e",
          3420 => x"83388152",
          3421 => x"7181faba",
          3422 => x"34800b87",
          3423 => x"c09e9008",
          3424 => x"70a08006",
          3425 => x"51525270",
          3426 => x"802e8338",
          3427 => x"81527181",
          3428 => x"fabb3487",
          3429 => x"c09e9008",
          3430 => x"70988006",
          3431 => x"708a2a51",
          3432 => x"51517081",
          3433 => x"fabc3480",
          3434 => x"0b87c09e",
          3435 => x"90087084",
          3436 => x"80065152",
          3437 => x"5270802e",
          3438 => x"83388152",
          3439 => x"7181fabd",
          3440 => x"3487c09e",
          3441 => x"90087083",
          3442 => x"f0067084",
          3443 => x"2a515151",
          3444 => x"7081fabe",
          3445 => x"34800b87",
          3446 => x"c09e9008",
          3447 => x"70880651",
          3448 => x"52527080",
          3449 => x"2e833881",
          3450 => x"527181fa",
          3451 => x"bf3487c0",
          3452 => x"9e900870",
          3453 => x"87065151",
          3454 => x"7081fac0",
          3455 => x"34833d0d",
          3456 => x"04fb3d0d",
          3457 => x"81e2ec51",
          3458 => x"8a9b3f81",
          3459 => x"fab03354",
          3460 => x"73802e88",
          3461 => x"3881e380",
          3462 => x"518a8a3f",
          3463 => x"81e39451",
          3464 => x"8a833f81",
          3465 => x"fab23354",
          3466 => x"73802e93",
          3467 => x"3881fa8c",
          3468 => x"0881fa90",
          3469 => x"08115452",
          3470 => x"81e3ac51",
          3471 => x"8fcb3f81",
          3472 => x"fab73354",
          3473 => x"73802e93",
          3474 => x"3881fa84",
          3475 => x"0881fa88",
          3476 => x"08115452",
          3477 => x"81e3c851",
          3478 => x"8faf3f81",
          3479 => x"fab43354",
          3480 => x"73802e93",
          3481 => x"3881f9ec",
          3482 => x"0881f9f0",
          3483 => x"08115452",
          3484 => x"81e3e451",
          3485 => x"8f933f81",
          3486 => x"fab53354",
          3487 => x"73802e93",
          3488 => x"3881f9f4",
          3489 => x"0881f9f8",
          3490 => x"08115452",
          3491 => x"81e48051",
          3492 => x"8ef73f81",
          3493 => x"fab63354",
          3494 => x"73802e93",
          3495 => x"3881f9fc",
          3496 => x"0881fa80",
          3497 => x"08115452",
          3498 => x"81e49c51",
          3499 => x"8edb3f81",
          3500 => x"fabb3354",
          3501 => x"73802e8d",
          3502 => x"3881fabc",
          3503 => x"335281e4",
          3504 => x"b8518ec5",
          3505 => x"3f81fabf",
          3506 => x"33547380",
          3507 => x"2e8d3881",
          3508 => x"fac03352",
          3509 => x"81e4d851",
          3510 => x"8eaf3f81",
          3511 => x"fabd3354",
          3512 => x"73802e8d",
          3513 => x"3881fabe",
          3514 => x"335281e4",
          3515 => x"f8518e99",
          3516 => x"3f81fab1",
          3517 => x"33547380",
          3518 => x"2e883881",
          3519 => x"e5985188",
          3520 => x"a43f81fa",
          3521 => x"b3335473",
          3522 => x"802e8838",
          3523 => x"81e5ac51",
          3524 => x"88933f81",
          3525 => x"fab83354",
          3526 => x"73802e88",
          3527 => x"3881e5b8",
          3528 => x"5188823f",
          3529 => x"81fab933",
          3530 => x"5473802e",
          3531 => x"883881e5",
          3532 => x"c45187f1",
          3533 => x"3f81faba",
          3534 => x"33547380",
          3535 => x"2e883881",
          3536 => x"e5d05187",
          3537 => x"e03f81e5",
          3538 => x"dc5187d9",
          3539 => x"3f81fa94",
          3540 => x"085281e5",
          3541 => x"e8518db1",
          3542 => x"3f81fa98",
          3543 => x"085281e6",
          3544 => x"90518da5",
          3545 => x"3f81fa9c",
          3546 => x"085281e6",
          3547 => x"b8518d99",
          3548 => x"3f81e6e0",
          3549 => x"5187ae3f",
          3550 => x"81faa022",
          3551 => x"5281e6e8",
          3552 => x"518d863f",
          3553 => x"81faa408",
          3554 => x"56bd84c0",
          3555 => x"527551e4",
          3556 => x"9a3f81fe",
          3557 => x"f008bd84",
          3558 => x"c0297671",
          3559 => x"31545481",
          3560 => x"fef00852",
          3561 => x"81e79051",
          3562 => x"8cdf3f81",
          3563 => x"fab73354",
          3564 => x"73802ea8",
          3565 => x"3881faa8",
          3566 => x"0856bd84",
          3567 => x"c0527551",
          3568 => x"e3e93f81",
          3569 => x"fef008bd",
          3570 => x"84c02976",
          3571 => x"71315454",
          3572 => x"81fef008",
          3573 => x"5281e7bc",
          3574 => x"518cae3f",
          3575 => x"81fab233",
          3576 => x"5473802e",
          3577 => x"a83881fa",
          3578 => x"ac0856bd",
          3579 => x"84c05275",
          3580 => x"51e3b83f",
          3581 => x"81fef008",
          3582 => x"bd84c029",
          3583 => x"76713154",
          3584 => x"5481fef0",
          3585 => x"085281e7",
          3586 => x"e8518bfd",
          3587 => x"3f81f5e4",
          3588 => x"5186923f",
          3589 => x"873d0d04",
          3590 => x"fe3d0d02",
          3591 => x"920533ff",
          3592 => x"05527184",
          3593 => x"26aa3871",
          3594 => x"842981e1",
          3595 => x"c0055271",
          3596 => x"080481e8",
          3597 => x"94519d39",
          3598 => x"81e89c51",
          3599 => x"973981e8",
          3600 => x"a4519139",
          3601 => x"81e8ac51",
          3602 => x"8b3981e8",
          3603 => x"b0518539",
          3604 => x"81e8b851",
          3605 => x"85cf3f84",
          3606 => x"3d0d0471",
          3607 => x"88800c04",
          3608 => x"ff3d0d87",
          3609 => x"c0968470",
          3610 => x"08525280",
          3611 => x"720c7074",
          3612 => x"077081fa",
          3613 => x"c40c720c",
          3614 => x"833d0d04",
          3615 => x"ff3d0d87",
          3616 => x"c0968470",
          3617 => x"0881fac4",
          3618 => x"0c528072",
          3619 => x"0c730970",
          3620 => x"81fac408",
          3621 => x"067081fa",
          3622 => x"c40c730c",
          3623 => x"51833d0d",
          3624 => x"04800b87",
          3625 => x"c096840c",
          3626 => x"0481fac4",
          3627 => x"0887c096",
          3628 => x"840c04fe",
          3629 => x"3d0d81ff",
          3630 => x"80088938",
          3631 => x"8296b00b",
          3632 => x"81ff800c",
          3633 => x"81ff8008",
          3634 => x"75115252",
          3635 => x"ff537083",
          3636 => x"b7f82688",
          3637 => x"387081ff",
          3638 => x"800c7153",
          3639 => x"7281fef0",
          3640 => x"0c843d0d",
          3641 => x"04f93d0d",
          3642 => x"797b8412",
          3643 => x"08a01290",
          3644 => x"14089415",
          3645 => x"0890165e",
          3646 => x"5a585459",
          3647 => x"57537077",
          3648 => x"26ba3875",
          3649 => x"13881408",
          3650 => x"53518171",
          3651 => x"0c767631",
          3652 => x"84120c80",
          3653 => x"730c7584",
          3654 => x"140c728c",
          3655 => x"120c7188",
          3656 => x"120c708c",
          3657 => x"130c7088",
          3658 => x"140c7390",
          3659 => x"120c7494",
          3660 => x"120c7094",
          3661 => x"150c7090",
          3662 => x"160c8c39",
          3663 => x"80730c73",
          3664 => x"90160c74",
          3665 => x"94150c77",
          3666 => x"81fef00c",
          3667 => x"893d0d04",
          3668 => x"fc3d0d76",
          3669 => x"8c110888",
          3670 => x"12085653",
          3671 => x"53710881",
          3672 => x"2e098106",
          3673 => x"a3388412",
          3674 => x"08701352",
          3675 => x"5570732e",
          3676 => x"09810694",
          3677 => x"38841308",
          3678 => x"1584130c",
          3679 => x"7388130c",
          3680 => x"718c150c",
          3681 => x"71539f39",
          3682 => x"81730c81",
          3683 => x"fad80890",
          3684 => x"140c81fa",
          3685 => x"c80b9414",
          3686 => x"0c7281fa",
          3687 => x"d80c9013",
          3688 => x"08739412",
          3689 => x"0c517308",
          3690 => x"812e0981",
          3691 => x"06b33884",
          3692 => x"13087014",
          3693 => x"52527074",
          3694 => x"2e098106",
          3695 => x"a4388414",
          3696 => x"08128414",
          3697 => x"0c941408",
          3698 => x"90150870",
          3699 => x"90130c52",
          3700 => x"94120c8c",
          3701 => x"14088815",
          3702 => x"08708813",
          3703 => x"0c528c12",
          3704 => x"0c7281fe",
          3705 => x"f00c863d",
          3706 => x"0d04f93d",
          3707 => x"0d797055",
          3708 => x"5776802e",
          3709 => x"81b5389f",
          3710 => x"17f00681",
          3711 => x"fad80857",
          3712 => x"57750882",
          3713 => x"2e8f3884",
          3714 => x"16087727",
          3715 => x"80c73890",
          3716 => x"160856ed",
          3717 => x"3983ffff",
          3718 => x"17fc8080",
          3719 => x"06705258",
          3720 => x"fd913f81",
          3721 => x"fef00881",
          3722 => x"fef00830",
          3723 => x"7081fef0",
          3724 => x"08078025",
          3725 => x"81fef008",
          3726 => x"09703070",
          3727 => x"72078025",
          3728 => x"73075358",
          3729 => x"58515456",
          3730 => x"80547274",
          3731 => x"2e098106",
          3732 => x"80d93888",
          3733 => x"39765275",
          3734 => x"5180c839",
          3735 => x"810b81fe",
          3736 => x"f0080c77",
          3737 => x"81fef008",
          3738 => x"84050c81",
          3739 => x"fad40853",
          3740 => x"7208822e",
          3741 => x"8c387573",
          3742 => x"2687388c",
          3743 => x"130853f0",
          3744 => x"39881308",
          3745 => x"88170c72",
          3746 => x"8c170c75",
          3747 => x"88140c88",
          3748 => x"1608768c",
          3749 => x"120c5375",
          3750 => x"51fdb53f",
          3751 => x"765281fe",
          3752 => x"f00851fc",
          3753 => x"c03f81fe",
          3754 => x"f0085473",
          3755 => x"81fef00c",
          3756 => x"893d0d04",
          3757 => x"ff3d0d73",
          3758 => x"5271802e",
          3759 => x"8738f012",
          3760 => x"51fd8d3f",
          3761 => x"833d0d04",
          3762 => x"fe3d0d02",
          3763 => x"93053353",
          3764 => x"728a2e09",
          3765 => x"81068538",
          3766 => x"8d51ed3f",
          3767 => x"81ff8c08",
          3768 => x"5271802e",
          3769 => x"90387272",
          3770 => x"3481ff8c",
          3771 => x"08810581",
          3772 => x"ff8c0c8f",
          3773 => x"3981ff84",
          3774 => x"08527180",
          3775 => x"2e853872",
          3776 => x"51712d84",
          3777 => x"3d0d04fe",
          3778 => x"3d0d0297",
          3779 => x"053381ff",
          3780 => x"84087681",
          3781 => x"ff840c54",
          3782 => x"51ffad3f",
          3783 => x"7281ff84",
          3784 => x"0c843d0d",
          3785 => x"04fd3d0d",
          3786 => x"75547333",
          3787 => x"7081ff06",
          3788 => x"53537180",
          3789 => x"2e8e3872",
          3790 => x"81ff0651",
          3791 => x"811454ff",
          3792 => x"873fe739",
          3793 => x"853d0d04",
          3794 => x"fc3d0d77",
          3795 => x"81ff8408",
          3796 => x"7881ff84",
          3797 => x"0c565473",
          3798 => x"337081ff",
          3799 => x"06535371",
          3800 => x"802e8e38",
          3801 => x"7281ff06",
          3802 => x"51811454",
          3803 => x"feda3fe7",
          3804 => x"397481ff",
          3805 => x"840c863d",
          3806 => x"0d04ec3d",
          3807 => x"0d666859",
          3808 => x"59787081",
          3809 => x"055a3356",
          3810 => x"75802e84",
          3811 => x"f83875a5",
          3812 => x"2e098106",
          3813 => x"82de3880",
          3814 => x"707a7081",
          3815 => x"055c3358",
          3816 => x"5b5b75b0",
          3817 => x"2e098106",
          3818 => x"8538815a",
          3819 => x"8b3975ad",
          3820 => x"2e098106",
          3821 => x"8a38825a",
          3822 => x"78708105",
          3823 => x"5a335675",
          3824 => x"aa2e0981",
          3825 => x"06923877",
          3826 => x"84197108",
          3827 => x"7b708105",
          3828 => x"5d33595d",
          3829 => x"59539d39",
          3830 => x"d0165372",
          3831 => x"89269538",
          3832 => x"7a88297b",
          3833 => x"10057605",
          3834 => x"d0057970",
          3835 => x"81055b33",
          3836 => x"575be539",
          3837 => x"7580ec32",
          3838 => x"70307072",
          3839 => x"07802578",
          3840 => x"80cc3270",
          3841 => x"30707207",
          3842 => x"80257307",
          3843 => x"53545851",
          3844 => x"55537380",
          3845 => x"2e8c3879",
          3846 => x"84077970",
          3847 => x"81055b33",
          3848 => x"575a7580",
          3849 => x"2e83de38",
          3850 => x"755480e0",
          3851 => x"76278938",
          3852 => x"e0167081",
          3853 => x"ff065553",
          3854 => x"7380cf2e",
          3855 => x"81aa3873",
          3856 => x"80cf24a2",
          3857 => x"387380c3",
          3858 => x"2e818e38",
          3859 => x"7380c324",
          3860 => x"8b387380",
          3861 => x"c22e818c",
          3862 => x"38819939",
          3863 => x"7380c42e",
          3864 => x"818a3881",
          3865 => x"8f397380",
          3866 => x"d52e8180",
          3867 => x"387380d5",
          3868 => x"248a3873",
          3869 => x"80d32e8e",
          3870 => x"3880f939",
          3871 => x"7380d82e",
          3872 => x"80ee3880",
          3873 => x"ef397784",
          3874 => x"19710856",
          3875 => x"59538074",
          3876 => x"33545572",
          3877 => x"752e8d38",
          3878 => x"81157015",
          3879 => x"70335154",
          3880 => x"5572f538",
          3881 => x"79812a56",
          3882 => x"90397481",
          3883 => x"16565372",
          3884 => x"7b278f38",
          3885 => x"a051fc90",
          3886 => x"3f758106",
          3887 => x"5372802e",
          3888 => x"e9387351",
          3889 => x"fcdf3f74",
          3890 => x"81165653",
          3891 => x"727b27fd",
          3892 => x"b038a051",
          3893 => x"fbf23fef",
          3894 => x"39778419",
          3895 => x"83123353",
          3896 => x"59539339",
          3897 => x"825c9539",
          3898 => x"885c9139",
          3899 => x"8a5c8d39",
          3900 => x"905c8939",
          3901 => x"7551fbd0",
          3902 => x"3ffd8639",
          3903 => x"79822a70",
          3904 => x"81065153",
          3905 => x"72802e88",
          3906 => x"38778419",
          3907 => x"59538639",
          3908 => x"84187854",
          3909 => x"58720874",
          3910 => x"80c43270",
          3911 => x"30707207",
          3912 => x"80255155",
          3913 => x"55557480",
          3914 => x"258d3872",
          3915 => x"802e8838",
          3916 => x"74307a90",
          3917 => x"075b5580",
          3918 => x"0b8f3d5e",
          3919 => x"577b5274",
          3920 => x"51d99b3f",
          3921 => x"81fef008",
          3922 => x"81ff067c",
          3923 => x"53755254",
          3924 => x"d8d93f81",
          3925 => x"fef00855",
          3926 => x"89742792",
          3927 => x"38a71453",
          3928 => x"7580f82e",
          3929 => x"84388714",
          3930 => x"537281ff",
          3931 => x"0654b014",
          3932 => x"53727d70",
          3933 => x"81055f34",
          3934 => x"81177530",
          3935 => x"7077079f",
          3936 => x"2a515457",
          3937 => x"769f2685",
          3938 => x"3872ffb1",
          3939 => x"3879842a",
          3940 => x"70810651",
          3941 => x"5372802e",
          3942 => x"8e38963d",
          3943 => x"7705e005",
          3944 => x"53ad7334",
          3945 => x"81175776",
          3946 => x"7a810654",
          3947 => x"55b05472",
          3948 => x"8338a054",
          3949 => x"79812a70",
          3950 => x"81065456",
          3951 => x"729f3881",
          3952 => x"1755767b",
          3953 => x"27973873",
          3954 => x"51f9fd3f",
          3955 => x"75810653",
          3956 => x"728b3874",
          3957 => x"81165653",
          3958 => x"7a7326eb",
          3959 => x"38963d77",
          3960 => x"05e00553",
          3961 => x"ff17ff14",
          3962 => x"70335354",
          3963 => x"57f9d93f",
          3964 => x"76f23874",
          3965 => x"81165653",
          3966 => x"727b27fb",
          3967 => x"8438a051",
          3968 => x"f9c63fef",
          3969 => x"39963d0d",
          3970 => x"04fd3d0d",
          3971 => x"863d7070",
          3972 => x"84055208",
          3973 => x"55527351",
          3974 => x"fae03f85",
          3975 => x"3d0d04fe",
          3976 => x"3d0d7481",
          3977 => x"ff8c0c85",
          3978 => x"3d880552",
          3979 => x"7551faca",
          3980 => x"3f81ff8c",
          3981 => x"08538073",
          3982 => x"34800b81",
          3983 => x"ff8c0c84",
          3984 => x"3d0d04fd",
          3985 => x"3d0d81ff",
          3986 => x"84087681",
          3987 => x"ff840c87",
          3988 => x"3d880553",
          3989 => x"775253fa",
          3990 => x"a13f7281",
          3991 => x"ff840c85",
          3992 => x"3d0d04fb",
          3993 => x"3d0d7779",
          3994 => x"81ff8808",
          3995 => x"70565457",
          3996 => x"55805471",
          3997 => x"802e80e0",
          3998 => x"3881ff88",
          3999 => x"0852712d",
          4000 => x"81fef008",
          4001 => x"81ff0653",
          4002 => x"72802e80",
          4003 => x"cb38728d",
          4004 => x"2eb93872",
          4005 => x"88327030",
          4006 => x"70802551",
          4007 => x"51527380",
          4008 => x"2e8b3871",
          4009 => x"802e8638",
          4010 => x"ff145497",
          4011 => x"399f7325",
          4012 => x"c838ff16",
          4013 => x"52737225",
          4014 => x"c0387414",
          4015 => x"52727234",
          4016 => x"81145472",
          4017 => x"51f8813f",
          4018 => x"ffaf3973",
          4019 => x"15528072",
          4020 => x"348a51f7",
          4021 => x"f33f8153",
          4022 => x"7281fef0",
          4023 => x"0c873d0d",
          4024 => x"04fe3d0d",
          4025 => x"81ff8808",
          4026 => x"7581ff88",
          4027 => x"0c775376",
          4028 => x"5253feef",
          4029 => x"3f7281ff",
          4030 => x"880c843d",
          4031 => x"0d04f83d",
          4032 => x"0d7a7c5a",
          4033 => x"5680707a",
          4034 => x"0c587508",
          4035 => x"70335553",
          4036 => x"73a02e09",
          4037 => x"81068738",
          4038 => x"8113760c",
          4039 => x"ed3973ad",
          4040 => x"2e098106",
          4041 => x"8e388176",
          4042 => x"0811770c",
          4043 => x"76087033",
          4044 => x"56545873",
          4045 => x"b02e0981",
          4046 => x"0680c238",
          4047 => x"75088105",
          4048 => x"760c7508",
          4049 => x"70335553",
          4050 => x"7380e22e",
          4051 => x"8b389057",
          4052 => x"7380f82e",
          4053 => x"85388f39",
          4054 => x"82578113",
          4055 => x"760c7508",
          4056 => x"70335553",
          4057 => x"ac398155",
          4058 => x"a0742780",
          4059 => x"fa38d014",
          4060 => x"53805588",
          4061 => x"57897327",
          4062 => x"983880eb",
          4063 => x"39d01453",
          4064 => x"80557289",
          4065 => x"2680e038",
          4066 => x"86398055",
          4067 => x"80d9398a",
          4068 => x"578055a0",
          4069 => x"742780c2",
          4070 => x"3880e074",
          4071 => x"278938e0",
          4072 => x"147081ff",
          4073 => x"065553d0",
          4074 => x"147081ff",
          4075 => x"06555390",
          4076 => x"74278e38",
          4077 => x"f9147081",
          4078 => x"ff065553",
          4079 => x"897427ca",
          4080 => x"38737727",
          4081 => x"c5387477",
          4082 => x"29147608",
          4083 => x"8105770c",
          4084 => x"76087033",
          4085 => x"565455ff",
          4086 => x"ba397780",
          4087 => x"2e843874",
          4088 => x"30557479",
          4089 => x"0c815574",
          4090 => x"81fef00c",
          4091 => x"8a3d0d04",
          4092 => x"f83d0d7a",
          4093 => x"7c5a5680",
          4094 => x"707a0c58",
          4095 => x"75087033",
          4096 => x"555373a0",
          4097 => x"2e098106",
          4098 => x"87388113",
          4099 => x"760ced39",
          4100 => x"73ad2e09",
          4101 => x"81068e38",
          4102 => x"81760811",
          4103 => x"770c7608",
          4104 => x"70335654",
          4105 => x"5873b02e",
          4106 => x"09810680",
          4107 => x"c2387508",
          4108 => x"8105760c",
          4109 => x"75087033",
          4110 => x"55537380",
          4111 => x"e22e8b38",
          4112 => x"90577380",
          4113 => x"f82e8538",
          4114 => x"8f398257",
          4115 => x"8113760c",
          4116 => x"75087033",
          4117 => x"5553ac39",
          4118 => x"8155a074",
          4119 => x"2780fa38",
          4120 => x"d0145380",
          4121 => x"55885789",
          4122 => x"73279838",
          4123 => x"80eb39d0",
          4124 => x"14538055",
          4125 => x"72892680",
          4126 => x"e0388639",
          4127 => x"805580d9",
          4128 => x"398a5780",
          4129 => x"55a07427",
          4130 => x"80c23880",
          4131 => x"e0742789",
          4132 => x"38e01470",
          4133 => x"81ff0655",
          4134 => x"53d01470",
          4135 => x"81ff0655",
          4136 => x"53907427",
          4137 => x"8e38f914",
          4138 => x"7081ff06",
          4139 => x"55538974",
          4140 => x"27ca3873",
          4141 => x"7727c538",
          4142 => x"74772914",
          4143 => x"76088105",
          4144 => x"770c7608",
          4145 => x"70335654",
          4146 => x"55ffba39",
          4147 => x"77802e84",
          4148 => x"38743055",
          4149 => x"74790c81",
          4150 => x"557481fe",
          4151 => x"f00c8a3d",
          4152 => x"0d04fd3d",
          4153 => x"0d76982b",
          4154 => x"70982c79",
          4155 => x"982b7098",
          4156 => x"2c721013",
          4157 => x"70822b51",
          4158 => x"53515451",
          4159 => x"51800b81",
          4160 => x"e9cc1233",
          4161 => x"55537174",
          4162 => x"259c3881",
          4163 => x"e9c81108",
          4164 => x"12028405",
          4165 => x"97053371",
          4166 => x"33525252",
          4167 => x"70722e09",
          4168 => x"81068338",
          4169 => x"81537281",
          4170 => x"fef00c85",
          4171 => x"3d0d04fc",
          4172 => x"3d0d7802",
          4173 => x"84059f05",
          4174 => x"33713354",
          4175 => x"55537180",
          4176 => x"2e9f3888",
          4177 => x"51f3813f",
          4178 => x"a051f2fc",
          4179 => x"3f8851f2",
          4180 => x"f73f7233",
          4181 => x"ff055271",
          4182 => x"73347181",
          4183 => x"ff0652de",
          4184 => x"397651f3",
          4185 => x"c03f7373",
          4186 => x"34863d0d",
          4187 => x"04f63d0d",
          4188 => x"7c028405",
          4189 => x"b7053302",
          4190 => x"8805bb05",
          4191 => x"3381fbbc",
          4192 => x"33708429",
          4193 => x"81fae405",
          4194 => x"70085159",
          4195 => x"595a5859",
          4196 => x"74802e86",
          4197 => x"387451f2",
          4198 => x"9b3f81fb",
          4199 => x"bc337084",
          4200 => x"2981fae4",
          4201 => x"05811970",
          4202 => x"5458565a",
          4203 => x"f0bc3f81",
          4204 => x"fef00875",
          4205 => x"0c81fbbc",
          4206 => x"33708429",
          4207 => x"81fae405",
          4208 => x"70085156",
          4209 => x"5a74802e",
          4210 => x"a6387553",
          4211 => x"78527451",
          4212 => x"d5e03f81",
          4213 => x"fbbc3381",
          4214 => x"05557481",
          4215 => x"fbbc3474",
          4216 => x"81ff0655",
          4217 => x"93752787",
          4218 => x"38800b81",
          4219 => x"fbbc3477",
          4220 => x"802eb638",
          4221 => x"81fbb808",
          4222 => x"5675802e",
          4223 => x"ac3881fb",
          4224 => x"b4335574",
          4225 => x"a4388c3d",
          4226 => x"fc055476",
          4227 => x"53785275",
          4228 => x"5180c891",
          4229 => x"3f81fbb8",
          4230 => x"08528a51",
          4231 => x"80fd9e3f",
          4232 => x"81fbb808",
          4233 => x"5180cbee",
          4234 => x"3f8c3d0d",
          4235 => x"04dc3d0d",
          4236 => x"81578052",
          4237 => x"81fbb808",
          4238 => x"5180d287",
          4239 => x"3f81fef0",
          4240 => x"0880d138",
          4241 => x"81fbb808",
          4242 => x"5380f852",
          4243 => x"883d7052",
          4244 => x"5680fad5",
          4245 => x"3f81fef0",
          4246 => x"08802eb8",
          4247 => x"387551d7",
          4248 => x"ec3f81fe",
          4249 => x"f0085580",
          4250 => x"0b81fef0",
          4251 => x"08259c38",
          4252 => x"81fef008",
          4253 => x"ff057017",
          4254 => x"55558074",
          4255 => x"34755376",
          4256 => x"52811781",
          4257 => x"e8e05257",
          4258 => x"f6ff3f74",
          4259 => x"ff2e0981",
          4260 => x"06ffb138",
          4261 => x"a63d0d04",
          4262 => x"d93d0daa",
          4263 => x"3d08ad3d",
          4264 => x"085a5a81",
          4265 => x"70585880",
          4266 => x"5281fbb8",
          4267 => x"085180d1",
          4268 => x"923f81fe",
          4269 => x"f0088191",
          4270 => x"38ff0b81",
          4271 => x"fbb80854",
          4272 => x"5580f852",
          4273 => x"8b3d7052",
          4274 => x"5680f9dd",
          4275 => x"3f81fef0",
          4276 => x"08802ea4",
          4277 => x"387551d6",
          4278 => x"f43f81fe",
          4279 => x"f0088118",
          4280 => x"5855800b",
          4281 => x"81fef008",
          4282 => x"258e3881",
          4283 => x"fef008ff",
          4284 => x"05701755",
          4285 => x"55807434",
          4286 => x"74097030",
          4287 => x"7072079f",
          4288 => x"2a515555",
          4289 => x"78772e85",
          4290 => x"3873ffad",
          4291 => x"3881fbb8",
          4292 => x"088c1108",
          4293 => x"535180d0",
          4294 => x"aa3f81fe",
          4295 => x"f008802e",
          4296 => x"883881e8",
          4297 => x"ec51effd",
          4298 => x"3f78772e",
          4299 => x"09810699",
          4300 => x"38755279",
          4301 => x"51d5a73f",
          4302 => x"7951d691",
          4303 => x"3fab3d08",
          4304 => x"5481fef0",
          4305 => x"08743480",
          4306 => x"587781fe",
          4307 => x"f00ca93d",
          4308 => x"0d04f63d",
          4309 => x"0d7c7e71",
          4310 => x"5c717233",
          4311 => x"57595a58",
          4312 => x"73a02e09",
          4313 => x"8106a238",
          4314 => x"78337805",
          4315 => x"56777627",
          4316 => x"98388117",
          4317 => x"705b7071",
          4318 => x"33565855",
          4319 => x"73a02e09",
          4320 => x"81068638",
          4321 => x"757526ea",
          4322 => x"38805473",
          4323 => x"882981fb",
          4324 => x"c0057008",
          4325 => x"5255d5b5",
          4326 => x"3f81fef0",
          4327 => x"08537952",
          4328 => x"740851d6",
          4329 => x"893f81fe",
          4330 => x"f00880c4",
          4331 => x"38841533",
          4332 => x"5574812e",
          4333 => x"88387482",
          4334 => x"2e8838b4",
          4335 => x"39fcee3f",
          4336 => x"ab39811a",
          4337 => x"5a8c3dfc",
          4338 => x"1153f805",
          4339 => x"51f6af3f",
          4340 => x"81fef008",
          4341 => x"802e9938",
          4342 => x"7a537852",
          4343 => x"7751fdb8",
          4344 => x"3f81fef0",
          4345 => x"0881ff06",
          4346 => x"55748538",
          4347 => x"74549139",
          4348 => x"81147081",
          4349 => x"ff065154",
          4350 => x"827427ff",
          4351 => x"8e388054",
          4352 => x"7381fef0",
          4353 => x"0c8c3d0d",
          4354 => x"04d33d0d",
          4355 => x"b03d0802",
          4356 => x"840581c3",
          4357 => x"05335f5a",
          4358 => x"800baf3d",
          4359 => x"3481fbbc",
          4360 => x"335b81fb",
          4361 => x"b80881a3",
          4362 => x"3881fbb4",
          4363 => x"33547381",
          4364 => x"9a38a851",
          4365 => x"ebb43f81",
          4366 => x"fef00881",
          4367 => x"fbb80c81",
          4368 => x"fef00880",
          4369 => x"2e80fe38",
          4370 => x"935381fa",
          4371 => x"e0085281",
          4372 => x"fef00851",
          4373 => x"bbed3f81",
          4374 => x"fef00880",
          4375 => x"2e8b3881",
          4376 => x"e99851f3",
          4377 => x"a43f80e3",
          4378 => x"3981fbb8",
          4379 => x"085380f8",
          4380 => x"52903d70",
          4381 => x"525480f6",
          4382 => x"b03f81fe",
          4383 => x"f0085681",
          4384 => x"fef00874",
          4385 => x"2e098106",
          4386 => x"80c13881",
          4387 => x"fef00851",
          4388 => x"d3bb3f81",
          4389 => x"fef00855",
          4390 => x"800b81fe",
          4391 => x"f008259a",
          4392 => x"3881fef0",
          4393 => x"08ff0570",
          4394 => x"17555580",
          4395 => x"74348053",
          4396 => x"7481ff06",
          4397 => x"527551f9",
          4398 => x"b43f74ff",
          4399 => x"2e098106",
          4400 => x"ffa73887",
          4401 => x"39810b81",
          4402 => x"fbb4348f",
          4403 => x"3d5ddd8d",
          4404 => x"3f81fef0",
          4405 => x"08982b70",
          4406 => x"982c5159",
          4407 => x"78ff2eee",
          4408 => x"387881ff",
          4409 => x"0681ff94",
          4410 => x"3370982b",
          4411 => x"70982c81",
          4412 => x"ff903370",
          4413 => x"982b7097",
          4414 => x"2c71982c",
          4415 => x"05708429",
          4416 => x"81e9c805",
          4417 => x"70081570",
          4418 => x"33515151",
          4419 => x"51595951",
          4420 => x"595d5881",
          4421 => x"5673782e",
          4422 => x"80e93877",
          4423 => x"7427b438",
          4424 => x"7481800a",
          4425 => x"2981ff0a",
          4426 => x"0570982c",
          4427 => x"51558075",
          4428 => x"2480ce38",
          4429 => x"76537452",
          4430 => x"7751f7a6",
          4431 => x"3f81fef0",
          4432 => x"0881ff06",
          4433 => x"5473802e",
          4434 => x"d7387481",
          4435 => x"ff903481",
          4436 => x"56b13974",
          4437 => x"81800a29",
          4438 => x"81800a05",
          4439 => x"70982c70",
          4440 => x"81ff0656",
          4441 => x"5155738a",
          4442 => x"26973876",
          4443 => x"53745277",
          4444 => x"51f6ef3f",
          4445 => x"81fef008",
          4446 => x"81ff0654",
          4447 => x"73cc38d3",
          4448 => x"39805675",
          4449 => x"802e80ca",
          4450 => x"38811c55",
          4451 => x"7481ff94",
          4452 => x"3474982b",
          4453 => x"70982c81",
          4454 => x"ff903370",
          4455 => x"982b7098",
          4456 => x"2c701011",
          4457 => x"70822b81",
          4458 => x"e9cc1133",
          4459 => x"5e515151",
          4460 => x"57585155",
          4461 => x"74772e09",
          4462 => x"8106fe92",
          4463 => x"3881e9d0",
          4464 => x"14087d0c",
          4465 => x"800b81ff",
          4466 => x"9434800b",
          4467 => x"81ff9034",
          4468 => x"92397581",
          4469 => x"ff943475",
          4470 => x"81ff9034",
          4471 => x"78af3d34",
          4472 => x"757d0c7e",
          4473 => x"54738b26",
          4474 => x"fde13873",
          4475 => x"842981e1",
          4476 => x"d4055473",
          4477 => x"080481ff",
          4478 => x"9c335473",
          4479 => x"7e2efdcb",
          4480 => x"3881ff98",
          4481 => x"33557375",
          4482 => x"27ab3874",
          4483 => x"982b7098",
          4484 => x"2c515573",
          4485 => x"75249e38",
          4486 => x"741a5473",
          4487 => x"33811534",
          4488 => x"7481800a",
          4489 => x"2981ff0a",
          4490 => x"0570982c",
          4491 => x"81ff9c33",
          4492 => x"565155df",
          4493 => x"3981ff9c",
          4494 => x"33811156",
          4495 => x"547481ff",
          4496 => x"9c34731a",
          4497 => x"54ae3d33",
          4498 => x"743481ff",
          4499 => x"98335473",
          4500 => x"7e278938",
          4501 => x"81145473",
          4502 => x"81ff9834",
          4503 => x"81ff9c33",
          4504 => x"7081800a",
          4505 => x"2981ff0a",
          4506 => x"0570982c",
          4507 => x"81ff9833",
          4508 => x"5a515656",
          4509 => x"747725a2",
          4510 => x"38741a70",
          4511 => x"335254e8",
          4512 => x"c73f7481",
          4513 => x"800a2981",
          4514 => x"800a0570",
          4515 => x"982c81ff",
          4516 => x"98335651",
          4517 => x"55737524",
          4518 => x"e03881ff",
          4519 => x"9c337098",
          4520 => x"2b70982c",
          4521 => x"81ff9833",
          4522 => x"5a515656",
          4523 => x"747725fc",
          4524 => x"9a388851",
          4525 => x"e8923f74",
          4526 => x"81800a29",
          4527 => x"81800a05",
          4528 => x"70982c81",
          4529 => x"ff983356",
          4530 => x"51557375",
          4531 => x"24e438fb",
          4532 => x"fa3981ff",
          4533 => x"9c337081",
          4534 => x"ff065555",
          4535 => x"73802efb",
          4536 => x"ea3881ff",
          4537 => x"9833ff05",
          4538 => x"547381ff",
          4539 => x"9834ff15",
          4540 => x"547381ff",
          4541 => x"9c348851",
          4542 => x"e7ce3f81",
          4543 => x"ff9c3370",
          4544 => x"982b7098",
          4545 => x"2c81ff98",
          4546 => x"33575156",
          4547 => x"57747425",
          4548 => x"a738741a",
          4549 => x"54811433",
          4550 => x"74347333",
          4551 => x"51e7a93f",
          4552 => x"7481800a",
          4553 => x"2981800a",
          4554 => x"0570982c",
          4555 => x"81ff9833",
          4556 => x"58515575",
          4557 => x"7524db38",
          4558 => x"a051e78c",
          4559 => x"3f81ff9c",
          4560 => x"3370982b",
          4561 => x"70982c81",
          4562 => x"ff983357",
          4563 => x"51565774",
          4564 => x"7424faf7",
          4565 => x"388851e6",
          4566 => x"ef3f7481",
          4567 => x"800a2981",
          4568 => x"800a0570",
          4569 => x"982c81ff",
          4570 => x"98335851",
          4571 => x"55757525",
          4572 => x"e438fad7",
          4573 => x"3981ff98",
          4574 => x"337a0554",
          4575 => x"8074348a",
          4576 => x"51e6c53f",
          4577 => x"81ff9852",
          4578 => x"7951f7c6",
          4579 => x"3f81fef0",
          4580 => x"0881ff06",
          4581 => x"54739838",
          4582 => x"81ff9833",
          4583 => x"5473802e",
          4584 => x"84c93881",
          4585 => x"53735279",
          4586 => x"51f3c23f",
          4587 => x"84bd3980",
          4588 => x"7a3484b7",
          4589 => x"3981ff9c",
          4590 => x"33547380",
          4591 => x"2efa8c38",
          4592 => x"8851e684",
          4593 => x"3f81ff9c",
          4594 => x"33ff0554",
          4595 => x"7381ff9c",
          4596 => x"347381ff",
          4597 => x"0654e339",
          4598 => x"81ff9c33",
          4599 => x"81ff9833",
          4600 => x"55557375",
          4601 => x"2ef9e438",
          4602 => x"ff145473",
          4603 => x"81ff9834",
          4604 => x"74982b70",
          4605 => x"982c7581",
          4606 => x"ff065651",
          4607 => x"55747425",
          4608 => x"a738741a",
          4609 => x"54811433",
          4610 => x"74347333",
          4611 => x"51e5b93f",
          4612 => x"7481800a",
          4613 => x"2981800a",
          4614 => x"0570982c",
          4615 => x"81ff9833",
          4616 => x"58515575",
          4617 => x"7524db38",
          4618 => x"a051e59c",
          4619 => x"3f81ff9c",
          4620 => x"3370982b",
          4621 => x"70982c81",
          4622 => x"ff983357",
          4623 => x"51565774",
          4624 => x"7424f987",
          4625 => x"388851e4",
          4626 => x"ff3f7481",
          4627 => x"800a2981",
          4628 => x"800a0570",
          4629 => x"982c81ff",
          4630 => x"98335851",
          4631 => x"55757525",
          4632 => x"e438f8e7",
          4633 => x"3981ff9c",
          4634 => x"337081ff",
          4635 => x"0681ff98",
          4636 => x"33595654",
          4637 => x"747727f8",
          4638 => x"d2388114",
          4639 => x"547381ff",
          4640 => x"9c34741a",
          4641 => x"70335254",
          4642 => x"e4be3f81",
          4643 => x"ff9c3370",
          4644 => x"81ff0681",
          4645 => x"ff983358",
          4646 => x"56547575",
          4647 => x"26dc38f8",
          4648 => x"aa397aae",
          4649 => x"3881fbb0",
          4650 => x"08557480",
          4651 => x"2ea43874",
          4652 => x"51cb9a3f",
          4653 => x"81fef008",
          4654 => x"81ff9834",
          4655 => x"81fef008",
          4656 => x"81ff0681",
          4657 => x"05537452",
          4658 => x"7951c7e6",
          4659 => x"3f935b81",
          4660 => x"c1397a84",
          4661 => x"2981fae4",
          4662 => x"05fc1108",
          4663 => x"56547480",
          4664 => x"2ea53874",
          4665 => x"51cae63f",
          4666 => x"81fef008",
          4667 => x"81ff9834",
          4668 => x"81fef008",
          4669 => x"81ff0681",
          4670 => x"05537452",
          4671 => x"7951c7b2",
          4672 => x"3fff1b54",
          4673 => x"80de3973",
          4674 => x"08557480",
          4675 => x"2ef7bc38",
          4676 => x"7451cab9",
          4677 => x"3f80e239",
          4678 => x"7a932e09",
          4679 => x"81069338",
          4680 => x"81fae408",
          4681 => x"5574802e",
          4682 => x"89387451",
          4683 => x"ca9f3f80",
          4684 => x"c8397a84",
          4685 => x"2981fae4",
          4686 => x"05841108",
          4687 => x"56547480",
          4688 => x"2ea93874",
          4689 => x"51ca863f",
          4690 => x"81fef008",
          4691 => x"81ff9834",
          4692 => x"81fef008",
          4693 => x"81ff0681",
          4694 => x"05537452",
          4695 => x"7951c6d2",
          4696 => x"3f811b54",
          4697 => x"7381ff06",
          4698 => x"5ba83973",
          4699 => x"08557480",
          4700 => x"2ef6d838",
          4701 => x"7451c9d5",
          4702 => x"3f81fef0",
          4703 => x"0881ff98",
          4704 => x"3481fef0",
          4705 => x"0881ff06",
          4706 => x"81055374",
          4707 => x"527951c6",
          4708 => x"a13f81ff",
          4709 => x"9c5381ff",
          4710 => x"98335279",
          4711 => x"51ef903f",
          4712 => x"f6a93981",
          4713 => x"ff9c3370",
          4714 => x"81ff0681",
          4715 => x"ff983359",
          4716 => x"56547477",
          4717 => x"27f69438",
          4718 => x"81145473",
          4719 => x"81ff9c34",
          4720 => x"741a7033",
          4721 => x"5254e280",
          4722 => x"3ff68039",
          4723 => x"81ff9c33",
          4724 => x"5473802e",
          4725 => x"f5f53888",
          4726 => x"51e1ed3f",
          4727 => x"81ff9c33",
          4728 => x"ff055473",
          4729 => x"81ff9c34",
          4730 => x"f5e13980",
          4731 => x"0b81ff9c",
          4732 => x"34800b81",
          4733 => x"ff983479",
          4734 => x"81fef00c",
          4735 => x"af3d0d04",
          4736 => x"ff3d0d02",
          4737 => x"8f053351",
          4738 => x"81527072",
          4739 => x"26873881",
          4740 => x"fbd81133",
          4741 => x"527181fe",
          4742 => x"f00c833d",
          4743 => x"0d04fc3d",
          4744 => x"0d029b05",
          4745 => x"33028405",
          4746 => x"9f053356",
          4747 => x"53835172",
          4748 => x"812680e0",
          4749 => x"3872842b",
          4750 => x"87c0928c",
          4751 => x"11535188",
          4752 => x"5474802e",
          4753 => x"84388188",
          4754 => x"5473720c",
          4755 => x"87c0928c",
          4756 => x"11518171",
          4757 => x"0c850b87",
          4758 => x"c0988c0c",
          4759 => x"70527108",
          4760 => x"70820651",
          4761 => x"5170802e",
          4762 => x"8a3887c0",
          4763 => x"988c0851",
          4764 => x"70ec3871",
          4765 => x"08fc8080",
          4766 => x"06527192",
          4767 => x"3887c098",
          4768 => x"8c085170",
          4769 => x"802e8738",
          4770 => x"7181fbd8",
          4771 => x"143481fb",
          4772 => x"d8133351",
          4773 => x"7081fef0",
          4774 => x"0c863d0d",
          4775 => x"04f33d0d",
          4776 => x"60626402",
          4777 => x"8c05bf05",
          4778 => x"33574058",
          4779 => x"5b837452",
          4780 => x"5afecd3f",
          4781 => x"81fef008",
          4782 => x"81067a54",
          4783 => x"527181be",
          4784 => x"38717275",
          4785 => x"842b87c0",
          4786 => x"92801187",
          4787 => x"c0928c12",
          4788 => x"87c09284",
          4789 => x"13415a40",
          4790 => x"575a5885",
          4791 => x"0b87c098",
          4792 => x"8c0c767d",
          4793 => x"0c84760c",
          4794 => x"75087085",
          4795 => x"2a708106",
          4796 => x"51535471",
          4797 => x"802e8e38",
          4798 => x"7b085271",
          4799 => x"7b708105",
          4800 => x"5d348119",
          4801 => x"598074a2",
          4802 => x"06535371",
          4803 => x"732e8338",
          4804 => x"81537883",
          4805 => x"ff268f38",
          4806 => x"72802e8a",
          4807 => x"3887c098",
          4808 => x"8c085271",
          4809 => x"c33887c0",
          4810 => x"988c0852",
          4811 => x"71802e87",
          4812 => x"38788480",
          4813 => x"2e993881",
          4814 => x"760c87c0",
          4815 => x"928c1553",
          4816 => x"72087082",
          4817 => x"06515271",
          4818 => x"f738ff1a",
          4819 => x"5a8d3984",
          4820 => x"80178119",
          4821 => x"7081ff06",
          4822 => x"5a535779",
          4823 => x"802e9038",
          4824 => x"73fc8080",
          4825 => x"06527187",
          4826 => x"387d7826",
          4827 => x"feed3873",
          4828 => x"fc808006",
          4829 => x"5271802e",
          4830 => x"83388152",
          4831 => x"71537281",
          4832 => x"fef00c8f",
          4833 => x"3d0d04f3",
          4834 => x"3d0d6062",
          4835 => x"64028c05",
          4836 => x"bf053357",
          4837 => x"40585b83",
          4838 => x"59807452",
          4839 => x"58fce13f",
          4840 => x"81fef008",
          4841 => x"81067954",
          4842 => x"5271782e",
          4843 => x"09810681",
          4844 => x"b1387774",
          4845 => x"842b87c0",
          4846 => x"92801187",
          4847 => x"c0928c12",
          4848 => x"87c09284",
          4849 => x"1340595f",
          4850 => x"565a850b",
          4851 => x"87c0988c",
          4852 => x"0c767d0c",
          4853 => x"82760c80",
          4854 => x"58750870",
          4855 => x"842a7081",
          4856 => x"06515354",
          4857 => x"71802e8c",
          4858 => x"387a7081",
          4859 => x"055c337c",
          4860 => x"0c811858",
          4861 => x"73812a70",
          4862 => x"81065152",
          4863 => x"71802e8a",
          4864 => x"3887c098",
          4865 => x"8c085271",
          4866 => x"d03887c0",
          4867 => x"988c0852",
          4868 => x"71802e87",
          4869 => x"38778480",
          4870 => x"2e993881",
          4871 => x"760c87c0",
          4872 => x"928c1553",
          4873 => x"72087082",
          4874 => x"06515271",
          4875 => x"f738ff19",
          4876 => x"598d3981",
          4877 => x"1a7081ff",
          4878 => x"06848019",
          4879 => x"595b5278",
          4880 => x"802e9038",
          4881 => x"73fc8080",
          4882 => x"06527187",
          4883 => x"387d7a26",
          4884 => x"fef83873",
          4885 => x"fc808006",
          4886 => x"5271802e",
          4887 => x"83388152",
          4888 => x"71537281",
          4889 => x"fef00c8f",
          4890 => x"3d0d04fa",
          4891 => x"3d0d7a02",
          4892 => x"8405a305",
          4893 => x"33028805",
          4894 => x"a7053371",
          4895 => x"54545657",
          4896 => x"fafe3f81",
          4897 => x"fef00881",
          4898 => x"06538354",
          4899 => x"7280fe38",
          4900 => x"850b87c0",
          4901 => x"988c0c81",
          4902 => x"5671762e",
          4903 => x"80dc3871",
          4904 => x"76249338",
          4905 => x"74842b87",
          4906 => x"c0928c11",
          4907 => x"54547180",
          4908 => x"2e8d3880",
          4909 => x"d4397183",
          4910 => x"2e80c638",
          4911 => x"80cb3972",
          4912 => x"0870812a",
          4913 => x"70810651",
          4914 => x"51527180",
          4915 => x"2e8a3887",
          4916 => x"c0988c08",
          4917 => x"5271e838",
          4918 => x"87c0988c",
          4919 => x"08527196",
          4920 => x"3881730c",
          4921 => x"87c0928c",
          4922 => x"14537208",
          4923 => x"70820651",
          4924 => x"5271f738",
          4925 => x"96398056",
          4926 => x"92398880",
          4927 => x"0a770c85",
          4928 => x"39818077",
          4929 => x"0c725683",
          4930 => x"39845675",
          4931 => x"547381fe",
          4932 => x"f00c883d",
          4933 => x"0d04fe3d",
          4934 => x"0d748111",
          4935 => x"33713371",
          4936 => x"882b0781",
          4937 => x"fef00c53",
          4938 => x"51843d0d",
          4939 => x"04fd3d0d",
          4940 => x"75831133",
          4941 => x"82123371",
          4942 => x"902b7188",
          4943 => x"2b078114",
          4944 => x"33707207",
          4945 => x"882b7533",
          4946 => x"710781fe",
          4947 => x"f00c5253",
          4948 => x"54565452",
          4949 => x"853d0d04",
          4950 => x"ff3d0d73",
          4951 => x"02840592",
          4952 => x"05225252",
          4953 => x"70727081",
          4954 => x"05543470",
          4955 => x"882a5170",
          4956 => x"7234833d",
          4957 => x"0d04ff3d",
          4958 => x"0d737552",
          4959 => x"52707270",
          4960 => x"81055434",
          4961 => x"70882a51",
          4962 => x"70727081",
          4963 => x"05543470",
          4964 => x"882a5170",
          4965 => x"72708105",
          4966 => x"54347088",
          4967 => x"2a517072",
          4968 => x"34833d0d",
          4969 => x"04fe3d0d",
          4970 => x"76757754",
          4971 => x"54517080",
          4972 => x"2e923871",
          4973 => x"70810553",
          4974 => x"33737081",
          4975 => x"055534ff",
          4976 => x"1151eb39",
          4977 => x"843d0d04",
          4978 => x"fe3d0d75",
          4979 => x"77765452",
          4980 => x"53727270",
          4981 => x"81055434",
          4982 => x"ff115170",
          4983 => x"f438843d",
          4984 => x"0d04fc3d",
          4985 => x"0d787779",
          4986 => x"56565374",
          4987 => x"70810556",
          4988 => x"33747081",
          4989 => x"05563371",
          4990 => x"7131ff16",
          4991 => x"56525252",
          4992 => x"72802e86",
          4993 => x"3871802e",
          4994 => x"e2387181",
          4995 => x"fef00c86",
          4996 => x"3d0d04fe",
          4997 => x"3d0d7476",
          4998 => x"54518939",
          4999 => x"71732e8a",
          5000 => x"38811151",
          5001 => x"70335271",
          5002 => x"f3387033",
          5003 => x"81fef00c",
          5004 => x"843d0d04",
          5005 => x"800b81fe",
          5006 => x"f00c0480",
          5007 => x"0b81fef0",
          5008 => x"0c04f73d",
          5009 => x"0d7b5680",
          5010 => x"0b831733",
          5011 => x"565a747a",
          5012 => x"2e80d638",
          5013 => x"8154b016",
          5014 => x"0853b416",
          5015 => x"70538117",
          5016 => x"335259fa",
          5017 => x"a23f81fe",
          5018 => x"f0087a2e",
          5019 => x"098106b7",
          5020 => x"3881fef0",
          5021 => x"08831734",
          5022 => x"b0160870",
          5023 => x"a4180831",
          5024 => x"9c180859",
          5025 => x"56587477",
          5026 => x"279f3882",
          5027 => x"16335574",
          5028 => x"822e0981",
          5029 => x"06933881",
          5030 => x"54761853",
          5031 => x"78528116",
          5032 => x"3351f9e3",
          5033 => x"3f833981",
          5034 => x"5a7981fe",
          5035 => x"f00c8b3d",
          5036 => x"0d04fa3d",
          5037 => x"0d787a56",
          5038 => x"56805774",
          5039 => x"b017082e",
          5040 => x"af387551",
          5041 => x"fefc3f81",
          5042 => x"fef00857",
          5043 => x"81fef008",
          5044 => x"9f388154",
          5045 => x"7453b416",
          5046 => x"52811633",
          5047 => x"51f7be3f",
          5048 => x"81fef008",
          5049 => x"802e8538",
          5050 => x"ff558157",
          5051 => x"74b0170c",
          5052 => x"7681fef0",
          5053 => x"0c883d0d",
          5054 => x"04f83d0d",
          5055 => x"7a705257",
          5056 => x"fec03f81",
          5057 => x"fef00858",
          5058 => x"81fef008",
          5059 => x"81913876",
          5060 => x"33557483",
          5061 => x"2e098106",
          5062 => x"80f03884",
          5063 => x"17335978",
          5064 => x"812e0981",
          5065 => x"0680e338",
          5066 => x"84805381",
          5067 => x"fef00852",
          5068 => x"b4177052",
          5069 => x"56fd913f",
          5070 => x"82d4d552",
          5071 => x"84b21751",
          5072 => x"fc963f84",
          5073 => x"8b85a4d2",
          5074 => x"527551fc",
          5075 => x"a93f868a",
          5076 => x"85e4f252",
          5077 => x"84981751",
          5078 => x"fc9c3f90",
          5079 => x"17085284",
          5080 => x"9c1751fc",
          5081 => x"913f8c17",
          5082 => x"085284a0",
          5083 => x"1751fc86",
          5084 => x"3fa01708",
          5085 => x"810570b0",
          5086 => x"190c7955",
          5087 => x"53755281",
          5088 => x"173351f8",
          5089 => x"823f7784",
          5090 => x"18348053",
          5091 => x"80528117",
          5092 => x"3351f9d7",
          5093 => x"3f81fef0",
          5094 => x"08802e83",
          5095 => x"38815877",
          5096 => x"81fef00c",
          5097 => x"8a3d0d04",
          5098 => x"fb3d0d77",
          5099 => x"fe1a9812",
          5100 => x"08fe0555",
          5101 => x"56548056",
          5102 => x"7473278d",
          5103 => x"388a1422",
          5104 => x"757129ac",
          5105 => x"16080557",
          5106 => x"537581fe",
          5107 => x"f00c873d",
          5108 => x"0d04f93d",
          5109 => x"0d7a7a70",
          5110 => x"08565457",
          5111 => x"81772781",
          5112 => x"df387698",
          5113 => x"15082781",
          5114 => x"d738ff74",
          5115 => x"33545872",
          5116 => x"822e80f5",
          5117 => x"38728224",
          5118 => x"89387281",
          5119 => x"2e8d3881",
          5120 => x"bf397283",
          5121 => x"2e818e38",
          5122 => x"81b63976",
          5123 => x"812a1770",
          5124 => x"892aa416",
          5125 => x"08055374",
          5126 => x"5255fd96",
          5127 => x"3f81fef0",
          5128 => x"08819f38",
          5129 => x"7483ff06",
          5130 => x"14b41133",
          5131 => x"81177089",
          5132 => x"2aa41808",
          5133 => x"05557654",
          5134 => x"575753fc",
          5135 => x"f53f81fe",
          5136 => x"f00880fe",
          5137 => x"387483ff",
          5138 => x"0614b411",
          5139 => x"3370882b",
          5140 => x"78077981",
          5141 => x"0671842a",
          5142 => x"5c525851",
          5143 => x"537280e2",
          5144 => x"38759fff",
          5145 => x"065880da",
          5146 => x"3976882a",
          5147 => x"a4150805",
          5148 => x"527351fc",
          5149 => x"bd3f81fe",
          5150 => x"f00880c6",
          5151 => x"38761083",
          5152 => x"fe067405",
          5153 => x"b40551f9",
          5154 => x"8d3f81fe",
          5155 => x"f00883ff",
          5156 => x"ff0658ae",
          5157 => x"3976872a",
          5158 => x"a4150805",
          5159 => x"527351fc",
          5160 => x"913f81fe",
          5161 => x"f0089b38",
          5162 => x"76822b83",
          5163 => x"fc067405",
          5164 => x"b40551f8",
          5165 => x"f83f81fe",
          5166 => x"f008f00a",
          5167 => x"06588339",
          5168 => x"81587781",
          5169 => x"fef00c89",
          5170 => x"3d0d04f8",
          5171 => x"3d0d7a7c",
          5172 => x"7e5a5856",
          5173 => x"82598177",
          5174 => x"27829e38",
          5175 => x"76981708",
          5176 => x"27829638",
          5177 => x"75335372",
          5178 => x"792e819d",
          5179 => x"38727924",
          5180 => x"89387281",
          5181 => x"2e8d3882",
          5182 => x"80397283",
          5183 => x"2e81b838",
          5184 => x"81f73976",
          5185 => x"812a1770",
          5186 => x"892aa418",
          5187 => x"08055376",
          5188 => x"5255fb9e",
          5189 => x"3f81fef0",
          5190 => x"085981fe",
          5191 => x"f00881d9",
          5192 => x"387483ff",
          5193 => x"0616b405",
          5194 => x"81167881",
          5195 => x"06595654",
          5196 => x"77537680",
          5197 => x"2e8f3877",
          5198 => x"842b9ff0",
          5199 => x"0674338f",
          5200 => x"06710751",
          5201 => x"53727434",
          5202 => x"810b8317",
          5203 => x"3474892a",
          5204 => x"a4170805",
          5205 => x"527551fa",
          5206 => x"d93f81fe",
          5207 => x"f0085981",
          5208 => x"fef00881",
          5209 => x"94387483",
          5210 => x"ff0616b4",
          5211 => x"0578842a",
          5212 => x"5454768f",
          5213 => x"3877882a",
          5214 => x"743381f0",
          5215 => x"06718f06",
          5216 => x"07515372",
          5217 => x"743480ec",
          5218 => x"3976882a",
          5219 => x"a4170805",
          5220 => x"527551fa",
          5221 => x"9d3f81fe",
          5222 => x"f0085981",
          5223 => x"fef00880",
          5224 => x"d8387783",
          5225 => x"ffff0652",
          5226 => x"761083fe",
          5227 => x"067605b4",
          5228 => x"0551f7a4",
          5229 => x"3fbe3976",
          5230 => x"872aa417",
          5231 => x"08055275",
          5232 => x"51f9ef3f",
          5233 => x"81fef008",
          5234 => x"5981fef0",
          5235 => x"08ab3877",
          5236 => x"f00a0677",
          5237 => x"822b83fc",
          5238 => x"067018b4",
          5239 => x"05705451",
          5240 => x"5454f6c9",
          5241 => x"3f81fef0",
          5242 => x"088f0a06",
          5243 => x"74075272",
          5244 => x"51f7833f",
          5245 => x"810b8317",
          5246 => x"347881fe",
          5247 => x"f00c8a3d",
          5248 => x"0d04f83d",
          5249 => x"0d7a7c7e",
          5250 => x"72085956",
          5251 => x"56598175",
          5252 => x"27a43874",
          5253 => x"98170827",
          5254 => x"9d387380",
          5255 => x"2eaa38ff",
          5256 => x"53735275",
          5257 => x"51fda43f",
          5258 => x"81fef008",
          5259 => x"5481fef0",
          5260 => x"0880f238",
          5261 => x"93398254",
          5262 => x"80eb3981",
          5263 => x"5480e639",
          5264 => x"81fef008",
          5265 => x"5480de39",
          5266 => x"74527851",
          5267 => x"fb843f81",
          5268 => x"fef00858",
          5269 => x"81fef008",
          5270 => x"802e80c7",
          5271 => x"3881fef0",
          5272 => x"08812ed2",
          5273 => x"3881fef0",
          5274 => x"08ff2ecf",
          5275 => x"38805374",
          5276 => x"527551fc",
          5277 => x"d63f81fe",
          5278 => x"f008c538",
          5279 => x"981608fe",
          5280 => x"11901808",
          5281 => x"57555774",
          5282 => x"74279038",
          5283 => x"81159017",
          5284 => x"0c841633",
          5285 => x"81075473",
          5286 => x"84173477",
          5287 => x"55767826",
          5288 => x"ffa63880",
          5289 => x"547381fe",
          5290 => x"f00c8a3d",
          5291 => x"0d04f63d",
          5292 => x"0d7c7e71",
          5293 => x"08595b5b",
          5294 => x"7995388c",
          5295 => x"17085877",
          5296 => x"802e8838",
          5297 => x"98170878",
          5298 => x"26b23881",
          5299 => x"58ae3979",
          5300 => x"527a51f9",
          5301 => x"fd3f8155",
          5302 => x"7481fef0",
          5303 => x"082782e0",
          5304 => x"3881fef0",
          5305 => x"085581fe",
          5306 => x"f008ff2e",
          5307 => x"82d23898",
          5308 => x"170881fe",
          5309 => x"f0082682",
          5310 => x"c7387958",
          5311 => x"90170870",
          5312 => x"56547380",
          5313 => x"2e82b938",
          5314 => x"777a2e09",
          5315 => x"810680e2",
          5316 => x"38811a56",
          5317 => x"98170876",
          5318 => x"26833882",
          5319 => x"5675527a",
          5320 => x"51f9af3f",
          5321 => x"805981fe",
          5322 => x"f008812e",
          5323 => x"09810686",
          5324 => x"3881fef0",
          5325 => x"085981fe",
          5326 => x"f0080970",
          5327 => x"30707207",
          5328 => x"8025707c",
          5329 => x"0781fef0",
          5330 => x"08545151",
          5331 => x"55557381",
          5332 => x"ef3881fe",
          5333 => x"f008802e",
          5334 => x"95388c17",
          5335 => x"08548174",
          5336 => x"27903873",
          5337 => x"98180827",
          5338 => x"89387358",
          5339 => x"85397580",
          5340 => x"db387756",
          5341 => x"81165698",
          5342 => x"17087626",
          5343 => x"89388256",
          5344 => x"75782681",
          5345 => x"ac387552",
          5346 => x"7a51f8c6",
          5347 => x"3f81fef0",
          5348 => x"08802eb8",
          5349 => x"38805981",
          5350 => x"fef00881",
          5351 => x"2e098106",
          5352 => x"863881fe",
          5353 => x"f0085981",
          5354 => x"fef00809",
          5355 => x"70307072",
          5356 => x"07802570",
          5357 => x"7c075151",
          5358 => x"55557380",
          5359 => x"f8387578",
          5360 => x"2e098106",
          5361 => x"ffae3873",
          5362 => x"5580f539",
          5363 => x"ff537552",
          5364 => x"7651f9f7",
          5365 => x"3f81fef0",
          5366 => x"0881fef0",
          5367 => x"08307081",
          5368 => x"fef00807",
          5369 => x"80255155",
          5370 => x"5579802e",
          5371 => x"94387380",
          5372 => x"2e8f3875",
          5373 => x"53795276",
          5374 => x"51f9d03f",
          5375 => x"81fef008",
          5376 => x"5574a538",
          5377 => x"758c180c",
          5378 => x"981708fe",
          5379 => x"05901808",
          5380 => x"56547474",
          5381 => x"268638ff",
          5382 => x"1590180c",
          5383 => x"84173381",
          5384 => x"07547384",
          5385 => x"18349739",
          5386 => x"ff567481",
          5387 => x"2e90388c",
          5388 => x"3980558c",
          5389 => x"3981fef0",
          5390 => x"08558539",
          5391 => x"81567555",
          5392 => x"7481fef0",
          5393 => x"0c8c3d0d",
          5394 => x"04f83d0d",
          5395 => x"7a705255",
          5396 => x"f3f03f81",
          5397 => x"fef00858",
          5398 => x"815681fe",
          5399 => x"f00880d8",
          5400 => x"387b5274",
          5401 => x"51f6c13f",
          5402 => x"81fef008",
          5403 => x"81fef008",
          5404 => x"b0170c59",
          5405 => x"84805377",
          5406 => x"52b41570",
          5407 => x"5257f2c8",
          5408 => x"3f775684",
          5409 => x"39811656",
          5410 => x"8a152258",
          5411 => x"75782797",
          5412 => x"38815475",
          5413 => x"19537652",
          5414 => x"81153351",
          5415 => x"ede93f81",
          5416 => x"fef00880",
          5417 => x"2edf388a",
          5418 => x"15227632",
          5419 => x"70307072",
          5420 => x"07709f2a",
          5421 => x"53515656",
          5422 => x"7581fef0",
          5423 => x"0c8a3d0d",
          5424 => x"04f83d0d",
          5425 => x"7a7c7108",
          5426 => x"58565774",
          5427 => x"f0800a26",
          5428 => x"80f13874",
          5429 => x"9f065372",
          5430 => x"80e93874",
          5431 => x"90180c88",
          5432 => x"17085473",
          5433 => x"aa387533",
          5434 => x"53827327",
          5435 => x"8838a816",
          5436 => x"0854739b",
          5437 => x"3874852a",
          5438 => x"53820b88",
          5439 => x"17225a58",
          5440 => x"72792780",
          5441 => x"fe38a816",
          5442 => x"0898180c",
          5443 => x"80cd398a",
          5444 => x"16227089",
          5445 => x"2b545872",
          5446 => x"7526b238",
          5447 => x"73527651",
          5448 => x"f5b03f81",
          5449 => x"fef00854",
          5450 => x"81fef008",
          5451 => x"ff2ebd38",
          5452 => x"810b81fe",
          5453 => x"f008278b",
          5454 => x"38981608",
          5455 => x"81fef008",
          5456 => x"26853882",
          5457 => x"58bd3974",
          5458 => x"733155cb",
          5459 => x"39735275",
          5460 => x"51f4d53f",
          5461 => x"81fef008",
          5462 => x"98180c73",
          5463 => x"94180c98",
          5464 => x"17085382",
          5465 => x"5872802e",
          5466 => x"9a388539",
          5467 => x"81589439",
          5468 => x"74892a13",
          5469 => x"98180c74",
          5470 => x"83ff0616",
          5471 => x"b4059c18",
          5472 => x"0c805877",
          5473 => x"81fef00c",
          5474 => x"8a3d0d04",
          5475 => x"f83d0d7a",
          5476 => x"70089012",
          5477 => x"08a00559",
          5478 => x"5754f080",
          5479 => x"0a772786",
          5480 => x"38800b98",
          5481 => x"150c9814",
          5482 => x"08538455",
          5483 => x"72802e81",
          5484 => x"cb387683",
          5485 => x"ff065877",
          5486 => x"81b53881",
          5487 => x"1398150c",
          5488 => x"94140855",
          5489 => x"74923876",
          5490 => x"852a8817",
          5491 => x"22565374",
          5492 => x"7326819b",
          5493 => x"3880c039",
          5494 => x"8a1622ff",
          5495 => x"0577892a",
          5496 => x"06537281",
          5497 => x"8a387452",
          5498 => x"7351f3e6",
          5499 => x"3f81fef0",
          5500 => x"08538255",
          5501 => x"810b81fe",
          5502 => x"f0082780",
          5503 => x"ff388155",
          5504 => x"81fef008",
          5505 => x"ff2e80f4",
          5506 => x"38981608",
          5507 => x"81fef008",
          5508 => x"2680ca38",
          5509 => x"7b8a3877",
          5510 => x"98150c84",
          5511 => x"5580dd39",
          5512 => x"94140852",
          5513 => x"7351f986",
          5514 => x"3f81fef0",
          5515 => x"08538755",
          5516 => x"81fef008",
          5517 => x"802e80c4",
          5518 => x"38825581",
          5519 => x"fef00881",
          5520 => x"2eba3881",
          5521 => x"5581fef0",
          5522 => x"08ff2eb0",
          5523 => x"3881fef0",
          5524 => x"08527551",
          5525 => x"fbf33f81",
          5526 => x"fef008a0",
          5527 => x"38729415",
          5528 => x"0c725275",
          5529 => x"51f2c13f",
          5530 => x"81fef008",
          5531 => x"98150c76",
          5532 => x"90150c77",
          5533 => x"16b4059c",
          5534 => x"150c8055",
          5535 => x"7481fef0",
          5536 => x"0c8a3d0d",
          5537 => x"04f73d0d",
          5538 => x"7b7d7108",
          5539 => x"5b5b5780",
          5540 => x"527651fc",
          5541 => x"ac3f81fe",
          5542 => x"f0085481",
          5543 => x"fef00880",
          5544 => x"ec3881fe",
          5545 => x"f0085698",
          5546 => x"17085278",
          5547 => x"51f0833f",
          5548 => x"81fef008",
          5549 => x"5481fef0",
          5550 => x"0880d238",
          5551 => x"81fef008",
          5552 => x"9c180870",
          5553 => x"33515458",
          5554 => x"7281e52e",
          5555 => x"09810683",
          5556 => x"38815881",
          5557 => x"fef00855",
          5558 => x"72833881",
          5559 => x"55777507",
          5560 => x"5372802e",
          5561 => x"8e388116",
          5562 => x"56757a2e",
          5563 => x"09810688",
          5564 => x"38a53981",
          5565 => x"fef00856",
          5566 => x"81527651",
          5567 => x"fd8e3f81",
          5568 => x"fef00854",
          5569 => x"81fef008",
          5570 => x"802eff9b",
          5571 => x"3873842e",
          5572 => x"09810683",
          5573 => x"38875473",
          5574 => x"81fef00c",
          5575 => x"8b3d0d04",
          5576 => x"fd3d0d76",
          5577 => x"9a115254",
          5578 => x"ebec3f81",
          5579 => x"fef00883",
          5580 => x"ffff0676",
          5581 => x"70335153",
          5582 => x"5371832e",
          5583 => x"09810690",
          5584 => x"38941451",
          5585 => x"ebd03f81",
          5586 => x"fef00890",
          5587 => x"2b730753",
          5588 => x"7281fef0",
          5589 => x"0c853d0d",
          5590 => x"04fc3d0d",
          5591 => x"77797083",
          5592 => x"ffff0654",
          5593 => x"9a125355",
          5594 => x"55ebed3f",
          5595 => x"76703351",
          5596 => x"5372832e",
          5597 => x"0981068b",
          5598 => x"3873902a",
          5599 => x"52941551",
          5600 => x"ebd63f86",
          5601 => x"3d0d04f7",
          5602 => x"3d0d7b7d",
          5603 => x"5b558475",
          5604 => x"085a5898",
          5605 => x"1508802e",
          5606 => x"818a3898",
          5607 => x"15085278",
          5608 => x"51ee8f3f",
          5609 => x"81fef008",
          5610 => x"5881fef0",
          5611 => x"0880f538",
          5612 => x"9c150870",
          5613 => x"33555373",
          5614 => x"86388458",
          5615 => x"80e6398b",
          5616 => x"133370bf",
          5617 => x"067081ff",
          5618 => x"06585153",
          5619 => x"72861634",
          5620 => x"81fef008",
          5621 => x"537381e5",
          5622 => x"2e833881",
          5623 => x"5373ae2e",
          5624 => x"a9388170",
          5625 => x"74065457",
          5626 => x"72802e9e",
          5627 => x"38758f2e",
          5628 => x"993881fe",
          5629 => x"f00876df",
          5630 => x"06545472",
          5631 => x"882e0981",
          5632 => x"06833876",
          5633 => x"54737a2e",
          5634 => x"a0388052",
          5635 => x"7451fafc",
          5636 => x"3f81fef0",
          5637 => x"085881fe",
          5638 => x"f0088938",
          5639 => x"981508fe",
          5640 => x"fa388639",
          5641 => x"800b9816",
          5642 => x"0c7781fe",
          5643 => x"f00c8b3d",
          5644 => x"0d04fb3d",
          5645 => x"0d777008",
          5646 => x"57548152",
          5647 => x"7351fcc5",
          5648 => x"3f81fef0",
          5649 => x"085581fe",
          5650 => x"f008b438",
          5651 => x"98140852",
          5652 => x"7551ecde",
          5653 => x"3f81fef0",
          5654 => x"085581fe",
          5655 => x"f008a038",
          5656 => x"a05381fe",
          5657 => x"f008529c",
          5658 => x"140851ea",
          5659 => x"db3f8b53",
          5660 => x"a014529c",
          5661 => x"140851ea",
          5662 => x"ac3f810b",
          5663 => x"83173474",
          5664 => x"81fef00c",
          5665 => x"873d0d04",
          5666 => x"fd3d0d75",
          5667 => x"70089812",
          5668 => x"08547053",
          5669 => x"5553ec9a",
          5670 => x"3f81fef0",
          5671 => x"088d389c",
          5672 => x"130853e5",
          5673 => x"7334810b",
          5674 => x"83153485",
          5675 => x"3d0d04fa",
          5676 => x"3d0d787a",
          5677 => x"5757800b",
          5678 => x"89173498",
          5679 => x"1708802e",
          5680 => x"81823880",
          5681 => x"70891855",
          5682 => x"55559c17",
          5683 => x"08147033",
          5684 => x"81165651",
          5685 => x"5271a02e",
          5686 => x"a8387185",
          5687 => x"2e098106",
          5688 => x"843881e5",
          5689 => x"5273892e",
          5690 => x"0981068b",
          5691 => x"38ae7370",
          5692 => x"81055534",
          5693 => x"81155571",
          5694 => x"73708105",
          5695 => x"55348115",
          5696 => x"558a7427",
          5697 => x"c5387515",
          5698 => x"88055280",
          5699 => x"0b811334",
          5700 => x"9c170852",
          5701 => x"8b123388",
          5702 => x"17349c17",
          5703 => x"089c1152",
          5704 => x"52e88a3f",
          5705 => x"81fef008",
          5706 => x"760c9612",
          5707 => x"51e7e73f",
          5708 => x"81fef008",
          5709 => x"86172398",
          5710 => x"1251e7da",
          5711 => x"3f81fef0",
          5712 => x"08841723",
          5713 => x"883d0d04",
          5714 => x"f33d0d7f",
          5715 => x"70085e5b",
          5716 => x"80617033",
          5717 => x"51555573",
          5718 => x"af2e8338",
          5719 => x"81557380",
          5720 => x"dc2e9138",
          5721 => x"74802e8c",
          5722 => x"38941d08",
          5723 => x"881c0caa",
          5724 => x"39811541",
          5725 => x"80617033",
          5726 => x"56565673",
          5727 => x"af2e0981",
          5728 => x"06833881",
          5729 => x"567380dc",
          5730 => x"32703070",
          5731 => x"80257807",
          5732 => x"51515473",
          5733 => x"dc387388",
          5734 => x"1c0c6070",
          5735 => x"33515473",
          5736 => x"9f269638",
          5737 => x"ff800bab",
          5738 => x"1c348052",
          5739 => x"7a51f691",
          5740 => x"3f81fef0",
          5741 => x"08558598",
          5742 => x"39913d61",
          5743 => x"a01d5c5a",
          5744 => x"5e8b53a0",
          5745 => x"527951e7",
          5746 => x"ff3f8070",
          5747 => x"59578879",
          5748 => x"33555c73",
          5749 => x"ae2e0981",
          5750 => x"0680d438",
          5751 => x"78187033",
          5752 => x"811a71ae",
          5753 => x"32703070",
          5754 => x"9f2a7382",
          5755 => x"26075151",
          5756 => x"535a5754",
          5757 => x"738c3879",
          5758 => x"17547574",
          5759 => x"34811757",
          5760 => x"db3975af",
          5761 => x"32703070",
          5762 => x"9f2a5151",
          5763 => x"547580dc",
          5764 => x"2e8c3873",
          5765 => x"802e8738",
          5766 => x"75a02682",
          5767 => x"bd387719",
          5768 => x"7e0ca454",
          5769 => x"a0762782",
          5770 => x"bd38a054",
          5771 => x"82b83978",
          5772 => x"18703381",
          5773 => x"1a5a5754",
          5774 => x"a0762781",
          5775 => x"fc3875af",
          5776 => x"32703077",
          5777 => x"80dc3270",
          5778 => x"30728025",
          5779 => x"71802507",
          5780 => x"51515651",
          5781 => x"5573802e",
          5782 => x"ac388439",
          5783 => x"81185880",
          5784 => x"781a7033",
          5785 => x"51555573",
          5786 => x"af2e0981",
          5787 => x"06833881",
          5788 => x"557380dc",
          5789 => x"32703070",
          5790 => x"80257707",
          5791 => x"51515473",
          5792 => x"db3881b5",
          5793 => x"3975ae2e",
          5794 => x"09810683",
          5795 => x"38815476",
          5796 => x"7c277407",
          5797 => x"5473802e",
          5798 => x"a2387b8b",
          5799 => x"32703077",
          5800 => x"ae327030",
          5801 => x"72802571",
          5802 => x"9f2a0753",
          5803 => x"51565155",
          5804 => x"7481a738",
          5805 => x"88578b5c",
          5806 => x"fef53975",
          5807 => x"982b5473",
          5808 => x"80258c38",
          5809 => x"7580ff06",
          5810 => x"81ebdc11",
          5811 => x"33575475",
          5812 => x"51e6e13f",
          5813 => x"81fef008",
          5814 => x"802eb238",
          5815 => x"78187033",
          5816 => x"811a7154",
          5817 => x"5a5654e6",
          5818 => x"d23f81fe",
          5819 => x"f008802e",
          5820 => x"80e838ff",
          5821 => x"1c547674",
          5822 => x"2780df38",
          5823 => x"79175475",
          5824 => x"74348117",
          5825 => x"7a115557",
          5826 => x"747434a7",
          5827 => x"39755281",
          5828 => x"eafc51e5",
          5829 => x"fe3f81fe",
          5830 => x"f008bf38",
          5831 => x"ff9f1654",
          5832 => x"73992689",
          5833 => x"38e01670",
          5834 => x"81ff0657",
          5835 => x"54791754",
          5836 => x"75743481",
          5837 => x"1757fdf7",
          5838 => x"3977197e",
          5839 => x"0c76802e",
          5840 => x"99387933",
          5841 => x"547381e5",
          5842 => x"2e098106",
          5843 => x"8438857a",
          5844 => x"348454a0",
          5845 => x"76278f38",
          5846 => x"8b398655",
          5847 => x"81f23984",
          5848 => x"5680f339",
          5849 => x"8054738b",
          5850 => x"1b34807b",
          5851 => x"0858527a",
          5852 => x"51f2ce3f",
          5853 => x"81fef008",
          5854 => x"5681fef0",
          5855 => x"0880d738",
          5856 => x"981b0852",
          5857 => x"7651e6aa",
          5858 => x"3f81fef0",
          5859 => x"085681fe",
          5860 => x"f00880c2",
          5861 => x"389c1b08",
          5862 => x"70335555",
          5863 => x"73802eff",
          5864 => x"be388b15",
          5865 => x"33bf0654",
          5866 => x"73861c34",
          5867 => x"8b153370",
          5868 => x"832a7081",
          5869 => x"06515558",
          5870 => x"7392388b",
          5871 => x"53795274",
          5872 => x"51e49f3f",
          5873 => x"81fef008",
          5874 => x"802e8b38",
          5875 => x"75527a51",
          5876 => x"f3ba3fff",
          5877 => x"9f3975ab",
          5878 => x"1c335755",
          5879 => x"74802ebb",
          5880 => x"3874842e",
          5881 => x"09810680",
          5882 => x"e7387585",
          5883 => x"2a708106",
          5884 => x"77822a58",
          5885 => x"51547380",
          5886 => x"2e963875",
          5887 => x"81065473",
          5888 => x"802efbb5",
          5889 => x"38ff800b",
          5890 => x"ab1c3480",
          5891 => x"5580c139",
          5892 => x"75810654",
          5893 => x"73ba3885",
          5894 => x"55b63975",
          5895 => x"822a7081",
          5896 => x"06515473",
          5897 => x"ab38861b",
          5898 => x"3370842a",
          5899 => x"70810651",
          5900 => x"55557380",
          5901 => x"2ee13890",
          5902 => x"1b0883ff",
          5903 => x"061db405",
          5904 => x"527c51f5",
          5905 => x"db3f81fe",
          5906 => x"f008881c",
          5907 => x"0cfaea39",
          5908 => x"7481fef0",
          5909 => x"0c8f3d0d",
          5910 => x"04f63d0d",
          5911 => x"7c5bff7b",
          5912 => x"08707173",
          5913 => x"55595c55",
          5914 => x"5973802e",
          5915 => x"81c63875",
          5916 => x"70810557",
          5917 => x"3370a026",
          5918 => x"525271ba",
          5919 => x"2e8d3870",
          5920 => x"ee3871ba",
          5921 => x"2e098106",
          5922 => x"81a53873",
          5923 => x"33d01170",
          5924 => x"81ff0651",
          5925 => x"52537089",
          5926 => x"26913882",
          5927 => x"147381ff",
          5928 => x"06d00556",
          5929 => x"5271762e",
          5930 => x"80f73880",
          5931 => x"0b81ebcc",
          5932 => x"59557708",
          5933 => x"7a555776",
          5934 => x"70810558",
          5935 => x"33747081",
          5936 => x"055633ff",
          5937 => x"9f125353",
          5938 => x"53709926",
          5939 => x"8938e013",
          5940 => x"7081ff06",
          5941 => x"5451ff9f",
          5942 => x"12517099",
          5943 => x"268938e0",
          5944 => x"127081ff",
          5945 => x"06535172",
          5946 => x"30709f2a",
          5947 => x"51517272",
          5948 => x"2e098106",
          5949 => x"853870ff",
          5950 => x"be387230",
          5951 => x"74773270",
          5952 => x"30707207",
          5953 => x"9f2a739f",
          5954 => x"2a075354",
          5955 => x"54517080",
          5956 => x"2e8f3881",
          5957 => x"15841959",
          5958 => x"55837525",
          5959 => x"ff94388b",
          5960 => x"39748324",
          5961 => x"86387476",
          5962 => x"7c0c5978",
          5963 => x"51863981",
          5964 => x"ffb43351",
          5965 => x"7081fef0",
          5966 => x"0c8c3d0d",
          5967 => x"04fa3d0d",
          5968 => x"7856800b",
          5969 => x"831734ff",
          5970 => x"0bb0170c",
          5971 => x"79527551",
          5972 => x"e2e03f84",
          5973 => x"5581fef0",
          5974 => x"08818038",
          5975 => x"84b21651",
          5976 => x"dfb43f81",
          5977 => x"fef00883",
          5978 => x"ffff0654",
          5979 => x"83557382",
          5980 => x"d4d52e09",
          5981 => x"810680e3",
          5982 => x"38800bb4",
          5983 => x"17335657",
          5984 => x"7481e92e",
          5985 => x"09810683",
          5986 => x"38815774",
          5987 => x"81eb3270",
          5988 => x"30708025",
          5989 => x"79075151",
          5990 => x"54738a38",
          5991 => x"7481e82e",
          5992 => x"098106b5",
          5993 => x"38835381",
          5994 => x"eb8c5280",
          5995 => x"ea1651e0",
          5996 => x"b13f81fe",
          5997 => x"f0085581",
          5998 => x"fef00880",
          5999 => x"2e9d3885",
          6000 => x"5381eb90",
          6001 => x"52818616",
          6002 => x"51e0973f",
          6003 => x"81fef008",
          6004 => x"5581fef0",
          6005 => x"08802e83",
          6006 => x"38825574",
          6007 => x"81fef00c",
          6008 => x"883d0d04",
          6009 => x"f23d0d61",
          6010 => x"02840580",
          6011 => x"cb053358",
          6012 => x"5580750c",
          6013 => x"6051fce1",
          6014 => x"3f81fef0",
          6015 => x"08588b56",
          6016 => x"800b81fe",
          6017 => x"f0082486",
          6018 => x"fc3881fe",
          6019 => x"f0088429",
          6020 => x"81ffa005",
          6021 => x"70085553",
          6022 => x"8c567380",
          6023 => x"2e86e638",
          6024 => x"73750c76",
          6025 => x"81fe0674",
          6026 => x"33545772",
          6027 => x"802eae38",
          6028 => x"81143351",
          6029 => x"d7ca3f81",
          6030 => x"fef00881",
          6031 => x"ff067081",
          6032 => x"06545572",
          6033 => x"98387680",
          6034 => x"2e86b838",
          6035 => x"74822a70",
          6036 => x"81065153",
          6037 => x"8a567286",
          6038 => x"ac3886a7",
          6039 => x"39807434",
          6040 => x"77811534",
          6041 => x"81528114",
          6042 => x"3351d7b2",
          6043 => x"3f81fef0",
          6044 => x"0881ff06",
          6045 => x"70810654",
          6046 => x"55835672",
          6047 => x"86873876",
          6048 => x"802e8f38",
          6049 => x"74822a70",
          6050 => x"81065153",
          6051 => x"8a567285",
          6052 => x"f4388070",
          6053 => x"5374525b",
          6054 => x"fda33f81",
          6055 => x"fef00881",
          6056 => x"ff065776",
          6057 => x"822e0981",
          6058 => x"0680e238",
          6059 => x"8c3d7456",
          6060 => x"58835683",
          6061 => x"f6153370",
          6062 => x"58537280",
          6063 => x"2e8d3883",
          6064 => x"fa1551dc",
          6065 => x"e83f81fe",
          6066 => x"f0085776",
          6067 => x"78708405",
          6068 => x"5a0cff16",
          6069 => x"90165656",
          6070 => x"758025d7",
          6071 => x"38800b8d",
          6072 => x"3d545672",
          6073 => x"70840554",
          6074 => x"085b8357",
          6075 => x"7a802e95",
          6076 => x"387a5273",
          6077 => x"51fcc63f",
          6078 => x"81fef008",
          6079 => x"81ff0657",
          6080 => x"81772789",
          6081 => x"38811656",
          6082 => x"837627d7",
          6083 => x"38815676",
          6084 => x"842e84f1",
          6085 => x"388d5676",
          6086 => x"812684e9",
          6087 => x"38bf1451",
          6088 => x"dbf43f81",
          6089 => x"fef00883",
          6090 => x"ffff0653",
          6091 => x"7284802e",
          6092 => x"09810684",
          6093 => x"d03880ca",
          6094 => x"1451dbda",
          6095 => x"3f81fef0",
          6096 => x"0883ffff",
          6097 => x"0658778d",
          6098 => x"3880d814",
          6099 => x"51dbde3f",
          6100 => x"81fef008",
          6101 => x"58779c15",
          6102 => x"0c80c414",
          6103 => x"33821534",
          6104 => x"80c41433",
          6105 => x"ff117081",
          6106 => x"ff065154",
          6107 => x"558d5672",
          6108 => x"81268491",
          6109 => x"387481ff",
          6110 => x"06787129",
          6111 => x"80c11633",
          6112 => x"52595372",
          6113 => x"8a152372",
          6114 => x"802e8b38",
          6115 => x"ff137306",
          6116 => x"5372802e",
          6117 => x"86388d56",
          6118 => x"83eb3980",
          6119 => x"c51451da",
          6120 => x"f53f81fe",
          6121 => x"f0085381",
          6122 => x"fef00888",
          6123 => x"1523728f",
          6124 => x"06578d56",
          6125 => x"7683ce38",
          6126 => x"80c71451",
          6127 => x"dad83f81",
          6128 => x"fef00883",
          6129 => x"ffff0655",
          6130 => x"748d3880",
          6131 => x"d41451da",
          6132 => x"dc3f81fe",
          6133 => x"f0085580",
          6134 => x"c21451da",
          6135 => x"b93f81fe",
          6136 => x"f00883ff",
          6137 => x"ff06538d",
          6138 => x"5672802e",
          6139 => x"83973888",
          6140 => x"14227814",
          6141 => x"71842a05",
          6142 => x"5a5a7875",
          6143 => x"26838638",
          6144 => x"8a142252",
          6145 => x"74793151",
          6146 => x"ff93a03f",
          6147 => x"81fef008",
          6148 => x"5581fef0",
          6149 => x"08802e82",
          6150 => x"ec3881fe",
          6151 => x"f00880ff",
          6152 => x"fffff526",
          6153 => x"83388357",
          6154 => x"7483fff5",
          6155 => x"26833882",
          6156 => x"57749ff5",
          6157 => x"26853881",
          6158 => x"5789398d",
          6159 => x"5676802e",
          6160 => x"82c33882",
          6161 => x"15709816",
          6162 => x"0c7ba016",
          6163 => x"0c731c70",
          6164 => x"a4170c7a",
          6165 => x"1dac170c",
          6166 => x"54557683",
          6167 => x"2e098106",
          6168 => x"af3880de",
          6169 => x"1451d9ae",
          6170 => x"3f81fef0",
          6171 => x"0883ffff",
          6172 => x"06538d56",
          6173 => x"72828e38",
          6174 => x"79828a38",
          6175 => x"80e01451",
          6176 => x"d9ab3f81",
          6177 => x"fef008a8",
          6178 => x"150c7482",
          6179 => x"2b53a239",
          6180 => x"8d567980",
          6181 => x"2e81ee38",
          6182 => x"7713a815",
          6183 => x"0c741553",
          6184 => x"76822e8d",
          6185 => x"38741015",
          6186 => x"70812a76",
          6187 => x"81060551",
          6188 => x"5383ff13",
          6189 => x"892a538d",
          6190 => x"56729c15",
          6191 => x"082681c5",
          6192 => x"38ff0b90",
          6193 => x"150cff0b",
          6194 => x"8c150cff",
          6195 => x"800b8415",
          6196 => x"3476832e",
          6197 => x"09810681",
          6198 => x"923880e4",
          6199 => x"1451d8b6",
          6200 => x"3f81fef0",
          6201 => x"0883ffff",
          6202 => x"06537281",
          6203 => x"2e098106",
          6204 => x"80f93881",
          6205 => x"1b527351",
          6206 => x"dbb83f81",
          6207 => x"fef00880",
          6208 => x"ea3881fe",
          6209 => x"f0088415",
          6210 => x"3484b214",
          6211 => x"51d8873f",
          6212 => x"81fef008",
          6213 => x"83ffff06",
          6214 => x"537282d4",
          6215 => x"d52e0981",
          6216 => x"0680c838",
          6217 => x"b41451d8",
          6218 => x"843f81fe",
          6219 => x"f008848b",
          6220 => x"85a4d22e",
          6221 => x"098106b3",
          6222 => x"38849814",
          6223 => x"51d7ee3f",
          6224 => x"81fef008",
          6225 => x"868a85e4",
          6226 => x"f22e0981",
          6227 => x"069d3884",
          6228 => x"9c1451d7",
          6229 => x"d83f81fe",
          6230 => x"f0089015",
          6231 => x"0c84a014",
          6232 => x"51d7ca3f",
          6233 => x"81fef008",
          6234 => x"8c150c76",
          6235 => x"743481ff",
          6236 => x"b0228105",
          6237 => x"537281ff",
          6238 => x"b0237286",
          6239 => x"1523800b",
          6240 => x"94150c80",
          6241 => x"567581fe",
          6242 => x"f00c903d",
          6243 => x"0d04fb3d",
          6244 => x"0d775489",
          6245 => x"5573802e",
          6246 => x"b9387308",
          6247 => x"5372802e",
          6248 => x"b1387233",
          6249 => x"5271802e",
          6250 => x"a9388613",
          6251 => x"22841522",
          6252 => x"57527176",
          6253 => x"2e098106",
          6254 => x"99388113",
          6255 => x"3351d0c0",
          6256 => x"3f81fef0",
          6257 => x"08810652",
          6258 => x"71883871",
          6259 => x"74085455",
          6260 => x"83398053",
          6261 => x"7873710c",
          6262 => x"527481fe",
          6263 => x"f00c873d",
          6264 => x"0d04fa3d",
          6265 => x"0d02ab05",
          6266 => x"337a5889",
          6267 => x"3dfc0552",
          6268 => x"56f4e63f",
          6269 => x"8b54800b",
          6270 => x"81fef008",
          6271 => x"24bc3881",
          6272 => x"fef00884",
          6273 => x"2981ffa0",
          6274 => x"05700855",
          6275 => x"5573802e",
          6276 => x"84388074",
          6277 => x"34785473",
          6278 => x"802e8438",
          6279 => x"80743478",
          6280 => x"750c7554",
          6281 => x"75802e92",
          6282 => x"38805389",
          6283 => x"3d705384",
          6284 => x"0551f7b0",
          6285 => x"3f81fef0",
          6286 => x"08547381",
          6287 => x"fef00c88",
          6288 => x"3d0d04eb",
          6289 => x"3d0d6702",
          6290 => x"840580e7",
          6291 => x"05335959",
          6292 => x"89547880",
          6293 => x"2e84c838",
          6294 => x"77bf0670",
          6295 => x"54983dd0",
          6296 => x"0553993d",
          6297 => x"84055258",
          6298 => x"f6fa3f81",
          6299 => x"fef00855",
          6300 => x"81fef008",
          6301 => x"84a4387a",
          6302 => x"5c68528c",
          6303 => x"3d705256",
          6304 => x"edc63f81",
          6305 => x"fef00855",
          6306 => x"81fef008",
          6307 => x"92380280",
          6308 => x"d7053370",
          6309 => x"982b5557",
          6310 => x"73802583",
          6311 => x"38865577",
          6312 => x"9c065473",
          6313 => x"802e81ab",
          6314 => x"3874802e",
          6315 => x"95387484",
          6316 => x"2e098106",
          6317 => x"aa387551",
          6318 => x"eaf83f81",
          6319 => x"fef00855",
          6320 => x"9e3902b2",
          6321 => x"05339106",
          6322 => x"547381b8",
          6323 => x"3877822a",
          6324 => x"70810651",
          6325 => x"5473802e",
          6326 => x"8e388855",
          6327 => x"83bc3977",
          6328 => x"88075874",
          6329 => x"83b43877",
          6330 => x"832a7081",
          6331 => x"06515473",
          6332 => x"802e81af",
          6333 => x"3862527a",
          6334 => x"51e8a53f",
          6335 => x"81fef008",
          6336 => x"568288b2",
          6337 => x"0a52628e",
          6338 => x"0551d4ea",
          6339 => x"3f6254a0",
          6340 => x"0b8b1534",
          6341 => x"80536252",
          6342 => x"7a51e8bd",
          6343 => x"3f805262",
          6344 => x"9c0551d4",
          6345 => x"d13f7a54",
          6346 => x"810b8315",
          6347 => x"3475802e",
          6348 => x"80f1387a",
          6349 => x"b0110851",
          6350 => x"54805375",
          6351 => x"52973dd4",
          6352 => x"0551ddbe",
          6353 => x"3f81fef0",
          6354 => x"085581fe",
          6355 => x"f00882ca",
          6356 => x"38b73974",
          6357 => x"82c43802",
          6358 => x"b2053370",
          6359 => x"842a7081",
          6360 => x"06515556",
          6361 => x"73802e86",
          6362 => x"38845582",
          6363 => x"ad397781",
          6364 => x"2a708106",
          6365 => x"51547380",
          6366 => x"2ea93875",
          6367 => x"81065473",
          6368 => x"802ea038",
          6369 => x"87558292",
          6370 => x"3973527a",
          6371 => x"51d6a33f",
          6372 => x"81fef008",
          6373 => x"7bff188c",
          6374 => x"120c5555",
          6375 => x"81fef008",
          6376 => x"81f83877",
          6377 => x"832a7081",
          6378 => x"06515473",
          6379 => x"802e8638",
          6380 => x"7780c007",
          6381 => x"587ab011",
          6382 => x"08a01b0c",
          6383 => x"63a41b0c",
          6384 => x"63537052",
          6385 => x"57e6d93f",
          6386 => x"81fef008",
          6387 => x"81fef008",
          6388 => x"881b0c63",
          6389 => x"9c05525a",
          6390 => x"d2d33f81",
          6391 => x"fef00881",
          6392 => x"fef0088c",
          6393 => x"1b0c777a",
          6394 => x"0c568617",
          6395 => x"22841a23",
          6396 => x"77901a34",
          6397 => x"800b911a",
          6398 => x"34800b9c",
          6399 => x"1a0c800b",
          6400 => x"941a0c77",
          6401 => x"852a7081",
          6402 => x"06515473",
          6403 => x"802e818d",
          6404 => x"3881fef0",
          6405 => x"08802e81",
          6406 => x"843881fe",
          6407 => x"f008941a",
          6408 => x"0c8a1722",
          6409 => x"70892b7b",
          6410 => x"525957a8",
          6411 => x"39765278",
          6412 => x"51d79f3f",
          6413 => x"81fef008",
          6414 => x"5781fef0",
          6415 => x"08812683",
          6416 => x"38825581",
          6417 => x"fef008ff",
          6418 => x"2e098106",
          6419 => x"83387955",
          6420 => x"75783156",
          6421 => x"74307076",
          6422 => x"07802551",
          6423 => x"54777627",
          6424 => x"8a388170",
          6425 => x"7506555a",
          6426 => x"73c33876",
          6427 => x"981a0c74",
          6428 => x"a9387583",
          6429 => x"ff065473",
          6430 => x"802ea238",
          6431 => x"76527a51",
          6432 => x"d6a63f81",
          6433 => x"fef00885",
          6434 => x"3882558e",
          6435 => x"3975892a",
          6436 => x"81fef008",
          6437 => x"059c1a0c",
          6438 => x"84398079",
          6439 => x"0c745473",
          6440 => x"81fef00c",
          6441 => x"973d0d04",
          6442 => x"f23d0d60",
          6443 => x"63656440",
          6444 => x"405d5980",
          6445 => x"7e0c903d",
          6446 => x"fc055278",
          6447 => x"51f9cf3f",
          6448 => x"81fef008",
          6449 => x"5581fef0",
          6450 => x"088a3891",
          6451 => x"19335574",
          6452 => x"802e8638",
          6453 => x"745682c4",
          6454 => x"39901933",
          6455 => x"81065587",
          6456 => x"5674802e",
          6457 => x"82b63895",
          6458 => x"39820b91",
          6459 => x"1a348256",
          6460 => x"82aa3981",
          6461 => x"0b911a34",
          6462 => x"815682a0",
          6463 => x"398c1908",
          6464 => x"941a0831",
          6465 => x"55747c27",
          6466 => x"8338745c",
          6467 => x"7b802e82",
          6468 => x"89389419",
          6469 => x"087083ff",
          6470 => x"06565674",
          6471 => x"81b2387e",
          6472 => x"8a1122ff",
          6473 => x"0577892a",
          6474 => x"065b5579",
          6475 => x"a8387587",
          6476 => x"38881908",
          6477 => x"558f3998",
          6478 => x"19085278",
          6479 => x"51d5933f",
          6480 => x"81fef008",
          6481 => x"55817527",
          6482 => x"ff9f3874",
          6483 => x"ff2effa3",
          6484 => x"3874981a",
          6485 => x"0c981908",
          6486 => x"527e51d4",
          6487 => x"cb3f81fe",
          6488 => x"f008802e",
          6489 => x"ff833881",
          6490 => x"fef0081a",
          6491 => x"7c892a59",
          6492 => x"5777802e",
          6493 => x"80d63877",
          6494 => x"1a7f8a11",
          6495 => x"22585c55",
          6496 => x"75752785",
          6497 => x"38757a31",
          6498 => x"58775476",
          6499 => x"537c5281",
          6500 => x"1b3351ca",
          6501 => x"883f81fe",
          6502 => x"f008fed7",
          6503 => x"387e8311",
          6504 => x"33565674",
          6505 => x"802e9f38",
          6506 => x"b0160877",
          6507 => x"31557478",
          6508 => x"27943884",
          6509 => x"8053b416",
          6510 => x"52b01608",
          6511 => x"7731892b",
          6512 => x"7d0551cf",
          6513 => x"e03f7789",
          6514 => x"2b56b939",
          6515 => x"769c1a0c",
          6516 => x"94190883",
          6517 => x"ff068480",
          6518 => x"71315755",
          6519 => x"7b762783",
          6520 => x"387b569c",
          6521 => x"1908527e",
          6522 => x"51d1c73f",
          6523 => x"81fef008",
          6524 => x"fe813875",
          6525 => x"53941908",
          6526 => x"83ff061f",
          6527 => x"b405527c",
          6528 => x"51cfa23f",
          6529 => x"7b76317e",
          6530 => x"08177f0c",
          6531 => x"761e941b",
          6532 => x"0818941c",
          6533 => x"0c5e5cfd",
          6534 => x"f3398056",
          6535 => x"7581fef0",
          6536 => x"0c903d0d",
          6537 => x"04f23d0d",
          6538 => x"60636564",
          6539 => x"40405d58",
          6540 => x"807e0c90",
          6541 => x"3dfc0552",
          6542 => x"7751f6d2",
          6543 => x"3f81fef0",
          6544 => x"085581fe",
          6545 => x"f0088a38",
          6546 => x"91183355",
          6547 => x"74802e86",
          6548 => x"38745683",
          6549 => x"b8399018",
          6550 => x"3370812a",
          6551 => x"70810651",
          6552 => x"56568756",
          6553 => x"74802e83",
          6554 => x"a4389539",
          6555 => x"820b9119",
          6556 => x"34825683",
          6557 => x"9839810b",
          6558 => x"91193481",
          6559 => x"56838e39",
          6560 => x"9418087c",
          6561 => x"11565674",
          6562 => x"76278438",
          6563 => x"75095c7b",
          6564 => x"802e82ec",
          6565 => x"38941808",
          6566 => x"7083ff06",
          6567 => x"56567481",
          6568 => x"fd387e8a",
          6569 => x"1122ff05",
          6570 => x"77892a06",
          6571 => x"5c557abf",
          6572 => x"38758c38",
          6573 => x"88180855",
          6574 => x"749c387a",
          6575 => x"52853998",
          6576 => x"18085277",
          6577 => x"51d7e73f",
          6578 => x"81fef008",
          6579 => x"5581fef0",
          6580 => x"08802e82",
          6581 => x"ab387481",
          6582 => x"2eff9138",
          6583 => x"74ff2eff",
          6584 => x"95387498",
          6585 => x"190c8818",
          6586 => x"08853874",
          6587 => x"88190c7e",
          6588 => x"55b01508",
          6589 => x"9c19082e",
          6590 => x"0981068d",
          6591 => x"387451ce",
          6592 => x"c13f81fe",
          6593 => x"f008feee",
          6594 => x"38981808",
          6595 => x"527e51d1",
          6596 => x"973f81fe",
          6597 => x"f008802e",
          6598 => x"fed23881",
          6599 => x"fef0081b",
          6600 => x"7c892a5a",
          6601 => x"5778802e",
          6602 => x"80d53878",
          6603 => x"1b7f8a11",
          6604 => x"22585b55",
          6605 => x"75752785",
          6606 => x"38757b31",
          6607 => x"59785476",
          6608 => x"537c5281",
          6609 => x"1a3351c8",
          6610 => x"be3f81fe",
          6611 => x"f008fea6",
          6612 => x"387eb011",
          6613 => x"08783156",
          6614 => x"56747927",
          6615 => x"9b388480",
          6616 => x"53b01608",
          6617 => x"7731892b",
          6618 => x"7d0552b4",
          6619 => x"1651ccb5",
          6620 => x"3f7e5580",
          6621 => x"0b831634",
          6622 => x"78892b56",
          6623 => x"80db398c",
          6624 => x"18089419",
          6625 => x"08269338",
          6626 => x"7e51cdb6",
          6627 => x"3f81fef0",
          6628 => x"08fde338",
          6629 => x"7e77b012",
          6630 => x"0c55769c",
          6631 => x"190c9418",
          6632 => x"0883ff06",
          6633 => x"84807131",
          6634 => x"57557b76",
          6635 => x"2783387b",
          6636 => x"569c1808",
          6637 => x"527e51cd",
          6638 => x"f93f81fe",
          6639 => x"f008fdb6",
          6640 => x"3875537c",
          6641 => x"52941808",
          6642 => x"83ff061f",
          6643 => x"b40551cb",
          6644 => x"d43f7e55",
          6645 => x"810b8316",
          6646 => x"347b7631",
          6647 => x"7e08177f",
          6648 => x"0c761e94",
          6649 => x"1a081870",
          6650 => x"941c0c8c",
          6651 => x"1b085858",
          6652 => x"5e5c7476",
          6653 => x"27833875",
          6654 => x"55748c19",
          6655 => x"0cfd9039",
          6656 => x"90183380",
          6657 => x"c0075574",
          6658 => x"90193480",
          6659 => x"567581fe",
          6660 => x"f00c903d",
          6661 => x"0d04f83d",
          6662 => x"0d7a8b3d",
          6663 => x"fc055370",
          6664 => x"5256f2ea",
          6665 => x"3f81fef0",
          6666 => x"085781fe",
          6667 => x"f00880fb",
          6668 => x"38901633",
          6669 => x"70862a70",
          6670 => x"81065155",
          6671 => x"5573802e",
          6672 => x"80e938a0",
          6673 => x"16085278",
          6674 => x"51cce73f",
          6675 => x"81fef008",
          6676 => x"5781fef0",
          6677 => x"0880d438",
          6678 => x"a416088b",
          6679 => x"1133a007",
          6680 => x"5555738b",
          6681 => x"16348816",
          6682 => x"08537452",
          6683 => x"750851dd",
          6684 => x"e83f8c16",
          6685 => x"08529c15",
          6686 => x"51c9fb3f",
          6687 => x"8288b20a",
          6688 => x"52961551",
          6689 => x"c9f03f76",
          6690 => x"52921551",
          6691 => x"c9ca3f78",
          6692 => x"54810b83",
          6693 => x"15347851",
          6694 => x"ccdf3f81",
          6695 => x"fef00890",
          6696 => x"173381bf",
          6697 => x"06555773",
          6698 => x"90173476",
          6699 => x"81fef00c",
          6700 => x"8a3d0d04",
          6701 => x"fc3d0d76",
          6702 => x"705254fe",
          6703 => x"d93f81fe",
          6704 => x"f0085381",
          6705 => x"fef0089c",
          6706 => x"38863dfc",
          6707 => x"05527351",
          6708 => x"f1bc3f81",
          6709 => x"fef00853",
          6710 => x"81fef008",
          6711 => x"873881fe",
          6712 => x"f008740c",
          6713 => x"7281fef0",
          6714 => x"0c863d0d",
          6715 => x"04ff3d0d",
          6716 => x"843d51e6",
          6717 => x"e43f8b52",
          6718 => x"800b81fe",
          6719 => x"f008248b",
          6720 => x"3881fef0",
          6721 => x"0881ffb4",
          6722 => x"34805271",
          6723 => x"81fef00c",
          6724 => x"833d0d04",
          6725 => x"ef3d0d80",
          6726 => x"53933dd0",
          6727 => x"0552943d",
          6728 => x"51e9c13f",
          6729 => x"81fef008",
          6730 => x"5581fef0",
          6731 => x"0880e038",
          6732 => x"76586352",
          6733 => x"933dd405",
          6734 => x"51e08d3f",
          6735 => x"81fef008",
          6736 => x"5581fef0",
          6737 => x"08bc3802",
          6738 => x"80c70533",
          6739 => x"70982b55",
          6740 => x"56738025",
          6741 => x"8938767a",
          6742 => x"94120c54",
          6743 => x"b23902a2",
          6744 => x"05337084",
          6745 => x"2a708106",
          6746 => x"51555673",
          6747 => x"802e9e38",
          6748 => x"767f5370",
          6749 => x"5254dba8",
          6750 => x"3f81fef0",
          6751 => x"0894150c",
          6752 => x"8e3981fe",
          6753 => x"f008842e",
          6754 => x"09810683",
          6755 => x"38855574",
          6756 => x"81fef00c",
          6757 => x"933d0d04",
          6758 => x"e43d0d6f",
          6759 => x"6f5b5b80",
          6760 => x"7a348053",
          6761 => x"9e3dffb8",
          6762 => x"05529f3d",
          6763 => x"51e8b53f",
          6764 => x"81fef008",
          6765 => x"5781fef0",
          6766 => x"0882fc38",
          6767 => x"7b437a7c",
          6768 => x"94110847",
          6769 => x"55586454",
          6770 => x"73802e81",
          6771 => x"ed38a052",
          6772 => x"933d7052",
          6773 => x"55d5ea3f",
          6774 => x"81fef008",
          6775 => x"5781fef0",
          6776 => x"0882d438",
          6777 => x"68527b51",
          6778 => x"c9c83f81",
          6779 => x"fef00857",
          6780 => x"81fef008",
          6781 => x"82c13869",
          6782 => x"527b51da",
          6783 => x"a33f81fe",
          6784 => x"f0084576",
          6785 => x"527451d5",
          6786 => x"b83f81fe",
          6787 => x"f0085781",
          6788 => x"fef00882",
          6789 => x"a2388052",
          6790 => x"7451daeb",
          6791 => x"3f81fef0",
          6792 => x"085781fe",
          6793 => x"f008a438",
          6794 => x"69527b51",
          6795 => x"d9f23f73",
          6796 => x"81fef008",
          6797 => x"2ea63876",
          6798 => x"527451d6",
          6799 => x"cf3f81fe",
          6800 => x"f0085781",
          6801 => x"fef00880",
          6802 => x"2ecc3876",
          6803 => x"842e0981",
          6804 => x"06863882",
          6805 => x"5781e039",
          6806 => x"7681dc38",
          6807 => x"9e3dffbc",
          6808 => x"05527451",
          6809 => x"dcc93f76",
          6810 => x"903d7811",
          6811 => x"81113351",
          6812 => x"565a5673",
          6813 => x"802e9138",
          6814 => x"02b90555",
          6815 => x"81168116",
          6816 => x"70335656",
          6817 => x"5673f538",
          6818 => x"81165473",
          6819 => x"78268190",
          6820 => x"3875802e",
          6821 => x"99387816",
          6822 => x"810555ff",
          6823 => x"186f11ff",
          6824 => x"18ff1858",
          6825 => x"58555874",
          6826 => x"33743475",
          6827 => x"ee38ff18",
          6828 => x"6f115558",
          6829 => x"af7434fe",
          6830 => x"8d39777b",
          6831 => x"2e098106",
          6832 => x"8a38ff18",
          6833 => x"6f115558",
          6834 => x"af743480",
          6835 => x"0b81ffb4",
          6836 => x"33708429",
          6837 => x"81ebcc05",
          6838 => x"70087033",
          6839 => x"525c5656",
          6840 => x"5673762e",
          6841 => x"8d388116",
          6842 => x"701a7033",
          6843 => x"51555673",
          6844 => x"f5388216",
          6845 => x"54737826",
          6846 => x"a7388055",
          6847 => x"74762791",
          6848 => x"38741954",
          6849 => x"73337a70",
          6850 => x"81055c34",
          6851 => x"811555ec",
          6852 => x"39ba7a70",
          6853 => x"81055c34",
          6854 => x"74ff2e09",
          6855 => x"81068538",
          6856 => x"91579439",
          6857 => x"6e188119",
          6858 => x"59547333",
          6859 => x"7a708105",
          6860 => x"5c347a78",
          6861 => x"26ee3880",
          6862 => x"7a347681",
          6863 => x"fef00c9e",
          6864 => x"3d0d04f7",
          6865 => x"3d0d7b7d",
          6866 => x"8d3dfc05",
          6867 => x"54715357",
          6868 => x"55ecbb3f",
          6869 => x"81fef008",
          6870 => x"5381fef0",
          6871 => x"0882fa38",
          6872 => x"91153353",
          6873 => x"7282f238",
          6874 => x"8c150854",
          6875 => x"73762792",
          6876 => x"38901533",
          6877 => x"70812a70",
          6878 => x"81065154",
          6879 => x"57728338",
          6880 => x"73569415",
          6881 => x"08548070",
          6882 => x"94170c58",
          6883 => x"75782e82",
          6884 => x"9738798a",
          6885 => x"11227089",
          6886 => x"2b595153",
          6887 => x"73782eb7",
          6888 => x"387652ff",
          6889 => x"1651fefc",
          6890 => x"823f81fe",
          6891 => x"f008ff15",
          6892 => x"78547053",
          6893 => x"5553fefb",
          6894 => x"f23f81fe",
          6895 => x"f0087326",
          6896 => x"96387630",
          6897 => x"70750670",
          6898 => x"94180c77",
          6899 => x"71319818",
          6900 => x"08575851",
          6901 => x"53b13988",
          6902 => x"15085473",
          6903 => x"a6387352",
          6904 => x"7451cdca",
          6905 => x"3f81fef0",
          6906 => x"085481fe",
          6907 => x"f008812e",
          6908 => x"819a3881",
          6909 => x"fef008ff",
          6910 => x"2e819b38",
          6911 => x"81fef008",
          6912 => x"88160c73",
          6913 => x"98160c73",
          6914 => x"802e819c",
          6915 => x"38767627",
          6916 => x"80dc3875",
          6917 => x"77319416",
          6918 => x"08189417",
          6919 => x"0c901633",
          6920 => x"70812a70",
          6921 => x"81065155",
          6922 => x"5a567280",
          6923 => x"2e9a3873",
          6924 => x"527451cc",
          6925 => x"f93f81fe",
          6926 => x"f0085481",
          6927 => x"fef00894",
          6928 => x"3881fef0",
          6929 => x"0856a739",
          6930 => x"73527451",
          6931 => x"c7843f81",
          6932 => x"fef00854",
          6933 => x"73ff2ebe",
          6934 => x"38817427",
          6935 => x"af387953",
          6936 => x"73981408",
          6937 => x"27a63873",
          6938 => x"98160cff",
          6939 => x"a0399415",
          6940 => x"08169416",
          6941 => x"0c7583ff",
          6942 => x"06537280",
          6943 => x"2eaa3873",
          6944 => x"527951c6",
          6945 => x"a33f81fe",
          6946 => x"f0089438",
          6947 => x"820b9116",
          6948 => x"34825380",
          6949 => x"c439810b",
          6950 => x"91163481",
          6951 => x"53bb3975",
          6952 => x"892a81fe",
          6953 => x"f0080558",
          6954 => x"94150854",
          6955 => x"8c150874",
          6956 => x"27903873",
          6957 => x"8c160c90",
          6958 => x"153380c0",
          6959 => x"07537290",
          6960 => x"16347383",
          6961 => x"ff065372",
          6962 => x"802e8c38",
          6963 => x"779c1608",
          6964 => x"2e853877",
          6965 => x"9c160c80",
          6966 => x"537281fe",
          6967 => x"f00c8b3d",
          6968 => x"0d04f93d",
          6969 => x"0d795689",
          6970 => x"5475802e",
          6971 => x"818a3880",
          6972 => x"53893dfc",
          6973 => x"05528a3d",
          6974 => x"840551e1",
          6975 => x"e73f81fe",
          6976 => x"f0085581",
          6977 => x"fef00880",
          6978 => x"ea387776",
          6979 => x"0c7a5275",
          6980 => x"51d8b53f",
          6981 => x"81fef008",
          6982 => x"5581fef0",
          6983 => x"0880c338",
          6984 => x"ab163370",
          6985 => x"982b5557",
          6986 => x"807424a2",
          6987 => x"38861633",
          6988 => x"70842a70",
          6989 => x"81065155",
          6990 => x"5773802e",
          6991 => x"ad389c16",
          6992 => x"08527751",
          6993 => x"d3da3f81",
          6994 => x"fef00888",
          6995 => x"170c7754",
          6996 => x"86142284",
          6997 => x"17237452",
          6998 => x"7551cee5",
          6999 => x"3f81fef0",
          7000 => x"08557484",
          7001 => x"2e098106",
          7002 => x"85388555",
          7003 => x"86397480",
          7004 => x"2e843880",
          7005 => x"760c7454",
          7006 => x"7381fef0",
          7007 => x"0c893d0d",
          7008 => x"04fc3d0d",
          7009 => x"76873dfc",
          7010 => x"05537052",
          7011 => x"53e7ff3f",
          7012 => x"81fef008",
          7013 => x"873881fe",
          7014 => x"f008730c",
          7015 => x"863d0d04",
          7016 => x"fb3d0d77",
          7017 => x"79893dfc",
          7018 => x"05547153",
          7019 => x"5654e7de",
          7020 => x"3f81fef0",
          7021 => x"085381fe",
          7022 => x"f00880df",
          7023 => x"38749338",
          7024 => x"81fef008",
          7025 => x"527351cd",
          7026 => x"f83f81fe",
          7027 => x"f0085380",
          7028 => x"ca3981fe",
          7029 => x"f0085273",
          7030 => x"51d3ac3f",
          7031 => x"81fef008",
          7032 => x"5381fef0",
          7033 => x"08842e09",
          7034 => x"81068538",
          7035 => x"80538739",
          7036 => x"81fef008",
          7037 => x"a6387452",
          7038 => x"7351d5b3",
          7039 => x"3f725273",
          7040 => x"51cf893f",
          7041 => x"81fef008",
          7042 => x"84327030",
          7043 => x"7072079f",
          7044 => x"2c7081fe",
          7045 => x"f0080651",
          7046 => x"51545472",
          7047 => x"81fef00c",
          7048 => x"873d0d04",
          7049 => x"ee3d0d65",
          7050 => x"57805389",
          7051 => x"3d705396",
          7052 => x"3d5256df",
          7053 => x"af3f81fe",
          7054 => x"f0085581",
          7055 => x"fef008b2",
          7056 => x"38645275",
          7057 => x"51d6813f",
          7058 => x"81fef008",
          7059 => x"5581fef0",
          7060 => x"08a03802",
          7061 => x"80cb0533",
          7062 => x"70982b55",
          7063 => x"58738025",
          7064 => x"85388655",
          7065 => x"8d397680",
          7066 => x"2e883876",
          7067 => x"527551d4",
          7068 => x"be3f7481",
          7069 => x"fef00c94",
          7070 => x"3d0d04f0",
          7071 => x"3d0d6365",
          7072 => x"555c8053",
          7073 => x"923dec05",
          7074 => x"52933d51",
          7075 => x"ded63f81",
          7076 => x"fef0085b",
          7077 => x"81fef008",
          7078 => x"8280387c",
          7079 => x"740c7308",
          7080 => x"981108fe",
          7081 => x"11901308",
          7082 => x"59565855",
          7083 => x"75742691",
          7084 => x"38757c0c",
          7085 => x"81e43981",
          7086 => x"5b81cc39",
          7087 => x"825b81c7",
          7088 => x"3981fef0",
          7089 => x"08753355",
          7090 => x"5973812e",
          7091 => x"098106bf",
          7092 => x"3882755f",
          7093 => x"57765292",
          7094 => x"3df00551",
          7095 => x"c1f43f81",
          7096 => x"fef008ff",
          7097 => x"2ed13881",
          7098 => x"fef00881",
          7099 => x"2ece3881",
          7100 => x"fef00830",
          7101 => x"7081fef0",
          7102 => x"08078025",
          7103 => x"7a058119",
          7104 => x"7f53595a",
          7105 => x"54981408",
          7106 => x"7726ca38",
          7107 => x"80f939a4",
          7108 => x"150881fe",
          7109 => x"f0085758",
          7110 => x"75983877",
          7111 => x"5281187d",
          7112 => x"5258ffbf",
          7113 => x"8d3f81fe",
          7114 => x"f0085b81",
          7115 => x"fef00880",
          7116 => x"d6387c70",
          7117 => x"337712ff",
          7118 => x"1a5d5256",
          7119 => x"5474822e",
          7120 => x"0981069e",
          7121 => x"38b41451",
          7122 => x"ffbbcb3f",
          7123 => x"81fef008",
          7124 => x"83ffff06",
          7125 => x"70307080",
          7126 => x"251b8219",
          7127 => x"595b5154",
          7128 => x"9b39b414",
          7129 => x"51ffbbc5",
          7130 => x"3f81fef0",
          7131 => x"08f00a06",
          7132 => x"70307080",
          7133 => x"251b8419",
          7134 => x"595b5154",
          7135 => x"7583ff06",
          7136 => x"7a585679",
          7137 => x"ff923878",
          7138 => x"7c0c7c79",
          7139 => x"90120c84",
          7140 => x"11338107",
          7141 => x"56547484",
          7142 => x"15347a81",
          7143 => x"fef00c92",
          7144 => x"3d0d04f9",
          7145 => x"3d0d798a",
          7146 => x"3dfc0553",
          7147 => x"705257e3",
          7148 => x"dd3f81fe",
          7149 => x"f0085681",
          7150 => x"fef00881",
          7151 => x"a8389117",
          7152 => x"33567581",
          7153 => x"a0389017",
          7154 => x"3370812a",
          7155 => x"70810651",
          7156 => x"55558755",
          7157 => x"73802e81",
          7158 => x"8e389417",
          7159 => x"0854738c",
          7160 => x"18082781",
          7161 => x"8038739b",
          7162 => x"3881fef0",
          7163 => x"08538817",
          7164 => x"08527651",
          7165 => x"c48c3f81",
          7166 => x"fef00874",
          7167 => x"88190c56",
          7168 => x"80c93998",
          7169 => x"17085276",
          7170 => x"51ffbfc6",
          7171 => x"3f81fef0",
          7172 => x"08ff2e09",
          7173 => x"81068338",
          7174 => x"815681fe",
          7175 => x"f008812e",
          7176 => x"09810685",
          7177 => x"388256a3",
          7178 => x"3975a038",
          7179 => x"775481fe",
          7180 => x"f0089815",
          7181 => x"08279438",
          7182 => x"98170853",
          7183 => x"81fef008",
          7184 => x"527651c3",
          7185 => x"bd3f81fe",
          7186 => x"f0085694",
          7187 => x"17088c18",
          7188 => x"0c901733",
          7189 => x"80c00754",
          7190 => x"73901834",
          7191 => x"75802e85",
          7192 => x"38759118",
          7193 => x"34755574",
          7194 => x"81fef00c",
          7195 => x"893d0d04",
          7196 => x"e23d0d82",
          7197 => x"53a03dff",
          7198 => x"a40552a1",
          7199 => x"3d51dae4",
          7200 => x"3f81fef0",
          7201 => x"085581fe",
          7202 => x"f00881f5",
          7203 => x"387845a1",
          7204 => x"3d085295",
          7205 => x"3d705258",
          7206 => x"d1ae3f81",
          7207 => x"fef00855",
          7208 => x"81fef008",
          7209 => x"81db3802",
          7210 => x"80fb0533",
          7211 => x"70852a70",
          7212 => x"81065155",
          7213 => x"56865573",
          7214 => x"81c73875",
          7215 => x"982b5480",
          7216 => x"742481bd",
          7217 => x"380280d6",
          7218 => x"05337081",
          7219 => x"06585487",
          7220 => x"557681ad",
          7221 => x"386b5278",
          7222 => x"51ccc53f",
          7223 => x"81fef008",
          7224 => x"74842a70",
          7225 => x"81065155",
          7226 => x"5673802e",
          7227 => x"80d43878",
          7228 => x"5481fef0",
          7229 => x"08941508",
          7230 => x"2e818638",
          7231 => x"735a81fe",
          7232 => x"f0085c76",
          7233 => x"528a3d70",
          7234 => x"5254c7b5",
          7235 => x"3f81fef0",
          7236 => x"085581fe",
          7237 => x"f00880e9",
          7238 => x"3881fef0",
          7239 => x"08527351",
          7240 => x"cce53f81",
          7241 => x"fef00855",
          7242 => x"81fef008",
          7243 => x"86388755",
          7244 => x"80cf3981",
          7245 => x"fef00884",
          7246 => x"2e883881",
          7247 => x"fef00880",
          7248 => x"c0387751",
          7249 => x"cec23f81",
          7250 => x"fef00881",
          7251 => x"fef00830",
          7252 => x"7081fef0",
          7253 => x"08078025",
          7254 => x"51555575",
          7255 => x"802e9438",
          7256 => x"73802e8f",
          7257 => x"38805375",
          7258 => x"527751c1",
          7259 => x"953f81fe",
          7260 => x"f0085574",
          7261 => x"8c387851",
          7262 => x"ffbafe3f",
          7263 => x"81fef008",
          7264 => x"557481fe",
          7265 => x"f00ca03d",
          7266 => x"0d04e93d",
          7267 => x"0d825399",
          7268 => x"3dc00552",
          7269 => x"9a3d51d8",
          7270 => x"cb3f81fe",
          7271 => x"f0085481",
          7272 => x"fef00882",
          7273 => x"b038785e",
          7274 => x"69528e3d",
          7275 => x"705258cf",
          7276 => x"973f81fe",
          7277 => x"f0085481",
          7278 => x"fef00886",
          7279 => x"38885482",
          7280 => x"943981fe",
          7281 => x"f008842e",
          7282 => x"09810682",
          7283 => x"88380280",
          7284 => x"df053370",
          7285 => x"852a8106",
          7286 => x"51558654",
          7287 => x"7481f638",
          7288 => x"785a7452",
          7289 => x"8a3d7052",
          7290 => x"57c1c33f",
          7291 => x"81fef008",
          7292 => x"75555681",
          7293 => x"fef00883",
          7294 => x"38875481",
          7295 => x"fef00881",
          7296 => x"2e098106",
          7297 => x"83388254",
          7298 => x"81fef008",
          7299 => x"ff2e0981",
          7300 => x"06863881",
          7301 => x"5481b439",
          7302 => x"7381b038",
          7303 => x"81fef008",
          7304 => x"527851c4",
          7305 => x"a43f81fe",
          7306 => x"f0085481",
          7307 => x"fef00881",
          7308 => x"9a388b53",
          7309 => x"a052b419",
          7310 => x"51ffb78c",
          7311 => x"3f7854ae",
          7312 => x"0bb41534",
          7313 => x"7854900b",
          7314 => x"bf153482",
          7315 => x"88b20a52",
          7316 => x"80ca1951",
          7317 => x"ffb69f3f",
          7318 => x"755378b4",
          7319 => x"115351c9",
          7320 => x"f83fa053",
          7321 => x"78b41153",
          7322 => x"80d40551",
          7323 => x"ffb6b63f",
          7324 => x"7854ae0b",
          7325 => x"80d51534",
          7326 => x"7f537880",
          7327 => x"d4115351",
          7328 => x"c9d73f78",
          7329 => x"54810b83",
          7330 => x"15347751",
          7331 => x"cba43f81",
          7332 => x"fef00854",
          7333 => x"81fef008",
          7334 => x"b2388288",
          7335 => x"b20a5264",
          7336 => x"960551ff",
          7337 => x"b5d03f75",
          7338 => x"53645278",
          7339 => x"51c9aa3f",
          7340 => x"6454900b",
          7341 => x"8b153478",
          7342 => x"54810b83",
          7343 => x"15347851",
          7344 => x"ffb8b63f",
          7345 => x"81fef008",
          7346 => x"548b3980",
          7347 => x"53755276",
          7348 => x"51ffbeae",
          7349 => x"3f7381fe",
          7350 => x"f00c993d",
          7351 => x"0d04da3d",
          7352 => x"0da93d84",
          7353 => x"0551d2f1",
          7354 => x"3f8253a8",
          7355 => x"3dff8405",
          7356 => x"52a93d51",
          7357 => x"d5ee3f81",
          7358 => x"fef00855",
          7359 => x"81fef008",
          7360 => x"82d33878",
          7361 => x"4da93d08",
          7362 => x"529d3d70",
          7363 => x"5258ccb8",
          7364 => x"3f81fef0",
          7365 => x"085581fe",
          7366 => x"f00882b9",
          7367 => x"3802819b",
          7368 => x"053381a0",
          7369 => x"06548655",
          7370 => x"7382aa38",
          7371 => x"a053a43d",
          7372 => x"0852a83d",
          7373 => x"ff880551",
          7374 => x"ffb4ea3f",
          7375 => x"ac537752",
          7376 => x"923d7052",
          7377 => x"54ffb4dd",
          7378 => x"3faa3d08",
          7379 => x"527351cb",
          7380 => x"f73f81fe",
          7381 => x"f0085581",
          7382 => x"fef00895",
          7383 => x"38636f2e",
          7384 => x"09810688",
          7385 => x"3865a23d",
          7386 => x"082e9238",
          7387 => x"885581e5",
          7388 => x"3981fef0",
          7389 => x"08842e09",
          7390 => x"810681b8",
          7391 => x"387351c9",
          7392 => x"b13f81fe",
          7393 => x"f0085581",
          7394 => x"fef00881",
          7395 => x"c8386856",
          7396 => x"9353a83d",
          7397 => x"ff950552",
          7398 => x"8d1651ff",
          7399 => x"b4873f02",
          7400 => x"af05338b",
          7401 => x"17348b16",
          7402 => x"3370842a",
          7403 => x"70810651",
          7404 => x"55557389",
          7405 => x"3874a007",
          7406 => x"54738b17",
          7407 => x"34785481",
          7408 => x"0b831534",
          7409 => x"8b163370",
          7410 => x"842a7081",
          7411 => x"06515555",
          7412 => x"73802e80",
          7413 => x"e5386e64",
          7414 => x"2e80df38",
          7415 => x"75527851",
          7416 => x"c6be3f81",
          7417 => x"fef00852",
          7418 => x"7851ffb7",
          7419 => x"bb3f8255",
          7420 => x"81fef008",
          7421 => x"802e80dd",
          7422 => x"3881fef0",
          7423 => x"08527851",
          7424 => x"ffb5af3f",
          7425 => x"81fef008",
          7426 => x"7980d411",
          7427 => x"58585581",
          7428 => x"fef00880",
          7429 => x"c0388116",
          7430 => x"335473ae",
          7431 => x"2e098106",
          7432 => x"99386353",
          7433 => x"75527651",
          7434 => x"c6af3f78",
          7435 => x"54810b83",
          7436 => x"15348739",
          7437 => x"81fef008",
          7438 => x"9c387751",
          7439 => x"c8ca3f81",
          7440 => x"fef00855",
          7441 => x"81fef008",
          7442 => x"8c387851",
          7443 => x"ffb5aa3f",
          7444 => x"81fef008",
          7445 => x"557481fe",
          7446 => x"f00ca83d",
          7447 => x"0d04ed3d",
          7448 => x"0d0280db",
          7449 => x"05330284",
          7450 => x"0580df05",
          7451 => x"33575782",
          7452 => x"53953dd0",
          7453 => x"0552963d",
          7454 => x"51d2e93f",
          7455 => x"81fef008",
          7456 => x"5581fef0",
          7457 => x"0880cf38",
          7458 => x"785a6552",
          7459 => x"953dd405",
          7460 => x"51c9b53f",
          7461 => x"81fef008",
          7462 => x"5581fef0",
          7463 => x"08b83802",
          7464 => x"80cf0533",
          7465 => x"81a00654",
          7466 => x"865573aa",
          7467 => x"3875a706",
          7468 => x"6171098b",
          7469 => x"12337106",
          7470 => x"7a740607",
          7471 => x"51575556",
          7472 => x"748b1534",
          7473 => x"7854810b",
          7474 => x"83153478",
          7475 => x"51ffb4a9",
          7476 => x"3f81fef0",
          7477 => x"08557481",
          7478 => x"fef00c95",
          7479 => x"3d0d04ef",
          7480 => x"3d0d6456",
          7481 => x"8253933d",
          7482 => x"d0055294",
          7483 => x"3d51d1f4",
          7484 => x"3f81fef0",
          7485 => x"085581fe",
          7486 => x"f00880cb",
          7487 => x"38765863",
          7488 => x"52933dd4",
          7489 => x"0551c8c0",
          7490 => x"3f81fef0",
          7491 => x"085581fe",
          7492 => x"f008b438",
          7493 => x"0280c705",
          7494 => x"3381a006",
          7495 => x"54865573",
          7496 => x"a6388416",
          7497 => x"22861722",
          7498 => x"71902b07",
          7499 => x"5354961f",
          7500 => x"51ffb0c2",
          7501 => x"3f765481",
          7502 => x"0b831534",
          7503 => x"7651ffb3",
          7504 => x"b83f81fe",
          7505 => x"f0085574",
          7506 => x"81fef00c",
          7507 => x"933d0d04",
          7508 => x"ea3d0d69",
          7509 => x"6b5c5a80",
          7510 => x"53983dd0",
          7511 => x"0552993d",
          7512 => x"51d1813f",
          7513 => x"81fef008",
          7514 => x"81fef008",
          7515 => x"307081fe",
          7516 => x"f0080780",
          7517 => x"25515557",
          7518 => x"79802e81",
          7519 => x"85388170",
          7520 => x"75065555",
          7521 => x"73802e80",
          7522 => x"f9387b5d",
          7523 => x"805f8052",
          7524 => x"8d3d7052",
          7525 => x"54ffbea9",
          7526 => x"3f81fef0",
          7527 => x"085781fe",
          7528 => x"f00880d1",
          7529 => x"38745273",
          7530 => x"51c3dc3f",
          7531 => x"81fef008",
          7532 => x"5781fef0",
          7533 => x"08bf3881",
          7534 => x"fef00881",
          7535 => x"fef00865",
          7536 => x"5b595678",
          7537 => x"1881197b",
          7538 => x"18565955",
          7539 => x"74337434",
          7540 => x"8116568a",
          7541 => x"7827ec38",
          7542 => x"8b56751a",
          7543 => x"54807434",
          7544 => x"75802e9e",
          7545 => x"38ff1670",
          7546 => x"1b703351",
          7547 => x"555673a0",
          7548 => x"2ee8388e",
          7549 => x"3976842e",
          7550 => x"09810686",
          7551 => x"38807a34",
          7552 => x"80577630",
          7553 => x"70780780",
          7554 => x"2551547a",
          7555 => x"802e80c1",
          7556 => x"3873802e",
          7557 => x"bc387ba0",
          7558 => x"11085351",
          7559 => x"ffb1933f",
          7560 => x"81fef008",
          7561 => x"5781fef0",
          7562 => x"08a7387b",
          7563 => x"70335555",
          7564 => x"80c35673",
          7565 => x"832e8b38",
          7566 => x"80e45673",
          7567 => x"842e8338",
          7568 => x"a7567515",
          7569 => x"b40551ff",
          7570 => x"ade33f81",
          7571 => x"fef0087b",
          7572 => x"0c7681fe",
          7573 => x"f00c983d",
          7574 => x"0d04e63d",
          7575 => x"0d82539c",
          7576 => x"3dffb805",
          7577 => x"529d3d51",
          7578 => x"cefa3f81",
          7579 => x"fef00881",
          7580 => x"fef00856",
          7581 => x"5481fef0",
          7582 => x"08839838",
          7583 => x"8b53a052",
          7584 => x"8b3d7052",
          7585 => x"59ffaec0",
          7586 => x"3f736d70",
          7587 => x"337081ff",
          7588 => x"06525755",
          7589 => x"579f7427",
          7590 => x"81bc3878",
          7591 => x"587481ff",
          7592 => x"066d8105",
          7593 => x"4e705255",
          7594 => x"ffaf893f",
          7595 => x"81fef008",
          7596 => x"802ea538",
          7597 => x"6c703370",
          7598 => x"535754ff",
          7599 => x"aefd3f81",
          7600 => x"fef00880",
          7601 => x"2e8d3874",
          7602 => x"882b7607",
          7603 => x"6d81054e",
          7604 => x"55863981",
          7605 => x"fef00855",
          7606 => x"ff9f1570",
          7607 => x"83ffff06",
          7608 => x"51547399",
          7609 => x"268a38e0",
          7610 => x"157083ff",
          7611 => x"ff065654",
          7612 => x"80ff7527",
          7613 => x"873881ea",
          7614 => x"dc153355",
          7615 => x"74802ea3",
          7616 => x"38745281",
          7617 => x"ecdc51ff",
          7618 => x"ae893f81",
          7619 => x"fef00893",
          7620 => x"3881ff75",
          7621 => x"27883876",
          7622 => x"89268838",
          7623 => x"8b398a77",
          7624 => x"27863886",
          7625 => x"5581ec39",
          7626 => x"81ff7527",
          7627 => x"8f387488",
          7628 => x"2a547378",
          7629 => x"7081055a",
          7630 => x"34811757",
          7631 => x"74787081",
          7632 => x"055a3481",
          7633 => x"176d7033",
          7634 => x"7081ff06",
          7635 => x"52575557",
          7636 => x"739f26fe",
          7637 => x"c8388b3d",
          7638 => x"33548655",
          7639 => x"7381e52e",
          7640 => x"81b13876",
          7641 => x"802e9938",
          7642 => x"02a70555",
          7643 => x"76157033",
          7644 => x"515473a0",
          7645 => x"2e098106",
          7646 => x"8738ff17",
          7647 => x"5776ed38",
          7648 => x"79418043",
          7649 => x"8052913d",
          7650 => x"705255ff",
          7651 => x"bab33f81",
          7652 => x"fef00854",
          7653 => x"81fef008",
          7654 => x"80f73881",
          7655 => x"527451ff",
          7656 => x"bfe53f81",
          7657 => x"fef00854",
          7658 => x"81fef008",
          7659 => x"8d387680",
          7660 => x"c4386754",
          7661 => x"e5743480",
          7662 => x"c63981fe",
          7663 => x"f008842e",
          7664 => x"09810680",
          7665 => x"cc388054",
          7666 => x"76742e80",
          7667 => x"c4388152",
          7668 => x"7451ffbd",
          7669 => x"b03f81fe",
          7670 => x"f0085481",
          7671 => x"fef008b1",
          7672 => x"38a05381",
          7673 => x"fef00852",
          7674 => x"6751ffab",
          7675 => x"db3f6754",
          7676 => x"880b8b15",
          7677 => x"348b5378",
          7678 => x"526751ff",
          7679 => x"aba73f79",
          7680 => x"54810b83",
          7681 => x"15347951",
          7682 => x"ffadee3f",
          7683 => x"81fef008",
          7684 => x"54735574",
          7685 => x"81fef00c",
          7686 => x"9c3d0d04",
          7687 => x"f23d0d60",
          7688 => x"62028805",
          7689 => x"80cb0533",
          7690 => x"933dfc05",
          7691 => x"55725440",
          7692 => x"5e5ad2da",
          7693 => x"3f81fef0",
          7694 => x"085881fe",
          7695 => x"f00882bd",
          7696 => x"38911a33",
          7697 => x"587782b5",
          7698 => x"387c802e",
          7699 => x"97388c1a",
          7700 => x"08597890",
          7701 => x"38901a33",
          7702 => x"70812a70",
          7703 => x"81065155",
          7704 => x"55739038",
          7705 => x"87548297",
          7706 => x"39825882",
          7707 => x"90398158",
          7708 => x"828b397e",
          7709 => x"8a112270",
          7710 => x"892b7055",
          7711 => x"7f545656",
          7712 => x"56fee2a7",
          7713 => x"3fff147d",
          7714 => x"06703070",
          7715 => x"72079f2a",
          7716 => x"81fef008",
          7717 => x"058c1908",
          7718 => x"7c405a5d",
          7719 => x"55558177",
          7720 => x"27883898",
          7721 => x"16087726",
          7722 => x"83388257",
          7723 => x"76775659",
          7724 => x"80567452",
          7725 => x"7951ffae",
          7726 => x"993f8115",
          7727 => x"7f555598",
          7728 => x"14087526",
          7729 => x"83388255",
          7730 => x"81fef008",
          7731 => x"812eff99",
          7732 => x"3881fef0",
          7733 => x"08ff2eff",
          7734 => x"953881fe",
          7735 => x"f0088e38",
          7736 => x"81165675",
          7737 => x"7b2e0981",
          7738 => x"06873893",
          7739 => x"39745980",
          7740 => x"5674772e",
          7741 => x"098106ff",
          7742 => x"b9388758",
          7743 => x"80ff397d",
          7744 => x"802eba38",
          7745 => x"787b5555",
          7746 => x"7a802eb4",
          7747 => x"38811556",
          7748 => x"73812e09",
          7749 => x"81068338",
          7750 => x"ff567553",
          7751 => x"74527e51",
          7752 => x"ffafa83f",
          7753 => x"81fef008",
          7754 => x"5881fef0",
          7755 => x"0880ce38",
          7756 => x"748116ff",
          7757 => x"1656565c",
          7758 => x"73d33884",
          7759 => x"39ff195c",
          7760 => x"7e7c8c12",
          7761 => x"0c557d80",
          7762 => x"2eb33878",
          7763 => x"881b0c7c",
          7764 => x"8c1b0c90",
          7765 => x"1a3380c0",
          7766 => x"07547390",
          7767 => x"1b349815",
          7768 => x"08fe0590",
          7769 => x"16085754",
          7770 => x"75742691",
          7771 => x"38757b31",
          7772 => x"90160c84",
          7773 => x"15338107",
          7774 => x"54738416",
          7775 => x"34775473",
          7776 => x"81fef00c",
          7777 => x"903d0d04",
          7778 => x"e93d0d6b",
          7779 => x"6d028805",
          7780 => x"80eb0533",
          7781 => x"9d3d545a",
          7782 => x"5c59c5bd",
          7783 => x"3f8b5680",
          7784 => x"0b81fef0",
          7785 => x"08248bf8",
          7786 => x"3881fef0",
          7787 => x"08842981",
          7788 => x"ffa00570",
          7789 => x"08515574",
          7790 => x"802e8438",
          7791 => x"80753481",
          7792 => x"fef00881",
          7793 => x"ff065f81",
          7794 => x"527e51ff",
          7795 => x"a0d03f81",
          7796 => x"fef00881",
          7797 => x"ff067081",
          7798 => x"06565783",
          7799 => x"56748bc0",
          7800 => x"3876822a",
          7801 => x"70810651",
          7802 => x"558a5674",
          7803 => x"8bb23899",
          7804 => x"3dfc0553",
          7805 => x"83527e51",
          7806 => x"ffa4f03f",
          7807 => x"81fef008",
          7808 => x"99386755",
          7809 => x"74802e92",
          7810 => x"38748280",
          7811 => x"80268b38",
          7812 => x"ff157506",
          7813 => x"5574802e",
          7814 => x"83388148",
          7815 => x"78802e87",
          7816 => x"38848079",
          7817 => x"26923878",
          7818 => x"81800a26",
          7819 => x"8b38ff19",
          7820 => x"79065574",
          7821 => x"802e8638",
          7822 => x"93568ae4",
          7823 => x"3978892a",
          7824 => x"6e892a70",
          7825 => x"892b7759",
          7826 => x"4843597a",
          7827 => x"83388156",
          7828 => x"61307080",
          7829 => x"25770751",
          7830 => x"55915674",
          7831 => x"8ac23899",
          7832 => x"3df80553",
          7833 => x"81527e51",
          7834 => x"ffa4803f",
          7835 => x"815681fe",
          7836 => x"f0088aac",
          7837 => x"3877832a",
          7838 => x"70770681",
          7839 => x"fef00843",
          7840 => x"56457483",
          7841 => x"38bf4166",
          7842 => x"558e5660",
          7843 => x"75268a90",
          7844 => x"38746131",
          7845 => x"70485580",
          7846 => x"ff75278a",
          7847 => x"83389356",
          7848 => x"78818026",
          7849 => x"89fa3877",
          7850 => x"812a7081",
          7851 => x"06564374",
          7852 => x"802e9538",
          7853 => x"77870655",
          7854 => x"74822e83",
          7855 => x"8d387781",
          7856 => x"06557480",
          7857 => x"2e838338",
          7858 => x"77810655",
          7859 => x"9356825e",
          7860 => x"74802e89",
          7861 => x"cb38785a",
          7862 => x"7d832e09",
          7863 => x"810680e1",
          7864 => x"3878ae38",
          7865 => x"66912a57",
          7866 => x"810b81ed",
          7867 => x"8022565a",
          7868 => x"74802e9d",
          7869 => x"38747726",
          7870 => x"983881ed",
          7871 => x"80567910",
          7872 => x"82177022",
          7873 => x"57575a74",
          7874 => x"802e8638",
          7875 => x"767527ee",
          7876 => x"38795266",
          7877 => x"51fedd93",
          7878 => x"3f81fef0",
          7879 => x"08842984",
          7880 => x"87057089",
          7881 => x"2a5e55a0",
          7882 => x"5c800b81",
          7883 => x"fef008fc",
          7884 => x"808a0556",
          7885 => x"44fdfff0",
          7886 => x"0a752780",
          7887 => x"ec3888d3",
          7888 => x"3978ae38",
          7889 => x"668c2a57",
          7890 => x"810b81ec",
          7891 => x"f022565a",
          7892 => x"74802e9d",
          7893 => x"38747726",
          7894 => x"983881ec",
          7895 => x"f0567910",
          7896 => x"82177022",
          7897 => x"57575a74",
          7898 => x"802e8638",
          7899 => x"767527ee",
          7900 => x"38795266",
          7901 => x"51fedcb3",
          7902 => x"3f81fef0",
          7903 => x"08108405",
          7904 => x"5781fef0",
          7905 => x"089ff526",
          7906 => x"9638810b",
          7907 => x"81fef008",
          7908 => x"1081fef0",
          7909 => x"08057111",
          7910 => x"722a8305",
          7911 => x"59565e83",
          7912 => x"ff17892a",
          7913 => x"5d815ca0",
          7914 => x"44601c7d",
          7915 => x"11650569",
          7916 => x"7012ff05",
          7917 => x"71307072",
          7918 => x"0674315c",
          7919 => x"52595759",
          7920 => x"407d832e",
          7921 => x"09810689",
          7922 => x"38761c60",
          7923 => x"18415c84",
          7924 => x"39761d5d",
          7925 => x"79902918",
          7926 => x"70623168",
          7927 => x"58515574",
          7928 => x"762687af",
          7929 => x"38757c31",
          7930 => x"7d317a53",
          7931 => x"70653152",
          7932 => x"55fedbb7",
          7933 => x"3f81fef0",
          7934 => x"08587d83",
          7935 => x"2e098106",
          7936 => x"9b3881fe",
          7937 => x"f00883ff",
          7938 => x"f52680dd",
          7939 => x"38788783",
          7940 => x"3879812a",
          7941 => x"5978fdbe",
          7942 => x"3886f839",
          7943 => x"7d822e09",
          7944 => x"810680c5",
          7945 => x"3883fff5",
          7946 => x"0b81fef0",
          7947 => x"0827a038",
          7948 => x"788f3879",
          7949 => x"1a557480",
          7950 => x"c0268638",
          7951 => x"7459fd96",
          7952 => x"39628106",
          7953 => x"5574802e",
          7954 => x"8f38835e",
          7955 => x"fd883981",
          7956 => x"fef0089f",
          7957 => x"f5269238",
          7958 => x"7886b838",
          7959 => x"791a5981",
          7960 => x"807927fc",
          7961 => x"f13886ab",
          7962 => x"3980557d",
          7963 => x"812e0981",
          7964 => x"0683387d",
          7965 => x"559ff578",
          7966 => x"278b3874",
          7967 => x"8106558e",
          7968 => x"5674869c",
          7969 => x"38848053",
          7970 => x"80527a51",
          7971 => x"ffa2b93f",
          7972 => x"8b5381eb",
          7973 => x"98527a51",
          7974 => x"ffa28a3f",
          7975 => x"8480528b",
          7976 => x"1b51ffa1",
          7977 => x"b33f798d",
          7978 => x"1c347b83",
          7979 => x"ffff0652",
          7980 => x"8e1b51ff",
          7981 => x"a1a23f81",
          7982 => x"0b901c34",
          7983 => x"7d833270",
          7984 => x"3070962a",
          7985 => x"84800654",
          7986 => x"5155911b",
          7987 => x"51ffa188",
          7988 => x"3f665574",
          7989 => x"83ffff26",
          7990 => x"90387483",
          7991 => x"ffff0652",
          7992 => x"931b51ff",
          7993 => x"a0f23f8a",
          7994 => x"397452a0",
          7995 => x"1b51ffa1",
          7996 => x"853ff80b",
          7997 => x"951c34bf",
          7998 => x"52981b51",
          7999 => x"ffa0d93f",
          8000 => x"81ff529a",
          8001 => x"1b51ffa0",
          8002 => x"cf3f6052",
          8003 => x"9c1b51ff",
          8004 => x"a0e43f7d",
          8005 => x"832e0981",
          8006 => x"0680cb38",
          8007 => x"8288b20a",
          8008 => x"5280c31b",
          8009 => x"51ffa0ce",
          8010 => x"3f7c52a4",
          8011 => x"1b51ffa0",
          8012 => x"c53f8252",
          8013 => x"ac1b51ff",
          8014 => x"a0bc3f81",
          8015 => x"52b01b51",
          8016 => x"ffa0953f",
          8017 => x"8652b21b",
          8018 => x"51ffa08c",
          8019 => x"3fff800b",
          8020 => x"80c01c34",
          8021 => x"a90b80c2",
          8022 => x"1c349353",
          8023 => x"81eba452",
          8024 => x"80c71b51",
          8025 => x"ae398288",
          8026 => x"b20a52a7",
          8027 => x"1b51ffa0",
          8028 => x"853f7c83",
          8029 => x"ffff0652",
          8030 => x"961b51ff",
          8031 => x"9fda3fff",
          8032 => x"800ba41c",
          8033 => x"34a90ba6",
          8034 => x"1c349353",
          8035 => x"81ebb852",
          8036 => x"ab1b51ff",
          8037 => x"a08f3f82",
          8038 => x"d4d55283",
          8039 => x"fe1b7052",
          8040 => x"59ff9fb4",
          8041 => x"3f815460",
          8042 => x"537a527e",
          8043 => x"51ff9bd7",
          8044 => x"3f815681",
          8045 => x"fef00883",
          8046 => x"e7387d83",
          8047 => x"2e098106",
          8048 => x"80ee3875",
          8049 => x"54608605",
          8050 => x"537a527e",
          8051 => x"51ff9bb7",
          8052 => x"3f848053",
          8053 => x"80527a51",
          8054 => x"ff9fed3f",
          8055 => x"848b85a4",
          8056 => x"d2527a51",
          8057 => x"ff9f8f3f",
          8058 => x"868a85e4",
          8059 => x"f25283e4",
          8060 => x"1b51ff9f",
          8061 => x"813fff18",
          8062 => x"5283e81b",
          8063 => x"51ff9ef6",
          8064 => x"3f825283",
          8065 => x"ec1b51ff",
          8066 => x"9eec3f82",
          8067 => x"d4d55278",
          8068 => x"51ff9ec4",
          8069 => x"3f755460",
          8070 => x"8705537a",
          8071 => x"527e51ff",
          8072 => x"9ae53f75",
          8073 => x"54601653",
          8074 => x"7a527e51",
          8075 => x"ff9ad83f",
          8076 => x"65538052",
          8077 => x"7a51ff9f",
          8078 => x"8f3f7f56",
          8079 => x"80587d83",
          8080 => x"2e098106",
          8081 => x"9a38f852",
          8082 => x"7a51ff9e",
          8083 => x"a93fff52",
          8084 => x"841b51ff",
          8085 => x"9ea03ff0",
          8086 => x"0a52881b",
          8087 => x"51913987",
          8088 => x"fffff855",
          8089 => x"7d812e83",
          8090 => x"38f85574",
          8091 => x"527a51ff",
          8092 => x"9e843f7c",
          8093 => x"55615774",
          8094 => x"62268338",
          8095 => x"74577654",
          8096 => x"75537a52",
          8097 => x"7e51ff99",
          8098 => x"fe3f81fe",
          8099 => x"f0088287",
          8100 => x"38848053",
          8101 => x"81fef008",
          8102 => x"527a51ff",
          8103 => x"9eaa3f76",
          8104 => x"16757831",
          8105 => x"565674cd",
          8106 => x"38811858",
          8107 => x"77802eff",
          8108 => x"8d387955",
          8109 => x"7d832e83",
          8110 => x"38635561",
          8111 => x"57746226",
          8112 => x"83387457",
          8113 => x"76547553",
          8114 => x"7a527e51",
          8115 => x"ff99b83f",
          8116 => x"81fef008",
          8117 => x"81c13876",
          8118 => x"16757831",
          8119 => x"565674db",
          8120 => x"388c567d",
          8121 => x"832e9338",
          8122 => x"86566683",
          8123 => x"ffff268a",
          8124 => x"3884567d",
          8125 => x"822e8338",
          8126 => x"81566481",
          8127 => x"06587780",
          8128 => x"fe388480",
          8129 => x"5377527a",
          8130 => x"51ff9dbc",
          8131 => x"3f82d4d5",
          8132 => x"527851ff",
          8133 => x"9cc23f83",
          8134 => x"be1b5577",
          8135 => x"7534810b",
          8136 => x"81163481",
          8137 => x"0b821634",
          8138 => x"77831634",
          8139 => x"75841634",
          8140 => x"60670556",
          8141 => x"80fdc152",
          8142 => x"7551fed4",
          8143 => x"ee3ffe0b",
          8144 => x"85163481",
          8145 => x"fef00882",
          8146 => x"2abf0756",
          8147 => x"75861634",
          8148 => x"81fef008",
          8149 => x"87163460",
          8150 => x"5283c61b",
          8151 => x"51ff9c96",
          8152 => x"3f665283",
          8153 => x"ca1b51ff",
          8154 => x"9c8c3f81",
          8155 => x"5477537a",
          8156 => x"527e51ff",
          8157 => x"98913f81",
          8158 => x"5681fef0",
          8159 => x"08a23880",
          8160 => x"5380527e",
          8161 => x"51ff99e3",
          8162 => x"3f815681",
          8163 => x"fef00890",
          8164 => x"3889398e",
          8165 => x"568a3981",
          8166 => x"56863981",
          8167 => x"fef00856",
          8168 => x"7581fef0",
          8169 => x"0c993d0d",
          8170 => x"04f53d0d",
          8171 => x"7d605b59",
          8172 => x"807960ff",
          8173 => x"055a5757",
          8174 => x"767825b4",
          8175 => x"388d3df8",
          8176 => x"11555581",
          8177 => x"53fc1552",
          8178 => x"7951c9dc",
          8179 => x"3f7a812e",
          8180 => x"0981069c",
          8181 => x"388c3d33",
          8182 => x"55748d2e",
          8183 => x"db387476",
          8184 => x"70810558",
          8185 => x"34811757",
          8186 => x"748a2e09",
          8187 => x"8106c938",
          8188 => x"80763478",
          8189 => x"55768338",
          8190 => x"76557481",
          8191 => x"fef00c8d",
          8192 => x"3d0d04f7",
          8193 => x"3d0d7b02",
          8194 => x"8405b305",
          8195 => x"33595777",
          8196 => x"8a2e0981",
          8197 => x"0687388d",
          8198 => x"527651e7",
          8199 => x"3f841708",
          8200 => x"56807624",
          8201 => x"be388817",
          8202 => x"0877178c",
          8203 => x"05565977",
          8204 => x"75348116",
          8205 => x"56bb7625",
          8206 => x"a1388b3d",
          8207 => x"fc055475",
          8208 => x"538c1752",
          8209 => x"760851cb",
          8210 => x"dc3f7976",
          8211 => x"32703070",
          8212 => x"72079f2a",
          8213 => x"70305351",
          8214 => x"56567584",
          8215 => x"180c8119",
          8216 => x"88180c8b",
          8217 => x"3d0d04f9",
          8218 => x"3d0d7984",
          8219 => x"11085656",
          8220 => x"807524a7",
          8221 => x"38893dfc",
          8222 => x"05547453",
          8223 => x"8c165275",
          8224 => x"0851cba1",
          8225 => x"3f81fef0",
          8226 => x"08913884",
          8227 => x"1608782e",
          8228 => x"09810687",
          8229 => x"38881608",
          8230 => x"558339ff",
          8231 => x"557481fe",
          8232 => x"f00c893d",
          8233 => x"0d04fd3d",
          8234 => x"0d755480",
          8235 => x"cc538052",
          8236 => x"7351ff9a",
          8237 => x"933f7674",
          8238 => x"0c853d0d",
          8239 => x"04ea3d0d",
          8240 => x"0280e305",
          8241 => x"336a5386",
          8242 => x"3d705354",
          8243 => x"54d83f73",
          8244 => x"527251fe",
          8245 => x"ae3f7251",
          8246 => x"ff8d3f98",
          8247 => x"3d0d04f8",
          8248 => x"3d0d7a70",
          8249 => x"08705656",
          8250 => x"5974802e",
          8251 => x"80e1388c",
          8252 => x"39771579",
          8253 => x"0c851633",
          8254 => x"5480d439",
          8255 => x"74335473",
          8256 => x"a02e0981",
          8257 => x"06863881",
          8258 => x"1555f139",
          8259 => x"80577690",
          8260 => x"2981fbe0",
          8261 => x"05700852",
          8262 => x"56fedab1",
          8263 => x"3f81fef0",
          8264 => x"0881fef0",
          8265 => x"08547553",
          8266 => x"76085258",
          8267 => x"fedaff3f",
          8268 => x"81fef008",
          8269 => x"8b388416",
          8270 => x"33547381",
          8271 => x"2effb238",
          8272 => x"81177081",
          8273 => x"ff065854",
          8274 => x"987727c2",
          8275 => x"38ff5473",
          8276 => x"81fef00c",
          8277 => x"8a3d0d04",
          8278 => x"ff3d0d73",
          8279 => x"52719326",
          8280 => x"818e3871",
          8281 => x"842981e2",
          8282 => x"84055271",
          8283 => x"080481ee",
          8284 => x"b8518180",
          8285 => x"3981eec4",
          8286 => x"5180f939",
          8287 => x"81eed851",
          8288 => x"80f23981",
          8289 => x"eeec5180",
          8290 => x"eb3981ee",
          8291 => x"fc5180e4",
          8292 => x"3981ef8c",
          8293 => x"5180dd39",
          8294 => x"81efa051",
          8295 => x"80d63981",
          8296 => x"efb05180",
          8297 => x"cf3981ef",
          8298 => x"c85180c8",
          8299 => x"3981efe0",
          8300 => x"5180c139",
          8301 => x"81eff851",
          8302 => x"bb3981f0",
          8303 => x"9451b539",
          8304 => x"81f0a851",
          8305 => x"af3981f0",
          8306 => x"d451a939",
          8307 => x"81f0e851",
          8308 => x"a33981f1",
          8309 => x"88519d39",
          8310 => x"81f19c51",
          8311 => x"973981f1",
          8312 => x"b4519139",
          8313 => x"81f1cc51",
          8314 => x"8b3981f1",
          8315 => x"e4518539",
          8316 => x"81f1f051",
          8317 => x"fef2ae3f",
          8318 => x"833d0d04",
          8319 => x"fb3d0d77",
          8320 => x"79565674",
          8321 => x"87e7268a",
          8322 => x"38745275",
          8323 => x"87e82951",
          8324 => x"913987e8",
          8325 => x"527451fe",
          8326 => x"cf913f81",
          8327 => x"fef00852",
          8328 => x"7551fecf",
          8329 => x"863f81fe",
          8330 => x"f0085479",
          8331 => x"53755281",
          8332 => x"f28051fe",
          8333 => x"f7d33f87",
          8334 => x"3d0d04ec",
          8335 => x"3d0d6602",
          8336 => x"840580e3",
          8337 => x"05335b57",
          8338 => x"80687830",
          8339 => x"707a0773",
          8340 => x"25515759",
          8341 => x"59785677",
          8342 => x"87ff2683",
          8343 => x"38815674",
          8344 => x"76077081",
          8345 => x"ff065155",
          8346 => x"93567481",
          8347 => x"80388153",
          8348 => x"76528c3d",
          8349 => x"705256ff",
          8350 => x"bfc93f81",
          8351 => x"fef00857",
          8352 => x"81fef008",
          8353 => x"b83881fe",
          8354 => x"f00887c0",
          8355 => x"98880c81",
          8356 => x"fef00859",
          8357 => x"963dd405",
          8358 => x"54848053",
          8359 => x"77527551",
          8360 => x"c4863f81",
          8361 => x"fef00857",
          8362 => x"81fef008",
          8363 => x"90387a55",
          8364 => x"74802e89",
          8365 => x"38741975",
          8366 => x"195959d8",
          8367 => x"39963dd8",
          8368 => x"0551cbf0",
          8369 => x"3f763070",
          8370 => x"78078025",
          8371 => x"7b30709f",
          8372 => x"2a720651",
          8373 => x"57515674",
          8374 => x"802e9038",
          8375 => x"81f2a453",
          8376 => x"87c09888",
          8377 => x"08527851",
          8378 => x"fe923f76",
          8379 => x"567581fe",
          8380 => x"f00c963d",
          8381 => x"0d04f93d",
          8382 => x"0d7b0284",
          8383 => x"05b30533",
          8384 => x"5758ff57",
          8385 => x"80537a52",
          8386 => x"7951feaf",
          8387 => x"3f81fef0",
          8388 => x"08a43875",
          8389 => x"802e8838",
          8390 => x"75812e98",
          8391 => x"38983960",
          8392 => x"557f5481",
          8393 => x"fef0537e",
          8394 => x"527d5177",
          8395 => x"2d81fef0",
          8396 => x"08578339",
          8397 => x"77047681",
          8398 => x"fef00c89",
          8399 => x"3d0d04f3",
          8400 => x"3d0d7f61",
          8401 => x"63028c05",
          8402 => x"80cf0533",
          8403 => x"73731568",
          8404 => x"415f5c5c",
          8405 => x"5e5e5e7a",
          8406 => x"5281f2ac",
          8407 => x"51fef5a9",
          8408 => x"3f81f2b4",
          8409 => x"51feefbd",
          8410 => x"3f805574",
          8411 => x"792780fc",
          8412 => x"387b902e",
          8413 => x"89387ba0",
          8414 => x"2ea73880",
          8415 => x"c6397418",
          8416 => x"53727a27",
          8417 => x"8e387222",
          8418 => x"5281f2b8",
          8419 => x"51fef4f9",
          8420 => x"3f893981",
          8421 => x"f2c451fe",
          8422 => x"ef8b3f82",
          8423 => x"155580c3",
          8424 => x"39741853",
          8425 => x"727a278e",
          8426 => x"38720852",
          8427 => x"81f2ac51",
          8428 => x"fef4d63f",
          8429 => x"893981f2",
          8430 => x"c051feee",
          8431 => x"e83f8415",
          8432 => x"55a13974",
          8433 => x"1853727a",
          8434 => x"278e3872",
          8435 => x"335281f2",
          8436 => x"cc51fef4",
          8437 => x"b43f8939",
          8438 => x"81f2d451",
          8439 => x"feeec63f",
          8440 => x"811555a0",
          8441 => x"51feede0",
          8442 => x"3fff8039",
          8443 => x"81f2d851",
          8444 => x"feeeb23f",
          8445 => x"80557479",
          8446 => x"27bc3874",
          8447 => x"18703355",
          8448 => x"53805672",
          8449 => x"7a278338",
          8450 => x"81568053",
          8451 => x"9f742783",
          8452 => x"38815375",
          8453 => x"73067081",
          8454 => x"ff065153",
          8455 => x"72802e8b",
          8456 => x"387380fe",
          8457 => x"26853873",
          8458 => x"518339a0",
          8459 => x"51feed98",
          8460 => x"3f811555",
          8461 => x"c13981f2",
          8462 => x"dc51feed",
          8463 => x"e83f7818",
          8464 => x"791c5c58",
          8465 => x"fede963f",
          8466 => x"81fef008",
          8467 => x"982b7098",
          8468 => x"2c515776",
          8469 => x"a02e0981",
          8470 => x"06ab38fe",
          8471 => x"ddff3f81",
          8472 => x"fef00898",
          8473 => x"2b70982c",
          8474 => x"70a03270",
          8475 => x"30729b32",
          8476 => x"70307072",
          8477 => x"07737507",
          8478 => x"06515858",
          8479 => x"59575157",
          8480 => x"807324d7",
          8481 => x"38769b2e",
          8482 => x"09810685",
          8483 => x"3880538c",
          8484 => x"397c1e53",
          8485 => x"727826fd",
          8486 => x"be38ff53",
          8487 => x"7281fef0",
          8488 => x"0c8f3d0d",
          8489 => x"04fc3d0d",
          8490 => x"029b0533",
          8491 => x"81f2e053",
          8492 => x"81f2e852",
          8493 => x"55fef2d1",
          8494 => x"3f81faa0",
          8495 => x"2251fee6",
          8496 => x"d73f81f2",
          8497 => x"f45481f3",
          8498 => x"805381fa",
          8499 => x"a1335281",
          8500 => x"f38851fe",
          8501 => x"f2b33f74",
          8502 => x"802e8538",
          8503 => x"fee2a23f",
          8504 => x"863d0d04",
          8505 => x"fe3d0d87",
          8506 => x"c0968008",
          8507 => x"53fee7b1",
          8508 => x"3f8151fe",
          8509 => x"d8fb3f81",
          8510 => x"f3a451fe",
          8511 => x"daf33f80",
          8512 => x"51fed8ed",
          8513 => x"3f72812a",
          8514 => x"70810651",
          8515 => x"5271802e",
          8516 => x"95388151",
          8517 => x"fed8da3f",
          8518 => x"81f3c051",
          8519 => x"fedad23f",
          8520 => x"8051fed8",
          8521 => x"cc3f7282",
          8522 => x"2a708106",
          8523 => x"51527180",
          8524 => x"2e953881",
          8525 => x"51fed8b9",
          8526 => x"3f81f3d4",
          8527 => x"51fedab1",
          8528 => x"3f8051fe",
          8529 => x"d8ab3f72",
          8530 => x"832a7081",
          8531 => x"06515271",
          8532 => x"802e9538",
          8533 => x"8151fed8",
          8534 => x"983f81f3",
          8535 => x"e451feda",
          8536 => x"903f8051",
          8537 => x"fed88a3f",
          8538 => x"72842a70",
          8539 => x"81065152",
          8540 => x"71802e95",
          8541 => x"388151fe",
          8542 => x"d7f73f81",
          8543 => x"f3f851fe",
          8544 => x"d9ef3f80",
          8545 => x"51fed7e9",
          8546 => x"3f72852a",
          8547 => x"70810651",
          8548 => x"5271802e",
          8549 => x"95388151",
          8550 => x"fed7d63f",
          8551 => x"81f48c51",
          8552 => x"fed9ce3f",
          8553 => x"8051fed7",
          8554 => x"c83f7286",
          8555 => x"2a708106",
          8556 => x"51527180",
          8557 => x"2e953881",
          8558 => x"51fed7b5",
          8559 => x"3f81f4a0",
          8560 => x"51fed9ad",
          8561 => x"3f8051fe",
          8562 => x"d7a73f72",
          8563 => x"872a7081",
          8564 => x"06515271",
          8565 => x"802e9538",
          8566 => x"8151fed7",
          8567 => x"943f81f4",
          8568 => x"b451fed9",
          8569 => x"8c3f8051",
          8570 => x"fed7863f",
          8571 => x"72882a70",
          8572 => x"81065152",
          8573 => x"71802e95",
          8574 => x"388151fe",
          8575 => x"d6f33f81",
          8576 => x"f4c851fe",
          8577 => x"d8eb3f80",
          8578 => x"51fed6e5",
          8579 => x"3ffee599",
          8580 => x"3f843d0d",
          8581 => x"04fb3d0d",
          8582 => x"77028405",
          8583 => x"a3053370",
          8584 => x"55565680",
          8585 => x"527551fe",
          8586 => x"cea33f81",
          8587 => x"fbdc3354",
          8588 => x"73a73881",
          8589 => x"5381f588",
          8590 => x"52829688",
          8591 => x"51ffb883",
          8592 => x"3f81fef0",
          8593 => x"08307081",
          8594 => x"fef00807",
          8595 => x"80258271",
          8596 => x"31515154",
          8597 => x"7381fbdc",
          8598 => x"3481fbdc",
          8599 => x"33547381",
          8600 => x"2e098106",
          8601 => x"ac388296",
          8602 => x"88537452",
          8603 => x"7551f2b9",
          8604 => x"3f81fef0",
          8605 => x"08802e8c",
          8606 => x"3881fef0",
          8607 => x"0851fee9",
          8608 => x"a43f8e39",
          8609 => x"82968851",
          8610 => x"c4aa3f82",
          8611 => x"0b81fbdc",
          8612 => x"3481fbdc",
          8613 => x"33547382",
          8614 => x"2e098106",
          8615 => x"89387452",
          8616 => x"7551fefa",
          8617 => x"e43f800b",
          8618 => x"81fef00c",
          8619 => x"873d0d04",
          8620 => x"ce3d0d80",
          8621 => x"70718296",
          8622 => x"840c5f5d",
          8623 => x"81527c51",
          8624 => x"ff86db3f",
          8625 => x"81fef008",
          8626 => x"81ff0659",
          8627 => x"787d2e09",
          8628 => x"8106a238",
          8629 => x"81f59852",
          8630 => x"963d7052",
          8631 => x"59feeebf",
          8632 => x"3f7c5378",
          8633 => x"528280b4",
          8634 => x"51ffb5f6",
          8635 => x"3f81fef0",
          8636 => x"087d2e88",
          8637 => x"3881f59c",
          8638 => x"5191fe39",
          8639 => x"81705f5d",
          8640 => x"81f5d451",
          8641 => x"fee89e3f",
          8642 => x"963d7046",
          8643 => x"5a80f852",
          8644 => x"7951fe81",
          8645 => x"3fb43dff",
          8646 => x"840551f3",
          8647 => x"c23f81fe",
          8648 => x"f008902b",
          8649 => x"70902c51",
          8650 => x"597880c1",
          8651 => x"2e89f138",
          8652 => x"7880c124",
          8653 => x"80d93878",
          8654 => x"ab2e83c0",
          8655 => x"3878ab24",
          8656 => x"a4387882",
          8657 => x"2e81b338",
          8658 => x"7882248a",
          8659 => x"3878802e",
          8660 => x"ffae388f",
          8661 => x"a5397884",
          8662 => x"2e828638",
          8663 => x"78942e82",
          8664 => x"b1388f96",
          8665 => x"3978bd2e",
          8666 => x"858c3878",
          8667 => x"bd249038",
          8668 => x"78b02e83",
          8669 => x"af3878bc",
          8670 => x"2e849138",
          8671 => x"8efc3978",
          8672 => x"bf2e85d7",
          8673 => x"387880c0",
          8674 => x"2e86d238",
          8675 => x"8eec3978",
          8676 => x"80d52e8d",
          8677 => x"c2387880",
          8678 => x"d524b038",
          8679 => x"7880d02e",
          8680 => x"8cf63878",
          8681 => x"80d02492",
          8682 => x"387880c2",
          8683 => x"2e8a9938",
          8684 => x"7880c32e",
          8685 => x"8bc2388e",
          8686 => x"c1397880",
          8687 => x"d12e8ce9",
          8688 => x"387880d4",
          8689 => x"2e8cf338",
          8690 => x"8eb03978",
          8691 => x"81822e8e",
          8692 => x"86387881",
          8693 => x"82249238",
          8694 => x"7880f82e",
          8695 => x"8d963878",
          8696 => x"80f92e8d",
          8697 => x"b4388e92",
          8698 => x"39788183",
          8699 => x"2e8df738",
          8700 => x"7881852e",
          8701 => x"8dfd388e",
          8702 => x"8139b43d",
          8703 => x"ff801153",
          8704 => x"ff840551",
          8705 => x"feedf73f",
          8706 => x"81fef008",
          8707 => x"883881f5",
          8708 => x"d8518fe5",
          8709 => x"39b43dfe",
          8710 => x"fc1153ff",
          8711 => x"840551fe",
          8712 => x"eddc3f81",
          8713 => x"fef00880",
          8714 => x"2e883881",
          8715 => x"63258338",
          8716 => x"80430280",
          8717 => x"cb053352",
          8718 => x"0280cf05",
          8719 => x"3351ff83",
          8720 => x"dd3f81fe",
          8721 => x"f00881ff",
          8722 => x"0659788e",
          8723 => x"3881f5e8",
          8724 => x"51fee5d1",
          8725 => x"3f815efd",
          8726 => x"a73981f5",
          8727 => x"f85187b9",
          8728 => x"39b43dff",
          8729 => x"801153ff",
          8730 => x"840551fe",
          8731 => x"ed903f81",
          8732 => x"fef00880",
          8733 => x"2efd8938",
          8734 => x"80538052",
          8735 => x"0280cf05",
          8736 => x"3351ff87",
          8737 => x"e63f81fe",
          8738 => x"f0085281",
          8739 => x"f690518c",
          8740 => x"bf39b43d",
          8741 => x"ff801153",
          8742 => x"ff840551",
          8743 => x"feecdf3f",
          8744 => x"81fef008",
          8745 => x"802e8738",
          8746 => x"638926fc",
          8747 => x"d338b43d",
          8748 => x"fefc1153",
          8749 => x"ff840551",
          8750 => x"feecc33f",
          8751 => x"81fef008",
          8752 => x"863881fe",
          8753 => x"f0084363",
          8754 => x"5381f698",
          8755 => x"527951fe",
          8756 => x"eacd3f02",
          8757 => x"80cb0533",
          8758 => x"53795263",
          8759 => x"84b42982",
          8760 => x"80b40551",
          8761 => x"ffb1fb3f",
          8762 => x"81fef008",
          8763 => x"81933881",
          8764 => x"f5e851fe",
          8765 => x"e4af3f81",
          8766 => x"5dfc8539",
          8767 => x"b43dff84",
          8768 => x"0551fecd",
          8769 => x"9d3f81fe",
          8770 => x"f008b53d",
          8771 => x"ff840552",
          8772 => x"5bfecdf0",
          8773 => x"3f815381",
          8774 => x"fef00852",
          8775 => x"7a51f29b",
          8776 => x"3f80d539",
          8777 => x"b43dff84",
          8778 => x"0551fecc",
          8779 => x"f53f81fe",
          8780 => x"f008b53d",
          8781 => x"ff840552",
          8782 => x"5bfecdc8",
          8783 => x"3f81fef0",
          8784 => x"08b53dff",
          8785 => x"8405525a",
          8786 => x"fecdb93f",
          8787 => x"81fef008",
          8788 => x"b53dff84",
          8789 => x"055259fe",
          8790 => x"cdaa3f81",
          8791 => x"f9ec5881",
          8792 => x"ffb85780",
          8793 => x"56805581",
          8794 => x"fef00881",
          8795 => x"ff065478",
          8796 => x"5379527a",
          8797 => x"51f2ff3f",
          8798 => x"81fef008",
          8799 => x"802efb80",
          8800 => x"3881fef0",
          8801 => x"0851efd0",
          8802 => x"3ffaf539",
          8803 => x"b43dff80",
          8804 => x"1153ff84",
          8805 => x"0551feea",
          8806 => x"e53f81fe",
          8807 => x"f008802e",
          8808 => x"fade38b4",
          8809 => x"3dfefc11",
          8810 => x"53ff8405",
          8811 => x"51feeace",
          8812 => x"3f81fef0",
          8813 => x"08802efa",
          8814 => x"c738b43d",
          8815 => x"fef81153",
          8816 => x"ff840551",
          8817 => x"feeab73f",
          8818 => x"81fef008",
          8819 => x"863881fe",
          8820 => x"f0084281",
          8821 => x"f69c51fe",
          8822 => x"e2cb3f63",
          8823 => x"635c5a79",
          8824 => x"7b2781f2",
          8825 => x"38615978",
          8826 => x"7a708405",
          8827 => x"5c0c7a7a",
          8828 => x"26f53881",
          8829 => x"e139b43d",
          8830 => x"ff801153",
          8831 => x"ff840551",
          8832 => x"fee9fb3f",
          8833 => x"81fef008",
          8834 => x"802ef9f4",
          8835 => x"38b43dfe",
          8836 => x"fc1153ff",
          8837 => x"840551fe",
          8838 => x"e9e43f81",
          8839 => x"fef00880",
          8840 => x"2ef9dd38",
          8841 => x"b43dfef8",
          8842 => x"1153ff84",
          8843 => x"0551fee9",
          8844 => x"cd3f81fe",
          8845 => x"f008802e",
          8846 => x"f9c63881",
          8847 => x"f6ac51fe",
          8848 => x"e1e33f63",
          8849 => x"5a796327",
          8850 => x"818c3861",
          8851 => x"59797081",
          8852 => x"055b3379",
          8853 => x"34618105",
          8854 => x"42eb39b4",
          8855 => x"3dff8011",
          8856 => x"53ff8405",
          8857 => x"51fee996",
          8858 => x"3f81fef0",
          8859 => x"08802ef9",
          8860 => x"8f38b43d",
          8861 => x"fefc1153",
          8862 => x"ff840551",
          8863 => x"fee8ff3f",
          8864 => x"81fef008",
          8865 => x"802ef8f8",
          8866 => x"38b43dfe",
          8867 => x"f81153ff",
          8868 => x"840551fe",
          8869 => x"e8e83f81",
          8870 => x"fef00880",
          8871 => x"2ef8e138",
          8872 => x"81f6b851",
          8873 => x"fee0fe3f",
          8874 => x"635a7963",
          8875 => x"27a83861",
          8876 => x"70337b33",
          8877 => x"5e5a5b78",
          8878 => x"7c2e9238",
          8879 => x"78557a54",
          8880 => x"79335379",
          8881 => x"5281f6c8",
          8882 => x"51fee6bd",
          8883 => x"3f811a62",
          8884 => x"8105435a",
          8885 => x"d53981f5",
          8886 => x"e45182bd",
          8887 => x"39b43dff",
          8888 => x"801153ff",
          8889 => x"840551fe",
          8890 => x"e8943f81",
          8891 => x"fef00880",
          8892 => x"df3881fa",
          8893 => x"b4335978",
          8894 => x"802e8938",
          8895 => x"81f9ec08",
          8896 => x"4480cd39",
          8897 => x"81fab533",
          8898 => x"5978802e",
          8899 => x"883881f9",
          8900 => x"f40844bc",
          8901 => x"3981fab6",
          8902 => x"33597880",
          8903 => x"2e883881",
          8904 => x"f9fc0844",
          8905 => x"ab3981fa",
          8906 => x"b7335978",
          8907 => x"802e8838",
          8908 => x"81fa8408",
          8909 => x"449a3981",
          8910 => x"fab23359",
          8911 => x"78802e88",
          8912 => x"3881fa8c",
          8913 => x"08448939",
          8914 => x"81fa9c08",
          8915 => x"fc800544",
          8916 => x"b43dfefc",
          8917 => x"1153ff84",
          8918 => x"0551fee7",
          8919 => x"a13f81fe",
          8920 => x"f00880de",
          8921 => x"3881fab4",
          8922 => x"33597880",
          8923 => x"2e893881",
          8924 => x"f9f00843",
          8925 => x"80cc3981",
          8926 => x"fab53359",
          8927 => x"78802e88",
          8928 => x"3881f9f8",
          8929 => x"0843bb39",
          8930 => x"81fab633",
          8931 => x"5978802e",
          8932 => x"883881fa",
          8933 => x"800843aa",
          8934 => x"3981fab7",
          8935 => x"33597880",
          8936 => x"2e883881",
          8937 => x"fa880843",
          8938 => x"993981fa",
          8939 => x"b2335978",
          8940 => x"802e8838",
          8941 => x"81fa9008",
          8942 => x"43883981",
          8943 => x"fa9c0888",
          8944 => x"0543b43d",
          8945 => x"fef81153",
          8946 => x"ff840551",
          8947 => x"fee6af3f",
          8948 => x"81fef008",
          8949 => x"802ea738",
          8950 => x"80625c5c",
          8951 => x"7a882e83",
          8952 => x"38815c7a",
          8953 => x"90327030",
          8954 => x"7072079f",
          8955 => x"2a707f06",
          8956 => x"51515a5a",
          8957 => x"78802e88",
          8958 => x"387aa02e",
          8959 => x"83388842",
          8960 => x"81f6e451",
          8961 => x"fede9e3f",
          8962 => x"a0556354",
          8963 => x"61536252",
          8964 => x"6351eeab",
          8965 => x"3f81f6f4",
          8966 => x"51fede89",
          8967 => x"3ff5e139",
          8968 => x"b43dff80",
          8969 => x"1153ff84",
          8970 => x"0551fee5",
          8971 => x"d13f81fe",
          8972 => x"f008802e",
          8973 => x"f5ca38b4",
          8974 => x"3dfefc11",
          8975 => x"53ff8405",
          8976 => x"51fee5ba",
          8977 => x"3f81fef0",
          8978 => x"08802ea5",
          8979 => x"38635902",
          8980 => x"80cb0533",
          8981 => x"79346381",
          8982 => x"0544b43d",
          8983 => x"fefc1153",
          8984 => x"ff840551",
          8985 => x"fee5973f",
          8986 => x"81fef008",
          8987 => x"e038f590",
          8988 => x"39637033",
          8989 => x"545281f7",
          8990 => x"8051fee3",
          8991 => x"8c3f80f8",
          8992 => x"527951fe",
          8993 => x"e3dd3f79",
          8994 => x"45793359",
          8995 => x"78ae2ef4",
          8996 => x"ef389f79",
          8997 => x"27a038b4",
          8998 => x"3dfefc11",
          8999 => x"53ff8405",
          9000 => x"51fee4da",
          9001 => x"3f81fef0",
          9002 => x"08802e91",
          9003 => x"38635902",
          9004 => x"80cb0533",
          9005 => x"79346381",
          9006 => x"0544ffb5",
          9007 => x"3981f78c",
          9008 => x"51fedce1",
          9009 => x"3fffaa39",
          9010 => x"b43dfef4",
          9011 => x"1153ff84",
          9012 => x"0551fee6",
          9013 => x"9b3f81fe",
          9014 => x"f008802e",
          9015 => x"f4a238b4",
          9016 => x"3dfef011",
          9017 => x"53ff8405",
          9018 => x"51fee684",
          9019 => x"3f81fef0",
          9020 => x"08802ea6",
          9021 => x"38605902",
          9022 => x"be052279",
          9023 => x"7082055b",
          9024 => x"237841b4",
          9025 => x"3dfef011",
          9026 => x"53ff8405",
          9027 => x"51fee5e0",
          9028 => x"3f81fef0",
          9029 => x"08df38f3",
          9030 => x"e7396070",
          9031 => x"22545281",
          9032 => x"f79451fe",
          9033 => x"e1e33f80",
          9034 => x"f8527951",
          9035 => x"fee2b43f",
          9036 => x"79457933",
          9037 => x"5978ae2e",
          9038 => x"f3c63878",
          9039 => x"9f268738",
          9040 => x"60820541",
          9041 => x"d539b43d",
          9042 => x"fef01153",
          9043 => x"ff840551",
          9044 => x"fee59d3f",
          9045 => x"81fef008",
          9046 => x"802e9238",
          9047 => x"605902be",
          9048 => x"05227970",
          9049 => x"82055b23",
          9050 => x"7841ffae",
          9051 => x"3981f78c",
          9052 => x"51fedbb1",
          9053 => x"3fffa339",
          9054 => x"b43dfef4",
          9055 => x"1153ff84",
          9056 => x"0551fee4",
          9057 => x"eb3f81fe",
          9058 => x"f008802e",
          9059 => x"f2f238b4",
          9060 => x"3dfef011",
          9061 => x"53ff8405",
          9062 => x"51fee4d4",
          9063 => x"3f81fef0",
          9064 => x"08802ea1",
          9065 => x"38606071",
          9066 => x"0c596084",
          9067 => x"0541b43d",
          9068 => x"fef01153",
          9069 => x"ff840551",
          9070 => x"fee4b53f",
          9071 => x"81fef008",
          9072 => x"e438f2bc",
          9073 => x"39607008",
          9074 => x"545281f7",
          9075 => x"a051fee0",
          9076 => x"b83f80f8",
          9077 => x"527951fe",
          9078 => x"e1893f79",
          9079 => x"45793359",
          9080 => x"78ae2ef2",
          9081 => x"9b389f79",
          9082 => x"279c38b4",
          9083 => x"3dfef011",
          9084 => x"53ff8405",
          9085 => x"51fee3f8",
          9086 => x"3f81fef0",
          9087 => x"08802e8d",
          9088 => x"38606071",
          9089 => x"0c596084",
          9090 => x"0541ffb9",
          9091 => x"3981f78c",
          9092 => x"51feda91",
          9093 => x"3fffae39",
          9094 => x"81f7ac51",
          9095 => x"feda863f",
          9096 => x"8251fed4",
          9097 => x"d73ff1d8",
          9098 => x"3981f7c4",
          9099 => x"51fed9f5",
          9100 => x"3fa251fe",
          9101 => x"d4aa3ff1",
          9102 => x"c73981f7",
          9103 => x"dc51fed9",
          9104 => x"e43f8480",
          9105 => x"810b87c0",
          9106 => x"94840c84",
          9107 => x"80810b87",
          9108 => x"c094940c",
          9109 => x"f1aa3981",
          9110 => x"f7f051fe",
          9111 => x"d9c73f8c",
          9112 => x"80830b87",
          9113 => x"c094840c",
          9114 => x"8c80830b",
          9115 => x"87c09494",
          9116 => x"0cf18d39",
          9117 => x"b43dff80",
          9118 => x"1153ff84",
          9119 => x"0551fee0",
          9120 => x"fd3f81fe",
          9121 => x"f008802e",
          9122 => x"f0f63863",
          9123 => x"5281f884",
          9124 => x"51fedef5",
          9125 => x"3f635978",
          9126 => x"04b43dff",
          9127 => x"801153ff",
          9128 => x"840551fe",
          9129 => x"e0d83f81",
          9130 => x"fef00880",
          9131 => x"2ef0d138",
          9132 => x"635281f8",
          9133 => x"a051fede",
          9134 => x"d03f6359",
          9135 => x"782d81fe",
          9136 => x"f008802e",
          9137 => x"f0ba3881",
          9138 => x"fef00852",
          9139 => x"81f8bc51",
          9140 => x"fedeb63f",
          9141 => x"f0aa3981",
          9142 => x"f8d851fe",
          9143 => x"d8c73ffe",
          9144 => x"b5aa3ff0",
          9145 => x"9b3981f8",
          9146 => x"f451fed8",
          9147 => x"b83f8059",
          9148 => x"ffa539fe",
          9149 => x"ce8b3ff0",
          9150 => x"87397945",
          9151 => x"79335978",
          9152 => x"802eeffc",
          9153 => x"387d7d06",
          9154 => x"5978802e",
          9155 => x"81d338b4",
          9156 => x"3dff8405",
          9157 => x"51fec18a",
          9158 => x"3f81fef0",
          9159 => x"085b815c",
          9160 => x"7b822eb2",
          9161 => x"387b8224",
          9162 => x"89387b81",
          9163 => x"2e8c3880",
          9164 => x"cd397b83",
          9165 => x"2eb03880",
          9166 => x"c53981f9",
          9167 => x"88567a55",
          9168 => x"81f98c54",
          9169 => x"805381f9",
          9170 => x"9052b43d",
          9171 => x"ffb00551",
          9172 => x"feddcc3f",
          9173 => x"bb3981f9",
          9174 => x"b052b43d",
          9175 => x"ffb00551",
          9176 => x"feddbc3f",
          9177 => x"ab397a55",
          9178 => x"81f98c54",
          9179 => x"805381f9",
          9180 => x"a052b43d",
          9181 => x"ffb00551",
          9182 => x"fedda43f",
          9183 => x"93397a54",
          9184 => x"805381f9",
          9185 => x"ac52b43d",
          9186 => x"ffb00551",
          9187 => x"fedd903f",
          9188 => x"81f9ec58",
          9189 => x"81ffb857",
          9190 => x"80566455",
          9191 => x"80548380",
          9192 => x"80538380",
          9193 => x"8052b43d",
          9194 => x"ffb00551",
          9195 => x"e6c83f81",
          9196 => x"fef00881",
          9197 => x"fef00809",
          9198 => x"70307072",
          9199 => x"07802551",
          9200 => x"5b5b5f80",
          9201 => x"5a7b8326",
          9202 => x"8338815a",
          9203 => x"787a0659",
          9204 => x"78802e8d",
          9205 => x"38811c70",
          9206 => x"81ff065d",
          9207 => x"597bfec0",
          9208 => x"387d8132",
          9209 => x"7d813207",
          9210 => x"59788a38",
          9211 => x"7eff2e09",
          9212 => x"8106ee8c",
          9213 => x"3881f9b4",
          9214 => x"51fedc8d",
          9215 => x"3fee8139",
          9216 => x"fc3d0d80",
          9217 => x"0b81ffb8",
          9218 => x"3487c094",
          9219 => x"8c700854",
          9220 => x"55878480",
          9221 => x"527251fe",
          9222 => x"b3913f81",
          9223 => x"fef00890",
          9224 => x"2b750855",
          9225 => x"53878480",
          9226 => x"527351fe",
          9227 => x"b2fd3f72",
          9228 => x"81fef008",
          9229 => x"07750c87",
          9230 => x"c0949c70",
          9231 => x"08545587",
          9232 => x"84805272",
          9233 => x"51feb2e3",
          9234 => x"3f81fef0",
          9235 => x"08902b75",
          9236 => x"08555387",
          9237 => x"84805273",
          9238 => x"51feb2cf",
          9239 => x"3f7281fe",
          9240 => x"f0080775",
          9241 => x"0c8c8083",
          9242 => x"0b87c094",
          9243 => x"840c8c80",
          9244 => x"830b87c0",
          9245 => x"94940ca3",
          9246 => x"8b0b81ff",
          9247 => x"840ca68c",
          9248 => x"0b81ff88",
          9249 => x"0cfec6ad",
          9250 => x"3ffed095",
          9251 => x"3f81f9c4",
          9252 => x"51fed591",
          9253 => x"3f81f9d0",
          9254 => x"51fed589",
          9255 => x"3f81c9e4",
          9256 => x"51fecfb7",
          9257 => x"3f8151e7",
          9258 => x"fc3fec84",
          9259 => x"3f800400",
          9260 => x"00ffffff",
          9261 => x"ff00ffff",
          9262 => x"ffff00ff",
          9263 => x"ffffff00",
          9264 => x"00001832",
          9265 => x"00001838",
          9266 => x"0000183e",
          9267 => x"00001844",
          9268 => x"0000184a",
          9269 => x"000025f6",
          9270 => x"000026d2",
          9271 => x"00002775",
          9272 => x"000027b5",
          9273 => x"000027d8",
          9274 => x"00002865",
          9275 => x"000024cb",
          9276 => x"000024cb",
          9277 => x"000028a2",
          9278 => x"00002918",
          9279 => x"000029a3",
          9280 => x"000029cc",
          9281 => x"000061ea",
          9282 => x"0000616e",
          9283 => x"00006175",
          9284 => x"0000617c",
          9285 => x"00006183",
          9286 => x"0000618a",
          9287 => x"00006191",
          9288 => x"00006198",
          9289 => x"0000619f",
          9290 => x"000061a6",
          9291 => x"000061ad",
          9292 => x"000061b4",
          9293 => x"000061ba",
          9294 => x"000061c0",
          9295 => x"000061c6",
          9296 => x"000061cc",
          9297 => x"000061d2",
          9298 => x"000061d8",
          9299 => x"000061de",
          9300 => x"000061e4",
          9301 => x"25642f25",
          9302 => x"642f2564",
          9303 => x"2025643a",
          9304 => x"25643a25",
          9305 => x"642e2564",
          9306 => x"25640a00",
          9307 => x"536f4320",
          9308 => x"436f6e66",
          9309 => x"69677572",
          9310 => x"6174696f",
          9311 => x"6e000000",
          9312 => x"20286672",
          9313 => x"6f6d2053",
          9314 => x"6f432063",
          9315 => x"6f6e6669",
          9316 => x"67290000",
          9317 => x"3a0a4465",
          9318 => x"76696365",
          9319 => x"7320696d",
          9320 => x"706c656d",
          9321 => x"656e7465",
          9322 => x"643a0a00",
          9323 => x"20202020",
          9324 => x"57422053",
          9325 => x"4452414d",
          9326 => x"20202825",
          9327 => x"3038583a",
          9328 => x"25303858",
          9329 => x"292e0a00",
          9330 => x"20202020",
          9331 => x"53445241",
          9332 => x"4d202020",
          9333 => x"20202825",
          9334 => x"3038583a",
          9335 => x"25303858",
          9336 => x"292e0a00",
          9337 => x"20202020",
          9338 => x"494e534e",
          9339 => x"20425241",
          9340 => x"4d202825",
          9341 => x"3038583a",
          9342 => x"25303858",
          9343 => x"292e0a00",
          9344 => x"20202020",
          9345 => x"4252414d",
          9346 => x"20202020",
          9347 => x"20202825",
          9348 => x"3038583a",
          9349 => x"25303858",
          9350 => x"292e0a00",
          9351 => x"20202020",
          9352 => x"52414d20",
          9353 => x"20202020",
          9354 => x"20202825",
          9355 => x"3038583a",
          9356 => x"25303858",
          9357 => x"292e0a00",
          9358 => x"20202020",
          9359 => x"53442043",
          9360 => x"41524420",
          9361 => x"20202844",
          9362 => x"65766963",
          9363 => x"6573203d",
          9364 => x"25303264",
          9365 => x"292e0a00",
          9366 => x"20202020",
          9367 => x"54494d45",
          9368 => x"52312020",
          9369 => x"20202854",
          9370 => x"696d6572",
          9371 => x"7320203d",
          9372 => x"25303264",
          9373 => x"292e0a00",
          9374 => x"20202020",
          9375 => x"494e5452",
          9376 => x"20435452",
          9377 => x"4c202843",
          9378 => x"68616e6e",
          9379 => x"656c733d",
          9380 => x"25303264",
          9381 => x"292e0a00",
          9382 => x"20202020",
          9383 => x"57495348",
          9384 => x"424f4e45",
          9385 => x"20425553",
          9386 => x"0a000000",
          9387 => x"20202020",
          9388 => x"57422049",
          9389 => x"32430a00",
          9390 => x"20202020",
          9391 => x"494f4354",
          9392 => x"4c0a0000",
          9393 => x"20202020",
          9394 => x"5053320a",
          9395 => x"00000000",
          9396 => x"20202020",
          9397 => x"5350490a",
          9398 => x"00000000",
          9399 => x"41646472",
          9400 => x"65737365",
          9401 => x"733a0a00",
          9402 => x"20202020",
          9403 => x"43505520",
          9404 => x"52657365",
          9405 => x"74205665",
          9406 => x"63746f72",
          9407 => x"20416464",
          9408 => x"72657373",
          9409 => x"203d2025",
          9410 => x"3038580a",
          9411 => x"00000000",
          9412 => x"20202020",
          9413 => x"43505520",
          9414 => x"4d656d6f",
          9415 => x"72792053",
          9416 => x"74617274",
          9417 => x"20416464",
          9418 => x"72657373",
          9419 => x"203d2025",
          9420 => x"3038580a",
          9421 => x"00000000",
          9422 => x"20202020",
          9423 => x"53746163",
          9424 => x"6b205374",
          9425 => x"61727420",
          9426 => x"41646472",
          9427 => x"65737320",
          9428 => x"20202020",
          9429 => x"203d2025",
          9430 => x"3038580a",
          9431 => x"00000000",
          9432 => x"4d697363",
          9433 => x"3a0a0000",
          9434 => x"20202020",
          9435 => x"5a505520",
          9436 => x"49642020",
          9437 => x"20202020",
          9438 => x"20202020",
          9439 => x"20202020",
          9440 => x"20202020",
          9441 => x"203d2025",
          9442 => x"3034580a",
          9443 => x"00000000",
          9444 => x"20202020",
          9445 => x"53797374",
          9446 => x"656d2043",
          9447 => x"6c6f636b",
          9448 => x"20467265",
          9449 => x"71202020",
          9450 => x"20202020",
          9451 => x"203d2025",
          9452 => x"642e2530",
          9453 => x"34644d48",
          9454 => x"7a0a0000",
          9455 => x"20202020",
          9456 => x"53445241",
          9457 => x"4d20436c",
          9458 => x"6f636b20",
          9459 => x"46726571",
          9460 => x"20202020",
          9461 => x"20202020",
          9462 => x"203d2025",
          9463 => x"642e2530",
          9464 => x"34644d48",
          9465 => x"7a0a0000",
          9466 => x"20202020",
          9467 => x"57697368",
          9468 => x"626f6e65",
          9469 => x"20534452",
          9470 => x"414d2043",
          9471 => x"6c6f636b",
          9472 => x"20467265",
          9473 => x"713d2025",
          9474 => x"642e2530",
          9475 => x"34644d48",
          9476 => x"7a0a0000",
          9477 => x"536d616c",
          9478 => x"6c000000",
          9479 => x"4d656469",
          9480 => x"756d0000",
          9481 => x"466c6578",
          9482 => x"00000000",
          9483 => x"45564f00",
          9484 => x"45564f6d",
          9485 => x"696e0000",
          9486 => x"556e6b6e",
          9487 => x"6f776e00",
          9488 => x"68697374",
          9489 => x"6f72792e",
          9490 => x"74787400",
          9491 => x"68697374",
          9492 => x"6f727900",
          9493 => x"68697374",
          9494 => x"00000000",
          9495 => x"21000000",
          9496 => x"25303464",
          9497 => x"20202573",
          9498 => x"0a000000",
          9499 => x"4661696c",
          9500 => x"65642074",
          9501 => x"6f207265",
          9502 => x"73657420",
          9503 => x"74686520",
          9504 => x"68697374",
          9505 => x"6f727920",
          9506 => x"66696c65",
          9507 => x"20746f20",
          9508 => x"454f462e",
          9509 => x"0a000000",
          9510 => x"43616e6e",
          9511 => x"6f74206f",
          9512 => x"70656e2f",
          9513 => x"63726561",
          9514 => x"74652068",
          9515 => x"6973746f",
          9516 => x"72792066",
          9517 => x"696c652c",
          9518 => x"20646973",
          9519 => x"61626c69",
          9520 => x"6e672e0a",
          9521 => x"00000000",
          9522 => x"00007574",
          9523 => x"01000000",
          9524 => x"00000001",
          9525 => x"00007570",
          9526 => x"01000000",
          9527 => x"00000002",
          9528 => x"0000756c",
          9529 => x"04000000",
          9530 => x"00000003",
          9531 => x"00007568",
          9532 => x"04000000",
          9533 => x"00000004",
          9534 => x"00007564",
          9535 => x"04000000",
          9536 => x"00000005",
          9537 => x"00007560",
          9538 => x"04000000",
          9539 => x"00000006",
          9540 => x"0000755c",
          9541 => x"04000000",
          9542 => x"00000007",
          9543 => x"00007558",
          9544 => x"03000000",
          9545 => x"00000008",
          9546 => x"00007554",
          9547 => x"03000000",
          9548 => x"00000009",
          9549 => x"00007550",
          9550 => x"03000000",
          9551 => x"0000000a",
          9552 => x"0000754c",
          9553 => x"03000000",
          9554 => x"0000000b",
          9555 => x"1b5b4400",
          9556 => x"1b5b4300",
          9557 => x"1b5b4200",
          9558 => x"1b5b4100",
          9559 => x"1b5b367e",
          9560 => x"1b5b357e",
          9561 => x"1b5b347e",
          9562 => x"1b5b337e",
          9563 => x"1b5b317e",
          9564 => x"0d000000",
          9565 => x"08000000",
          9566 => x"53440000",
          9567 => x"222a2b2c",
          9568 => x"3a3b3c3d",
          9569 => x"3e3f5b5d",
          9570 => x"7c7f0000",
          9571 => x"46415400",
          9572 => x"46415433",
          9573 => x"32000000",
          9574 => x"ebfe904d",
          9575 => x"53444f53",
          9576 => x"352e3000",
          9577 => x"4e4f204e",
          9578 => x"414d4520",
          9579 => x"20202046",
          9580 => x"41543332",
          9581 => x"20202000",
          9582 => x"4e4f204e",
          9583 => x"414d4520",
          9584 => x"20202046",
          9585 => x"41542020",
          9586 => x"20202000",
          9587 => x"00007578",
          9588 => x"00000000",
          9589 => x"00000000",
          9590 => x"00000000",
          9591 => x"809a4541",
          9592 => x"8e418f80",
          9593 => x"45454549",
          9594 => x"49498e8f",
          9595 => x"9092924f",
          9596 => x"994f5555",
          9597 => x"59999a9b",
          9598 => x"9c9d9e9f",
          9599 => x"41494f55",
          9600 => x"a5a5a6a7",
          9601 => x"a8a9aaab",
          9602 => x"acadaeaf",
          9603 => x"b0b1b2b3",
          9604 => x"b4b5b6b7",
          9605 => x"b8b9babb",
          9606 => x"bcbdbebf",
          9607 => x"c0c1c2c3",
          9608 => x"c4c5c6c7",
          9609 => x"c8c9cacb",
          9610 => x"cccdcecf",
          9611 => x"d0d1d2d3",
          9612 => x"d4d5d6d7",
          9613 => x"d8d9dadb",
          9614 => x"dcdddedf",
          9615 => x"e0e1e2e3",
          9616 => x"e4e5e6e7",
          9617 => x"e8e9eaeb",
          9618 => x"ecedeeef",
          9619 => x"f0f1f2f3",
          9620 => x"f4f5f6f7",
          9621 => x"f8f9fafb",
          9622 => x"fcfdfeff",
          9623 => x"2b2e2c3b",
          9624 => x"3d5b5d2f",
          9625 => x"5c222a3a",
          9626 => x"3c3e3f7c",
          9627 => x"7f000000",
          9628 => x"00010004",
          9629 => x"00100040",
          9630 => x"01000200",
          9631 => x"00000000",
          9632 => x"00010002",
          9633 => x"00040008",
          9634 => x"00100020",
          9635 => x"00000000",
          9636 => x"64696e69",
          9637 => x"74000000",
          9638 => x"64696f63",
          9639 => x"746c0000",
          9640 => x"66696e69",
          9641 => x"74000000",
          9642 => x"666c6f61",
          9643 => x"64000000",
          9644 => x"66657865",
          9645 => x"63000000",
          9646 => x"6d636c65",
          9647 => x"61720000",
          9648 => x"6d636f70",
          9649 => x"79000000",
          9650 => x"6d646966",
          9651 => x"66000000",
          9652 => x"6d64756d",
          9653 => x"70000000",
          9654 => x"6d656200",
          9655 => x"6d656800",
          9656 => x"6d657700",
          9657 => x"68696400",
          9658 => x"68696500",
          9659 => x"68666400",
          9660 => x"68666500",
          9661 => x"63616c6c",
          9662 => x"00000000",
          9663 => x"6a6d7000",
          9664 => x"72657374",
          9665 => x"61727400",
          9666 => x"72657365",
          9667 => x"74000000",
          9668 => x"696e666f",
          9669 => x"00000000",
          9670 => x"74657374",
          9671 => x"00000000",
          9672 => x"74626173",
          9673 => x"69630000",
          9674 => x"6d626173",
          9675 => x"69630000",
          9676 => x"6b696c6f",
          9677 => x"00000000",
          9678 => x"4469736b",
          9679 => x"20457272",
          9680 => x"6f720a00",
          9681 => x"496e7465",
          9682 => x"726e616c",
          9683 => x"20657272",
          9684 => x"6f722e0a",
          9685 => x"00000000",
          9686 => x"4469736b",
          9687 => x"206e6f74",
          9688 => x"20726561",
          9689 => x"64792e0a",
          9690 => x"00000000",
          9691 => x"4e6f2066",
          9692 => x"696c6520",
          9693 => x"666f756e",
          9694 => x"642e0a00",
          9695 => x"4e6f2070",
          9696 => x"61746820",
          9697 => x"666f756e",
          9698 => x"642e0a00",
          9699 => x"496e7661",
          9700 => x"6c696420",
          9701 => x"66696c65",
          9702 => x"6e616d65",
          9703 => x"2e0a0000",
          9704 => x"41636365",
          9705 => x"73732064",
          9706 => x"656e6965",
          9707 => x"642e0a00",
          9708 => x"46696c65",
          9709 => x"20616c72",
          9710 => x"65616479",
          9711 => x"20657869",
          9712 => x"7374732e",
          9713 => x"0a000000",
          9714 => x"46696c65",
          9715 => x"2068616e",
          9716 => x"646c6520",
          9717 => x"696e7661",
          9718 => x"6c69642e",
          9719 => x"0a000000",
          9720 => x"53442069",
          9721 => x"73207772",
          9722 => x"69746520",
          9723 => x"70726f74",
          9724 => x"65637465",
          9725 => x"642e0a00",
          9726 => x"44726976",
          9727 => x"65206e75",
          9728 => x"6d626572",
          9729 => x"20697320",
          9730 => x"696e7661",
          9731 => x"6c69642e",
          9732 => x"0a000000",
          9733 => x"4469736b",
          9734 => x"206e6f74",
          9735 => x"20656e61",
          9736 => x"626c6564",
          9737 => x"2e0a0000",
          9738 => x"4e6f2063",
          9739 => x"6f6d7061",
          9740 => x"7469626c",
          9741 => x"65206669",
          9742 => x"6c657379",
          9743 => x"7374656d",
          9744 => x"20666f75",
          9745 => x"6e64206f",
          9746 => x"6e206469",
          9747 => x"736b2e0a",
          9748 => x"00000000",
          9749 => x"466f726d",
          9750 => x"61742061",
          9751 => x"626f7274",
          9752 => x"65642e0a",
          9753 => x"00000000",
          9754 => x"54696d65",
          9755 => x"6f75742c",
          9756 => x"206f7065",
          9757 => x"72617469",
          9758 => x"6f6e2063",
          9759 => x"616e6365",
          9760 => x"6c6c6564",
          9761 => x"2e0a0000",
          9762 => x"46696c65",
          9763 => x"20697320",
          9764 => x"6c6f636b",
          9765 => x"65642e0a",
          9766 => x"00000000",
          9767 => x"496e7375",
          9768 => x"66666963",
          9769 => x"69656e74",
          9770 => x"206d656d",
          9771 => x"6f72792e",
          9772 => x"0a000000",
          9773 => x"546f6f20",
          9774 => x"6d616e79",
          9775 => x"206f7065",
          9776 => x"6e206669",
          9777 => x"6c65732e",
          9778 => x"0a000000",
          9779 => x"50617261",
          9780 => x"6d657465",
          9781 => x"72732069",
          9782 => x"6e636f72",
          9783 => x"72656374",
          9784 => x"2e0a0000",
          9785 => x"53756363",
          9786 => x"6573732e",
          9787 => x"0a000000",
          9788 => x"556e6b6e",
          9789 => x"6f776e20",
          9790 => x"6572726f",
          9791 => x"722e0a00",
          9792 => x"0a256c75",
          9793 => x"20627974",
          9794 => x"65732025",
          9795 => x"73206174",
          9796 => x"20256c75",
          9797 => x"20627974",
          9798 => x"65732f73",
          9799 => x"65632e0a",
          9800 => x"00000000",
          9801 => x"72656164",
          9802 => x"00000000",
          9803 => x"25303858",
          9804 => x"00000000",
          9805 => x"3a202000",
          9806 => x"25303458",
          9807 => x"00000000",
          9808 => x"20202020",
          9809 => x"20202020",
          9810 => x"00000000",
          9811 => x"25303258",
          9812 => x"00000000",
          9813 => x"20200000",
          9814 => x"207c0000",
          9815 => x"7c0d0a00",
          9816 => x"5a505554",
          9817 => x"41000000",
          9818 => x"0a2a2a20",
          9819 => x"25732028",
          9820 => x"00000000",
          9821 => x"32312f30",
          9822 => x"342f3230",
          9823 => x"32300000",
          9824 => x"76312e35",
          9825 => x"31000000",
          9826 => x"205a5055",
          9827 => x"2c207265",
          9828 => x"76202530",
          9829 => x"32782920",
          9830 => x"25732025",
          9831 => x"73202a2a",
          9832 => x"0a0a0000",
          9833 => x"5a505554",
          9834 => x"4120496e",
          9835 => x"74657272",
          9836 => x"75707420",
          9837 => x"48616e64",
          9838 => x"6c65720a",
          9839 => x"00000000",
          9840 => x"54696d65",
          9841 => x"7220696e",
          9842 => x"74657272",
          9843 => x"7570740a",
          9844 => x"00000000",
          9845 => x"50533220",
          9846 => x"696e7465",
          9847 => x"72727570",
          9848 => x"740a0000",
          9849 => x"494f4354",
          9850 => x"4c205244",
          9851 => x"20696e74",
          9852 => x"65727275",
          9853 => x"70740a00",
          9854 => x"494f4354",
          9855 => x"4c205752",
          9856 => x"20696e74",
          9857 => x"65727275",
          9858 => x"70740a00",
          9859 => x"55415254",
          9860 => x"30205258",
          9861 => x"20696e74",
          9862 => x"65727275",
          9863 => x"70740a00",
          9864 => x"55415254",
          9865 => x"30205458",
          9866 => x"20696e74",
          9867 => x"65727275",
          9868 => x"70740a00",
          9869 => x"55415254",
          9870 => x"31205258",
          9871 => x"20696e74",
          9872 => x"65727275",
          9873 => x"70740a00",
          9874 => x"55415254",
          9875 => x"31205458",
          9876 => x"20696e74",
          9877 => x"65727275",
          9878 => x"70740a00",
          9879 => x"53657474",
          9880 => x"696e6720",
          9881 => x"75702074",
          9882 => x"696d6572",
          9883 => x"2e2e2e0a",
          9884 => x"00000000",
          9885 => x"456e6162",
          9886 => x"6c696e67",
          9887 => x"2074696d",
          9888 => x"65722e2e",
          9889 => x"2e0a0000",
          9890 => x"6175746f",
          9891 => x"65786563",
          9892 => x"2e626174",
          9893 => x"00000000",
          9894 => x"303a0000",
          9895 => x"4661696c",
          9896 => x"65642074",
          9897 => x"6f20696e",
          9898 => x"69746961",
          9899 => x"6c697365",
          9900 => x"20736420",
          9901 => x"63617264",
          9902 => x"20302c20",
          9903 => x"706c6561",
          9904 => x"73652069",
          9905 => x"6e697420",
          9906 => x"6d616e75",
          9907 => x"616c6c79",
          9908 => x"2e0a0000",
          9909 => x"2a200000",
          9910 => x"42616420",
          9911 => x"6469736b",
          9912 => x"20696421",
          9913 => x"0a000000",
          9914 => x"496e6974",
          9915 => x"69616c69",
          9916 => x"7365642e",
          9917 => x"0a000000",
          9918 => x"4661696c",
          9919 => x"65642074",
          9920 => x"6f20696e",
          9921 => x"69746961",
          9922 => x"6c697365",
          9923 => x"2e0a0000",
          9924 => x"72633d25",
          9925 => x"640a0000",
          9926 => x"25753a00",
          9927 => x"436c6561",
          9928 => x"72696e67",
          9929 => x"2e2e2e2e",
          9930 => x"00000000",
          9931 => x"436f7079",
          9932 => x"696e672e",
          9933 => x"2e2e0000",
          9934 => x"436f6d70",
          9935 => x"6172696e",
          9936 => x"672e2e2e",
          9937 => x"00000000",
          9938 => x"2530386c",
          9939 => x"78282530",
          9940 => x"3878292d",
          9941 => x"3e253038",
          9942 => x"6c782825",
          9943 => x"30387829",
          9944 => x"0a000000",
          9945 => x"44756d70",
          9946 => x"204d656d",
          9947 => x"6f72790a",
          9948 => x"00000000",
          9949 => x"0a436f6d",
          9950 => x"706c6574",
          9951 => x"652e0a00",
          9952 => x"25303858",
          9953 => x"20253032",
          9954 => x"582d0000",
          9955 => x"3f3f3f0a",
          9956 => x"00000000",
          9957 => x"25303858",
          9958 => x"20253034",
          9959 => x"582d0000",
          9960 => x"25303858",
          9961 => x"20253038",
          9962 => x"582d0000",
          9963 => x"44697361",
          9964 => x"626c696e",
          9965 => x"6720696e",
          9966 => x"74657272",
          9967 => x"75707473",
          9968 => x"0a000000",
          9969 => x"456e6162",
          9970 => x"6c696e67",
          9971 => x"20696e74",
          9972 => x"65727275",
          9973 => x"7074730a",
          9974 => x"00000000",
          9975 => x"44697361",
          9976 => x"626c6564",
          9977 => x"20756172",
          9978 => x"74206669",
          9979 => x"666f0a00",
          9980 => x"456e6162",
          9981 => x"6c696e67",
          9982 => x"20756172",
          9983 => x"74206669",
          9984 => x"666f0a00",
          9985 => x"45786563",
          9986 => x"7574696e",
          9987 => x"6720636f",
          9988 => x"64652040",
          9989 => x"20253038",
          9990 => x"78202e2e",
          9991 => x"2e0a0000",
          9992 => x"43616c6c",
          9993 => x"696e6720",
          9994 => x"636f6465",
          9995 => x"20402025",
          9996 => x"30387820",
          9997 => x"2e2e2e0a",
          9998 => x"00000000",
          9999 => x"43616c6c",
         10000 => x"20726574",
         10001 => x"75726e65",
         10002 => x"6420636f",
         10003 => x"64652028",
         10004 => x"2564292e",
         10005 => x"0a000000",
         10006 => x"52657374",
         10007 => x"61727469",
         10008 => x"6e672061",
         10009 => x"70706c69",
         10010 => x"63617469",
         10011 => x"6f6e2e2e",
         10012 => x"2e0a0000",
         10013 => x"436f6c64",
         10014 => x"20726562",
         10015 => x"6f6f7469",
         10016 => x"6e672e2e",
         10017 => x"2e0a0000",
         10018 => x"5a505500",
         10019 => x"62696e00",
         10020 => x"25643a5c",
         10021 => x"25735c25",
         10022 => x"732e2573",
         10023 => x"00000000",
         10024 => x"25643a5c",
         10025 => x"25735c25",
         10026 => x"73000000",
         10027 => x"25643a5c",
         10028 => x"25730000",
         10029 => x"42616420",
         10030 => x"636f6d6d",
         10031 => x"616e642e",
         10032 => x"0a000000",
         10033 => x"52756e6e",
         10034 => x"696e672e",
         10035 => x"2e2e0a00",
         10036 => x"456e6162",
         10037 => x"6c696e67",
         10038 => x"20696e74",
         10039 => x"65727275",
         10040 => x"7074732e",
         10041 => x"2e2e0a00",
         10042 => x"00000000",
         10043 => x"00000000",
         10044 => x"00007fff",
         10045 => x"00000000",
         10046 => x"00007fff",
         10047 => x"00010000",
         10048 => x"00007fff",
         10049 => x"00010000",
         10050 => x"00810000",
         10051 => x"01000000",
         10052 => x"017fffff",
         10053 => x"00000000",
         10054 => x"00000000",
         10055 => x"00007800",
         10056 => x"00000000",
         10057 => x"05f5e100",
         10058 => x"05f5e100",
         10059 => x"05f5e100",
         10060 => x"00000000",
         10061 => x"01010101",
         10062 => x"01010101",
         10063 => x"01011001",
         10064 => x"01000000",
         10065 => x"00000000",
         10066 => x"00000002",
         10067 => x"00000000",
         10068 => x"00007d48",
         10069 => x"00007d48",
         10070 => x"00007d48",
         10071 => x"00007d48",
         10072 => x"00007440",
         10073 => x"00000000",
         10074 => x"00000000",
         10075 => x"00000000",
         10076 => x"00000000",
         10077 => x"00000000",
         10078 => x"00000000",
         10079 => x"00000000",
         10080 => x"00000000",
         10081 => x"00000000",
         10082 => x"00000000",
         10083 => x"00000000",
         10084 => x"00000000",
         10085 => x"00000000",
         10086 => x"00000000",
         10087 => x"00000000",
         10088 => x"00000000",
         10089 => x"00000000",
         10090 => x"00000000",
         10091 => x"00000000",
         10092 => x"00000000",
         10093 => x"00000000",
         10094 => x"00000000",
         10095 => x"00000000",
         10096 => x"0000744c",
         10097 => x"01000000",
         10098 => x"00007454",
         10099 => x"01000000",
         10100 => x"0000745c",
         10101 => x"02000000",
         10102 => x"01000000",
         10103 => x"00000000",
         10104 => x"00007690",
         10105 => x"01020100",
         10106 => x"00000000",
         10107 => x"00000000",
         10108 => x"00007698",
         10109 => x"01040100",
         10110 => x"00000000",
         10111 => x"00000000",
         10112 => x"000076a0",
         10113 => x"01140300",
         10114 => x"00000000",
         10115 => x"00000000",
         10116 => x"000076a8",
         10117 => x"012b0300",
         10118 => x"00000000",
         10119 => x"00000000",
         10120 => x"000076b0",
         10121 => x"01300300",
         10122 => x"00000000",
         10123 => x"00000000",
         10124 => x"000076b8",
         10125 => x"013c0400",
         10126 => x"00000000",
         10127 => x"00000000",
         10128 => x"000076c0",
         10129 => x"013d0400",
         10130 => x"00000000",
         10131 => x"00000000",
         10132 => x"000076c8",
         10133 => x"013f0400",
         10134 => x"00000000",
         10135 => x"00000000",
         10136 => x"000076d0",
         10137 => x"01400400",
         10138 => x"00000000",
         10139 => x"00000000",
         10140 => x"000076d8",
         10141 => x"01410400",
         10142 => x"00000000",
         10143 => x"00000000",
         10144 => x"000076dc",
         10145 => x"01420400",
         10146 => x"00000000",
         10147 => x"00000000",
         10148 => x"000076e0",
         10149 => x"01430400",
         10150 => x"00000000",
         10151 => x"00000000",
         10152 => x"000076e4",
         10153 => x"01500500",
         10154 => x"00000000",
         10155 => x"00000000",
         10156 => x"000076e8",
         10157 => x"01510500",
         10158 => x"00000000",
         10159 => x"00000000",
         10160 => x"000076ec",
         10161 => x"01540500",
         10162 => x"00000000",
         10163 => x"00000000",
         10164 => x"000076f0",
         10165 => x"01550500",
         10166 => x"00000000",
         10167 => x"00000000",
         10168 => x"000076f4",
         10169 => x"01790700",
         10170 => x"00000000",
         10171 => x"00000000",
         10172 => x"000076fc",
         10173 => x"01780700",
         10174 => x"00000000",
         10175 => x"00000000",
         10176 => x"00007700",
         10177 => x"01820800",
         10178 => x"00000000",
         10179 => x"00000000",
         10180 => x"00007708",
         10181 => x"01830800",
         10182 => x"00000000",
         10183 => x"00000000",
         10184 => x"00007710",
         10185 => x"01850800",
         10186 => x"00000000",
         10187 => x"00000000",
         10188 => x"00007718",
         10189 => x"01870800",
         10190 => x"00000000",
         10191 => x"00000000",
         10192 => x"00007720",
         10193 => x"018c0900",
         10194 => x"00000000",
         10195 => x"00000000",
         10196 => x"00007728",
         10197 => x"018d0900",
         10198 => x"00000000",
         10199 => x"00000000",
         10200 => x"00007730",
         10201 => x"018e0900",
         10202 => x"00000000",
         10203 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

