-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b83ff",
          2049 => x"f80d0b0b",
          2050 => x"0b93b904",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"9d040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b9380",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b8295",
          2210 => x"98738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93850400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b80c3",
          2219 => x"f42d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b80c5",
          2227 => x"e02d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"95040b0b",
          2317 => x"0b8ca404",
          2318 => x"0b0b0b8c",
          2319 => x"b3040b0b",
          2320 => x"0b8cc204",
          2321 => x"0b0b0b8c",
          2322 => x"d1040b0b",
          2323 => x"0b8ce004",
          2324 => x"0b0b0b8c",
          2325 => x"f0040b0b",
          2326 => x"0b8d8004",
          2327 => x"0b0b0b8d",
          2328 => x"8f040b0b",
          2329 => x"0b8d9e04",
          2330 => x"0b0b0b8d",
          2331 => x"ad040b0b",
          2332 => x"0b8dbd04",
          2333 => x"0b0b0b8d",
          2334 => x"cd040b0b",
          2335 => x"0b8ddd04",
          2336 => x"0b0b0b8d",
          2337 => x"ed040b0b",
          2338 => x"0b8dfd04",
          2339 => x"0b0b0b8e",
          2340 => x"8d040b0b",
          2341 => x"0b8e9d04",
          2342 => x"0b0b0b8e",
          2343 => x"ad040b0b",
          2344 => x"0b8ebd04",
          2345 => x"0b0b0b8e",
          2346 => x"cd040b0b",
          2347 => x"0b8edd04",
          2348 => x"0b0b0b8e",
          2349 => x"ed040b0b",
          2350 => x"0b8efd04",
          2351 => x"0b0b0b8f",
          2352 => x"8d040b0b",
          2353 => x"0b8f9d04",
          2354 => x"0b0b0b8f",
          2355 => x"ad040b0b",
          2356 => x"0b8fbd04",
          2357 => x"0b0b0b8f",
          2358 => x"cd040b0b",
          2359 => x"0b8fdd04",
          2360 => x"0b0b0b8f",
          2361 => x"ed040b0b",
          2362 => x"0b8ffd04",
          2363 => x"0b0b0b90",
          2364 => x"8d040b0b",
          2365 => x"0b909d04",
          2366 => x"0b0b0b90",
          2367 => x"ad040b0b",
          2368 => x"0b90bd04",
          2369 => x"0b0b0b90",
          2370 => x"cd040b0b",
          2371 => x"0b90dd04",
          2372 => x"0b0b0b90",
          2373 => x"ed040b0b",
          2374 => x"0b90fd04",
          2375 => x"0b0b0b91",
          2376 => x"8d040b0b",
          2377 => x"0b919d04",
          2378 => x"0b0b0b91",
          2379 => x"ad040b0b",
          2380 => x"0b91bd04",
          2381 => x"0b0b0b91",
          2382 => x"cd040b0b",
          2383 => x"0b91dd04",
          2384 => x"0b0b0b91",
          2385 => x"ed040b0b",
          2386 => x"0b91fd04",
          2387 => x"0b0b0b92",
          2388 => x"8d040b0b",
          2389 => x"0b929d04",
          2390 => x"0b0b0b92",
          2391 => x"ad040b0b",
          2392 => x"0b92bd04",
          2393 => x"0b0b0b92",
          2394 => x"cd04ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0482b5d4",
          2434 => x"0c80f4da",
          2435 => x"2d82b5d4",
          2436 => x"0882d090",
          2437 => x"0482b5d4",
          2438 => x"0cb3b22d",
          2439 => x"82b5d408",
          2440 => x"82d09004",
          2441 => x"82b5d40c",
          2442 => x"afe32d82",
          2443 => x"b5d40882",
          2444 => x"d0900482",
          2445 => x"b5d40caf",
          2446 => x"ad2d82b5",
          2447 => x"d40882d0",
          2448 => x"900482b5",
          2449 => x"d40c94ad",
          2450 => x"2d82b5d4",
          2451 => x"0882d090",
          2452 => x"0482b5d4",
          2453 => x"0cb1c22d",
          2454 => x"82b5d408",
          2455 => x"82d09004",
          2456 => x"82b5d40c",
          2457 => x"80cfcc2d",
          2458 => x"82b5d408",
          2459 => x"82d09004",
          2460 => x"82b5d40c",
          2461 => x"80c9fb2d",
          2462 => x"82b5d408",
          2463 => x"82d09004",
          2464 => x"82b5d40c",
          2465 => x"93d82d82",
          2466 => x"b5d40882",
          2467 => x"d0900482",
          2468 => x"b5d40c96",
          2469 => x"c02d82b5",
          2470 => x"d40882d0",
          2471 => x"900482b5",
          2472 => x"d40c97cd",
          2473 => x"2d82b5d4",
          2474 => x"0882d090",
          2475 => x"0482b5d4",
          2476 => x"0c80f884",
          2477 => x"2d82b5d4",
          2478 => x"0882d090",
          2479 => x"0482b5d4",
          2480 => x"0c80f8e2",
          2481 => x"2d82b5d4",
          2482 => x"0882d090",
          2483 => x"0482b5d4",
          2484 => x"0c80f09f",
          2485 => x"2d82b5d4",
          2486 => x"0882d090",
          2487 => x"0482b5d4",
          2488 => x"0c80f296",
          2489 => x"2d82b5d4",
          2490 => x"0882d090",
          2491 => x"0482b5d4",
          2492 => x"0c80f3c9",
          2493 => x"2d82b5d4",
          2494 => x"0882d090",
          2495 => x"0482b5d4",
          2496 => x"0c81d7fc",
          2497 => x"2d82b5d4",
          2498 => x"0882d090",
          2499 => x"0482b5d4",
          2500 => x"0c81e4ed",
          2501 => x"2d82b5d4",
          2502 => x"0882d090",
          2503 => x"0482b5d4",
          2504 => x"0c81dce1",
          2505 => x"2d82b5d4",
          2506 => x"0882d090",
          2507 => x"0482b5d4",
          2508 => x"0c81dfde",
          2509 => x"2d82b5d4",
          2510 => x"0882d090",
          2511 => x"0482b5d4",
          2512 => x"0c81e9fc",
          2513 => x"2d82b5d4",
          2514 => x"0882d090",
          2515 => x"0482b5d4",
          2516 => x"0c81f2dc",
          2517 => x"2d82b5d4",
          2518 => x"0882d090",
          2519 => x"0482b5d4",
          2520 => x"0c81e3cf",
          2521 => x"2d82b5d4",
          2522 => x"0882d090",
          2523 => x"0482b5d4",
          2524 => x"0c81ed9b",
          2525 => x"2d82b5d4",
          2526 => x"0882d090",
          2527 => x"0482b5d4",
          2528 => x"0c81eeba",
          2529 => x"2d82b5d4",
          2530 => x"0882d090",
          2531 => x"0482b5d4",
          2532 => x"0c81eed9",
          2533 => x"2d82b5d4",
          2534 => x"0882d090",
          2535 => x"0482b5d4",
          2536 => x"0c81f6c3",
          2537 => x"2d82b5d4",
          2538 => x"0882d090",
          2539 => x"0482b5d4",
          2540 => x"0c81f4a9",
          2541 => x"2d82b5d4",
          2542 => x"0882d090",
          2543 => x"0482b5d4",
          2544 => x"0c81f997",
          2545 => x"2d82b5d4",
          2546 => x"0882d090",
          2547 => x"0482b5d4",
          2548 => x"0c81efdd",
          2549 => x"2d82b5d4",
          2550 => x"0882d090",
          2551 => x"0482b5d4",
          2552 => x"0c81fc97",
          2553 => x"2d82b5d4",
          2554 => x"0882d090",
          2555 => x"0482b5d4",
          2556 => x"0c81fd98",
          2557 => x"2d82b5d4",
          2558 => x"0882d090",
          2559 => x"0482b5d4",
          2560 => x"0c81e5cd",
          2561 => x"2d82b5d4",
          2562 => x"0882d090",
          2563 => x"0482b5d4",
          2564 => x"0c81e5a6",
          2565 => x"2d82b5d4",
          2566 => x"0882d090",
          2567 => x"0482b5d4",
          2568 => x"0c81e6d1",
          2569 => x"2d82b5d4",
          2570 => x"0882d090",
          2571 => x"0482b5d4",
          2572 => x"0c81f0b4",
          2573 => x"2d82b5d4",
          2574 => x"0882d090",
          2575 => x"0482b5d4",
          2576 => x"0c81fe89",
          2577 => x"2d82b5d4",
          2578 => x"0882d090",
          2579 => x"0482b5d4",
          2580 => x"0c828093",
          2581 => x"2d82b5d4",
          2582 => x"0882d090",
          2583 => x"0482b5d4",
          2584 => x"0c8283d5",
          2585 => x"2d82b5d4",
          2586 => x"0882d090",
          2587 => x"0482b5d4",
          2588 => x"0c81d79b",
          2589 => x"2d82b5d4",
          2590 => x"0882d090",
          2591 => x"0482b5d4",
          2592 => x"0c8286c1",
          2593 => x"2d82b5d4",
          2594 => x"0882d090",
          2595 => x"0482b5d4",
          2596 => x"0c8294f6",
          2597 => x"2d82b5d4",
          2598 => x"0882d090",
          2599 => x"0482b5d4",
          2600 => x"0c8292e2",
          2601 => x"2d82b5d4",
          2602 => x"0882d090",
          2603 => x"0482b5d4",
          2604 => x"0c81a8d6",
          2605 => x"2d82b5d4",
          2606 => x"0882d090",
          2607 => x"0482b5d4",
          2608 => x"0c81aac0",
          2609 => x"2d82b5d4",
          2610 => x"0882d090",
          2611 => x"0482b5d4",
          2612 => x"0c81aca4",
          2613 => x"2d82b5d4",
          2614 => x"0882d090",
          2615 => x"0482b5d4",
          2616 => x"0c80f0c8",
          2617 => x"2d82b5d4",
          2618 => x"0882d090",
          2619 => x"0482b5d4",
          2620 => x"0c80f1ec",
          2621 => x"2d82b5d4",
          2622 => x"0882d090",
          2623 => x"0482b5d4",
          2624 => x"0c80f5cf",
          2625 => x"2d82b5d4",
          2626 => x"0882d090",
          2627 => x"0482b5d4",
          2628 => x"0c80d698",
          2629 => x"2d82b5d4",
          2630 => x"0882d090",
          2631 => x"0482b5d4",
          2632 => x"0c81a2ea",
          2633 => x"2d82b5d4",
          2634 => x"0882d090",
          2635 => x"0482b5d4",
          2636 => x"0c81a392",
          2637 => x"2d82b5d4",
          2638 => x"0882d090",
          2639 => x"0482b5d4",
          2640 => x"0c81a78a",
          2641 => x"2d82b5d4",
          2642 => x"0882d090",
          2643 => x"0482b5d4",
          2644 => x"0c819fd4",
          2645 => x"2d82b5d4",
          2646 => x"0882d090",
          2647 => x"043c0400",
          2648 => x"00101010",
          2649 => x"10101010",
          2650 => x"10101010",
          2651 => x"10101010",
          2652 => x"10101010",
          2653 => x"10101010",
          2654 => x"10101010",
          2655 => x"10101010",
          2656 => x"53510400",
          2657 => x"007381ff",
          2658 => x"06738306",
          2659 => x"09810583",
          2660 => x"05101010",
          2661 => x"2b0772fc",
          2662 => x"060c5151",
          2663 => x"04727280",
          2664 => x"728106ff",
          2665 => x"05097206",
          2666 => x"05711052",
          2667 => x"720a100a",
          2668 => x"5372ed38",
          2669 => x"51515351",
          2670 => x"0482b5c8",
          2671 => x"7082cda4",
          2672 => x"278e3880",
          2673 => x"71708405",
          2674 => x"530c0b0b",
          2675 => x"0b93bc04",
          2676 => x"8c815180",
          2677 => x"eee20400",
          2678 => x"82b5d408",
          2679 => x"0282b5d4",
          2680 => x"0cfb3d0d",
          2681 => x"82b5d408",
          2682 => x"8c057082",
          2683 => x"b5d408fc",
          2684 => x"050c82b5",
          2685 => x"d408fc05",
          2686 => x"085482b5",
          2687 => x"d4088805",
          2688 => x"085382cd",
          2689 => x"9c085254",
          2690 => x"849a3f82",
          2691 => x"b5c80870",
          2692 => x"82b5d408",
          2693 => x"f8050c82",
          2694 => x"b5d408f8",
          2695 => x"05087082",
          2696 => x"b5c80c51",
          2697 => x"54873d0d",
          2698 => x"82b5d40c",
          2699 => x"0482b5d4",
          2700 => x"080282b5",
          2701 => x"d40cfb3d",
          2702 => x"0d82b5d4",
          2703 => x"08900508",
          2704 => x"85113370",
          2705 => x"81327081",
          2706 => x"06515151",
          2707 => x"52718f38",
          2708 => x"800b82b5",
          2709 => x"d4088c05",
          2710 => x"08258338",
          2711 => x"8d39800b",
          2712 => x"82b5d408",
          2713 => x"f4050c81",
          2714 => x"c43982b5",
          2715 => x"d4088c05",
          2716 => x"08ff0582",
          2717 => x"b5d4088c",
          2718 => x"050c800b",
          2719 => x"82b5d408",
          2720 => x"f8050c82",
          2721 => x"b5d40888",
          2722 => x"050882b5",
          2723 => x"d408fc05",
          2724 => x"0c82b5d4",
          2725 => x"08f80508",
          2726 => x"8a2e80f6",
          2727 => x"38800b82",
          2728 => x"b5d4088c",
          2729 => x"05082580",
          2730 => x"e93882b5",
          2731 => x"d4089005",
          2732 => x"0851a090",
          2733 => x"3f82b5c8",
          2734 => x"087082b5",
          2735 => x"d408f805",
          2736 => x"0c5282b5",
          2737 => x"d408f805",
          2738 => x"08ff2e09",
          2739 => x"81068d38",
          2740 => x"800b82b5",
          2741 => x"d408f405",
          2742 => x"0c80d239",
          2743 => x"82b5d408",
          2744 => x"fc050882",
          2745 => x"b5d408f8",
          2746 => x"05085353",
          2747 => x"71733482",
          2748 => x"b5d4088c",
          2749 => x"0508ff05",
          2750 => x"82b5d408",
          2751 => x"8c050c82",
          2752 => x"b5d408fc",
          2753 => x"05088105",
          2754 => x"82b5d408",
          2755 => x"fc050cff",
          2756 => x"803982b5",
          2757 => x"d408fc05",
          2758 => x"08528072",
          2759 => x"3482b5d4",
          2760 => x"08880508",
          2761 => x"7082b5d4",
          2762 => x"08f4050c",
          2763 => x"5282b5d4",
          2764 => x"08f40508",
          2765 => x"82b5c80c",
          2766 => x"873d0d82",
          2767 => x"b5d40c04",
          2768 => x"82b5d408",
          2769 => x"0282b5d4",
          2770 => x"0cf43d0d",
          2771 => x"860b82b5",
          2772 => x"d408e505",
          2773 => x"3482b5d4",
          2774 => x"08880508",
          2775 => x"82b5d408",
          2776 => x"e0050cfe",
          2777 => x"0a0b82b5",
          2778 => x"d408e805",
          2779 => x"0c82b5d4",
          2780 => x"08900570",
          2781 => x"82b5d408",
          2782 => x"fc050c82",
          2783 => x"b5d408fc",
          2784 => x"05085482",
          2785 => x"b5d4088c",
          2786 => x"05085382",
          2787 => x"b5d408e0",
          2788 => x"05705351",
          2789 => x"54818d3f",
          2790 => x"82b5c808",
          2791 => x"7082b5d4",
          2792 => x"08dc050c",
          2793 => x"82b5d408",
          2794 => x"ec050882",
          2795 => x"b5d40888",
          2796 => x"05080551",
          2797 => x"54807434",
          2798 => x"82b5d408",
          2799 => x"dc050870",
          2800 => x"82b5c80c",
          2801 => x"548e3d0d",
          2802 => x"82b5d40c",
          2803 => x"0482b5d4",
          2804 => x"080282b5",
          2805 => x"d40cfb3d",
          2806 => x"0d82b5d4",
          2807 => x"08900570",
          2808 => x"82b5d408",
          2809 => x"fc050c82",
          2810 => x"b5d408fc",
          2811 => x"05085482",
          2812 => x"b5d4088c",
          2813 => x"05085382",
          2814 => x"b5d40888",
          2815 => x"05085254",
          2816 => x"a33f82b5",
          2817 => x"c8087082",
          2818 => x"b5d408f8",
          2819 => x"050c82b5",
          2820 => x"d408f805",
          2821 => x"087082b5",
          2822 => x"c80c5154",
          2823 => x"873d0d82",
          2824 => x"b5d40c04",
          2825 => x"82b5d408",
          2826 => x"0282b5d4",
          2827 => x"0ced3d0d",
          2828 => x"800b82b5",
          2829 => x"d408e405",
          2830 => x"2382b5d4",
          2831 => x"08880508",
          2832 => x"53800b8c",
          2833 => x"140c82b5",
          2834 => x"d4088805",
          2835 => x"08851133",
          2836 => x"70812a70",
          2837 => x"81327081",
          2838 => x"06515151",
          2839 => x"51537280",
          2840 => x"2e8d38ff",
          2841 => x"0b82b5d4",
          2842 => x"08e0050c",
          2843 => x"96ac3982",
          2844 => x"b5d4088c",
          2845 => x"05085372",
          2846 => x"33537282",
          2847 => x"b5d408f8",
          2848 => x"05347281",
          2849 => x"ff065372",
          2850 => x"802e95fa",
          2851 => x"3882b5d4",
          2852 => x"088c0508",
          2853 => x"810582b5",
          2854 => x"d4088c05",
          2855 => x"0c82b5d4",
          2856 => x"08e40522",
          2857 => x"70810651",
          2858 => x"5372802e",
          2859 => x"958b3882",
          2860 => x"b5d408f8",
          2861 => x"053353af",
          2862 => x"732781fc",
          2863 => x"3882b5d4",
          2864 => x"08f80533",
          2865 => x"5372b926",
          2866 => x"81ee3882",
          2867 => x"b5d408f8",
          2868 => x"05335372",
          2869 => x"b02e0981",
          2870 => x"0680c538",
          2871 => x"82b5d408",
          2872 => x"e8053370",
          2873 => x"982b7098",
          2874 => x"2c515153",
          2875 => x"72b23882",
          2876 => x"b5d408e4",
          2877 => x"05227083",
          2878 => x"2a708132",
          2879 => x"70810651",
          2880 => x"51515372",
          2881 => x"802e9938",
          2882 => x"82b5d408",
          2883 => x"e4052270",
          2884 => x"82800751",
          2885 => x"537282b5",
          2886 => x"d408e405",
          2887 => x"23fed039",
          2888 => x"82b5d408",
          2889 => x"e8053370",
          2890 => x"982b7098",
          2891 => x"2c707083",
          2892 => x"2b721173",
          2893 => x"11515151",
          2894 => x"53515553",
          2895 => x"7282b5d4",
          2896 => x"08e80534",
          2897 => x"82b5d408",
          2898 => x"e8053354",
          2899 => x"82b5d408",
          2900 => x"f8053370",
          2901 => x"15d01151",
          2902 => x"51537282",
          2903 => x"b5d408e8",
          2904 => x"053482b5",
          2905 => x"d408e805",
          2906 => x"3370982b",
          2907 => x"70982c51",
          2908 => x"51537280",
          2909 => x"258b3880",
          2910 => x"ff0b82b5",
          2911 => x"d408e805",
          2912 => x"3482b5d4",
          2913 => x"08e40522",
          2914 => x"70832a70",
          2915 => x"81065151",
          2916 => x"5372fddb",
          2917 => x"3882b5d4",
          2918 => x"08e80533",
          2919 => x"70882b70",
          2920 => x"902b7090",
          2921 => x"2c70882c",
          2922 => x"51515151",
          2923 => x"537282b5",
          2924 => x"d408ec05",
          2925 => x"23fdb839",
          2926 => x"82b5d408",
          2927 => x"e4052270",
          2928 => x"832a7081",
          2929 => x"06515153",
          2930 => x"72802e9d",
          2931 => x"3882b5d4",
          2932 => x"08e80533",
          2933 => x"70982b70",
          2934 => x"982c5151",
          2935 => x"53728a38",
          2936 => x"810b82b5",
          2937 => x"d408e805",
          2938 => x"3482b5d4",
          2939 => x"08f80533",
          2940 => x"e01182b5",
          2941 => x"d408c405",
          2942 => x"0c5382b5",
          2943 => x"d408c405",
          2944 => x"0880d826",
          2945 => x"92943882",
          2946 => x"b5d408c4",
          2947 => x"05087082",
          2948 => x"2b8296e4",
          2949 => x"11700851",
          2950 => x"51515372",
          2951 => x"0482b5d4",
          2952 => x"08e40522",
          2953 => x"70900751",
          2954 => x"537282b5",
          2955 => x"d408e405",
          2956 => x"2382b5d4",
          2957 => x"08e40522",
          2958 => x"70a00751",
          2959 => x"537282b5",
          2960 => x"d408e405",
          2961 => x"23fca839",
          2962 => x"82b5d408",
          2963 => x"e4052270",
          2964 => x"81800751",
          2965 => x"537282b5",
          2966 => x"d408e405",
          2967 => x"23fc9039",
          2968 => x"82b5d408",
          2969 => x"e4052270",
          2970 => x"80c00751",
          2971 => x"537282b5",
          2972 => x"d408e405",
          2973 => x"23fbf839",
          2974 => x"82b5d408",
          2975 => x"e4052270",
          2976 => x"88075153",
          2977 => x"7282b5d4",
          2978 => x"08e40523",
          2979 => x"800b82b5",
          2980 => x"d408e805",
          2981 => x"34fbd839",
          2982 => x"82b5d408",
          2983 => x"e4052270",
          2984 => x"84075153",
          2985 => x"7282b5d4",
          2986 => x"08e40523",
          2987 => x"fbc139bf",
          2988 => x"0b82b5d4",
          2989 => x"08fc0534",
          2990 => x"82b5d408",
          2991 => x"ec0522ff",
          2992 => x"11515372",
          2993 => x"82b5d408",
          2994 => x"ec052380",
          2995 => x"e30b82b5",
          2996 => x"d408f805",
          2997 => x"348da839",
          2998 => x"82b5d408",
          2999 => x"90050882",
          3000 => x"b5d40890",
          3001 => x"05088405",
          3002 => x"82b5d408",
          3003 => x"90050c70",
          3004 => x"08515372",
          3005 => x"82b5d408",
          3006 => x"fc053482",
          3007 => x"b5d408ec",
          3008 => x"0522ff11",
          3009 => x"51537282",
          3010 => x"b5d408ec",
          3011 => x"05238cef",
          3012 => x"3982b5d4",
          3013 => x"08900508",
          3014 => x"82b5d408",
          3015 => x"90050884",
          3016 => x"0582b5d4",
          3017 => x"0890050c",
          3018 => x"700882b5",
          3019 => x"d408fc05",
          3020 => x"0c82b5d4",
          3021 => x"08e40522",
          3022 => x"70832a70",
          3023 => x"81065151",
          3024 => x"51537280",
          3025 => x"2eab3882",
          3026 => x"b5d408e8",
          3027 => x"05337098",
          3028 => x"2b537298",
          3029 => x"2c5382b5",
          3030 => x"d408fc05",
          3031 => x"085253a2",
          3032 => x"d83f82b5",
          3033 => x"c8085372",
          3034 => x"82b5d408",
          3035 => x"f4052399",
          3036 => x"3982b5d4",
          3037 => x"08fc0508",
          3038 => x"519d8a3f",
          3039 => x"82b5c808",
          3040 => x"537282b5",
          3041 => x"d408f405",
          3042 => x"2382b5d4",
          3043 => x"08ec0522",
          3044 => x"5382b5d4",
          3045 => x"08f40522",
          3046 => x"73713154",
          3047 => x"547282b5",
          3048 => x"d408ec05",
          3049 => x"238bd839",
          3050 => x"82b5d408",
          3051 => x"90050882",
          3052 => x"b5d40890",
          3053 => x"05088405",
          3054 => x"82b5d408",
          3055 => x"90050c70",
          3056 => x"0882b5d4",
          3057 => x"08fc050c",
          3058 => x"82b5d408",
          3059 => x"e4052270",
          3060 => x"832a7081",
          3061 => x"06515151",
          3062 => x"5372802e",
          3063 => x"ab3882b5",
          3064 => x"d408e805",
          3065 => x"3370982b",
          3066 => x"5372982c",
          3067 => x"5382b5d4",
          3068 => x"08fc0508",
          3069 => x"5253a1c1",
          3070 => x"3f82b5c8",
          3071 => x"08537282",
          3072 => x"b5d408f4",
          3073 => x"05239939",
          3074 => x"82b5d408",
          3075 => x"fc050851",
          3076 => x"9bf33f82",
          3077 => x"b5c80853",
          3078 => x"7282b5d4",
          3079 => x"08f40523",
          3080 => x"82b5d408",
          3081 => x"ec052253",
          3082 => x"82b5d408",
          3083 => x"f4052273",
          3084 => x"71315454",
          3085 => x"7282b5d4",
          3086 => x"08ec0523",
          3087 => x"8ac13982",
          3088 => x"b5d408e4",
          3089 => x"05227082",
          3090 => x"2a708106",
          3091 => x"51515372",
          3092 => x"802ea438",
          3093 => x"82b5d408",
          3094 => x"90050882",
          3095 => x"b5d40890",
          3096 => x"05088405",
          3097 => x"82b5d408",
          3098 => x"90050c70",
          3099 => x"0882b5d4",
          3100 => x"08dc050c",
          3101 => x"53a23982",
          3102 => x"b5d40890",
          3103 => x"050882b5",
          3104 => x"d4089005",
          3105 => x"08840582",
          3106 => x"b5d40890",
          3107 => x"050c7008",
          3108 => x"82b5d408",
          3109 => x"dc050c53",
          3110 => x"82b5d408",
          3111 => x"dc050882",
          3112 => x"b5d408fc",
          3113 => x"050c82b5",
          3114 => x"d408fc05",
          3115 => x"088025a4",
          3116 => x"3882b5d4",
          3117 => x"08e40522",
          3118 => x"70820751",
          3119 => x"537282b5",
          3120 => x"d408e405",
          3121 => x"2382b5d4",
          3122 => x"08fc0508",
          3123 => x"3082b5d4",
          3124 => x"08fc050c",
          3125 => x"82b5d408",
          3126 => x"e4052270",
          3127 => x"ffbf0651",
          3128 => x"537282b5",
          3129 => x"d408e405",
          3130 => x"2381af39",
          3131 => x"880b82b5",
          3132 => x"d408f405",
          3133 => x"23a93982",
          3134 => x"b5d408e4",
          3135 => x"05227080",
          3136 => x"c0075153",
          3137 => x"7282b5d4",
          3138 => x"08e40523",
          3139 => x"80f80b82",
          3140 => x"b5d408f8",
          3141 => x"0534900b",
          3142 => x"82b5d408",
          3143 => x"f4052382",
          3144 => x"b5d408e4",
          3145 => x"05227082",
          3146 => x"2a708106",
          3147 => x"51515372",
          3148 => x"802ea438",
          3149 => x"82b5d408",
          3150 => x"90050882",
          3151 => x"b5d40890",
          3152 => x"05088405",
          3153 => x"82b5d408",
          3154 => x"90050c70",
          3155 => x"0882b5d4",
          3156 => x"08d8050c",
          3157 => x"53a23982",
          3158 => x"b5d40890",
          3159 => x"050882b5",
          3160 => x"d4089005",
          3161 => x"08840582",
          3162 => x"b5d40890",
          3163 => x"050c7008",
          3164 => x"82b5d408",
          3165 => x"d8050c53",
          3166 => x"82b5d408",
          3167 => x"d8050882",
          3168 => x"b5d408fc",
          3169 => x"050c82b5",
          3170 => x"d408e405",
          3171 => x"2270cf06",
          3172 => x"51537282",
          3173 => x"b5d408e4",
          3174 => x"052382b5",
          3175 => x"d80b82b5",
          3176 => x"d408f005",
          3177 => x"0c82b5d4",
          3178 => x"08f00508",
          3179 => x"82b5d408",
          3180 => x"f4052282",
          3181 => x"b5d408fc",
          3182 => x"05087155",
          3183 => x"70545654",
          3184 => x"55a3f33f",
          3185 => x"82b5c808",
          3186 => x"53727534",
          3187 => x"82b5d408",
          3188 => x"f0050882",
          3189 => x"b5d408d4",
          3190 => x"050c82b5",
          3191 => x"d408f005",
          3192 => x"08703351",
          3193 => x"53897327",
          3194 => x"a43882b5",
          3195 => x"d408f005",
          3196 => x"08537233",
          3197 => x"5482b5d4",
          3198 => x"08f80533",
          3199 => x"7015df11",
          3200 => x"51515372",
          3201 => x"82b5d408",
          3202 => x"d0053497",
          3203 => x"3982b5d4",
          3204 => x"08f00508",
          3205 => x"537233b0",
          3206 => x"11515372",
          3207 => x"82b5d408",
          3208 => x"d0053482",
          3209 => x"b5d408d4",
          3210 => x"05085382",
          3211 => x"b5d408d0",
          3212 => x"05337334",
          3213 => x"82b5d408",
          3214 => x"f0050881",
          3215 => x"0582b5d4",
          3216 => x"08f0050c",
          3217 => x"82b5d408",
          3218 => x"f4052270",
          3219 => x"5382b5d4",
          3220 => x"08fc0508",
          3221 => x"5253a2ab",
          3222 => x"3f82b5c8",
          3223 => x"087082b5",
          3224 => x"d408fc05",
          3225 => x"0c5382b5",
          3226 => x"d408fc05",
          3227 => x"08802e84",
          3228 => x"38feb239",
          3229 => x"82b5d408",
          3230 => x"f0050882",
          3231 => x"b5d85455",
          3232 => x"72547470",
          3233 => x"75315153",
          3234 => x"7282b5d4",
          3235 => x"08fc0534",
          3236 => x"82b5d408",
          3237 => x"e4052270",
          3238 => x"b2065153",
          3239 => x"72802e94",
          3240 => x"3882b5d4",
          3241 => x"08ec0522",
          3242 => x"ff115153",
          3243 => x"7282b5d4",
          3244 => x"08ec0523",
          3245 => x"82b5d408",
          3246 => x"e4052270",
          3247 => x"862a7081",
          3248 => x"06515153",
          3249 => x"72802e80",
          3250 => x"e73882b5",
          3251 => x"d408ec05",
          3252 => x"2270902b",
          3253 => x"82b5d408",
          3254 => x"cc050c82",
          3255 => x"b5d408cc",
          3256 => x"0508902c",
          3257 => x"82b5d408",
          3258 => x"cc050c82",
          3259 => x"b5d408f4",
          3260 => x"05225153",
          3261 => x"72902e09",
          3262 => x"81069538",
          3263 => x"82b5d408",
          3264 => x"cc0508fe",
          3265 => x"05537282",
          3266 => x"b5d408c8",
          3267 => x"05239339",
          3268 => x"82b5d408",
          3269 => x"cc0508ff",
          3270 => x"05537282",
          3271 => x"b5d408c8",
          3272 => x"052382b5",
          3273 => x"d408c805",
          3274 => x"2282b5d4",
          3275 => x"08ec0523",
          3276 => x"82b5d408",
          3277 => x"e4052270",
          3278 => x"832a7081",
          3279 => x"06515153",
          3280 => x"72802e80",
          3281 => x"d03882b5",
          3282 => x"d408e805",
          3283 => x"3370982b",
          3284 => x"70982c82",
          3285 => x"b5d408fc",
          3286 => x"05335751",
          3287 => x"51537274",
          3288 => x"24973882",
          3289 => x"b5d408e4",
          3290 => x"052270f7",
          3291 => x"06515372",
          3292 => x"82b5d408",
          3293 => x"e405239d",
          3294 => x"3982b5d4",
          3295 => x"08e80533",
          3296 => x"5382b5d4",
          3297 => x"08fc0533",
          3298 => x"73713154",
          3299 => x"547282b5",
          3300 => x"d408e805",
          3301 => x"3482b5d4",
          3302 => x"08e40522",
          3303 => x"70832a70",
          3304 => x"81065151",
          3305 => x"5372802e",
          3306 => x"b13882b5",
          3307 => x"d408e805",
          3308 => x"3370882b",
          3309 => x"70902b70",
          3310 => x"902c7088",
          3311 => x"2c515151",
          3312 => x"51537254",
          3313 => x"82b5d408",
          3314 => x"ec052270",
          3315 => x"75315153",
          3316 => x"7282b5d4",
          3317 => x"08ec0523",
          3318 => x"af3982b5",
          3319 => x"d408fc05",
          3320 => x"3370882b",
          3321 => x"70902b70",
          3322 => x"902c7088",
          3323 => x"2c515151",
          3324 => x"51537254",
          3325 => x"82b5d408",
          3326 => x"ec052270",
          3327 => x"75315153",
          3328 => x"7282b5d4",
          3329 => x"08ec0523",
          3330 => x"82b5d408",
          3331 => x"e4052270",
          3332 => x"83800651",
          3333 => x"5372b038",
          3334 => x"82b5d408",
          3335 => x"ec0522ff",
          3336 => x"11545472",
          3337 => x"82b5d408",
          3338 => x"ec052373",
          3339 => x"902b7090",
          3340 => x"2c515380",
          3341 => x"73259038",
          3342 => x"82b5d408",
          3343 => x"88050852",
          3344 => x"a0518aee",
          3345 => x"3fd23982",
          3346 => x"b5d408e4",
          3347 => x"05227081",
          3348 => x"2a708106",
          3349 => x"51515372",
          3350 => x"802e9138",
          3351 => x"82b5d408",
          3352 => x"88050852",
          3353 => x"ad518aca",
          3354 => x"3f80c739",
          3355 => x"82b5d408",
          3356 => x"e4052270",
          3357 => x"842a7081",
          3358 => x"06515153",
          3359 => x"72802e90",
          3360 => x"3882b5d4",
          3361 => x"08880508",
          3362 => x"52ab518a",
          3363 => x"a53fa339",
          3364 => x"82b5d408",
          3365 => x"e4052270",
          3366 => x"852a7081",
          3367 => x"06515153",
          3368 => x"72802e8e",
          3369 => x"3882b5d4",
          3370 => x"08880508",
          3371 => x"52a0518a",
          3372 => x"813f82b5",
          3373 => x"d408e405",
          3374 => x"2270862a",
          3375 => x"70810651",
          3376 => x"51537280",
          3377 => x"2eb13882",
          3378 => x"b5d40888",
          3379 => x"050852b0",
          3380 => x"5189df3f",
          3381 => x"82b5d408",
          3382 => x"f4052253",
          3383 => x"72902e09",
          3384 => x"81069438",
          3385 => x"82b5d408",
          3386 => x"88050852",
          3387 => x"82b5d408",
          3388 => x"f8053351",
          3389 => x"89bc3f82",
          3390 => x"b5d408e4",
          3391 => x"05227088",
          3392 => x"2a708106",
          3393 => x"51515372",
          3394 => x"802eb038",
          3395 => x"82b5d408",
          3396 => x"ec0522ff",
          3397 => x"11545472",
          3398 => x"82b5d408",
          3399 => x"ec052373",
          3400 => x"902b7090",
          3401 => x"2c515380",
          3402 => x"73259038",
          3403 => x"82b5d408",
          3404 => x"88050852",
          3405 => x"b05188fa",
          3406 => x"3fd23982",
          3407 => x"b5d408e4",
          3408 => x"05227083",
          3409 => x"2a708106",
          3410 => x"51515372",
          3411 => x"802eb038",
          3412 => x"82b5d408",
          3413 => x"e80533ff",
          3414 => x"11545472",
          3415 => x"82b5d408",
          3416 => x"e8053473",
          3417 => x"982b7098",
          3418 => x"2c515380",
          3419 => x"73259038",
          3420 => x"82b5d408",
          3421 => x"88050852",
          3422 => x"b05188b6",
          3423 => x"3fd23982",
          3424 => x"b5d408e4",
          3425 => x"05227087",
          3426 => x"2a708106",
          3427 => x"51515372",
          3428 => x"b03882b5",
          3429 => x"d408ec05",
          3430 => x"22ff1154",
          3431 => x"547282b5",
          3432 => x"d408ec05",
          3433 => x"2373902b",
          3434 => x"70902c51",
          3435 => x"53807325",
          3436 => x"903882b5",
          3437 => x"d4088805",
          3438 => x"0852a051",
          3439 => x"87f43fd2",
          3440 => x"3982b5d4",
          3441 => x"08f80533",
          3442 => x"537280e3",
          3443 => x"2e098106",
          3444 => x"973882b5",
          3445 => x"d4088805",
          3446 => x"085282b5",
          3447 => x"d408fc05",
          3448 => x"335187ce",
          3449 => x"3f81ee39",
          3450 => x"82b5d408",
          3451 => x"f8053353",
          3452 => x"7280f32e",
          3453 => x"09810680",
          3454 => x"cb3882b5",
          3455 => x"d408f405",
          3456 => x"22ff1151",
          3457 => x"537282b5",
          3458 => x"d408f405",
          3459 => x"237283ff",
          3460 => x"ff065372",
          3461 => x"83ffff2e",
          3462 => x"81bb3882",
          3463 => x"b5d40888",
          3464 => x"05085282",
          3465 => x"b5d408fc",
          3466 => x"05087033",
          3467 => x"5282b5d4",
          3468 => x"08fc0508",
          3469 => x"810582b5",
          3470 => x"d408fc05",
          3471 => x"0c5386f2",
          3472 => x"3fffb739",
          3473 => x"82b5d408",
          3474 => x"f8053353",
          3475 => x"7280d32e",
          3476 => x"09810680",
          3477 => x"cb3882b5",
          3478 => x"d408f405",
          3479 => x"22ff1151",
          3480 => x"537282b5",
          3481 => x"d408f405",
          3482 => x"237283ff",
          3483 => x"ff065372",
          3484 => x"83ffff2e",
          3485 => x"80df3882",
          3486 => x"b5d40888",
          3487 => x"05085282",
          3488 => x"b5d408fc",
          3489 => x"05087033",
          3490 => x"525386a6",
          3491 => x"3f82b5d4",
          3492 => x"08fc0508",
          3493 => x"810582b5",
          3494 => x"d408fc05",
          3495 => x"0cffb739",
          3496 => x"82b5d408",
          3497 => x"f0050882",
          3498 => x"b5d82ea9",
          3499 => x"3882b5d4",
          3500 => x"08880508",
          3501 => x"5282b5d4",
          3502 => x"08f00508",
          3503 => x"ff0582b5",
          3504 => x"d408f005",
          3505 => x"0c82b5d4",
          3506 => x"08f00508",
          3507 => x"70335253",
          3508 => x"85e03fcc",
          3509 => x"3982b5d4",
          3510 => x"08e40522",
          3511 => x"70872a70",
          3512 => x"81065151",
          3513 => x"5372802e",
          3514 => x"80c33882",
          3515 => x"b5d408ec",
          3516 => x"0522ff11",
          3517 => x"54547282",
          3518 => x"b5d408ec",
          3519 => x"05237390",
          3520 => x"2b70902c",
          3521 => x"51538073",
          3522 => x"25a33882",
          3523 => x"b5d40888",
          3524 => x"050852a0",
          3525 => x"51859b3f",
          3526 => x"d23982b5",
          3527 => x"d4088805",
          3528 => x"085282b5",
          3529 => x"d408f805",
          3530 => x"33518586",
          3531 => x"3f800b82",
          3532 => x"b5d408e4",
          3533 => x"0523eab7",
          3534 => x"3982b5d4",
          3535 => x"08f80533",
          3536 => x"5372a52e",
          3537 => x"098106a8",
          3538 => x"38810b82",
          3539 => x"b5d408e4",
          3540 => x"0523800b",
          3541 => x"82b5d408",
          3542 => x"ec052380",
          3543 => x"0b82b5d4",
          3544 => x"08e80534",
          3545 => x"8a0b82b5",
          3546 => x"d408f405",
          3547 => x"23ea8039",
          3548 => x"82b5d408",
          3549 => x"88050852",
          3550 => x"82b5d408",
          3551 => x"f8053351",
          3552 => x"84b03fe9",
          3553 => x"ea3982b5",
          3554 => x"d4088805",
          3555 => x"088c1108",
          3556 => x"7082b5d4",
          3557 => x"08e0050c",
          3558 => x"515382b5",
          3559 => x"d408e005",
          3560 => x"0882b5c8",
          3561 => x"0c953d0d",
          3562 => x"82b5d40c",
          3563 => x"0482b5d4",
          3564 => x"080282b5",
          3565 => x"d40cfd3d",
          3566 => x"0d82cd98",
          3567 => x"085382b5",
          3568 => x"d4088c05",
          3569 => x"085282b5",
          3570 => x"d4088805",
          3571 => x"0851e4dd",
          3572 => x"3f82b5c8",
          3573 => x"087082b5",
          3574 => x"c80c5485",
          3575 => x"3d0d82b5",
          3576 => x"d40c0482",
          3577 => x"b5d40802",
          3578 => x"82b5d40c",
          3579 => x"fb3d0d80",
          3580 => x"0b82b5d4",
          3581 => x"08f8050c",
          3582 => x"82cd9c08",
          3583 => x"85113370",
          3584 => x"812a7081",
          3585 => x"32708106",
          3586 => x"51515151",
          3587 => x"5372802e",
          3588 => x"8d38ff0b",
          3589 => x"82b5d408",
          3590 => x"f4050c81",
          3591 => x"923982b5",
          3592 => x"d4088805",
          3593 => x"08537233",
          3594 => x"82b5d408",
          3595 => x"88050881",
          3596 => x"0582b5d4",
          3597 => x"0888050c",
          3598 => x"537282b5",
          3599 => x"d408fc05",
          3600 => x"347281ff",
          3601 => x"06537280",
          3602 => x"2eb03882",
          3603 => x"cd9c0882",
          3604 => x"cd9c0853",
          3605 => x"82b5d408",
          3606 => x"fc053352",
          3607 => x"90110851",
          3608 => x"53722d82",
          3609 => x"b5c80853",
          3610 => x"72802eff",
          3611 => x"b138ff0b",
          3612 => x"82b5d408",
          3613 => x"f8050cff",
          3614 => x"a53982cd",
          3615 => x"9c0882cd",
          3616 => x"9c085353",
          3617 => x"8a519013",
          3618 => x"0853722d",
          3619 => x"82b5c808",
          3620 => x"5372802e",
          3621 => x"8a38ff0b",
          3622 => x"82b5d408",
          3623 => x"f8050c82",
          3624 => x"b5d408f8",
          3625 => x"05087082",
          3626 => x"b5d408f4",
          3627 => x"050c5382",
          3628 => x"b5d408f4",
          3629 => x"050882b5",
          3630 => x"c80c873d",
          3631 => x"0d82b5d4",
          3632 => x"0c0482b5",
          3633 => x"d4080282",
          3634 => x"b5d40cfb",
          3635 => x"3d0d800b",
          3636 => x"82b5d408",
          3637 => x"f8050c82",
          3638 => x"b5d4088c",
          3639 => x"05088511",
          3640 => x"3370812a",
          3641 => x"70813270",
          3642 => x"81065151",
          3643 => x"51515372",
          3644 => x"802e8d38",
          3645 => x"ff0b82b5",
          3646 => x"d408f405",
          3647 => x"0c80f339",
          3648 => x"82b5d408",
          3649 => x"88050853",
          3650 => x"723382b5",
          3651 => x"d4088805",
          3652 => x"08810582",
          3653 => x"b5d40888",
          3654 => x"050c5372",
          3655 => x"82b5d408",
          3656 => x"fc053472",
          3657 => x"81ff0653",
          3658 => x"72802eb6",
          3659 => x"3882b5d4",
          3660 => x"088c0508",
          3661 => x"82b5d408",
          3662 => x"8c050853",
          3663 => x"82b5d408",
          3664 => x"fc053352",
          3665 => x"90110851",
          3666 => x"53722d82",
          3667 => x"b5c80853",
          3668 => x"72802eff",
          3669 => x"ab38ff0b",
          3670 => x"82b5d408",
          3671 => x"f8050cff",
          3672 => x"9f3982b5",
          3673 => x"d408f805",
          3674 => x"087082b5",
          3675 => x"d408f405",
          3676 => x"0c5382b5",
          3677 => x"d408f405",
          3678 => x"0882b5c8",
          3679 => x"0c873d0d",
          3680 => x"82b5d40c",
          3681 => x"0482b5d4",
          3682 => x"080282b5",
          3683 => x"d40cfe3d",
          3684 => x"0d82cd9c",
          3685 => x"085282b5",
          3686 => x"d4088805",
          3687 => x"0851933f",
          3688 => x"82b5c808",
          3689 => x"7082b5c8",
          3690 => x"0c53843d",
          3691 => x"0d82b5d4",
          3692 => x"0c0482b5",
          3693 => x"d4080282",
          3694 => x"b5d40cfb",
          3695 => x"3d0d82b5",
          3696 => x"d4088c05",
          3697 => x"08851133",
          3698 => x"70812a70",
          3699 => x"81327081",
          3700 => x"06515151",
          3701 => x"51537280",
          3702 => x"2e8d38ff",
          3703 => x"0b82b5d4",
          3704 => x"08fc050c",
          3705 => x"81cb3982",
          3706 => x"b5d4088c",
          3707 => x"05088511",
          3708 => x"3370822a",
          3709 => x"70810651",
          3710 => x"51515372",
          3711 => x"802e80db",
          3712 => x"3882b5d4",
          3713 => x"088c0508",
          3714 => x"82b5d408",
          3715 => x"8c050854",
          3716 => x"548c1408",
          3717 => x"88140825",
          3718 => x"9f3882b5",
          3719 => x"d4088c05",
          3720 => x"08700870",
          3721 => x"82b5d408",
          3722 => x"88050852",
          3723 => x"57545472",
          3724 => x"75347308",
          3725 => x"8105740c",
          3726 => x"82b5d408",
          3727 => x"8c05088c",
          3728 => x"11088105",
          3729 => x"8c120c82",
          3730 => x"b5d40888",
          3731 => x"05087082",
          3732 => x"b5d408fc",
          3733 => x"050c5153",
          3734 => x"80d73982",
          3735 => x"b5d4088c",
          3736 => x"050882b5",
          3737 => x"d4088c05",
          3738 => x"085382b5",
          3739 => x"d4088805",
          3740 => x"087081ff",
          3741 => x"06539012",
          3742 => x"08515454",
          3743 => x"722d82b5",
          3744 => x"c8085372",
          3745 => x"a33882b5",
          3746 => x"d4088c05",
          3747 => x"088c1108",
          3748 => x"81058c12",
          3749 => x"0c82b5d4",
          3750 => x"08880508",
          3751 => x"7082b5d4",
          3752 => x"08fc050c",
          3753 => x"51538a39",
          3754 => x"ff0b82b5",
          3755 => x"d408fc05",
          3756 => x"0c82b5d4",
          3757 => x"08fc0508",
          3758 => x"82b5c80c",
          3759 => x"873d0d82",
          3760 => x"b5d40c04",
          3761 => x"82b5d408",
          3762 => x"0282b5d4",
          3763 => x"0cf93d0d",
          3764 => x"82b5d408",
          3765 => x"88050885",
          3766 => x"11337081",
          3767 => x"32708106",
          3768 => x"51515152",
          3769 => x"71802e8d",
          3770 => x"38ff0b82",
          3771 => x"b5d408f8",
          3772 => x"050c8394",
          3773 => x"3982b5d4",
          3774 => x"08880508",
          3775 => x"85113370",
          3776 => x"862a7081",
          3777 => x"06515151",
          3778 => x"5271802e",
          3779 => x"80c53882",
          3780 => x"b5d40888",
          3781 => x"050882b5",
          3782 => x"d4088805",
          3783 => x"08535385",
          3784 => x"123370ff",
          3785 => x"bf065152",
          3786 => x"71851434",
          3787 => x"82b5d408",
          3788 => x"8805088c",
          3789 => x"11088105",
          3790 => x"8c120c82",
          3791 => x"b5d40888",
          3792 => x"05088411",
          3793 => x"337082b5",
          3794 => x"d408f805",
          3795 => x"0c515152",
          3796 => x"82b63982",
          3797 => x"b5d40888",
          3798 => x"05088511",
          3799 => x"3370822a",
          3800 => x"70810651",
          3801 => x"51515271",
          3802 => x"802e80d7",
          3803 => x"3882b5d4",
          3804 => x"08880508",
          3805 => x"70087033",
          3806 => x"82b5d408",
          3807 => x"fc050c51",
          3808 => x"5282b5d4",
          3809 => x"08fc0508",
          3810 => x"a93882b5",
          3811 => x"d4088805",
          3812 => x"0882b5d4",
          3813 => x"08880508",
          3814 => x"53538512",
          3815 => x"3370a007",
          3816 => x"51527185",
          3817 => x"1434ff0b",
          3818 => x"82b5d408",
          3819 => x"f8050c81",
          3820 => x"d73982b5",
          3821 => x"d4088805",
          3822 => x"08700881",
          3823 => x"05710c52",
          3824 => x"81a13982",
          3825 => x"b5d40888",
          3826 => x"050882b5",
          3827 => x"d4088805",
          3828 => x"08529411",
          3829 => x"08515271",
          3830 => x"2d82b5c8",
          3831 => x"087082b5",
          3832 => x"d408fc05",
          3833 => x"0c5282b5",
          3834 => x"d408fc05",
          3835 => x"08802580",
          3836 => x"f23882b5",
          3837 => x"d4088805",
          3838 => x"0882b5d4",
          3839 => x"08f4050c",
          3840 => x"82b5d408",
          3841 => x"88050885",
          3842 => x"113382b5",
          3843 => x"d408f005",
          3844 => x"0c5282b5",
          3845 => x"d408fc05",
          3846 => x"08ff2e09",
          3847 => x"81069538",
          3848 => x"82b5d408",
          3849 => x"f0050890",
          3850 => x"07527182",
          3851 => x"b5d408ec",
          3852 => x"05349339",
          3853 => x"82b5d408",
          3854 => x"f00508a0",
          3855 => x"07527182",
          3856 => x"b5d408ec",
          3857 => x"053482b5",
          3858 => x"d408f405",
          3859 => x"085282b5",
          3860 => x"d408ec05",
          3861 => x"33851334",
          3862 => x"ff0b82b5",
          3863 => x"d408f805",
          3864 => x"0ca63982",
          3865 => x"b5d40888",
          3866 => x"05088c11",
          3867 => x"0881058c",
          3868 => x"120c82b5",
          3869 => x"d408fc05",
          3870 => x"087081ff",
          3871 => x"067082b5",
          3872 => x"d408f805",
          3873 => x"0c515152",
          3874 => x"82b5d408",
          3875 => x"f8050882",
          3876 => x"b5c80c89",
          3877 => x"3d0d82b5",
          3878 => x"d40c0482",
          3879 => x"b5d40802",
          3880 => x"82b5d40c",
          3881 => x"fd3d0d82",
          3882 => x"b5d40888",
          3883 => x"050882b5",
          3884 => x"d408fc05",
          3885 => x"0c82b5d4",
          3886 => x"088c0508",
          3887 => x"82b5d408",
          3888 => x"f8050c82",
          3889 => x"b5d40890",
          3890 => x"0508802e",
          3891 => x"82a23882",
          3892 => x"b5d408f8",
          3893 => x"050882b5",
          3894 => x"d408fc05",
          3895 => x"082681ac",
          3896 => x"3882b5d4",
          3897 => x"08f80508",
          3898 => x"82b5d408",
          3899 => x"90050805",
          3900 => x"5182b5d4",
          3901 => x"08fc0508",
          3902 => x"71278190",
          3903 => x"3882b5d4",
          3904 => x"08fc0508",
          3905 => x"82b5d408",
          3906 => x"90050805",
          3907 => x"82b5d408",
          3908 => x"fc050c82",
          3909 => x"b5d408f8",
          3910 => x"050882b5",
          3911 => x"d4089005",
          3912 => x"080582b5",
          3913 => x"d408f805",
          3914 => x"0c82b5d4",
          3915 => x"08900508",
          3916 => x"810582b5",
          3917 => x"d4089005",
          3918 => x"0c82b5d4",
          3919 => x"08900508",
          3920 => x"ff0582b5",
          3921 => x"d4089005",
          3922 => x"0c82b5d4",
          3923 => x"08900508",
          3924 => x"802e819c",
          3925 => x"3882b5d4",
          3926 => x"08fc0508",
          3927 => x"ff0582b5",
          3928 => x"d408fc05",
          3929 => x"0c82b5d4",
          3930 => x"08f80508",
          3931 => x"ff0582b5",
          3932 => x"d408f805",
          3933 => x"0c82b5d4",
          3934 => x"08fc0508",
          3935 => x"82b5d408",
          3936 => x"f8050853",
          3937 => x"51713371",
          3938 => x"34ffae39",
          3939 => x"82b5d408",
          3940 => x"90050881",
          3941 => x"0582b5d4",
          3942 => x"0890050c",
          3943 => x"82b5d408",
          3944 => x"900508ff",
          3945 => x"0582b5d4",
          3946 => x"0890050c",
          3947 => x"82b5d408",
          3948 => x"90050880",
          3949 => x"2eba3882",
          3950 => x"b5d408f8",
          3951 => x"05085170",
          3952 => x"3382b5d4",
          3953 => x"08f80508",
          3954 => x"810582b5",
          3955 => x"d408f805",
          3956 => x"0c82b5d4",
          3957 => x"08fc0508",
          3958 => x"52527171",
          3959 => x"3482b5d4",
          3960 => x"08fc0508",
          3961 => x"810582b5",
          3962 => x"d408fc05",
          3963 => x"0cffad39",
          3964 => x"82b5d408",
          3965 => x"88050870",
          3966 => x"82b5c80c",
          3967 => x"51853d0d",
          3968 => x"82b5d40c",
          3969 => x"0482b5d4",
          3970 => x"080282b5",
          3971 => x"d40cfe3d",
          3972 => x"0d82b5d4",
          3973 => x"08880508",
          3974 => x"82b5d408",
          3975 => x"fc050c82",
          3976 => x"b5d408fc",
          3977 => x"05085271",
          3978 => x"3382b5d4",
          3979 => x"08fc0508",
          3980 => x"810582b5",
          3981 => x"d408fc05",
          3982 => x"0c7081ff",
          3983 => x"06515170",
          3984 => x"802e8338",
          3985 => x"da3982b5",
          3986 => x"d408fc05",
          3987 => x"08ff0582",
          3988 => x"b5d408fc",
          3989 => x"050c82b5",
          3990 => x"d408fc05",
          3991 => x"0882b5d4",
          3992 => x"08880508",
          3993 => x"317082b5",
          3994 => x"c80c5184",
          3995 => x"3d0d82b5",
          3996 => x"d40c0482",
          3997 => x"b5d40802",
          3998 => x"82b5d40c",
          3999 => x"fe3d0d82",
          4000 => x"b5d40888",
          4001 => x"050882b5",
          4002 => x"d408fc05",
          4003 => x"0c82b5d4",
          4004 => x"088c0508",
          4005 => x"52713382",
          4006 => x"b5d4088c",
          4007 => x"05088105",
          4008 => x"82b5d408",
          4009 => x"8c050c82",
          4010 => x"b5d408fc",
          4011 => x"05085351",
          4012 => x"70723482",
          4013 => x"b5d408fc",
          4014 => x"05088105",
          4015 => x"82b5d408",
          4016 => x"fc050c70",
          4017 => x"81ff0651",
          4018 => x"70802e84",
          4019 => x"38ffbe39",
          4020 => x"82b5d408",
          4021 => x"88050870",
          4022 => x"82b5c80c",
          4023 => x"51843d0d",
          4024 => x"82b5d40c",
          4025 => x"0482b5d4",
          4026 => x"080282b5",
          4027 => x"d40cfd3d",
          4028 => x"0d82b5d4",
          4029 => x"08880508",
          4030 => x"82b5d408",
          4031 => x"fc050c82",
          4032 => x"b5d4088c",
          4033 => x"050882b5",
          4034 => x"d408f805",
          4035 => x"0c82b5d4",
          4036 => x"08900508",
          4037 => x"802e80e5",
          4038 => x"3882b5d4",
          4039 => x"08900508",
          4040 => x"810582b5",
          4041 => x"d4089005",
          4042 => x"0c82b5d4",
          4043 => x"08900508",
          4044 => x"ff0582b5",
          4045 => x"d4089005",
          4046 => x"0c82b5d4",
          4047 => x"08900508",
          4048 => x"802eba38",
          4049 => x"82b5d408",
          4050 => x"f8050851",
          4051 => x"703382b5",
          4052 => x"d408f805",
          4053 => x"08810582",
          4054 => x"b5d408f8",
          4055 => x"050c82b5",
          4056 => x"d408fc05",
          4057 => x"08525271",
          4058 => x"713482b5",
          4059 => x"d408fc05",
          4060 => x"08810582",
          4061 => x"b5d408fc",
          4062 => x"050cffad",
          4063 => x"3982b5d4",
          4064 => x"08880508",
          4065 => x"7082b5c8",
          4066 => x"0c51853d",
          4067 => x"0d82b5d4",
          4068 => x"0c0482b5",
          4069 => x"d4080282",
          4070 => x"b5d40cfd",
          4071 => x"3d0d82b5",
          4072 => x"d4089005",
          4073 => x"08802e81",
          4074 => x"f43882b5",
          4075 => x"d4088c05",
          4076 => x"08527133",
          4077 => x"82b5d408",
          4078 => x"8c050881",
          4079 => x"0582b5d4",
          4080 => x"088c050c",
          4081 => x"82b5d408",
          4082 => x"88050870",
          4083 => x"337281ff",
          4084 => x"06535454",
          4085 => x"5171712e",
          4086 => x"843880ce",
          4087 => x"3982b5d4",
          4088 => x"08880508",
          4089 => x"52713382",
          4090 => x"b5d40888",
          4091 => x"05088105",
          4092 => x"82b5d408",
          4093 => x"88050c70",
          4094 => x"81ff0651",
          4095 => x"51708d38",
          4096 => x"800b82b5",
          4097 => x"d408fc05",
          4098 => x"0c819b39",
          4099 => x"82b5d408",
          4100 => x"900508ff",
          4101 => x"0582b5d4",
          4102 => x"0890050c",
          4103 => x"82b5d408",
          4104 => x"90050880",
          4105 => x"2e8438ff",
          4106 => x"813982b5",
          4107 => x"d4089005",
          4108 => x"08802e80",
          4109 => x"e83882b5",
          4110 => x"d4088805",
          4111 => x"08703352",
          4112 => x"53708d38",
          4113 => x"ff0b82b5",
          4114 => x"d408fc05",
          4115 => x"0c80d739",
          4116 => x"82b5d408",
          4117 => x"8c0508ff",
          4118 => x"0582b5d4",
          4119 => x"088c050c",
          4120 => x"82b5d408",
          4121 => x"8c050870",
          4122 => x"33525270",
          4123 => x"8c38810b",
          4124 => x"82b5d408",
          4125 => x"fc050cae",
          4126 => x"3982b5d4",
          4127 => x"08880508",
          4128 => x"703382b5",
          4129 => x"d4088c05",
          4130 => x"08703372",
          4131 => x"71317082",
          4132 => x"b5d408fc",
          4133 => x"050c5355",
          4134 => x"5252538a",
          4135 => x"39800b82",
          4136 => x"b5d408fc",
          4137 => x"050c82b5",
          4138 => x"d408fc05",
          4139 => x"0882b5c8",
          4140 => x"0c853d0d",
          4141 => x"82b5d40c",
          4142 => x"0482b5d4",
          4143 => x"080282b5",
          4144 => x"d40cfd3d",
          4145 => x"0d82b5d4",
          4146 => x"08880508",
          4147 => x"82b5d408",
          4148 => x"f8050c82",
          4149 => x"b5d4088c",
          4150 => x"05088d38",
          4151 => x"800b82b5",
          4152 => x"d408fc05",
          4153 => x"0c80ec39",
          4154 => x"82b5d408",
          4155 => x"f8050852",
          4156 => x"713382b5",
          4157 => x"d408f805",
          4158 => x"08810582",
          4159 => x"b5d408f8",
          4160 => x"050c7081",
          4161 => x"ff065151",
          4162 => x"70802e9f",
          4163 => x"3882b5d4",
          4164 => x"088c0508",
          4165 => x"ff0582b5",
          4166 => x"d4088c05",
          4167 => x"0c82b5d4",
          4168 => x"088c0508",
          4169 => x"ff2e8438",
          4170 => x"ffbe3982",
          4171 => x"b5d408f8",
          4172 => x"0508ff05",
          4173 => x"82b5d408",
          4174 => x"f8050c82",
          4175 => x"b5d408f8",
          4176 => x"050882b5",
          4177 => x"d4088805",
          4178 => x"08317082",
          4179 => x"b5d408fc",
          4180 => x"050c5182",
          4181 => x"b5d408fc",
          4182 => x"050882b5",
          4183 => x"c80c853d",
          4184 => x"0d82b5d4",
          4185 => x"0c0482b5",
          4186 => x"d4080282",
          4187 => x"b5d40cfe",
          4188 => x"3d0d82b5",
          4189 => x"d4088805",
          4190 => x"0882b5d4",
          4191 => x"08fc050c",
          4192 => x"82b5d408",
          4193 => x"90050880",
          4194 => x"2e80d438",
          4195 => x"82b5d408",
          4196 => x"90050881",
          4197 => x"0582b5d4",
          4198 => x"0890050c",
          4199 => x"82b5d408",
          4200 => x"900508ff",
          4201 => x"0582b5d4",
          4202 => x"0890050c",
          4203 => x"82b5d408",
          4204 => x"90050880",
          4205 => x"2ea93882",
          4206 => x"b5d4088c",
          4207 => x"05085170",
          4208 => x"82b5d408",
          4209 => x"fc050852",
          4210 => x"52717134",
          4211 => x"82b5d408",
          4212 => x"fc050881",
          4213 => x"0582b5d4",
          4214 => x"08fc050c",
          4215 => x"ffbe3982",
          4216 => x"b5d40888",
          4217 => x"05087082",
          4218 => x"b5c80c51",
          4219 => x"843d0d82",
          4220 => x"b5d40c04",
          4221 => x"82b5d408",
          4222 => x"0282b5d4",
          4223 => x"0cf93d0d",
          4224 => x"800b82b5",
          4225 => x"d408fc05",
          4226 => x"0c82b5d4",
          4227 => x"08880508",
          4228 => x"8025b938",
          4229 => x"82b5d408",
          4230 => x"88050830",
          4231 => x"82b5d408",
          4232 => x"88050c80",
          4233 => x"0b82b5d4",
          4234 => x"08f4050c",
          4235 => x"82b5d408",
          4236 => x"fc05088a",
          4237 => x"38810b82",
          4238 => x"b5d408f4",
          4239 => x"050c82b5",
          4240 => x"d408f405",
          4241 => x"0882b5d4",
          4242 => x"08fc050c",
          4243 => x"82b5d408",
          4244 => x"8c050880",
          4245 => x"25b93882",
          4246 => x"b5d4088c",
          4247 => x"05083082",
          4248 => x"b5d4088c",
          4249 => x"050c800b",
          4250 => x"82b5d408",
          4251 => x"f0050c82",
          4252 => x"b5d408fc",
          4253 => x"05088a38",
          4254 => x"810b82b5",
          4255 => x"d408f005",
          4256 => x"0c82b5d4",
          4257 => x"08f00508",
          4258 => x"82b5d408",
          4259 => x"fc050c80",
          4260 => x"5382b5d4",
          4261 => x"088c0508",
          4262 => x"5282b5d4",
          4263 => x"08880508",
          4264 => x"5182c53f",
          4265 => x"82b5c808",
          4266 => x"7082b5d4",
          4267 => x"08f8050c",
          4268 => x"5482b5d4",
          4269 => x"08fc0508",
          4270 => x"802e9038",
          4271 => x"82b5d408",
          4272 => x"f8050830",
          4273 => x"82b5d408",
          4274 => x"f8050c82",
          4275 => x"b5d408f8",
          4276 => x"05087082",
          4277 => x"b5c80c54",
          4278 => x"893d0d82",
          4279 => x"b5d40c04",
          4280 => x"82b5d408",
          4281 => x"0282b5d4",
          4282 => x"0cfb3d0d",
          4283 => x"800b82b5",
          4284 => x"d408fc05",
          4285 => x"0c82b5d4",
          4286 => x"08880508",
          4287 => x"80259938",
          4288 => x"82b5d408",
          4289 => x"88050830",
          4290 => x"82b5d408",
          4291 => x"88050c81",
          4292 => x"0b82b5d4",
          4293 => x"08fc050c",
          4294 => x"82b5d408",
          4295 => x"8c050880",
          4296 => x"25903882",
          4297 => x"b5d4088c",
          4298 => x"05083082",
          4299 => x"b5d4088c",
          4300 => x"050c8153",
          4301 => x"82b5d408",
          4302 => x"8c050852",
          4303 => x"82b5d408",
          4304 => x"88050851",
          4305 => x"81a23f82",
          4306 => x"b5c80870",
          4307 => x"82b5d408",
          4308 => x"f8050c54",
          4309 => x"82b5d408",
          4310 => x"fc050880",
          4311 => x"2e903882",
          4312 => x"b5d408f8",
          4313 => x"05083082",
          4314 => x"b5d408f8",
          4315 => x"050c82b5",
          4316 => x"d408f805",
          4317 => x"087082b5",
          4318 => x"c80c5487",
          4319 => x"3d0d82b5",
          4320 => x"d40c0482",
          4321 => x"b5d40802",
          4322 => x"82b5d40c",
          4323 => x"fd3d0d80",
          4324 => x"5382b5d4",
          4325 => x"088c0508",
          4326 => x"5282b5d4",
          4327 => x"08880508",
          4328 => x"5180c53f",
          4329 => x"82b5c808",
          4330 => x"7082b5c8",
          4331 => x"0c54853d",
          4332 => x"0d82b5d4",
          4333 => x"0c0482b5",
          4334 => x"d4080282",
          4335 => x"b5d40cfd",
          4336 => x"3d0d8153",
          4337 => x"82b5d408",
          4338 => x"8c050852",
          4339 => x"82b5d408",
          4340 => x"88050851",
          4341 => x"933f82b5",
          4342 => x"c8087082",
          4343 => x"b5c80c54",
          4344 => x"853d0d82",
          4345 => x"b5d40c04",
          4346 => x"82b5d408",
          4347 => x"0282b5d4",
          4348 => x"0cfd3d0d",
          4349 => x"810b82b5",
          4350 => x"d408fc05",
          4351 => x"0c800b82",
          4352 => x"b5d408f8",
          4353 => x"050c82b5",
          4354 => x"d4088c05",
          4355 => x"0882b5d4",
          4356 => x"08880508",
          4357 => x"27b93882",
          4358 => x"b5d408fc",
          4359 => x"0508802e",
          4360 => x"ae38800b",
          4361 => x"82b5d408",
          4362 => x"8c050824",
          4363 => x"a23882b5",
          4364 => x"d4088c05",
          4365 => x"081082b5",
          4366 => x"d4088c05",
          4367 => x"0c82b5d4",
          4368 => x"08fc0508",
          4369 => x"1082b5d4",
          4370 => x"08fc050c",
          4371 => x"ffb83982",
          4372 => x"b5d408fc",
          4373 => x"0508802e",
          4374 => x"80e13882",
          4375 => x"b5d4088c",
          4376 => x"050882b5",
          4377 => x"d4088805",
          4378 => x"0826ad38",
          4379 => x"82b5d408",
          4380 => x"88050882",
          4381 => x"b5d4088c",
          4382 => x"05083182",
          4383 => x"b5d40888",
          4384 => x"050c82b5",
          4385 => x"d408f805",
          4386 => x"0882b5d4",
          4387 => x"08fc0508",
          4388 => x"0782b5d4",
          4389 => x"08f8050c",
          4390 => x"82b5d408",
          4391 => x"fc050881",
          4392 => x"2a82b5d4",
          4393 => x"08fc050c",
          4394 => x"82b5d408",
          4395 => x"8c050881",
          4396 => x"2a82b5d4",
          4397 => x"088c050c",
          4398 => x"ff953982",
          4399 => x"b5d40890",
          4400 => x"0508802e",
          4401 => x"933882b5",
          4402 => x"d4088805",
          4403 => x"087082b5",
          4404 => x"d408f405",
          4405 => x"0c519139",
          4406 => x"82b5d408",
          4407 => x"f8050870",
          4408 => x"82b5d408",
          4409 => x"f4050c51",
          4410 => x"82b5d408",
          4411 => x"f4050882",
          4412 => x"b5c80c85",
          4413 => x"3d0d82b5",
          4414 => x"d40c0482",
          4415 => x"b5d40802",
          4416 => x"82b5d40c",
          4417 => x"f73d0d80",
          4418 => x"0b82b5d4",
          4419 => x"08f00534",
          4420 => x"82b5d408",
          4421 => x"8c050853",
          4422 => x"80730c82",
          4423 => x"b5d40888",
          4424 => x"05087008",
          4425 => x"51537233",
          4426 => x"537282b5",
          4427 => x"d408f805",
          4428 => x"347281ff",
          4429 => x"065372a0",
          4430 => x"2e098106",
          4431 => x"913882b5",
          4432 => x"d4088805",
          4433 => x"08700881",
          4434 => x"05710c53",
          4435 => x"ce3982b5",
          4436 => x"d408f805",
          4437 => x"335372ad",
          4438 => x"2e098106",
          4439 => x"a438810b",
          4440 => x"82b5d408",
          4441 => x"f0053482",
          4442 => x"b5d40888",
          4443 => x"05087008",
          4444 => x"8105710c",
          4445 => x"70085153",
          4446 => x"723382b5",
          4447 => x"d408f805",
          4448 => x"3482b5d4",
          4449 => x"08f80533",
          4450 => x"5372b02e",
          4451 => x"09810681",
          4452 => x"dc3882b5",
          4453 => x"d4088805",
          4454 => x"08700881",
          4455 => x"05710c70",
          4456 => x"08515372",
          4457 => x"3382b5d4",
          4458 => x"08f80534",
          4459 => x"82b5d408",
          4460 => x"f8053382",
          4461 => x"b5d408e8",
          4462 => x"050c82b5",
          4463 => x"d408e805",
          4464 => x"0880e22e",
          4465 => x"b63882b5",
          4466 => x"d408e805",
          4467 => x"0880f82e",
          4468 => x"843880cd",
          4469 => x"39900b82",
          4470 => x"b5d408f4",
          4471 => x"053482b5",
          4472 => x"d4088805",
          4473 => x"08700881",
          4474 => x"05710c70",
          4475 => x"08515372",
          4476 => x"3382b5d4",
          4477 => x"08f80534",
          4478 => x"81a43982",
          4479 => x"0b82b5d4",
          4480 => x"08f40534",
          4481 => x"82b5d408",
          4482 => x"88050870",
          4483 => x"08810571",
          4484 => x"0c700851",
          4485 => x"53723382",
          4486 => x"b5d408f8",
          4487 => x"053480fe",
          4488 => x"3982b5d4",
          4489 => x"08f80533",
          4490 => x"5372a026",
          4491 => x"8d38810b",
          4492 => x"82b5d408",
          4493 => x"ec050c83",
          4494 => x"803982b5",
          4495 => x"d408f805",
          4496 => x"3353af73",
          4497 => x"27903882",
          4498 => x"b5d408f8",
          4499 => x"05335372",
          4500 => x"b9268338",
          4501 => x"8d39800b",
          4502 => x"82b5d408",
          4503 => x"ec050c82",
          4504 => x"d839880b",
          4505 => x"82b5d408",
          4506 => x"f40534b2",
          4507 => x"3982b5d4",
          4508 => x"08f80533",
          4509 => x"53af7327",
          4510 => x"903882b5",
          4511 => x"d408f805",
          4512 => x"335372b9",
          4513 => x"2683388d",
          4514 => x"39800b82",
          4515 => x"b5d408ec",
          4516 => x"050c82a5",
          4517 => x"398a0b82",
          4518 => x"b5d408f4",
          4519 => x"0534800b",
          4520 => x"82b5d408",
          4521 => x"fc050c82",
          4522 => x"b5d408f8",
          4523 => x"053353a0",
          4524 => x"732781cf",
          4525 => x"3882b5d4",
          4526 => x"08f80533",
          4527 => x"5380e073",
          4528 => x"27943882",
          4529 => x"b5d408f8",
          4530 => x"0533e011",
          4531 => x"51537282",
          4532 => x"b5d408f8",
          4533 => x"053482b5",
          4534 => x"d408f805",
          4535 => x"33d01151",
          4536 => x"537282b5",
          4537 => x"d408f805",
          4538 => x"3482b5d4",
          4539 => x"08f80533",
          4540 => x"53907327",
          4541 => x"ad3882b5",
          4542 => x"d408f805",
          4543 => x"33f91151",
          4544 => x"537282b5",
          4545 => x"d408f805",
          4546 => x"3482b5d4",
          4547 => x"08f80533",
          4548 => x"53728926",
          4549 => x"8d38800b",
          4550 => x"82b5d408",
          4551 => x"ec050c81",
          4552 => x"983982b5",
          4553 => x"d408f805",
          4554 => x"3382b5d4",
          4555 => x"08f40533",
          4556 => x"54547274",
          4557 => x"268d3880",
          4558 => x"0b82b5d4",
          4559 => x"08ec050c",
          4560 => x"80f73982",
          4561 => x"b5d408f4",
          4562 => x"05337082",
          4563 => x"b5d408fc",
          4564 => x"05082982",
          4565 => x"b5d408f8",
          4566 => x"05337012",
          4567 => x"82b5d408",
          4568 => x"fc050c82",
          4569 => x"b5d40888",
          4570 => x"05087008",
          4571 => x"8105710c",
          4572 => x"70085151",
          4573 => x"52555372",
          4574 => x"3382b5d4",
          4575 => x"08f80534",
          4576 => x"fea53982",
          4577 => x"b5d408f0",
          4578 => x"05335372",
          4579 => x"802e9038",
          4580 => x"82b5d408",
          4581 => x"fc050830",
          4582 => x"82b5d408",
          4583 => x"fc050c82",
          4584 => x"b5d4088c",
          4585 => x"050882b5",
          4586 => x"d408fc05",
          4587 => x"08710c53",
          4588 => x"810b82b5",
          4589 => x"d408ec05",
          4590 => x"0c82b5d4",
          4591 => x"08ec0508",
          4592 => x"82b5c80c",
          4593 => x"8b3d0d82",
          4594 => x"b5d40c04",
          4595 => x"82b5d408",
          4596 => x"0282b5d4",
          4597 => x"0cf73d0d",
          4598 => x"800b82b5",
          4599 => x"d408f005",
          4600 => x"3482b5d4",
          4601 => x"088c0508",
          4602 => x"5380730c",
          4603 => x"82b5d408",
          4604 => x"88050870",
          4605 => x"08515372",
          4606 => x"33537282",
          4607 => x"b5d408f8",
          4608 => x"05347281",
          4609 => x"ff065372",
          4610 => x"a02e0981",
          4611 => x"06913882",
          4612 => x"b5d40888",
          4613 => x"05087008",
          4614 => x"8105710c",
          4615 => x"53ce3982",
          4616 => x"b5d408f8",
          4617 => x"05335372",
          4618 => x"ad2e0981",
          4619 => x"06a43881",
          4620 => x"0b82b5d4",
          4621 => x"08f00534",
          4622 => x"82b5d408",
          4623 => x"88050870",
          4624 => x"08810571",
          4625 => x"0c700851",
          4626 => x"53723382",
          4627 => x"b5d408f8",
          4628 => x"053482b5",
          4629 => x"d408f805",
          4630 => x"335372b0",
          4631 => x"2e098106",
          4632 => x"81dc3882",
          4633 => x"b5d40888",
          4634 => x"05087008",
          4635 => x"8105710c",
          4636 => x"70085153",
          4637 => x"723382b5",
          4638 => x"d408f805",
          4639 => x"3482b5d4",
          4640 => x"08f80533",
          4641 => x"82b5d408",
          4642 => x"e8050c82",
          4643 => x"b5d408e8",
          4644 => x"050880e2",
          4645 => x"2eb63882",
          4646 => x"b5d408e8",
          4647 => x"050880f8",
          4648 => x"2e843880",
          4649 => x"cd39900b",
          4650 => x"82b5d408",
          4651 => x"f4053482",
          4652 => x"b5d40888",
          4653 => x"05087008",
          4654 => x"8105710c",
          4655 => x"70085153",
          4656 => x"723382b5",
          4657 => x"d408f805",
          4658 => x"3481a439",
          4659 => x"820b82b5",
          4660 => x"d408f405",
          4661 => x"3482b5d4",
          4662 => x"08880508",
          4663 => x"70088105",
          4664 => x"710c7008",
          4665 => x"51537233",
          4666 => x"82b5d408",
          4667 => x"f8053480",
          4668 => x"fe3982b5",
          4669 => x"d408f805",
          4670 => x"335372a0",
          4671 => x"268d3881",
          4672 => x"0b82b5d4",
          4673 => x"08ec050c",
          4674 => x"83803982",
          4675 => x"b5d408f8",
          4676 => x"053353af",
          4677 => x"73279038",
          4678 => x"82b5d408",
          4679 => x"f8053353",
          4680 => x"72b92683",
          4681 => x"388d3980",
          4682 => x"0b82b5d4",
          4683 => x"08ec050c",
          4684 => x"82d83988",
          4685 => x"0b82b5d4",
          4686 => x"08f40534",
          4687 => x"b23982b5",
          4688 => x"d408f805",
          4689 => x"3353af73",
          4690 => x"27903882",
          4691 => x"b5d408f8",
          4692 => x"05335372",
          4693 => x"b9268338",
          4694 => x"8d39800b",
          4695 => x"82b5d408",
          4696 => x"ec050c82",
          4697 => x"a5398a0b",
          4698 => x"82b5d408",
          4699 => x"f4053480",
          4700 => x"0b82b5d4",
          4701 => x"08fc050c",
          4702 => x"82b5d408",
          4703 => x"f8053353",
          4704 => x"a0732781",
          4705 => x"cf3882b5",
          4706 => x"d408f805",
          4707 => x"335380e0",
          4708 => x"73279438",
          4709 => x"82b5d408",
          4710 => x"f80533e0",
          4711 => x"11515372",
          4712 => x"82b5d408",
          4713 => x"f8053482",
          4714 => x"b5d408f8",
          4715 => x"0533d011",
          4716 => x"51537282",
          4717 => x"b5d408f8",
          4718 => x"053482b5",
          4719 => x"d408f805",
          4720 => x"33539073",
          4721 => x"27ad3882",
          4722 => x"b5d408f8",
          4723 => x"0533f911",
          4724 => x"51537282",
          4725 => x"b5d408f8",
          4726 => x"053482b5",
          4727 => x"d408f805",
          4728 => x"33537289",
          4729 => x"268d3880",
          4730 => x"0b82b5d4",
          4731 => x"08ec050c",
          4732 => x"81983982",
          4733 => x"b5d408f8",
          4734 => x"053382b5",
          4735 => x"d408f405",
          4736 => x"33545472",
          4737 => x"74268d38",
          4738 => x"800b82b5",
          4739 => x"d408ec05",
          4740 => x"0c80f739",
          4741 => x"82b5d408",
          4742 => x"f4053370",
          4743 => x"82b5d408",
          4744 => x"fc050829",
          4745 => x"82b5d408",
          4746 => x"f8053370",
          4747 => x"1282b5d4",
          4748 => x"08fc050c",
          4749 => x"82b5d408",
          4750 => x"88050870",
          4751 => x"08810571",
          4752 => x"0c700851",
          4753 => x"51525553",
          4754 => x"723382b5",
          4755 => x"d408f805",
          4756 => x"34fea539",
          4757 => x"82b5d408",
          4758 => x"f0053353",
          4759 => x"72802e90",
          4760 => x"3882b5d4",
          4761 => x"08fc0508",
          4762 => x"3082b5d4",
          4763 => x"08fc050c",
          4764 => x"82b5d408",
          4765 => x"8c050882",
          4766 => x"b5d408fc",
          4767 => x"0508710c",
          4768 => x"53810b82",
          4769 => x"b5d408ec",
          4770 => x"050c82b5",
          4771 => x"d408ec05",
          4772 => x"0882b5c8",
          4773 => x"0c8b3d0d",
          4774 => x"82b5d40c",
          4775 => x"04f93d0d",
          4776 => x"79700870",
          4777 => x"56565874",
          4778 => x"802e80e3",
          4779 => x"38953975",
          4780 => x"0851e6d1",
          4781 => x"3f82b5c8",
          4782 => x"0815780c",
          4783 => x"85163354",
          4784 => x"80cd3974",
          4785 => x"335473a0",
          4786 => x"2e098106",
          4787 => x"86388115",
          4788 => x"55f13980",
          4789 => x"57769029",
          4790 => x"82b0c805",
          4791 => x"70085256",
          4792 => x"e6a33f82",
          4793 => x"b5c80853",
          4794 => x"74527508",
          4795 => x"51e9a33f",
          4796 => x"82b5c808",
          4797 => x"8b388416",
          4798 => x"33547381",
          4799 => x"2effb038",
          4800 => x"81177081",
          4801 => x"ff065854",
          4802 => x"997727c9",
          4803 => x"38ff5473",
          4804 => x"82b5c80c",
          4805 => x"893d0d04",
          4806 => x"ff3d0d73",
          4807 => x"52719326",
          4808 => x"818e3871",
          4809 => x"84298295",
          4810 => x"a8055271",
          4811 => x"0804829a",
          4812 => x"f4518180",
          4813 => x"39829b80",
          4814 => x"5180f939",
          4815 => x"829b9051",
          4816 => x"80f23982",
          4817 => x"9ba05180",
          4818 => x"eb39829b",
          4819 => x"b05180e4",
          4820 => x"39829bc0",
          4821 => x"5180dd39",
          4822 => x"829bd451",
          4823 => x"80d63982",
          4824 => x"9be45180",
          4825 => x"cf39829b",
          4826 => x"fc5180c8",
          4827 => x"39829c94",
          4828 => x"5180c139",
          4829 => x"829cac51",
          4830 => x"bb39829c",
          4831 => x"c851b539",
          4832 => x"829cdc51",
          4833 => x"af39829d",
          4834 => x"8451a939",
          4835 => x"829d9451",
          4836 => x"a339829d",
          4837 => x"b4519d39",
          4838 => x"829dc451",
          4839 => x"9739829d",
          4840 => x"dc519139",
          4841 => x"829df451",
          4842 => x"8b39829e",
          4843 => x"8c518539",
          4844 => x"829e9851",
          4845 => x"d8ad3f83",
          4846 => x"3d0d04fb",
          4847 => x"3d0d7779",
          4848 => x"56567487",
          4849 => x"e7268a38",
          4850 => x"74527587",
          4851 => x"e8295190",
          4852 => x"3987e852",
          4853 => x"7451efab",
          4854 => x"3f82b5c8",
          4855 => x"08527551",
          4856 => x"efa13f82",
          4857 => x"b5c80854",
          4858 => x"79537552",
          4859 => x"829ea851",
          4860 => x"ffbbe53f",
          4861 => x"873d0d04",
          4862 => x"ec3d0d66",
          4863 => x"02840580",
          4864 => x"e305335b",
          4865 => x"57806878",
          4866 => x"30707a07",
          4867 => x"73255157",
          4868 => x"59597856",
          4869 => x"7787ff26",
          4870 => x"83388156",
          4871 => x"74760770",
          4872 => x"81ff0651",
          4873 => x"55935674",
          4874 => x"81823881",
          4875 => x"5376528c",
          4876 => x"3d705256",
          4877 => x"80ffc53f",
          4878 => x"82b5c808",
          4879 => x"5782b5c8",
          4880 => x"08b93882",
          4881 => x"b5c80887",
          4882 => x"c098880c",
          4883 => x"82b5c808",
          4884 => x"59963dd4",
          4885 => x"05548480",
          4886 => x"53775275",
          4887 => x"51818481",
          4888 => x"3f82b5c8",
          4889 => x"085782b5",
          4890 => x"c8089038",
          4891 => x"7a557480",
          4892 => x"2e893874",
          4893 => x"19751959",
          4894 => x"59d73996",
          4895 => x"3dd80551",
          4896 => x"818bea3f",
          4897 => x"76307078",
          4898 => x"0780257b",
          4899 => x"30709f2a",
          4900 => x"72065157",
          4901 => x"51567480",
          4902 => x"2e903882",
          4903 => x"9ecc5387",
          4904 => x"c0988808",
          4905 => x"527851fe",
          4906 => x"923f7656",
          4907 => x"7582b5c8",
          4908 => x"0c963d0d",
          4909 => x"04f83d0d",
          4910 => x"7c028405",
          4911 => x"b7053358",
          4912 => x"59ff5880",
          4913 => x"537b527a",
          4914 => x"51fead3f",
          4915 => x"82b5c808",
          4916 => x"a8387680",
          4917 => x"2e883876",
          4918 => x"812e9c38",
          4919 => x"9c3982cd",
          4920 => x"98566155",
          4921 => x"605482b5",
          4922 => x"c8537f52",
          4923 => x"7e51782d",
          4924 => x"82b5c808",
          4925 => x"58833978",
          4926 => x"047782b5",
          4927 => x"c80c8a3d",
          4928 => x"0d04f33d",
          4929 => x"0d7f6163",
          4930 => x"028c0580",
          4931 => x"cf053373",
          4932 => x"73156841",
          4933 => x"5f5c5c5e",
          4934 => x"5e5e7a52",
          4935 => x"829ed451",
          4936 => x"ffb9b53f",
          4937 => x"829edc51",
          4938 => x"ffb9ad3f",
          4939 => x"80557479",
          4940 => x"27818038",
          4941 => x"7b902e89",
          4942 => x"387ba02e",
          4943 => x"a73880c6",
          4944 => x"39741853",
          4945 => x"727a278e",
          4946 => x"38722252",
          4947 => x"829ee051",
          4948 => x"ffb9853f",
          4949 => x"8939829e",
          4950 => x"ec51ffb8",
          4951 => x"fb3f8215",
          4952 => x"5580c339",
          4953 => x"74185372",
          4954 => x"7a278e38",
          4955 => x"72085282",
          4956 => x"9ed451ff",
          4957 => x"b8e23f89",
          4958 => x"39829ee8",
          4959 => x"51ffb8d8",
          4960 => x"3f841555",
          4961 => x"a1397418",
          4962 => x"53727a27",
          4963 => x"8e387233",
          4964 => x"52829ef4",
          4965 => x"51ffb8c0",
          4966 => x"3f893982",
          4967 => x"9efc51ff",
          4968 => x"b8b63f81",
          4969 => x"155582cd",
          4970 => x"9c0852a0",
          4971 => x"51d8833f",
          4972 => x"fefc3982",
          4973 => x"9f8051ff",
          4974 => x"b89e3f80",
          4975 => x"55747927",
          4976 => x"80c63874",
          4977 => x"18703355",
          4978 => x"53805672",
          4979 => x"7a278338",
          4980 => x"81568053",
          4981 => x"9f742783",
          4982 => x"38815375",
          4983 => x"73067081",
          4984 => x"ff065153",
          4985 => x"72802e90",
          4986 => x"387380fe",
          4987 => x"268a3882",
          4988 => x"cd9c0852",
          4989 => x"73518839",
          4990 => x"82cd9c08",
          4991 => x"52a051d7",
          4992 => x"b13f8115",
          4993 => x"55ffb639",
          4994 => x"829f8451",
          4995 => x"d3d53f78",
          4996 => x"18791c5c",
          4997 => x"589ccb3f",
          4998 => x"82b5c808",
          4999 => x"982b7098",
          5000 => x"2c515776",
          5001 => x"a02e0981",
          5002 => x"06aa389c",
          5003 => x"b53f82b5",
          5004 => x"c808982b",
          5005 => x"70982c70",
          5006 => x"a0327030",
          5007 => x"729b3270",
          5008 => x"30707207",
          5009 => x"73750706",
          5010 => x"51585859",
          5011 => x"57515780",
          5012 => x"7324d838",
          5013 => x"769b2e09",
          5014 => x"81068538",
          5015 => x"80538c39",
          5016 => x"7c1e5372",
          5017 => x"7826fdb2",
          5018 => x"38ff5372",
          5019 => x"82b5c80c",
          5020 => x"8f3d0d04",
          5021 => x"fc3d0d02",
          5022 => x"9b053382",
          5023 => x"9f885382",
          5024 => x"9f8c5255",
          5025 => x"ffb6d13f",
          5026 => x"82b4a022",
          5027 => x"51a5a63f",
          5028 => x"829f9854",
          5029 => x"829fa453",
          5030 => x"82b4a133",
          5031 => x"52829fac",
          5032 => x"51ffb6b4",
          5033 => x"3f74802e",
          5034 => x"8438a0d8",
          5035 => x"3f863d0d",
          5036 => x"04fe3d0d",
          5037 => x"87c09680",
          5038 => x"0853a5c2",
          5039 => x"3f815198",
          5040 => x"8e3f829f",
          5041 => x"c85199a3",
          5042 => x"3f805198",
          5043 => x"823f7281",
          5044 => x"2a708106",
          5045 => x"51527180",
          5046 => x"2e923881",
          5047 => x"5197f03f",
          5048 => x"829fe051",
          5049 => x"99853f80",
          5050 => x"5197e43f",
          5051 => x"72822a70",
          5052 => x"81065152",
          5053 => x"71802e92",
          5054 => x"38815197",
          5055 => x"d23f829f",
          5056 => x"f05198e7",
          5057 => x"3f805197",
          5058 => x"c63f7283",
          5059 => x"2a708106",
          5060 => x"51527180",
          5061 => x"2e923881",
          5062 => x"5197b43f",
          5063 => x"82a08051",
          5064 => x"98c93f80",
          5065 => x"5197a83f",
          5066 => x"72842a70",
          5067 => x"81065152",
          5068 => x"71802e92",
          5069 => x"38815197",
          5070 => x"963f82a0",
          5071 => x"945198ab",
          5072 => x"3f805197",
          5073 => x"8a3f7285",
          5074 => x"2a708106",
          5075 => x"51527180",
          5076 => x"2e923881",
          5077 => x"5196f83f",
          5078 => x"82a0a851",
          5079 => x"988d3f80",
          5080 => x"5196ec3f",
          5081 => x"72862a70",
          5082 => x"81065152",
          5083 => x"71802e92",
          5084 => x"38815196",
          5085 => x"da3f82a0",
          5086 => x"bc5197ef",
          5087 => x"3f805196",
          5088 => x"ce3f7287",
          5089 => x"2a708106",
          5090 => x"51527180",
          5091 => x"2e923881",
          5092 => x"5196bc3f",
          5093 => x"82a0d051",
          5094 => x"97d13f80",
          5095 => x"5196b03f",
          5096 => x"72882a70",
          5097 => x"81065152",
          5098 => x"71802e92",
          5099 => x"38815196",
          5100 => x"9e3f82a0",
          5101 => x"e45197b3",
          5102 => x"3f805196",
          5103 => x"923fa3c6",
          5104 => x"3f843d0d",
          5105 => x"04fb3d0d",
          5106 => x"77028405",
          5107 => x"a3053370",
          5108 => x"55565680",
          5109 => x"527551e3",
          5110 => x"8d3f0b0b",
          5111 => x"82b0c433",
          5112 => x"5473a938",
          5113 => x"815382a1",
          5114 => x"a05282cc",
          5115 => x"c85180f8",
          5116 => x"8b3f82b5",
          5117 => x"c8083070",
          5118 => x"82b5c808",
          5119 => x"07802582",
          5120 => x"71315151",
          5121 => x"54730b0b",
          5122 => x"82b0c434",
          5123 => x"0b0b82b0",
          5124 => x"c4335473",
          5125 => x"812e0981",
          5126 => x"06af3882",
          5127 => x"ccc85374",
          5128 => x"52755181",
          5129 => x"b2bc3f82",
          5130 => x"b5c80880",
          5131 => x"2e8b3882",
          5132 => x"b5c80851",
          5133 => x"cfad3f91",
          5134 => x"3982ccc8",
          5135 => x"518184ad",
          5136 => x"3f820b0b",
          5137 => x"0b82b0c4",
          5138 => x"340b0b82",
          5139 => x"b0c43354",
          5140 => x"73822e09",
          5141 => x"81068c38",
          5142 => x"82a1b053",
          5143 => x"74527551",
          5144 => x"a9be3f80",
          5145 => x"0b82b5c8",
          5146 => x"0c873d0d",
          5147 => x"04ce3d0d",
          5148 => x"80707182",
          5149 => x"ccc40c5f",
          5150 => x"5d81527c",
          5151 => x"5180c6d7",
          5152 => x"3f82b5c8",
          5153 => x"0881ff06",
          5154 => x"59787d2e",
          5155 => x"098106a3",
          5156 => x"38963d59",
          5157 => x"835382a1",
          5158 => x"b8527851",
          5159 => x"dcc73f7c",
          5160 => x"53785282",
          5161 => x"b6f45180",
          5162 => x"f5f13f82",
          5163 => x"b5c8087d",
          5164 => x"2e883882",
          5165 => x"a1bc518d",
          5166 => x"a3398170",
          5167 => x"5f5d82a1",
          5168 => x"f451ffb2",
          5169 => x"933f963d",
          5170 => x"70465a80",
          5171 => x"f8527951",
          5172 => x"fdf33fb4",
          5173 => x"3dff8405",
          5174 => x"51f3c23f",
          5175 => x"82b5c808",
          5176 => x"902b7090",
          5177 => x"2c515978",
          5178 => x"80c22e87",
          5179 => x"a3387880",
          5180 => x"c224b238",
          5181 => x"78bd2e81",
          5182 => x"d23878bd",
          5183 => x"24903878",
          5184 => x"802effba",
          5185 => x"3878bc2e",
          5186 => x"80da388a",
          5187 => x"d4397880",
          5188 => x"c02e8399",
          5189 => x"387880c0",
          5190 => x"2485cd38",
          5191 => x"78bf2e82",
          5192 => x"8c388abd",
          5193 => x"397880f9",
          5194 => x"2e89d938",
          5195 => x"7880f924",
          5196 => x"92387880",
          5197 => x"c32e8888",
          5198 => x"387880f8",
          5199 => x"2e89a138",
          5200 => x"8a9f3978",
          5201 => x"81832e8a",
          5202 => x"86387881",
          5203 => x"83248b38",
          5204 => x"7881822e",
          5205 => x"89eb388a",
          5206 => x"88397881",
          5207 => x"852e89fb",
          5208 => x"3889fe39",
          5209 => x"b43dff80",
          5210 => x"1153ff84",
          5211 => x"0551ecdc",
          5212 => x"3f82b5c8",
          5213 => x"08802efe",
          5214 => x"c538b43d",
          5215 => x"fefc1153",
          5216 => x"ff840551",
          5217 => x"ecc63f82",
          5218 => x"b5c80880",
          5219 => x"2efeaf38",
          5220 => x"b43dfef8",
          5221 => x"1153ff84",
          5222 => x"0551ecb0",
          5223 => x"3f82b5c8",
          5224 => x"08863882",
          5225 => x"b5c80842",
          5226 => x"82a1f851",
          5227 => x"ffb0a93f",
          5228 => x"63635c5a",
          5229 => x"797b2781",
          5230 => x"ec386159",
          5231 => x"787a7084",
          5232 => x"055c0c7a",
          5233 => x"7a26f538",
          5234 => x"81db39b4",
          5235 => x"3dff8011",
          5236 => x"53ff8405",
          5237 => x"51ebf53f",
          5238 => x"82b5c808",
          5239 => x"802efdde",
          5240 => x"38b43dfe",
          5241 => x"fc1153ff",
          5242 => x"840551eb",
          5243 => x"df3f82b5",
          5244 => x"c808802e",
          5245 => x"fdc838b4",
          5246 => x"3dfef811",
          5247 => x"53ff8405",
          5248 => x"51ebc93f",
          5249 => x"82b5c808",
          5250 => x"802efdb2",
          5251 => x"3882a288",
          5252 => x"51ffafc4",
          5253 => x"3f635a79",
          5254 => x"63278189",
          5255 => x"38615979",
          5256 => x"7081055b",
          5257 => x"33793461",
          5258 => x"810542eb",
          5259 => x"39b43dff",
          5260 => x"801153ff",
          5261 => x"840551eb",
          5262 => x"933f82b5",
          5263 => x"c808802e",
          5264 => x"fcfc38b4",
          5265 => x"3dfefc11",
          5266 => x"53ff8405",
          5267 => x"51eafd3f",
          5268 => x"82b5c808",
          5269 => x"802efce6",
          5270 => x"38b43dfe",
          5271 => x"f81153ff",
          5272 => x"840551ea",
          5273 => x"e73f82b5",
          5274 => x"c808802e",
          5275 => x"fcd03882",
          5276 => x"a29451ff",
          5277 => x"aee23f63",
          5278 => x"5a796327",
          5279 => x"a8386170",
          5280 => x"337b335e",
          5281 => x"5a5b787c",
          5282 => x"2e923878",
          5283 => x"557a5479",
          5284 => x"33537952",
          5285 => x"82a2a451",
          5286 => x"ffaebd3f",
          5287 => x"811a6281",
          5288 => x"05435ad5",
          5289 => x"398a51cd",
          5290 => x"dc3ffc92",
          5291 => x"39b43dff",
          5292 => x"801153ff",
          5293 => x"840551ea",
          5294 => x"933f82b5",
          5295 => x"c80880df",
          5296 => x"3882b4b4",
          5297 => x"33597880",
          5298 => x"2e893882",
          5299 => x"b3ec0844",
          5300 => x"80cd3982",
          5301 => x"b4b53359",
          5302 => x"78802e88",
          5303 => x"3882b3f4",
          5304 => x"0844bc39",
          5305 => x"82b4b633",
          5306 => x"5978802e",
          5307 => x"883882b3",
          5308 => x"fc0844ab",
          5309 => x"3982b4b7",
          5310 => x"33597880",
          5311 => x"2e883882",
          5312 => x"b4840844",
          5313 => x"9a3982b4",
          5314 => x"b2335978",
          5315 => x"802e8838",
          5316 => x"82b48c08",
          5317 => x"44893982",
          5318 => x"b49c08fc",
          5319 => x"800544b4",
          5320 => x"3dfefc11",
          5321 => x"53ff8405",
          5322 => x"51e9a13f",
          5323 => x"82b5c808",
          5324 => x"80de3882",
          5325 => x"b4b43359",
          5326 => x"78802e89",
          5327 => x"3882b3f0",
          5328 => x"084380cc",
          5329 => x"3982b4b5",
          5330 => x"33597880",
          5331 => x"2e883882",
          5332 => x"b3f80843",
          5333 => x"bb3982b4",
          5334 => x"b6335978",
          5335 => x"802e8838",
          5336 => x"82b48008",
          5337 => x"43aa3982",
          5338 => x"b4b73359",
          5339 => x"78802e88",
          5340 => x"3882b488",
          5341 => x"08439939",
          5342 => x"82b4b233",
          5343 => x"5978802e",
          5344 => x"883882b4",
          5345 => x"90084388",
          5346 => x"3982b49c",
          5347 => x"08880543",
          5348 => x"b43dfef8",
          5349 => x"1153ff84",
          5350 => x"0551e8b0",
          5351 => x"3f82b5c8",
          5352 => x"08802ea7",
          5353 => x"3880625c",
          5354 => x"5c7a882e",
          5355 => x"8338815c",
          5356 => x"7a903270",
          5357 => x"30707207",
          5358 => x"9f2a707f",
          5359 => x"0651515a",
          5360 => x"5a78802e",
          5361 => x"88387aa0",
          5362 => x"2e833888",
          5363 => x"4282a2c0",
          5364 => x"51c8903f",
          5365 => x"a0556354",
          5366 => x"61536252",
          5367 => x"6351f2a2",
          5368 => x"3f82a2cc",
          5369 => x"5186f539",
          5370 => x"b43dff80",
          5371 => x"1153ff84",
          5372 => x"0551e7d8",
          5373 => x"3f82b5c8",
          5374 => x"08802ef9",
          5375 => x"c138b43d",
          5376 => x"fefc1153",
          5377 => x"ff840551",
          5378 => x"e7c23f82",
          5379 => x"b5c80880",
          5380 => x"2ea43863",
          5381 => x"590280cb",
          5382 => x"05337934",
          5383 => x"63810544",
          5384 => x"b43dfefc",
          5385 => x"1153ff84",
          5386 => x"0551e7a0",
          5387 => x"3f82b5c8",
          5388 => x"08e138f9",
          5389 => x"89396370",
          5390 => x"33545282",
          5391 => x"a2d851ff",
          5392 => x"ab963f82",
          5393 => x"cd980853",
          5394 => x"80f85279",
          5395 => x"51ffabdd",
          5396 => x"3f794579",
          5397 => x"335978ae",
          5398 => x"2ef8e338",
          5399 => x"9f79279f",
          5400 => x"38b43dfe",
          5401 => x"fc1153ff",
          5402 => x"840551e6",
          5403 => x"df3f82b5",
          5404 => x"c808802e",
          5405 => x"91386359",
          5406 => x"0280cb05",
          5407 => x"33793463",
          5408 => x"810544ff",
          5409 => x"b13982a2",
          5410 => x"e451c6d7",
          5411 => x"3fffa739",
          5412 => x"b43dfef4",
          5413 => x"1153ff84",
          5414 => x"0551e0df",
          5415 => x"3f82b5c8",
          5416 => x"08802ef8",
          5417 => x"9938b43d",
          5418 => x"fef01153",
          5419 => x"ff840551",
          5420 => x"e0c93f82",
          5421 => x"b5c80880",
          5422 => x"2ea53860",
          5423 => x"5902be05",
          5424 => x"22797082",
          5425 => x"055b2378",
          5426 => x"41b43dfe",
          5427 => x"f01153ff",
          5428 => x"840551e0",
          5429 => x"a63f82b5",
          5430 => x"c808e038",
          5431 => x"f7e03960",
          5432 => x"70225452",
          5433 => x"82a2e851",
          5434 => x"ffa9ed3f",
          5435 => x"82cd9808",
          5436 => x"5380f852",
          5437 => x"7951ffaa",
          5438 => x"b43f7945",
          5439 => x"79335978",
          5440 => x"ae2ef7ba",
          5441 => x"38789f26",
          5442 => x"87386082",
          5443 => x"0541d039",
          5444 => x"b43dfef0",
          5445 => x"1153ff84",
          5446 => x"0551dfdf",
          5447 => x"3f82b5c8",
          5448 => x"08802e92",
          5449 => x"38605902",
          5450 => x"be052279",
          5451 => x"7082055b",
          5452 => x"237841ff",
          5453 => x"aa3982a2",
          5454 => x"e451c5a7",
          5455 => x"3fffa039",
          5456 => x"b43dfef4",
          5457 => x"1153ff84",
          5458 => x"0551dfaf",
          5459 => x"3f82b5c8",
          5460 => x"08802ef6",
          5461 => x"e938b43d",
          5462 => x"fef01153",
          5463 => x"ff840551",
          5464 => x"df993f82",
          5465 => x"b5c80880",
          5466 => x"2ea03860",
          5467 => x"60710c59",
          5468 => x"60840541",
          5469 => x"b43dfef0",
          5470 => x"1153ff84",
          5471 => x"0551defb",
          5472 => x"3f82b5c8",
          5473 => x"08e538f6",
          5474 => x"b5396070",
          5475 => x"08545282",
          5476 => x"a2f451ff",
          5477 => x"a8c23f82",
          5478 => x"cd980853",
          5479 => x"80f85279",
          5480 => x"51ffa989",
          5481 => x"3f794579",
          5482 => x"335978ae",
          5483 => x"2ef68f38",
          5484 => x"9f79279b",
          5485 => x"38b43dfe",
          5486 => x"f01153ff",
          5487 => x"840551de",
          5488 => x"ba3f82b5",
          5489 => x"c808802e",
          5490 => x"8d386060",
          5491 => x"710c5960",
          5492 => x"840541ff",
          5493 => x"b53982a2",
          5494 => x"e451c487",
          5495 => x"3fffab39",
          5496 => x"b43dff80",
          5497 => x"1153ff84",
          5498 => x"0551e3e0",
          5499 => x"3f82b5c8",
          5500 => x"08802ef5",
          5501 => x"c9386352",
          5502 => x"82a38451",
          5503 => x"ffa7d93f",
          5504 => x"63597804",
          5505 => x"b43dff80",
          5506 => x"1153ff84",
          5507 => x"0551e3bc",
          5508 => x"3f82b5c8",
          5509 => x"08802ef5",
          5510 => x"a5386352",
          5511 => x"82a3a051",
          5512 => x"ffa7b53f",
          5513 => x"6359782d",
          5514 => x"82b5c808",
          5515 => x"802ef58e",
          5516 => x"3882b5c8",
          5517 => x"085282a3",
          5518 => x"bc51ffa7",
          5519 => x"9b3ff4fe",
          5520 => x"3982a3d8",
          5521 => x"51c39c3f",
          5522 => x"ffa6ee3f",
          5523 => x"f4f03982",
          5524 => x"a3f451c3",
          5525 => x"8e3f8059",
          5526 => x"ffa83991",
          5527 => x"a73ff4de",
          5528 => x"39794579",
          5529 => x"33597880",
          5530 => x"2ef4d338",
          5531 => x"7d7d0659",
          5532 => x"78802e81",
          5533 => x"cf38b43d",
          5534 => x"ff840551",
          5535 => x"83ca3f82",
          5536 => x"b5c8085c",
          5537 => x"815b7a82",
          5538 => x"2eb2387a",
          5539 => x"82248938",
          5540 => x"7a812e8c",
          5541 => x"3880ca39",
          5542 => x"7a832ead",
          5543 => x"3880c239",
          5544 => x"82a48856",
          5545 => x"7b5582a4",
          5546 => x"8c548053",
          5547 => x"82a49052",
          5548 => x"b43dffb0",
          5549 => x"0551ffa9",
          5550 => x"873fb839",
          5551 => x"7b52b43d",
          5552 => x"ffb00551",
          5553 => x"cfad3fab",
          5554 => x"397b5582",
          5555 => x"a48c5480",
          5556 => x"5382a4a0",
          5557 => x"52b43dff",
          5558 => x"b00551ff",
          5559 => x"a8e23f93",
          5560 => x"397b5480",
          5561 => x"5382a4ac",
          5562 => x"52b43dff",
          5563 => x"b00551ff",
          5564 => x"a8ce3f82",
          5565 => x"b3ec5882",
          5566 => x"b5f85780",
          5567 => x"56645580",
          5568 => x"5482d080",
          5569 => x"5382d080",
          5570 => x"52b43dff",
          5571 => x"b00551eb",
          5572 => x"a43f82b5",
          5573 => x"c80882b5",
          5574 => x"c8080970",
          5575 => x"30707207",
          5576 => x"8025515b",
          5577 => x"5b5f805a",
          5578 => x"7a832683",
          5579 => x"38815a78",
          5580 => x"7a065978",
          5581 => x"802e8d38",
          5582 => x"811b7081",
          5583 => x"ff065c59",
          5584 => x"7afec338",
          5585 => x"7d81327d",
          5586 => x"81320759",
          5587 => x"788a387e",
          5588 => x"ff2e0981",
          5589 => x"06f2e738",
          5590 => x"82a4b451",
          5591 => x"c1853ff2",
          5592 => x"dd39f53d",
          5593 => x"0d800b82",
          5594 => x"b5f83487",
          5595 => x"c0948c70",
          5596 => x"08545587",
          5597 => x"84805272",
          5598 => x"51d8883f",
          5599 => x"82b5c808",
          5600 => x"902b7508",
          5601 => x"55538784",
          5602 => x"80527351",
          5603 => x"d7f53f72",
          5604 => x"82b5c808",
          5605 => x"07750c87",
          5606 => x"c0949c70",
          5607 => x"08545587",
          5608 => x"84805272",
          5609 => x"51d7dc3f",
          5610 => x"82b5c808",
          5611 => x"902b7508",
          5612 => x"55538784",
          5613 => x"80527351",
          5614 => x"d7c93f72",
          5615 => x"82b5c808",
          5616 => x"07750c8c",
          5617 => x"80830b87",
          5618 => x"c094840c",
          5619 => x"8c80830b",
          5620 => x"87c09494",
          5621 => x"0c80f5e7",
          5622 => x"5a80f8d3",
          5623 => x"5b830284",
          5624 => x"05990534",
          5625 => x"805c82cd",
          5626 => x"980b873d",
          5627 => x"7088130c",
          5628 => x"70720c82",
          5629 => x"cd9c0c54",
          5630 => x"89be3f93",
          5631 => x"813f82a4",
          5632 => x"c451ffbf",
          5633 => x"de3f82a4",
          5634 => x"d051ffbf",
          5635 => x"d63f80dd",
          5636 => x"b15192e5",
          5637 => x"3f8151ec",
          5638 => x"db3ff0d1",
          5639 => x"3f8004fe",
          5640 => x"3d0d8052",
          5641 => x"83537188",
          5642 => x"2b5287d8",
          5643 => x"3f82b5c8",
          5644 => x"0881ff06",
          5645 => x"7207ff14",
          5646 => x"54527280",
          5647 => x"25e83871",
          5648 => x"82b5c80c",
          5649 => x"843d0d04",
          5650 => x"fc3d0d76",
          5651 => x"70085455",
          5652 => x"80735254",
          5653 => x"72742e81",
          5654 => x"8a387233",
          5655 => x"5170a02e",
          5656 => x"09810686",
          5657 => x"38811353",
          5658 => x"f1397233",
          5659 => x"5170a22e",
          5660 => x"09810686",
          5661 => x"38811353",
          5662 => x"81547252",
          5663 => x"73812e09",
          5664 => x"81069f38",
          5665 => x"84398112",
          5666 => x"52807233",
          5667 => x"525470a2",
          5668 => x"2e833881",
          5669 => x"5470802e",
          5670 => x"9d3873ea",
          5671 => x"38983981",
          5672 => x"12528072",
          5673 => x"33525470",
          5674 => x"a02e8338",
          5675 => x"81547080",
          5676 => x"2e843873",
          5677 => x"ea388072",
          5678 => x"33525470",
          5679 => x"a02e0981",
          5680 => x"06833881",
          5681 => x"5470a232",
          5682 => x"70307080",
          5683 => x"25760751",
          5684 => x"51517080",
          5685 => x"2e883880",
          5686 => x"72708105",
          5687 => x"54347175",
          5688 => x"0c725170",
          5689 => x"82b5c80c",
          5690 => x"863d0d04",
          5691 => x"fc3d0d76",
          5692 => x"53720880",
          5693 => x"2e913886",
          5694 => x"3dfc0552",
          5695 => x"7251d7fb",
          5696 => x"3f82b5c8",
          5697 => x"08853880",
          5698 => x"53833974",
          5699 => x"537282b5",
          5700 => x"c80c863d",
          5701 => x"0d04fc3d",
          5702 => x"0d768211",
          5703 => x"33ff0552",
          5704 => x"53815270",
          5705 => x"8b268198",
          5706 => x"38831333",
          5707 => x"ff055182",
          5708 => x"52709e26",
          5709 => x"818a3884",
          5710 => x"13335183",
          5711 => x"52709726",
          5712 => x"80fe3885",
          5713 => x"13335184",
          5714 => x"5270bb26",
          5715 => x"80f23886",
          5716 => x"13335185",
          5717 => x"5270bb26",
          5718 => x"80e63888",
          5719 => x"13225586",
          5720 => x"527487e7",
          5721 => x"2680d938",
          5722 => x"8a132254",
          5723 => x"87527387",
          5724 => x"e72680cc",
          5725 => x"38810b87",
          5726 => x"c0989c0c",
          5727 => x"722287c0",
          5728 => x"98bc0c82",
          5729 => x"133387c0",
          5730 => x"98b80c83",
          5731 => x"133387c0",
          5732 => x"98b40c84",
          5733 => x"133387c0",
          5734 => x"98b00c85",
          5735 => x"133387c0",
          5736 => x"98ac0c86",
          5737 => x"133387c0",
          5738 => x"98a80c74",
          5739 => x"87c098a4",
          5740 => x"0c7387c0",
          5741 => x"98a00c80",
          5742 => x"0b87c098",
          5743 => x"9c0c8052",
          5744 => x"7182b5c8",
          5745 => x"0c863d0d",
          5746 => x"04f33d0d",
          5747 => x"7f5b87c0",
          5748 => x"989c5d81",
          5749 => x"7d0c87c0",
          5750 => x"98bc085e",
          5751 => x"7d7b2387",
          5752 => x"c098b808",
          5753 => x"5a79821c",
          5754 => x"3487c098",
          5755 => x"b4085a79",
          5756 => x"831c3487",
          5757 => x"c098b008",
          5758 => x"5a79841c",
          5759 => x"3487c098",
          5760 => x"ac085a79",
          5761 => x"851c3487",
          5762 => x"c098a808",
          5763 => x"5a79861c",
          5764 => x"3487c098",
          5765 => x"a4085c7b",
          5766 => x"881c2387",
          5767 => x"c098a008",
          5768 => x"5a798a1c",
          5769 => x"23807d0c",
          5770 => x"7983ffff",
          5771 => x"06597b83",
          5772 => x"ffff0658",
          5773 => x"861b3357",
          5774 => x"851b3356",
          5775 => x"841b3355",
          5776 => x"831b3354",
          5777 => x"821b3353",
          5778 => x"7d83ffff",
          5779 => x"065282a4",
          5780 => x"e851ff9f",
          5781 => x"833f8f3d",
          5782 => x"0d04fb3d",
          5783 => x"0d029f05",
          5784 => x"3382b3e8",
          5785 => x"337081ff",
          5786 => x"06585555",
          5787 => x"87c09484",
          5788 => x"5175802e",
          5789 => x"863887c0",
          5790 => x"94945170",
          5791 => x"0870962a",
          5792 => x"70810653",
          5793 => x"54527080",
          5794 => x"2e8c3871",
          5795 => x"912a7081",
          5796 => x"06515170",
          5797 => x"d7387281",
          5798 => x"32708106",
          5799 => x"51517080",
          5800 => x"2e8d3871",
          5801 => x"932a7081",
          5802 => x"06515170",
          5803 => x"ffbe3873",
          5804 => x"81ff0651",
          5805 => x"87c09480",
          5806 => x"5270802e",
          5807 => x"863887c0",
          5808 => x"94905274",
          5809 => x"720c7482",
          5810 => x"b5c80c87",
          5811 => x"3d0d04ff",
          5812 => x"3d0d028f",
          5813 => x"05337030",
          5814 => x"709f2a51",
          5815 => x"52527082",
          5816 => x"b3e83483",
          5817 => x"3d0d04f9",
          5818 => x"3d0d02a7",
          5819 => x"05335877",
          5820 => x"8a2e0981",
          5821 => x"0687387a",
          5822 => x"528d51eb",
          5823 => x"3f82b3e8",
          5824 => x"337081ff",
          5825 => x"06585687",
          5826 => x"c0948453",
          5827 => x"76802e86",
          5828 => x"3887c094",
          5829 => x"94537208",
          5830 => x"70962a70",
          5831 => x"81065556",
          5832 => x"5472802e",
          5833 => x"8c387391",
          5834 => x"2a708106",
          5835 => x"515372d7",
          5836 => x"38748132",
          5837 => x"70810651",
          5838 => x"5372802e",
          5839 => x"8d387393",
          5840 => x"2a708106",
          5841 => x"515372ff",
          5842 => x"be387581",
          5843 => x"ff065387",
          5844 => x"c0948054",
          5845 => x"72802e86",
          5846 => x"3887c094",
          5847 => x"90547774",
          5848 => x"0c800b82",
          5849 => x"b5c80c89",
          5850 => x"3d0d04f9",
          5851 => x"3d0d7954",
          5852 => x"80743370",
          5853 => x"81ff0653",
          5854 => x"53577077",
          5855 => x"2e80fc38",
          5856 => x"7181ff06",
          5857 => x"811582b3",
          5858 => x"e8337081",
          5859 => x"ff065957",
          5860 => x"555887c0",
          5861 => x"94845175",
          5862 => x"802e8638",
          5863 => x"87c09494",
          5864 => x"51700870",
          5865 => x"962a7081",
          5866 => x"06535452",
          5867 => x"70802e8c",
          5868 => x"3871912a",
          5869 => x"70810651",
          5870 => x"5170d738",
          5871 => x"72813270",
          5872 => x"81065151",
          5873 => x"70802e8d",
          5874 => x"3871932a",
          5875 => x"70810651",
          5876 => x"5170ffbe",
          5877 => x"387481ff",
          5878 => x"065187c0",
          5879 => x"94805270",
          5880 => x"802e8638",
          5881 => x"87c09490",
          5882 => x"5277720c",
          5883 => x"81177433",
          5884 => x"7081ff06",
          5885 => x"53535770",
          5886 => x"ff863876",
          5887 => x"82b5c80c",
          5888 => x"893d0d04",
          5889 => x"fe3d0d82",
          5890 => x"b3e83370",
          5891 => x"81ff0654",
          5892 => x"5287c094",
          5893 => x"84517280",
          5894 => x"2e863887",
          5895 => x"c0949451",
          5896 => x"70087082",
          5897 => x"2a708106",
          5898 => x"51515170",
          5899 => x"802ee238",
          5900 => x"7181ff06",
          5901 => x"5187c094",
          5902 => x"80527080",
          5903 => x"2e863887",
          5904 => x"c0949052",
          5905 => x"71087081",
          5906 => x"ff0682b5",
          5907 => x"c80c5184",
          5908 => x"3d0d04ff",
          5909 => x"af3f82b5",
          5910 => x"c80881ff",
          5911 => x"0682b5c8",
          5912 => x"0c04fe3d",
          5913 => x"0d82b3e8",
          5914 => x"337081ff",
          5915 => x"06525387",
          5916 => x"c0948452",
          5917 => x"70802e86",
          5918 => x"3887c094",
          5919 => x"94527108",
          5920 => x"70822a70",
          5921 => x"81065151",
          5922 => x"51ff5270",
          5923 => x"802ea038",
          5924 => x"7281ff06",
          5925 => x"5187c094",
          5926 => x"80527080",
          5927 => x"2e863887",
          5928 => x"c0949052",
          5929 => x"71087098",
          5930 => x"2b70982c",
          5931 => x"51535171",
          5932 => x"82b5c80c",
          5933 => x"843d0d04",
          5934 => x"ff3d0d87",
          5935 => x"c09e8008",
          5936 => x"709c2a8a",
          5937 => x"06515170",
          5938 => x"802e84b4",
          5939 => x"3887c09e",
          5940 => x"a40882b3",
          5941 => x"ec0c87c0",
          5942 => x"9ea80882",
          5943 => x"b3f00c87",
          5944 => x"c09e9408",
          5945 => x"82b3f40c",
          5946 => x"87c09e98",
          5947 => x"0882b3f8",
          5948 => x"0c87c09e",
          5949 => x"9c0882b3",
          5950 => x"fc0c87c0",
          5951 => x"9ea00882",
          5952 => x"b4800c87",
          5953 => x"c09eac08",
          5954 => x"82b4840c",
          5955 => x"87c09eb0",
          5956 => x"0882b488",
          5957 => x"0c87c09e",
          5958 => x"b40882b4",
          5959 => x"8c0c87c0",
          5960 => x"9eb80882",
          5961 => x"b4900c87",
          5962 => x"c09ebc08",
          5963 => x"82b4940c",
          5964 => x"87c09ec0",
          5965 => x"0882b498",
          5966 => x"0c87c09e",
          5967 => x"c40882b4",
          5968 => x"9c0c87c0",
          5969 => x"9e800851",
          5970 => x"7082b4a0",
          5971 => x"2387c09e",
          5972 => x"840882b4",
          5973 => x"a40c87c0",
          5974 => x"9e880882",
          5975 => x"b4a80c87",
          5976 => x"c09e8c08",
          5977 => x"82b4ac0c",
          5978 => x"810b82b4",
          5979 => x"b034800b",
          5980 => x"87c09e90",
          5981 => x"08708480",
          5982 => x"0a065152",
          5983 => x"5270802e",
          5984 => x"83388152",
          5985 => x"7182b4b1",
          5986 => x"34800b87",
          5987 => x"c09e9008",
          5988 => x"7088800a",
          5989 => x"06515252",
          5990 => x"70802e83",
          5991 => x"38815271",
          5992 => x"82b4b234",
          5993 => x"800b87c0",
          5994 => x"9e900870",
          5995 => x"90800a06",
          5996 => x"51525270",
          5997 => x"802e8338",
          5998 => x"81527182",
          5999 => x"b4b33480",
          6000 => x"0b87c09e",
          6001 => x"90087088",
          6002 => x"80800651",
          6003 => x"52527080",
          6004 => x"2e833881",
          6005 => x"527182b4",
          6006 => x"b434800b",
          6007 => x"87c09e90",
          6008 => x"0870a080",
          6009 => x"80065152",
          6010 => x"5270802e",
          6011 => x"83388152",
          6012 => x"7182b4b5",
          6013 => x"34800b87",
          6014 => x"c09e9008",
          6015 => x"70908080",
          6016 => x"06515252",
          6017 => x"70802e83",
          6018 => x"38815271",
          6019 => x"82b4b634",
          6020 => x"800b87c0",
          6021 => x"9e900870",
          6022 => x"84808006",
          6023 => x"51525270",
          6024 => x"802e8338",
          6025 => x"81527182",
          6026 => x"b4b73480",
          6027 => x"0b87c09e",
          6028 => x"90087082",
          6029 => x"80800651",
          6030 => x"52527080",
          6031 => x"2e833881",
          6032 => x"527182b4",
          6033 => x"b834800b",
          6034 => x"87c09e90",
          6035 => x"08708180",
          6036 => x"80065152",
          6037 => x"5270802e",
          6038 => x"83388152",
          6039 => x"7182b4b9",
          6040 => x"34800b87",
          6041 => x"c09e9008",
          6042 => x"7080c080",
          6043 => x"06515252",
          6044 => x"70802e83",
          6045 => x"38815271",
          6046 => x"82b4ba34",
          6047 => x"800b87c0",
          6048 => x"9e900870",
          6049 => x"a0800651",
          6050 => x"52527080",
          6051 => x"2e833881",
          6052 => x"527182b4",
          6053 => x"bb3487c0",
          6054 => x"9e900870",
          6055 => x"98800670",
          6056 => x"8a2a5151",
          6057 => x"517082b4",
          6058 => x"bc34800b",
          6059 => x"87c09e90",
          6060 => x"08708480",
          6061 => x"06515252",
          6062 => x"70802e83",
          6063 => x"38815271",
          6064 => x"82b4bd34",
          6065 => x"87c09e90",
          6066 => x"087083f0",
          6067 => x"0670842a",
          6068 => x"51515170",
          6069 => x"82b4be34",
          6070 => x"800b87c0",
          6071 => x"9e900870",
          6072 => x"88065152",
          6073 => x"5270802e",
          6074 => x"83388152",
          6075 => x"7182b4bf",
          6076 => x"3487c09e",
          6077 => x"90087087",
          6078 => x"06515170",
          6079 => x"82b4c034",
          6080 => x"833d0d04",
          6081 => x"fb3d0d82",
          6082 => x"a58051ff",
          6083 => x"b1d53f82",
          6084 => x"b4b03354",
          6085 => x"73802e89",
          6086 => x"3882a594",
          6087 => x"51ffb1c3",
          6088 => x"3f82a5a8",
          6089 => x"51ffb1bb",
          6090 => x"3f82b4b2",
          6091 => x"33547380",
          6092 => x"2e943882",
          6093 => x"b48c0882",
          6094 => x"b4900811",
          6095 => x"545282a5",
          6096 => x"c051ff95",
          6097 => x"933f82b4",
          6098 => x"b7335473",
          6099 => x"802e9438",
          6100 => x"82b48408",
          6101 => x"82b48808",
          6102 => x"11545282",
          6103 => x"a5dc51ff",
          6104 => x"94f63f82",
          6105 => x"b4b43354",
          6106 => x"73802e94",
          6107 => x"3882b3ec",
          6108 => x"0882b3f0",
          6109 => x"08115452",
          6110 => x"82a5f851",
          6111 => x"ff94d93f",
          6112 => x"82b4b533",
          6113 => x"5473802e",
          6114 => x"943882b3",
          6115 => x"f40882b3",
          6116 => x"f8081154",
          6117 => x"5282a694",
          6118 => x"51ff94bc",
          6119 => x"3f82b4b6",
          6120 => x"33547380",
          6121 => x"2e943882",
          6122 => x"b3fc0882",
          6123 => x"b4800811",
          6124 => x"545282a6",
          6125 => x"b051ff94",
          6126 => x"9f3f82b4",
          6127 => x"bb335473",
          6128 => x"802e8e38",
          6129 => x"82b4bc33",
          6130 => x"5282a6cc",
          6131 => x"51ff9488",
          6132 => x"3f82b4bf",
          6133 => x"33547380",
          6134 => x"2e8e3882",
          6135 => x"b4c03352",
          6136 => x"82a6ec51",
          6137 => x"ff93f13f",
          6138 => x"82b4bd33",
          6139 => x"5473802e",
          6140 => x"8e3882b4",
          6141 => x"be335282",
          6142 => x"a78c51ff",
          6143 => x"93da3f82",
          6144 => x"b4b13354",
          6145 => x"73802e89",
          6146 => x"3882a7ac",
          6147 => x"51ffafd3",
          6148 => x"3f82b4b3",
          6149 => x"33547380",
          6150 => x"2e893882",
          6151 => x"a7c051ff",
          6152 => x"afc13f82",
          6153 => x"b4b83354",
          6154 => x"73802e89",
          6155 => x"3882a7cc",
          6156 => x"51ffafaf",
          6157 => x"3f82b4b9",
          6158 => x"33547380",
          6159 => x"2e893882",
          6160 => x"a7d851ff",
          6161 => x"af9d3f82",
          6162 => x"b4ba3354",
          6163 => x"73802e89",
          6164 => x"3882a7e4",
          6165 => x"51ffaf8b",
          6166 => x"3f82a7f0",
          6167 => x"51ffaf83",
          6168 => x"3f82b494",
          6169 => x"085282a7",
          6170 => x"fc51ff92",
          6171 => x"eb3f82b4",
          6172 => x"98085282",
          6173 => x"a8a451ff",
          6174 => x"92de3f82",
          6175 => x"b49c0852",
          6176 => x"82a8cc51",
          6177 => x"ff92d13f",
          6178 => x"82a8f451",
          6179 => x"ffaed43f",
          6180 => x"82b4a022",
          6181 => x"5282a8fc",
          6182 => x"51ff92bc",
          6183 => x"3f82b4a4",
          6184 => x"0856bd84",
          6185 => x"c0527551",
          6186 => x"c5d93f82",
          6187 => x"b5c808bd",
          6188 => x"84c02976",
          6189 => x"71315454",
          6190 => x"82b5c808",
          6191 => x"5282a9a4",
          6192 => x"51ff9294",
          6193 => x"3f82b4b7",
          6194 => x"33547380",
          6195 => x"2ea93882",
          6196 => x"b4a80856",
          6197 => x"bd84c052",
          6198 => x"7551c5a7",
          6199 => x"3f82b5c8",
          6200 => x"08bd84c0",
          6201 => x"29767131",
          6202 => x"545482b5",
          6203 => x"c8085282",
          6204 => x"a9d051ff",
          6205 => x"91e23f82",
          6206 => x"b4b23354",
          6207 => x"73802ea9",
          6208 => x"3882b4ac",
          6209 => x"0856bd84",
          6210 => x"c0527551",
          6211 => x"c4f53f82",
          6212 => x"b5c808bd",
          6213 => x"84c02976",
          6214 => x"71315454",
          6215 => x"82b5c808",
          6216 => x"5282a9fc",
          6217 => x"51ff91b0",
          6218 => x"3f82a2bc",
          6219 => x"51ffadb3",
          6220 => x"3f873d0d",
          6221 => x"04fe3d0d",
          6222 => x"02920533",
          6223 => x"ff055271",
          6224 => x"8426aa38",
          6225 => x"71842982",
          6226 => x"95f80552",
          6227 => x"71080482",
          6228 => x"aaa8519d",
          6229 => x"3982aab0",
          6230 => x"51973982",
          6231 => x"aab85191",
          6232 => x"3982aac0",
          6233 => x"518b3982",
          6234 => x"aac45185",
          6235 => x"3982aacc",
          6236 => x"51ffacef",
          6237 => x"3f843d0d",
          6238 => x"04718880",
          6239 => x"0c04800b",
          6240 => x"87c09684",
          6241 => x"0c0482b4",
          6242 => x"c40887c0",
          6243 => x"96840c04",
          6244 => x"fd3d0d76",
          6245 => x"982b7098",
          6246 => x"2c79982b",
          6247 => x"70982c72",
          6248 => x"10137082",
          6249 => x"2b515351",
          6250 => x"54515180",
          6251 => x"0b82aad8",
          6252 => x"12335553",
          6253 => x"7174259c",
          6254 => x"3882aad4",
          6255 => x"11081202",
          6256 => x"84059705",
          6257 => x"33713352",
          6258 => x"52527072",
          6259 => x"2e098106",
          6260 => x"83388153",
          6261 => x"7282b5c8",
          6262 => x"0c853d0d",
          6263 => x"04fb3d0d",
          6264 => x"79028405",
          6265 => x"a3053371",
          6266 => x"33555654",
          6267 => x"72802eb1",
          6268 => x"3882cd9c",
          6269 => x"08528851",
          6270 => x"ffafb73f",
          6271 => x"82cd9c08",
          6272 => x"52a051ff",
          6273 => x"afac3f82",
          6274 => x"cd9c0852",
          6275 => x"8851ffaf",
          6276 => x"a13f7333",
          6277 => x"ff055372",
          6278 => x"74347281",
          6279 => x"ff0653cc",
          6280 => x"397751ff",
          6281 => x"8fb23f74",
          6282 => x"7434873d",
          6283 => x"0d04f63d",
          6284 => x"0d7c0284",
          6285 => x"05b70533",
          6286 => x"028805bb",
          6287 => x"053382b5",
          6288 => x"a0337084",
          6289 => x"2982b4c8",
          6290 => x"05700851",
          6291 => x"59595a58",
          6292 => x"5974802e",
          6293 => x"86387451",
          6294 => x"9afa3f82",
          6295 => x"b5a03370",
          6296 => x"842982b4",
          6297 => x"c8058119",
          6298 => x"70545856",
          6299 => x"5a9dfb3f",
          6300 => x"82b5c808",
          6301 => x"750c82b5",
          6302 => x"a0337084",
          6303 => x"2982b4c8",
          6304 => x"05700851",
          6305 => x"565a7480",
          6306 => x"2ea73875",
          6307 => x"53785274",
          6308 => x"51ffb8d1",
          6309 => x"3f82b5a0",
          6310 => x"33810555",
          6311 => x"7482b5a0",
          6312 => x"347481ff",
          6313 => x"06559375",
          6314 => x"27873880",
          6315 => x"0b82b5a0",
          6316 => x"3477802e",
          6317 => x"b63882b5",
          6318 => x"9c085675",
          6319 => x"802eac38",
          6320 => x"82b59833",
          6321 => x"5574a438",
          6322 => x"8c3dfc05",
          6323 => x"54765378",
          6324 => x"52755180",
          6325 => x"da883f82",
          6326 => x"b59c0852",
          6327 => x"8a51818f",
          6328 => x"953f82b5",
          6329 => x"9c085180",
          6330 => x"dde53f8c",
          6331 => x"3d0d04fd",
          6332 => x"3d0d82b4",
          6333 => x"c8539354",
          6334 => x"72085271",
          6335 => x"802e8938",
          6336 => x"715199d0",
          6337 => x"3f80730c",
          6338 => x"ff148414",
          6339 => x"54547380",
          6340 => x"25e63880",
          6341 => x"0b82b5a0",
          6342 => x"3482b59c",
          6343 => x"08527180",
          6344 => x"2e953871",
          6345 => x"5180dec5",
          6346 => x"3f82b59c",
          6347 => x"085199a4",
          6348 => x"3f800b82",
          6349 => x"b59c0c85",
          6350 => x"3d0d04dc",
          6351 => x"3d0d8157",
          6352 => x"805282b5",
          6353 => x"9c085180",
          6354 => x"e3b23f82",
          6355 => x"b5c80880",
          6356 => x"d33882b5",
          6357 => x"9c085380",
          6358 => x"f852883d",
          6359 => x"70525681",
          6360 => x"8c803f82",
          6361 => x"b5c80880",
          6362 => x"2eba3875",
          6363 => x"51ffb595",
          6364 => x"3f82b5c8",
          6365 => x"0855800b",
          6366 => x"82b5c808",
          6367 => x"259d3882",
          6368 => x"b5c808ff",
          6369 => x"05701755",
          6370 => x"55807434",
          6371 => x"75537652",
          6372 => x"811782ad",
          6373 => x"c85257ff",
          6374 => x"8cbe3f74",
          6375 => x"ff2e0981",
          6376 => x"06ffaf38",
          6377 => x"a63d0d04",
          6378 => x"d93d0daa",
          6379 => x"3d08ad3d",
          6380 => x"085a5a81",
          6381 => x"70585880",
          6382 => x"5282b59c",
          6383 => x"085180e2",
          6384 => x"bb3f82b5",
          6385 => x"c8088195",
          6386 => x"38ff0b82",
          6387 => x"b59c0854",
          6388 => x"5580f852",
          6389 => x"8b3d7052",
          6390 => x"56818b86",
          6391 => x"3f82b5c8",
          6392 => x"08802ea5",
          6393 => x"387551ff",
          6394 => x"b49b3f82",
          6395 => x"b5c80881",
          6396 => x"18585580",
          6397 => x"0b82b5c8",
          6398 => x"08258e38",
          6399 => x"82b5c808",
          6400 => x"ff057017",
          6401 => x"55558074",
          6402 => x"34740970",
          6403 => x"30707207",
          6404 => x"9f2a5155",
          6405 => x"5578772e",
          6406 => x"853873ff",
          6407 => x"ac3882b5",
          6408 => x"9c088c11",
          6409 => x"08535180",
          6410 => x"e1d23f82",
          6411 => x"b5c80880",
          6412 => x"2e893882",
          6413 => x"add451ff",
          6414 => x"8b9e3f78",
          6415 => x"772e0981",
          6416 => x"069b3875",
          6417 => x"527951ff",
          6418 => x"b4a93f79",
          6419 => x"51ffb3b5",
          6420 => x"3fab3d08",
          6421 => x"5482b5c8",
          6422 => x"08743480",
          6423 => x"587782b5",
          6424 => x"c80ca93d",
          6425 => x"0d04f63d",
          6426 => x"0d7c7e71",
          6427 => x"5c717233",
          6428 => x"57595a58",
          6429 => x"73a02e09",
          6430 => x"8106a238",
          6431 => x"78337805",
          6432 => x"56777627",
          6433 => x"98388117",
          6434 => x"705b7071",
          6435 => x"33565855",
          6436 => x"73a02e09",
          6437 => x"81068638",
          6438 => x"757526ea",
          6439 => x"38805473",
          6440 => x"882982b5",
          6441 => x"a4057008",
          6442 => x"5255ffb2",
          6443 => x"d83f82b5",
          6444 => x"c8085379",
          6445 => x"52740851",
          6446 => x"ffb5d73f",
          6447 => x"82b5c808",
          6448 => x"80c53884",
          6449 => x"15335574",
          6450 => x"812e8838",
          6451 => x"74822e88",
          6452 => x"38b539fc",
          6453 => x"e63fac39",
          6454 => x"811a5a8c",
          6455 => x"3dfc1153",
          6456 => x"f80551c5",
          6457 => x"e73f82b5",
          6458 => x"c808802e",
          6459 => x"9a38ff1b",
          6460 => x"53785277",
          6461 => x"51fdb13f",
          6462 => x"82b5c808",
          6463 => x"81ff0655",
          6464 => x"74853874",
          6465 => x"54913981",
          6466 => x"147081ff",
          6467 => x"06515482",
          6468 => x"7427ff8b",
          6469 => x"38805473",
          6470 => x"82b5c80c",
          6471 => x"8c3d0d04",
          6472 => x"d33d0db0",
          6473 => x"3d08b23d",
          6474 => x"08b43d08",
          6475 => x"595f5a80",
          6476 => x"0baf3d34",
          6477 => x"82b5a033",
          6478 => x"82b59c08",
          6479 => x"555b7381",
          6480 => x"cb387382",
          6481 => x"b5983355",
          6482 => x"55738338",
          6483 => x"81557680",
          6484 => x"2e81bc38",
          6485 => x"81707606",
          6486 => x"55567380",
          6487 => x"2e81ad38",
          6488 => x"a8519886",
          6489 => x"3f82b5c8",
          6490 => x"0882b59c",
          6491 => x"0c82b5c8",
          6492 => x"08802e81",
          6493 => x"92389353",
          6494 => x"765282b5",
          6495 => x"c8085180",
          6496 => x"ccfa3f82",
          6497 => x"b5c80880",
          6498 => x"2e8c3882",
          6499 => x"ae8051ff",
          6500 => x"a4d13f80",
          6501 => x"f73982b5",
          6502 => x"c8085b82",
          6503 => x"b59c0853",
          6504 => x"80f85290",
          6505 => x"3d705254",
          6506 => x"8187b73f",
          6507 => x"82b5c808",
          6508 => x"5682b5c8",
          6509 => x"08742e09",
          6510 => x"810680d0",
          6511 => x"3882b5c8",
          6512 => x"0851ffb0",
          6513 => x"c03f82b5",
          6514 => x"c8085580",
          6515 => x"0b82b5c8",
          6516 => x"0825a938",
          6517 => x"82b5c808",
          6518 => x"ff057017",
          6519 => x"55558074",
          6520 => x"34805374",
          6521 => x"81ff0652",
          6522 => x"7551f8c2",
          6523 => x"3f811b70",
          6524 => x"81ff065c",
          6525 => x"54937b27",
          6526 => x"8338805b",
          6527 => x"74ff2e09",
          6528 => x"8106ff97",
          6529 => x"38863975",
          6530 => x"82b59834",
          6531 => x"768c3882",
          6532 => x"b59c0880",
          6533 => x"2e8438f9",
          6534 => x"d63f8f3d",
          6535 => x"5decc33f",
          6536 => x"82b5c808",
          6537 => x"982b7098",
          6538 => x"2c515978",
          6539 => x"ff2eee38",
          6540 => x"7881ff06",
          6541 => x"82ccf433",
          6542 => x"70982b70",
          6543 => x"982c82cc",
          6544 => x"f0337098",
          6545 => x"2b70972c",
          6546 => x"71982c05",
          6547 => x"70842982",
          6548 => x"aad40570",
          6549 => x"08157033",
          6550 => x"51515151",
          6551 => x"59595159",
          6552 => x"5d588156",
          6553 => x"73782e80",
          6554 => x"e9387774",
          6555 => x"27b43874",
          6556 => x"81800a29",
          6557 => x"81ff0a05",
          6558 => x"70982c51",
          6559 => x"55807524",
          6560 => x"80ce3876",
          6561 => x"53745277",
          6562 => x"51f6853f",
          6563 => x"82b5c808",
          6564 => x"81ff0654",
          6565 => x"73802ed7",
          6566 => x"387482cc",
          6567 => x"f0348156",
          6568 => x"b1397481",
          6569 => x"800a2981",
          6570 => x"800a0570",
          6571 => x"982c7081",
          6572 => x"ff065651",
          6573 => x"55739526",
          6574 => x"97387653",
          6575 => x"74527751",
          6576 => x"f5ce3f82",
          6577 => x"b5c80881",
          6578 => x"ff065473",
          6579 => x"cc38d339",
          6580 => x"80567580",
          6581 => x"2e80ca38",
          6582 => x"811c5574",
          6583 => x"82ccf434",
          6584 => x"74982b70",
          6585 => x"982c82cc",
          6586 => x"f0337098",
          6587 => x"2b70982c",
          6588 => x"70101170",
          6589 => x"822b82aa",
          6590 => x"d811335e",
          6591 => x"51515157",
          6592 => x"58515574",
          6593 => x"772e0981",
          6594 => x"06fe9238",
          6595 => x"82aadc14",
          6596 => x"087d0c80",
          6597 => x"0b82ccf4",
          6598 => x"34800b82",
          6599 => x"ccf03492",
          6600 => x"397582cc",
          6601 => x"f4347582",
          6602 => x"ccf03478",
          6603 => x"af3d3475",
          6604 => x"7d0c7e54",
          6605 => x"739526fd",
          6606 => x"e1387384",
          6607 => x"2982968c",
          6608 => x"05547308",
          6609 => x"0482ccfc",
          6610 => x"3354737e",
          6611 => x"2efdcb38",
          6612 => x"82ccf833",
          6613 => x"55737527",
          6614 => x"ab387498",
          6615 => x"2b70982c",
          6616 => x"51557375",
          6617 => x"249e3874",
          6618 => x"1a547333",
          6619 => x"81153474",
          6620 => x"81800a29",
          6621 => x"81ff0a05",
          6622 => x"70982c82",
          6623 => x"ccfc3356",
          6624 => x"5155df39",
          6625 => x"82ccfc33",
          6626 => x"81115654",
          6627 => x"7482ccfc",
          6628 => x"34731a54",
          6629 => x"ae3d3374",
          6630 => x"3482ccf8",
          6631 => x"3354737e",
          6632 => x"25893881",
          6633 => x"14547382",
          6634 => x"ccf83482",
          6635 => x"ccfc3370",
          6636 => x"81800a29",
          6637 => x"81ff0a05",
          6638 => x"70982c82",
          6639 => x"ccf8335a",
          6640 => x"51565674",
          6641 => x"7725a838",
          6642 => x"82cd9c08",
          6643 => x"52741a70",
          6644 => x"335254ff",
          6645 => x"a3dc3f74",
          6646 => x"81800a29",
          6647 => x"81800a05",
          6648 => x"70982c82",
          6649 => x"ccf83356",
          6650 => x"51557375",
          6651 => x"24da3882",
          6652 => x"ccfc3370",
          6653 => x"982b7098",
          6654 => x"2c82ccf8",
          6655 => x"335a5156",
          6656 => x"56747725",
          6657 => x"fc943882",
          6658 => x"cd9c0852",
          6659 => x"8851ffa3",
          6660 => x"a13f7481",
          6661 => x"800a2981",
          6662 => x"800a0570",
          6663 => x"982c82cc",
          6664 => x"f8335651",
          6665 => x"55737524",
          6666 => x"de38fbee",
          6667 => x"39837a34",
          6668 => x"800b811b",
          6669 => x"3482ccfc",
          6670 => x"53805282",
          6671 => x"9ec851f3",
          6672 => x"9c3f81fd",
          6673 => x"3982ccfc",
          6674 => x"337081ff",
          6675 => x"06555573",
          6676 => x"802efbc6",
          6677 => x"3882ccf8",
          6678 => x"33ff0554",
          6679 => x"7382ccf8",
          6680 => x"34ff1554",
          6681 => x"7382ccfc",
          6682 => x"3482cd9c",
          6683 => x"08528851",
          6684 => x"ffa2bf3f",
          6685 => x"82ccfc33",
          6686 => x"70982b70",
          6687 => x"982c82cc",
          6688 => x"f8335751",
          6689 => x"56577474",
          6690 => x"25ad3874",
          6691 => x"1a548114",
          6692 => x"33743482",
          6693 => x"cd9c0852",
          6694 => x"733351ff",
          6695 => x"a2943f74",
          6696 => x"81800a29",
          6697 => x"81800a05",
          6698 => x"70982c82",
          6699 => x"ccf83358",
          6700 => x"51557575",
          6701 => x"24d53882",
          6702 => x"cd9c0852",
          6703 => x"a051ffa1",
          6704 => x"f13f82cc",
          6705 => x"fc337098",
          6706 => x"2b70982c",
          6707 => x"82ccf833",
          6708 => x"57515657",
          6709 => x"747424fa",
          6710 => x"c13882cd",
          6711 => x"9c085288",
          6712 => x"51ffa1ce",
          6713 => x"3f748180",
          6714 => x"0a298180",
          6715 => x"0a057098",
          6716 => x"2c82ccf8",
          6717 => x"33585155",
          6718 => x"757525de",
          6719 => x"38fa9b39",
          6720 => x"82ccf833",
          6721 => x"7a055480",
          6722 => x"743482cd",
          6723 => x"9c08528a",
          6724 => x"51ffa19e",
          6725 => x"3f82ccf8",
          6726 => x"527951f6",
          6727 => x"c93f82b5",
          6728 => x"c80881ff",
          6729 => x"06547396",
          6730 => x"3882ccf8",
          6731 => x"33547380",
          6732 => x"2e8f3881",
          6733 => x"53735279",
          6734 => x"51f1f33f",
          6735 => x"8439807a",
          6736 => x"34800b82",
          6737 => x"ccfc3480",
          6738 => x"0b82ccf8",
          6739 => x"347982b5",
          6740 => x"c80caf3d",
          6741 => x"0d0482cc",
          6742 => x"fc335473",
          6743 => x"802ef9ba",
          6744 => x"3882cd9c",
          6745 => x"08528851",
          6746 => x"ffa0c73f",
          6747 => x"82ccfc33",
          6748 => x"ff055473",
          6749 => x"82ccfc34",
          6750 => x"7381ff06",
          6751 => x"54dd3982",
          6752 => x"ccfc3382",
          6753 => x"ccf83355",
          6754 => x"5573752e",
          6755 => x"f98c38ff",
          6756 => x"14547382",
          6757 => x"ccf83474",
          6758 => x"982b7098",
          6759 => x"2c7581ff",
          6760 => x"06565155",
          6761 => x"747425ad",
          6762 => x"38741a54",
          6763 => x"81143374",
          6764 => x"3482cd9c",
          6765 => x"08527333",
          6766 => x"51ff9ff6",
          6767 => x"3f748180",
          6768 => x"0a298180",
          6769 => x"0a057098",
          6770 => x"2c82ccf8",
          6771 => x"33585155",
          6772 => x"757524d5",
          6773 => x"3882cd9c",
          6774 => x"0852a051",
          6775 => x"ff9fd33f",
          6776 => x"82ccfc33",
          6777 => x"70982b70",
          6778 => x"982c82cc",
          6779 => x"f8335751",
          6780 => x"56577474",
          6781 => x"24f8a338",
          6782 => x"82cd9c08",
          6783 => x"528851ff",
          6784 => x"9fb03f74",
          6785 => x"81800a29",
          6786 => x"81800a05",
          6787 => x"70982c82",
          6788 => x"ccf83358",
          6789 => x"51557575",
          6790 => x"25de38f7",
          6791 => x"fd3982cc",
          6792 => x"fc337081",
          6793 => x"ff0682cc",
          6794 => x"f8335956",
          6795 => x"54747727",
          6796 => x"f7e83882",
          6797 => x"cd9c0852",
          6798 => x"81145473",
          6799 => x"82ccfc34",
          6800 => x"741a7033",
          6801 => x"5254ff9e",
          6802 => x"e93f82cc",
          6803 => x"fc337081",
          6804 => x"ff0682cc",
          6805 => x"f8335856",
          6806 => x"54757526",
          6807 => x"d638f7ba",
          6808 => x"3982ccfc",
          6809 => x"53805282",
          6810 => x"9ec851ee",
          6811 => x"f03f800b",
          6812 => x"82ccfc34",
          6813 => x"800b82cc",
          6814 => x"f834f79e",
          6815 => x"397ab038",
          6816 => x"82b59408",
          6817 => x"5574802e",
          6818 => x"a6387451",
          6819 => x"ffa6f63f",
          6820 => x"82b5c808",
          6821 => x"82ccf834",
          6822 => x"82b5c808",
          6823 => x"81ff0681",
          6824 => x"05537452",
          6825 => x"7951ffa8",
          6826 => x"bc3f935b",
          6827 => x"81c0397a",
          6828 => x"842982b4",
          6829 => x"c805fc11",
          6830 => x"08565474",
          6831 => x"802ea738",
          6832 => x"7451ffa6",
          6833 => x"c03f82b5",
          6834 => x"c80882cc",
          6835 => x"f83482b5",
          6836 => x"c80881ff",
          6837 => x"06810553",
          6838 => x"74527951",
          6839 => x"ffa8863f",
          6840 => x"ff1b5480",
          6841 => x"fa397308",
          6842 => x"5574802e",
          6843 => x"f6ac3874",
          6844 => x"51ffa691",
          6845 => x"3f99397a",
          6846 => x"932e0981",
          6847 => x"06ae3882",
          6848 => x"b4c80855",
          6849 => x"74802ea4",
          6850 => x"387451ff",
          6851 => x"a5f73f82",
          6852 => x"b5c80882",
          6853 => x"ccf83482",
          6854 => x"b5c80881",
          6855 => x"ff068105",
          6856 => x"53745279",
          6857 => x"51ffa7bd",
          6858 => x"3f80c339",
          6859 => x"7a842982",
          6860 => x"b4cc0570",
          6861 => x"08565474",
          6862 => x"802eab38",
          6863 => x"7451ffa5",
          6864 => x"c43f82b5",
          6865 => x"c80882cc",
          6866 => x"f83482b5",
          6867 => x"c80881ff",
          6868 => x"06810553",
          6869 => x"74527951",
          6870 => x"ffa78a3f",
          6871 => x"811b5473",
          6872 => x"81ff065b",
          6873 => x"89397482",
          6874 => x"ccf83474",
          6875 => x"7a3482cc",
          6876 => x"fc5382cc",
          6877 => x"f8335279",
          6878 => x"51ece23f",
          6879 => x"f59c3982",
          6880 => x"ccfc3370",
          6881 => x"81ff0682",
          6882 => x"ccf83359",
          6883 => x"56547477",
          6884 => x"27f58738",
          6885 => x"82cd9c08",
          6886 => x"52811454",
          6887 => x"7382ccfc",
          6888 => x"34741a70",
          6889 => x"335254ff",
          6890 => x"9c883ff4",
          6891 => x"ed3982cc",
          6892 => x"fc335473",
          6893 => x"802ef4e2",
          6894 => x"3882cd9c",
          6895 => x"08528851",
          6896 => x"ff9bef3f",
          6897 => x"82ccfc33",
          6898 => x"ff055473",
          6899 => x"82ccfc34",
          6900 => x"f4c839f9",
          6901 => x"3d0d83bf",
          6902 => x"f40b82b5",
          6903 => x"c00c8480",
          6904 => x"0b82b5bc",
          6905 => x"23a08053",
          6906 => x"805283bf",
          6907 => x"f451ffaa",
          6908 => x"f53f82b5",
          6909 => x"c0085480",
          6910 => x"58777434",
          6911 => x"81577681",
          6912 => x"153482b5",
          6913 => x"c0085477",
          6914 => x"84153476",
          6915 => x"85153482",
          6916 => x"b5c00854",
          6917 => x"77861534",
          6918 => x"76871534",
          6919 => x"82b5c008",
          6920 => x"82b5bc22",
          6921 => x"ff05fe80",
          6922 => x"80077083",
          6923 => x"ffff0670",
          6924 => x"882a5851",
          6925 => x"55567488",
          6926 => x"17347389",
          6927 => x"173482b5",
          6928 => x"bc227088",
          6929 => x"2982b5c0",
          6930 => x"0805f811",
          6931 => x"51555577",
          6932 => x"82153476",
          6933 => x"83153489",
          6934 => x"3d0d04ff",
          6935 => x"3d0d7352",
          6936 => x"81518472",
          6937 => x"278f38fb",
          6938 => x"12832a82",
          6939 => x"117083ff",
          6940 => x"ff065151",
          6941 => x"517082b5",
          6942 => x"c80c833d",
          6943 => x"0d04f93d",
          6944 => x"0d02a605",
          6945 => x"22028405",
          6946 => x"aa052271",
          6947 => x"0582b5c0",
          6948 => x"0871832b",
          6949 => x"71117483",
          6950 => x"2b731170",
          6951 => x"33811233",
          6952 => x"71882b07",
          6953 => x"02a405ae",
          6954 => x"05227181",
          6955 => x"ffff0607",
          6956 => x"70882a53",
          6957 => x"51525954",
          6958 => x"5b5b5753",
          6959 => x"54557177",
          6960 => x"34708118",
          6961 => x"3482b5c0",
          6962 => x"08147588",
          6963 => x"2a525470",
          6964 => x"82153474",
          6965 => x"83153482",
          6966 => x"b5c00870",
          6967 => x"17703381",
          6968 => x"12337188",
          6969 => x"2b077083",
          6970 => x"2b8ffff8",
          6971 => x"06515256",
          6972 => x"52710573",
          6973 => x"83ffff06",
          6974 => x"70882a54",
          6975 => x"54517182",
          6976 => x"12347281",
          6977 => x"ff065372",
          6978 => x"83123482",
          6979 => x"b5c00816",
          6980 => x"56717634",
          6981 => x"72811734",
          6982 => x"893d0d04",
          6983 => x"fb3d0d82",
          6984 => x"b5c00802",
          6985 => x"84059e05",
          6986 => x"2270832b",
          6987 => x"72118611",
          6988 => x"33871233",
          6989 => x"718b2b71",
          6990 => x"832b0758",
          6991 => x"5b595255",
          6992 => x"52720584",
          6993 => x"12338513",
          6994 => x"3371882b",
          6995 => x"0770882a",
          6996 => x"54565652",
          6997 => x"70841334",
          6998 => x"73851334",
          6999 => x"82b5c008",
          7000 => x"70148411",
          7001 => x"33851233",
          7002 => x"718b2b71",
          7003 => x"832b0756",
          7004 => x"59575272",
          7005 => x"05861233",
          7006 => x"87133371",
          7007 => x"882b0770",
          7008 => x"882a5456",
          7009 => x"56527086",
          7010 => x"13347387",
          7011 => x"133482b5",
          7012 => x"c0081370",
          7013 => x"33811233",
          7014 => x"71882b07",
          7015 => x"7081ffff",
          7016 => x"0670882a",
          7017 => x"53515353",
          7018 => x"53717334",
          7019 => x"70811434",
          7020 => x"873d0d04",
          7021 => x"fa3d0d02",
          7022 => x"a2052282",
          7023 => x"b5c00871",
          7024 => x"832b7111",
          7025 => x"70338112",
          7026 => x"3371882b",
          7027 => x"07708829",
          7028 => x"15703381",
          7029 => x"12337198",
          7030 => x"2b71902b",
          7031 => x"07535f53",
          7032 => x"55525a56",
          7033 => x"57535471",
          7034 => x"802580f6",
          7035 => x"387251fe",
          7036 => x"ab3f82b5",
          7037 => x"c0087016",
          7038 => x"70338112",
          7039 => x"33718b2b",
          7040 => x"71832b07",
          7041 => x"74117033",
          7042 => x"81123371",
          7043 => x"882b0770",
          7044 => x"832b8fff",
          7045 => x"f8065152",
          7046 => x"5451535a",
          7047 => x"58537205",
          7048 => x"74882a54",
          7049 => x"52728213",
          7050 => x"34738313",
          7051 => x"3482b5c0",
          7052 => x"08701670",
          7053 => x"33811233",
          7054 => x"718b2b71",
          7055 => x"832b0756",
          7056 => x"59575572",
          7057 => x"05703381",
          7058 => x"12337188",
          7059 => x"2b077081",
          7060 => x"ffff0670",
          7061 => x"882a5751",
          7062 => x"52585272",
          7063 => x"74347181",
          7064 => x"1534883d",
          7065 => x"0d04fb3d",
          7066 => x"0d82b5c0",
          7067 => x"08028405",
          7068 => x"9e052270",
          7069 => x"832b7211",
          7070 => x"82113383",
          7071 => x"1233718b",
          7072 => x"2b71832b",
          7073 => x"07595b59",
          7074 => x"52565273",
          7075 => x"05713381",
          7076 => x"13337188",
          7077 => x"2b07028c",
          7078 => x"05a20522",
          7079 => x"71077088",
          7080 => x"2a535153",
          7081 => x"53537173",
          7082 => x"34708114",
          7083 => x"3482b5c0",
          7084 => x"08701570",
          7085 => x"33811233",
          7086 => x"718b2b71",
          7087 => x"832b0756",
          7088 => x"59575272",
          7089 => x"05821233",
          7090 => x"83133371",
          7091 => x"882b0770",
          7092 => x"882a5455",
          7093 => x"56527082",
          7094 => x"13347283",
          7095 => x"133482b5",
          7096 => x"c0081482",
          7097 => x"11338312",
          7098 => x"3371882b",
          7099 => x"0782b5c8",
          7100 => x"0c525487",
          7101 => x"3d0d04f7",
          7102 => x"3d0d7b82",
          7103 => x"b5c00831",
          7104 => x"832a7083",
          7105 => x"ffff0670",
          7106 => x"535753fd",
          7107 => x"a73f82b5",
          7108 => x"c0087683",
          7109 => x"2b711182",
          7110 => x"11338312",
          7111 => x"33718b2b",
          7112 => x"71832b07",
          7113 => x"75117033",
          7114 => x"81123371",
          7115 => x"982b7190",
          7116 => x"2b075342",
          7117 => x"4051535b",
          7118 => x"58555954",
          7119 => x"7280258d",
          7120 => x"38828080",
          7121 => x"527551fe",
          7122 => x"9d3f8184",
          7123 => x"39841433",
          7124 => x"85153371",
          7125 => x"8b2b7183",
          7126 => x"2b077611",
          7127 => x"79882a53",
          7128 => x"51555855",
          7129 => x"76861434",
          7130 => x"7581ff06",
          7131 => x"56758714",
          7132 => x"3482b5c0",
          7133 => x"08701984",
          7134 => x"12338513",
          7135 => x"3371882b",
          7136 => x"0770882a",
          7137 => x"54575b56",
          7138 => x"53728416",
          7139 => x"34738516",
          7140 => x"3482b5c0",
          7141 => x"08185380",
          7142 => x"0b861434",
          7143 => x"800b8714",
          7144 => x"3482b5c0",
          7145 => x"08537684",
          7146 => x"14347585",
          7147 => x"143482b5",
          7148 => x"c0081870",
          7149 => x"33811233",
          7150 => x"71882b07",
          7151 => x"70828080",
          7152 => x"0770882a",
          7153 => x"53515556",
          7154 => x"54747434",
          7155 => x"72811534",
          7156 => x"8b3d0d04",
          7157 => x"ff3d0d73",
          7158 => x"5282b5c0",
          7159 => x"088438f7",
          7160 => x"f23f7180",
          7161 => x"2e863871",
          7162 => x"51fe8c3f",
          7163 => x"833d0d04",
          7164 => x"f53d0d80",
          7165 => x"7e5258f8",
          7166 => x"e23f82b5",
          7167 => x"c80883ff",
          7168 => x"ff0682b5",
          7169 => x"c0088411",
          7170 => x"33851233",
          7171 => x"71882b07",
          7172 => x"705f5956",
          7173 => x"585a81ff",
          7174 => x"ff597578",
          7175 => x"2e80cb38",
          7176 => x"75882917",
          7177 => x"70338112",
          7178 => x"3371882b",
          7179 => x"077081ff",
          7180 => x"ff067931",
          7181 => x"7083ffff",
          7182 => x"06707f27",
          7183 => x"52535156",
          7184 => x"59557779",
          7185 => x"278a3873",
          7186 => x"802e8538",
          7187 => x"75785a5b",
          7188 => x"84153385",
          7189 => x"16337188",
          7190 => x"2b075754",
          7191 => x"75c23878",
          7192 => x"81ffff2e",
          7193 => x"85387a79",
          7194 => x"59568076",
          7195 => x"832b82b5",
          7196 => x"c0081170",
          7197 => x"33811233",
          7198 => x"71882b07",
          7199 => x"7081ffff",
          7200 => x"0651525a",
          7201 => x"565c5573",
          7202 => x"752e8338",
          7203 => x"81558054",
          7204 => x"79782681",
          7205 => x"cc387454",
          7206 => x"74802e81",
          7207 => x"c438777a",
          7208 => x"2e098106",
          7209 => x"89387551",
          7210 => x"f8f23f81",
          7211 => x"ac398280",
          7212 => x"80537952",
          7213 => x"7551f7c6",
          7214 => x"3f82b5c0",
          7215 => x"08701c86",
          7216 => x"11338712",
          7217 => x"33718b2b",
          7218 => x"71832b07",
          7219 => x"535a5e55",
          7220 => x"74057a17",
          7221 => x"7083ffff",
          7222 => x"0670882a",
          7223 => x"5c595654",
          7224 => x"78841534",
          7225 => x"7681ff06",
          7226 => x"57768515",
          7227 => x"3482b5c0",
          7228 => x"0875832b",
          7229 => x"7111721e",
          7230 => x"86113387",
          7231 => x"12337188",
          7232 => x"2b077088",
          7233 => x"2a535b5e",
          7234 => x"535a5654",
          7235 => x"73861934",
          7236 => x"75871934",
          7237 => x"82b5c008",
          7238 => x"701c8411",
          7239 => x"33851233",
          7240 => x"718b2b71",
          7241 => x"832b0753",
          7242 => x"5d5a5574",
          7243 => x"05547886",
          7244 => x"15347687",
          7245 => x"153482b5",
          7246 => x"c0087016",
          7247 => x"711d8411",
          7248 => x"33851233",
          7249 => x"71882b07",
          7250 => x"70882a53",
          7251 => x"5a5f5256",
          7252 => x"54738416",
          7253 => x"34758516",
          7254 => x"3482b5c0",
          7255 => x"081b8405",
          7256 => x"547382b5",
          7257 => x"c80c8d3d",
          7258 => x"0d04fe3d",
          7259 => x"0d745282",
          7260 => x"b5c00884",
          7261 => x"38f4dc3f",
          7262 => x"71537180",
          7263 => x"2e8b3871",
          7264 => x"51fced3f",
          7265 => x"82b5c808",
          7266 => x"537282b5",
          7267 => x"c80c843d",
          7268 => x"0d04ee3d",
          7269 => x"0d646640",
          7270 => x"5c807042",
          7271 => x"4082b5c0",
          7272 => x"08602e09",
          7273 => x"81068438",
          7274 => x"f4a93f7b",
          7275 => x"8e387e51",
          7276 => x"ffb83f82",
          7277 => x"b5c80854",
          7278 => x"83c7397e",
          7279 => x"8b387b51",
          7280 => x"fc923f7e",
          7281 => x"5483ba39",
          7282 => x"7e51f58f",
          7283 => x"3f82b5c8",
          7284 => x"0883ffff",
          7285 => x"0682b5c0",
          7286 => x"087d7131",
          7287 => x"832a7083",
          7288 => x"ffff0670",
          7289 => x"832b7311",
          7290 => x"70338112",
          7291 => x"3371882b",
          7292 => x"07707531",
          7293 => x"7083ffff",
          7294 => x"06708829",
          7295 => x"fc057388",
          7296 => x"291a7033",
          7297 => x"81123371",
          7298 => x"882b0770",
          7299 => x"902b5344",
          7300 => x"4e534841",
          7301 => x"525c545b",
          7302 => x"415c565b",
          7303 => x"5b738025",
          7304 => x"8f387681",
          7305 => x"ffff0675",
          7306 => x"317083ff",
          7307 => x"ff064254",
          7308 => x"82163383",
          7309 => x"17337188",
          7310 => x"2b077088",
          7311 => x"291c7033",
          7312 => x"81123371",
          7313 => x"982b7190",
          7314 => x"2b075347",
          7315 => x"45525654",
          7316 => x"7380258b",
          7317 => x"38787531",
          7318 => x"7083ffff",
          7319 => x"06415477",
          7320 => x"7b2781fe",
          7321 => x"38601854",
          7322 => x"737b2e09",
          7323 => x"81068f38",
          7324 => x"7851f6c0",
          7325 => x"3f7a83ff",
          7326 => x"ff065881",
          7327 => x"e5397f8e",
          7328 => x"387a7424",
          7329 => x"89387851",
          7330 => x"f6aa3f81",
          7331 => x"a5397f18",
          7332 => x"557a7524",
          7333 => x"80c83879",
          7334 => x"1d821133",
          7335 => x"83123371",
          7336 => x"882b0753",
          7337 => x"5754f4f4",
          7338 => x"3f805278",
          7339 => x"51f7b73f",
          7340 => x"82b5c808",
          7341 => x"83ffff06",
          7342 => x"7e547c53",
          7343 => x"70832b82",
          7344 => x"b5c00811",
          7345 => x"84055355",
          7346 => x"59ff93cf",
          7347 => x"3f82b5c0",
          7348 => x"08148405",
          7349 => x"7583ffff",
          7350 => x"06595c81",
          7351 => x"85396015",
          7352 => x"547a7424",
          7353 => x"80d43878",
          7354 => x"51f5c93f",
          7355 => x"82b5c008",
          7356 => x"1d821133",
          7357 => x"83123371",
          7358 => x"882b0753",
          7359 => x"4354f49c",
          7360 => x"3f805278",
          7361 => x"51f6df3f",
          7362 => x"82b5c808",
          7363 => x"83ffff06",
          7364 => x"7e547c53",
          7365 => x"70832b82",
          7366 => x"b5c00811",
          7367 => x"84055355",
          7368 => x"59ff92f7",
          7369 => x"3f82b5c0",
          7370 => x"08148405",
          7371 => x"60620519",
          7372 => x"555c7383",
          7373 => x"ffff0658",
          7374 => x"a9397b7f",
          7375 => x"5254f9b0",
          7376 => x"3f82b5c8",
          7377 => x"085c82b5",
          7378 => x"c808802e",
          7379 => x"93387d53",
          7380 => x"735282b5",
          7381 => x"c80851ff",
          7382 => x"978b3f73",
          7383 => x"51f7983f",
          7384 => x"7a587a78",
          7385 => x"27993880",
          7386 => x"537a5278",
          7387 => x"51f28f3f",
          7388 => x"7a19832b",
          7389 => x"82b5c008",
          7390 => x"05840551",
          7391 => x"f6f93f7b",
          7392 => x"547382b5",
          7393 => x"c80c943d",
          7394 => x"0d04fc3d",
          7395 => x"0d777729",
          7396 => x"705254fb",
          7397 => x"d53f82b5",
          7398 => x"c8085582",
          7399 => x"b5c80880",
          7400 => x"2e8e3873",
          7401 => x"53805282",
          7402 => x"b5c80851",
          7403 => x"ff9bb73f",
          7404 => x"7482b5c8",
          7405 => x"0c863d0d",
          7406 => x"04ff3d0d",
          7407 => x"028f0533",
          7408 => x"51815270",
          7409 => x"72268738",
          7410 => x"82b5c411",
          7411 => x"33527182",
          7412 => x"b5c80c83",
          7413 => x"3d0d04fc",
          7414 => x"3d0d029b",
          7415 => x"05330284",
          7416 => x"059f0533",
          7417 => x"56538351",
          7418 => x"72812680",
          7419 => x"e0387284",
          7420 => x"2b87c092",
          7421 => x"8c115351",
          7422 => x"88547480",
          7423 => x"2e843881",
          7424 => x"88547372",
          7425 => x"0c87c092",
          7426 => x"8c115181",
          7427 => x"710c850b",
          7428 => x"87c0988c",
          7429 => x"0c705271",
          7430 => x"08708206",
          7431 => x"51517080",
          7432 => x"2e8a3887",
          7433 => x"c0988c08",
          7434 => x"5170ec38",
          7435 => x"7108fc80",
          7436 => x"80065271",
          7437 => x"923887c0",
          7438 => x"988c0851",
          7439 => x"70802e87",
          7440 => x"387182b5",
          7441 => x"c4143482",
          7442 => x"b5c41333",
          7443 => x"517082b5",
          7444 => x"c80c863d",
          7445 => x"0d04f33d",
          7446 => x"0d606264",
          7447 => x"028c05bf",
          7448 => x"05335740",
          7449 => x"585b8374",
          7450 => x"525afecd",
          7451 => x"3f82b5c8",
          7452 => x"0881067a",
          7453 => x"54527181",
          7454 => x"be387172",
          7455 => x"75842b87",
          7456 => x"c0928011",
          7457 => x"87c0928c",
          7458 => x"1287c092",
          7459 => x"8413415a",
          7460 => x"40575a58",
          7461 => x"850b87c0",
          7462 => x"988c0c76",
          7463 => x"7d0c8476",
          7464 => x"0c750870",
          7465 => x"852a7081",
          7466 => x"06515354",
          7467 => x"71802e8e",
          7468 => x"387b0852",
          7469 => x"717b7081",
          7470 => x"055d3481",
          7471 => x"19598074",
          7472 => x"a2065353",
          7473 => x"71732e83",
          7474 => x"38815378",
          7475 => x"83ff268f",
          7476 => x"3872802e",
          7477 => x"8a3887c0",
          7478 => x"988c0852",
          7479 => x"71c33887",
          7480 => x"c0988c08",
          7481 => x"5271802e",
          7482 => x"87387884",
          7483 => x"802e9938",
          7484 => x"81760c87",
          7485 => x"c0928c15",
          7486 => x"53720870",
          7487 => x"82065152",
          7488 => x"71f738ff",
          7489 => x"1a5a8d39",
          7490 => x"84801781",
          7491 => x"197081ff",
          7492 => x"065a5357",
          7493 => x"79802e90",
          7494 => x"3873fc80",
          7495 => x"80065271",
          7496 => x"87387d78",
          7497 => x"26feed38",
          7498 => x"73fc8080",
          7499 => x"06527180",
          7500 => x"2e833881",
          7501 => x"52715372",
          7502 => x"82b5c80c",
          7503 => x"8f3d0d04",
          7504 => x"f33d0d60",
          7505 => x"6264028c",
          7506 => x"05bf0533",
          7507 => x"5740585b",
          7508 => x"83598074",
          7509 => x"5258fce1",
          7510 => x"3f82b5c8",
          7511 => x"08810679",
          7512 => x"54527178",
          7513 => x"2e098106",
          7514 => x"81b13877",
          7515 => x"74842b87",
          7516 => x"c0928011",
          7517 => x"87c0928c",
          7518 => x"1287c092",
          7519 => x"84134059",
          7520 => x"5f565a85",
          7521 => x"0b87c098",
          7522 => x"8c0c767d",
          7523 => x"0c82760c",
          7524 => x"80587508",
          7525 => x"70842a70",
          7526 => x"81065153",
          7527 => x"5471802e",
          7528 => x"8c387a70",
          7529 => x"81055c33",
          7530 => x"7c0c8118",
          7531 => x"5873812a",
          7532 => x"70810651",
          7533 => x"5271802e",
          7534 => x"8a3887c0",
          7535 => x"988c0852",
          7536 => x"71d03887",
          7537 => x"c0988c08",
          7538 => x"5271802e",
          7539 => x"87387784",
          7540 => x"802e9938",
          7541 => x"81760c87",
          7542 => x"c0928c15",
          7543 => x"53720870",
          7544 => x"82065152",
          7545 => x"71f738ff",
          7546 => x"19598d39",
          7547 => x"811a7081",
          7548 => x"ff068480",
          7549 => x"19595b52",
          7550 => x"78802e90",
          7551 => x"3873fc80",
          7552 => x"80065271",
          7553 => x"87387d7a",
          7554 => x"26fef838",
          7555 => x"73fc8080",
          7556 => x"06527180",
          7557 => x"2e833881",
          7558 => x"52715372",
          7559 => x"82b5c80c",
          7560 => x"8f3d0d04",
          7561 => x"fa3d0d7a",
          7562 => x"028405a3",
          7563 => x"05330288",
          7564 => x"05a70533",
          7565 => x"71545456",
          7566 => x"57fafe3f",
          7567 => x"82b5c808",
          7568 => x"81065383",
          7569 => x"547280fe",
          7570 => x"38850b87",
          7571 => x"c0988c0c",
          7572 => x"81567176",
          7573 => x"2e80dc38",
          7574 => x"71762493",
          7575 => x"3874842b",
          7576 => x"87c0928c",
          7577 => x"11545471",
          7578 => x"802e8d38",
          7579 => x"80d43971",
          7580 => x"832e80c6",
          7581 => x"3880cb39",
          7582 => x"72087081",
          7583 => x"2a708106",
          7584 => x"51515271",
          7585 => x"802e8a38",
          7586 => x"87c0988c",
          7587 => x"085271e8",
          7588 => x"3887c098",
          7589 => x"8c085271",
          7590 => x"96388173",
          7591 => x"0c87c092",
          7592 => x"8c145372",
          7593 => x"08708206",
          7594 => x"515271f7",
          7595 => x"38963980",
          7596 => x"56923988",
          7597 => x"800a770c",
          7598 => x"85398180",
          7599 => x"770c7256",
          7600 => x"83398456",
          7601 => x"75547382",
          7602 => x"b5c80c88",
          7603 => x"3d0d04fe",
          7604 => x"3d0d7481",
          7605 => x"11337133",
          7606 => x"71882b07",
          7607 => x"82b5c80c",
          7608 => x"5351843d",
          7609 => x"0d04fd3d",
          7610 => x"0d758311",
          7611 => x"33821233",
          7612 => x"71902b71",
          7613 => x"882b0781",
          7614 => x"14337072",
          7615 => x"07882b75",
          7616 => x"33710782",
          7617 => x"b5c80c52",
          7618 => x"53545654",
          7619 => x"52853d0d",
          7620 => x"04ff3d0d",
          7621 => x"73028405",
          7622 => x"92052252",
          7623 => x"52707270",
          7624 => x"81055434",
          7625 => x"70882a51",
          7626 => x"70723483",
          7627 => x"3d0d04ff",
          7628 => x"3d0d7375",
          7629 => x"52527072",
          7630 => x"70810554",
          7631 => x"3470882a",
          7632 => x"51707270",
          7633 => x"81055434",
          7634 => x"70882a51",
          7635 => x"70727081",
          7636 => x"05543470",
          7637 => x"882a5170",
          7638 => x"7234833d",
          7639 => x"0d04fe3d",
          7640 => x"0d767577",
          7641 => x"54545170",
          7642 => x"802e9238",
          7643 => x"71708105",
          7644 => x"53337370",
          7645 => x"81055534",
          7646 => x"ff1151eb",
          7647 => x"39843d0d",
          7648 => x"04fe3d0d",
          7649 => x"75777654",
          7650 => x"52537272",
          7651 => x"70810554",
          7652 => x"34ff1151",
          7653 => x"70f43884",
          7654 => x"3d0d04fc",
          7655 => x"3d0d7877",
          7656 => x"79565653",
          7657 => x"74708105",
          7658 => x"56337470",
          7659 => x"81055633",
          7660 => x"717131ff",
          7661 => x"16565252",
          7662 => x"5272802e",
          7663 => x"86387180",
          7664 => x"2ee23871",
          7665 => x"82b5c80c",
          7666 => x"863d0d04",
          7667 => x"fe3d0d74",
          7668 => x"76545189",
          7669 => x"3971732e",
          7670 => x"8a388111",
          7671 => x"51703352",
          7672 => x"71f33870",
          7673 => x"3382b5c8",
          7674 => x"0c843d0d",
          7675 => x"04800b82",
          7676 => x"b5c80c04",
          7677 => x"800b82b5",
          7678 => x"c80c04f7",
          7679 => x"3d0d7b56",
          7680 => x"800b8317",
          7681 => x"33565a74",
          7682 => x"7a2e80d6",
          7683 => x"388154b0",
          7684 => x"160853b4",
          7685 => x"16705381",
          7686 => x"17335259",
          7687 => x"faa23f82",
          7688 => x"b5c8087a",
          7689 => x"2e098106",
          7690 => x"b73882b5",
          7691 => x"c8088317",
          7692 => x"34b01608",
          7693 => x"70a41808",
          7694 => x"319c1808",
          7695 => x"59565874",
          7696 => x"77279f38",
          7697 => x"82163355",
          7698 => x"74822e09",
          7699 => x"81069338",
          7700 => x"81547618",
          7701 => x"53785281",
          7702 => x"163351f9",
          7703 => x"e33f8339",
          7704 => x"815a7982",
          7705 => x"b5c80c8b",
          7706 => x"3d0d04fa",
          7707 => x"3d0d787a",
          7708 => x"56568057",
          7709 => x"74b01708",
          7710 => x"2eaf3875",
          7711 => x"51fefc3f",
          7712 => x"82b5c808",
          7713 => x"5782b5c8",
          7714 => x"089f3881",
          7715 => x"547453b4",
          7716 => x"16528116",
          7717 => x"3351f7be",
          7718 => x"3f82b5c8",
          7719 => x"08802e85",
          7720 => x"38ff5581",
          7721 => x"5774b017",
          7722 => x"0c7682b5",
          7723 => x"c80c883d",
          7724 => x"0d04f83d",
          7725 => x"0d7a7052",
          7726 => x"57fec03f",
          7727 => x"82b5c808",
          7728 => x"5882b5c8",
          7729 => x"08819138",
          7730 => x"76335574",
          7731 => x"832e0981",
          7732 => x"0680f038",
          7733 => x"84173359",
          7734 => x"78812e09",
          7735 => x"810680e3",
          7736 => x"38848053",
          7737 => x"82b5c808",
          7738 => x"52b41770",
          7739 => x"5256fd91",
          7740 => x"3f82d4d5",
          7741 => x"5284b217",
          7742 => x"51fc963f",
          7743 => x"848b85a4",
          7744 => x"d2527551",
          7745 => x"fca93f86",
          7746 => x"8a85e4f2",
          7747 => x"52849817",
          7748 => x"51fc9c3f",
          7749 => x"90170852",
          7750 => x"849c1751",
          7751 => x"fc913f8c",
          7752 => x"17085284",
          7753 => x"a01751fc",
          7754 => x"863fa017",
          7755 => x"08810570",
          7756 => x"b0190c79",
          7757 => x"55537552",
          7758 => x"81173351",
          7759 => x"f8823f77",
          7760 => x"84183480",
          7761 => x"53805281",
          7762 => x"173351f9",
          7763 => x"d73f82b5",
          7764 => x"c808802e",
          7765 => x"83388158",
          7766 => x"7782b5c8",
          7767 => x"0c8a3d0d",
          7768 => x"04fb3d0d",
          7769 => x"77fe1a98",
          7770 => x"1208fe05",
          7771 => x"55565480",
          7772 => x"56747327",
          7773 => x"8d388a14",
          7774 => x"22757129",
          7775 => x"ac160805",
          7776 => x"57537582",
          7777 => x"b5c80c87",
          7778 => x"3d0d04f9",
          7779 => x"3d0d7a7a",
          7780 => x"70085654",
          7781 => x"57817727",
          7782 => x"81df3876",
          7783 => x"98150827",
          7784 => x"81d738ff",
          7785 => x"74335458",
          7786 => x"72822e80",
          7787 => x"f5387282",
          7788 => x"24893872",
          7789 => x"812e8d38",
          7790 => x"81bf3972",
          7791 => x"832e818e",
          7792 => x"3881b639",
          7793 => x"76812a17",
          7794 => x"70892aa4",
          7795 => x"16080553",
          7796 => x"745255fd",
          7797 => x"963f82b5",
          7798 => x"c808819f",
          7799 => x"387483ff",
          7800 => x"0614b411",
          7801 => x"33811770",
          7802 => x"892aa418",
          7803 => x"08055576",
          7804 => x"54575753",
          7805 => x"fcf53f82",
          7806 => x"b5c80880",
          7807 => x"fe387483",
          7808 => x"ff0614b4",
          7809 => x"11337088",
          7810 => x"2b780779",
          7811 => x"81067184",
          7812 => x"2a5c5258",
          7813 => x"51537280",
          7814 => x"e238759f",
          7815 => x"ff065880",
          7816 => x"da397688",
          7817 => x"2aa41508",
          7818 => x"05527351",
          7819 => x"fcbd3f82",
          7820 => x"b5c80880",
          7821 => x"c6387610",
          7822 => x"83fe0674",
          7823 => x"05b40551",
          7824 => x"f98d3f82",
          7825 => x"b5c80883",
          7826 => x"ffff0658",
          7827 => x"ae397687",
          7828 => x"2aa41508",
          7829 => x"05527351",
          7830 => x"fc913f82",
          7831 => x"b5c8089b",
          7832 => x"3876822b",
          7833 => x"83fc0674",
          7834 => x"05b40551",
          7835 => x"f8f83f82",
          7836 => x"b5c808f0",
          7837 => x"0a065883",
          7838 => x"39815877",
          7839 => x"82b5c80c",
          7840 => x"893d0d04",
          7841 => x"f83d0d7a",
          7842 => x"7c7e5a58",
          7843 => x"56825981",
          7844 => x"7727829e",
          7845 => x"38769817",
          7846 => x"08278296",
          7847 => x"38753353",
          7848 => x"72792e81",
          7849 => x"9d387279",
          7850 => x"24893872",
          7851 => x"812e8d38",
          7852 => x"82803972",
          7853 => x"832e81b8",
          7854 => x"3881f739",
          7855 => x"76812a17",
          7856 => x"70892aa4",
          7857 => x"18080553",
          7858 => x"765255fb",
          7859 => x"9e3f82b5",
          7860 => x"c8085982",
          7861 => x"b5c80881",
          7862 => x"d9387483",
          7863 => x"ff0616b4",
          7864 => x"05811678",
          7865 => x"81065956",
          7866 => x"54775376",
          7867 => x"802e8f38",
          7868 => x"77842b9f",
          7869 => x"f0067433",
          7870 => x"8f067107",
          7871 => x"51537274",
          7872 => x"34810b83",
          7873 => x"17347489",
          7874 => x"2aa41708",
          7875 => x"05527551",
          7876 => x"fad93f82",
          7877 => x"b5c80859",
          7878 => x"82b5c808",
          7879 => x"81943874",
          7880 => x"83ff0616",
          7881 => x"b4057884",
          7882 => x"2a545476",
          7883 => x"8f387788",
          7884 => x"2a743381",
          7885 => x"f006718f",
          7886 => x"06075153",
          7887 => x"72743480",
          7888 => x"ec397688",
          7889 => x"2aa41708",
          7890 => x"05527551",
          7891 => x"fa9d3f82",
          7892 => x"b5c80859",
          7893 => x"82b5c808",
          7894 => x"80d83877",
          7895 => x"83ffff06",
          7896 => x"52761083",
          7897 => x"fe067605",
          7898 => x"b40551f7",
          7899 => x"a43fbe39",
          7900 => x"76872aa4",
          7901 => x"17080552",
          7902 => x"7551f9ef",
          7903 => x"3f82b5c8",
          7904 => x"085982b5",
          7905 => x"c808ab38",
          7906 => x"77f00a06",
          7907 => x"77822b83",
          7908 => x"fc067018",
          7909 => x"b4057054",
          7910 => x"515454f6",
          7911 => x"c93f82b5",
          7912 => x"c8088f0a",
          7913 => x"06740752",
          7914 => x"7251f783",
          7915 => x"3f810b83",
          7916 => x"17347882",
          7917 => x"b5c80c8a",
          7918 => x"3d0d04f8",
          7919 => x"3d0d7a7c",
          7920 => x"7e720859",
          7921 => x"56565981",
          7922 => x"7527a438",
          7923 => x"74981708",
          7924 => x"279d3873",
          7925 => x"802eaa38",
          7926 => x"ff537352",
          7927 => x"7551fda4",
          7928 => x"3f82b5c8",
          7929 => x"085482b5",
          7930 => x"c80880f2",
          7931 => x"38933982",
          7932 => x"5480eb39",
          7933 => x"815480e6",
          7934 => x"3982b5c8",
          7935 => x"085480de",
          7936 => x"39745278",
          7937 => x"51fb843f",
          7938 => x"82b5c808",
          7939 => x"5882b5c8",
          7940 => x"08802e80",
          7941 => x"c73882b5",
          7942 => x"c808812e",
          7943 => x"d23882b5",
          7944 => x"c808ff2e",
          7945 => x"cf388053",
          7946 => x"74527551",
          7947 => x"fcd63f82",
          7948 => x"b5c808c5",
          7949 => x"38981608",
          7950 => x"fe119018",
          7951 => x"08575557",
          7952 => x"74742790",
          7953 => x"38811590",
          7954 => x"170c8416",
          7955 => x"33810754",
          7956 => x"73841734",
          7957 => x"77557678",
          7958 => x"26ffa638",
          7959 => x"80547382",
          7960 => x"b5c80c8a",
          7961 => x"3d0d04f6",
          7962 => x"3d0d7c7e",
          7963 => x"7108595b",
          7964 => x"5b799538",
          7965 => x"8c170858",
          7966 => x"77802e88",
          7967 => x"38981708",
          7968 => x"7826b238",
          7969 => x"8158ae39",
          7970 => x"79527a51",
          7971 => x"f9fd3f81",
          7972 => x"557482b5",
          7973 => x"c8082782",
          7974 => x"e03882b5",
          7975 => x"c8085582",
          7976 => x"b5c808ff",
          7977 => x"2e82d238",
          7978 => x"98170882",
          7979 => x"b5c80826",
          7980 => x"82c73879",
          7981 => x"58901708",
          7982 => x"70565473",
          7983 => x"802e82b9",
          7984 => x"38777a2e",
          7985 => x"09810680",
          7986 => x"e238811a",
          7987 => x"56981708",
          7988 => x"76268338",
          7989 => x"82567552",
          7990 => x"7a51f9af",
          7991 => x"3f805982",
          7992 => x"b5c80881",
          7993 => x"2e098106",
          7994 => x"863882b5",
          7995 => x"c8085982",
          7996 => x"b5c80809",
          7997 => x"70307072",
          7998 => x"07802570",
          7999 => x"7c0782b5",
          8000 => x"c8085451",
          8001 => x"51555573",
          8002 => x"81ef3882",
          8003 => x"b5c80880",
          8004 => x"2e95388c",
          8005 => x"17085481",
          8006 => x"74279038",
          8007 => x"73981808",
          8008 => x"27893873",
          8009 => x"58853975",
          8010 => x"80db3877",
          8011 => x"56811656",
          8012 => x"98170876",
          8013 => x"26893882",
          8014 => x"56757826",
          8015 => x"81ac3875",
          8016 => x"527a51f8",
          8017 => x"c63f82b5",
          8018 => x"c808802e",
          8019 => x"b8388059",
          8020 => x"82b5c808",
          8021 => x"812e0981",
          8022 => x"06863882",
          8023 => x"b5c80859",
          8024 => x"82b5c808",
          8025 => x"09703070",
          8026 => x"72078025",
          8027 => x"707c0751",
          8028 => x"51555573",
          8029 => x"80f83875",
          8030 => x"782e0981",
          8031 => x"06ffae38",
          8032 => x"735580f5",
          8033 => x"39ff5375",
          8034 => x"527651f9",
          8035 => x"f73f82b5",
          8036 => x"c80882b5",
          8037 => x"c8083070",
          8038 => x"82b5c808",
          8039 => x"07802551",
          8040 => x"55557980",
          8041 => x"2e943873",
          8042 => x"802e8f38",
          8043 => x"75537952",
          8044 => x"7651f9d0",
          8045 => x"3f82b5c8",
          8046 => x"085574a5",
          8047 => x"38758c18",
          8048 => x"0c981708",
          8049 => x"fe059018",
          8050 => x"08565474",
          8051 => x"74268638",
          8052 => x"ff159018",
          8053 => x"0c841733",
          8054 => x"81075473",
          8055 => x"84183497",
          8056 => x"39ff5674",
          8057 => x"812e9038",
          8058 => x"8c398055",
          8059 => x"8c3982b5",
          8060 => x"c8085585",
          8061 => x"39815675",
          8062 => x"557482b5",
          8063 => x"c80c8c3d",
          8064 => x"0d04f83d",
          8065 => x"0d7a7052",
          8066 => x"55f3f03f",
          8067 => x"82b5c808",
          8068 => x"58815682",
          8069 => x"b5c80880",
          8070 => x"d8387b52",
          8071 => x"7451f6c1",
          8072 => x"3f82b5c8",
          8073 => x"0882b5c8",
          8074 => x"08b0170c",
          8075 => x"59848053",
          8076 => x"7752b415",
          8077 => x"705257f2",
          8078 => x"c83f7756",
          8079 => x"84398116",
          8080 => x"568a1522",
          8081 => x"58757827",
          8082 => x"97388154",
          8083 => x"75195376",
          8084 => x"52811533",
          8085 => x"51ede93f",
          8086 => x"82b5c808",
          8087 => x"802edf38",
          8088 => x"8a152276",
          8089 => x"32703070",
          8090 => x"7207709f",
          8091 => x"2a535156",
          8092 => x"567582b5",
          8093 => x"c80c8a3d",
          8094 => x"0d04f83d",
          8095 => x"0d7a7c71",
          8096 => x"08585657",
          8097 => x"74f0800a",
          8098 => x"2680f138",
          8099 => x"749f0653",
          8100 => x"7280e938",
          8101 => x"7490180c",
          8102 => x"88170854",
          8103 => x"73aa3875",
          8104 => x"33538273",
          8105 => x"278838a8",
          8106 => x"16085473",
          8107 => x"9b387485",
          8108 => x"2a53820b",
          8109 => x"8817225a",
          8110 => x"58727927",
          8111 => x"80fe38a8",
          8112 => x"16089818",
          8113 => x"0c80cd39",
          8114 => x"8a162270",
          8115 => x"892b5458",
          8116 => x"727526b2",
          8117 => x"38735276",
          8118 => x"51f5b03f",
          8119 => x"82b5c808",
          8120 => x"5482b5c8",
          8121 => x"08ff2ebd",
          8122 => x"38810b82",
          8123 => x"b5c80827",
          8124 => x"8b389816",
          8125 => x"0882b5c8",
          8126 => x"08268538",
          8127 => x"8258bd39",
          8128 => x"74733155",
          8129 => x"cb397352",
          8130 => x"7551f4d5",
          8131 => x"3f82b5c8",
          8132 => x"0898180c",
          8133 => x"7394180c",
          8134 => x"98170853",
          8135 => x"82587280",
          8136 => x"2e9a3885",
          8137 => x"39815894",
          8138 => x"3974892a",
          8139 => x"1398180c",
          8140 => x"7483ff06",
          8141 => x"16b4059c",
          8142 => x"180c8058",
          8143 => x"7782b5c8",
          8144 => x"0c8a3d0d",
          8145 => x"04f83d0d",
          8146 => x"7a700890",
          8147 => x"1208a005",
          8148 => x"595754f0",
          8149 => x"800a7727",
          8150 => x"8638800b",
          8151 => x"98150c98",
          8152 => x"14085384",
          8153 => x"5572802e",
          8154 => x"81cb3876",
          8155 => x"83ff0658",
          8156 => x"7781b538",
          8157 => x"81139815",
          8158 => x"0c941408",
          8159 => x"55749238",
          8160 => x"76852a88",
          8161 => x"17225653",
          8162 => x"74732681",
          8163 => x"9b3880c0",
          8164 => x"398a1622",
          8165 => x"ff057789",
          8166 => x"2a065372",
          8167 => x"818a3874",
          8168 => x"527351f3",
          8169 => x"e63f82b5",
          8170 => x"c8085382",
          8171 => x"55810b82",
          8172 => x"b5c80827",
          8173 => x"80ff3881",
          8174 => x"5582b5c8",
          8175 => x"08ff2e80",
          8176 => x"f4389816",
          8177 => x"0882b5c8",
          8178 => x"082680ca",
          8179 => x"387b8a38",
          8180 => x"7798150c",
          8181 => x"845580dd",
          8182 => x"39941408",
          8183 => x"527351f9",
          8184 => x"863f82b5",
          8185 => x"c8085387",
          8186 => x"5582b5c8",
          8187 => x"08802e80",
          8188 => x"c4388255",
          8189 => x"82b5c808",
          8190 => x"812eba38",
          8191 => x"815582b5",
          8192 => x"c808ff2e",
          8193 => x"b03882b5",
          8194 => x"c8085275",
          8195 => x"51fbf33f",
          8196 => x"82b5c808",
          8197 => x"a0387294",
          8198 => x"150c7252",
          8199 => x"7551f2c1",
          8200 => x"3f82b5c8",
          8201 => x"0898150c",
          8202 => x"7690150c",
          8203 => x"7716b405",
          8204 => x"9c150c80",
          8205 => x"557482b5",
          8206 => x"c80c8a3d",
          8207 => x"0d04f73d",
          8208 => x"0d7b7d71",
          8209 => x"085b5b57",
          8210 => x"80527651",
          8211 => x"fcac3f82",
          8212 => x"b5c80854",
          8213 => x"82b5c808",
          8214 => x"80ec3882",
          8215 => x"b5c80856",
          8216 => x"98170852",
          8217 => x"7851f083",
          8218 => x"3f82b5c8",
          8219 => x"085482b5",
          8220 => x"c80880d2",
          8221 => x"3882b5c8",
          8222 => x"089c1808",
          8223 => x"70335154",
          8224 => x"587281e5",
          8225 => x"2e098106",
          8226 => x"83388158",
          8227 => x"82b5c808",
          8228 => x"55728338",
          8229 => x"81557775",
          8230 => x"07537280",
          8231 => x"2e8e3881",
          8232 => x"1656757a",
          8233 => x"2e098106",
          8234 => x"8838a539",
          8235 => x"82b5c808",
          8236 => x"56815276",
          8237 => x"51fd8e3f",
          8238 => x"82b5c808",
          8239 => x"5482b5c8",
          8240 => x"08802eff",
          8241 => x"9b387384",
          8242 => x"2e098106",
          8243 => x"83388754",
          8244 => x"7382b5c8",
          8245 => x"0c8b3d0d",
          8246 => x"04fd3d0d",
          8247 => x"769a1152",
          8248 => x"54ebec3f",
          8249 => x"82b5c808",
          8250 => x"83ffff06",
          8251 => x"76703351",
          8252 => x"53537183",
          8253 => x"2e098106",
          8254 => x"90389414",
          8255 => x"51ebd03f",
          8256 => x"82b5c808",
          8257 => x"902b7307",
          8258 => x"537282b5",
          8259 => x"c80c853d",
          8260 => x"0d04fc3d",
          8261 => x"0d777970",
          8262 => x"83ffff06",
          8263 => x"549a1253",
          8264 => x"5555ebed",
          8265 => x"3f767033",
          8266 => x"51537283",
          8267 => x"2e098106",
          8268 => x"8b387390",
          8269 => x"2a529415",
          8270 => x"51ebd63f",
          8271 => x"863d0d04",
          8272 => x"f73d0d7b",
          8273 => x"7d5b5584",
          8274 => x"75085a58",
          8275 => x"98150880",
          8276 => x"2e818a38",
          8277 => x"98150852",
          8278 => x"7851ee8f",
          8279 => x"3f82b5c8",
          8280 => x"085882b5",
          8281 => x"c80880f5",
          8282 => x"389c1508",
          8283 => x"70335553",
          8284 => x"73863884",
          8285 => x"5880e639",
          8286 => x"8b133370",
          8287 => x"bf067081",
          8288 => x"ff065851",
          8289 => x"53728616",
          8290 => x"3482b5c8",
          8291 => x"08537381",
          8292 => x"e52e8338",
          8293 => x"815373ae",
          8294 => x"2ea93881",
          8295 => x"70740654",
          8296 => x"5772802e",
          8297 => x"9e38758f",
          8298 => x"2e993882",
          8299 => x"b5c80876",
          8300 => x"df065454",
          8301 => x"72882e09",
          8302 => x"81068338",
          8303 => x"7654737a",
          8304 => x"2ea03880",
          8305 => x"527451fa",
          8306 => x"fc3f82b5",
          8307 => x"c8085882",
          8308 => x"b5c80889",
          8309 => x"38981508",
          8310 => x"fefa3886",
          8311 => x"39800b98",
          8312 => x"160c7782",
          8313 => x"b5c80c8b",
          8314 => x"3d0d04fb",
          8315 => x"3d0d7770",
          8316 => x"08575481",
          8317 => x"527351fc",
          8318 => x"c53f82b5",
          8319 => x"c8085582",
          8320 => x"b5c808b4",
          8321 => x"38981408",
          8322 => x"527551ec",
          8323 => x"de3f82b5",
          8324 => x"c8085582",
          8325 => x"b5c808a0",
          8326 => x"38a05382",
          8327 => x"b5c80852",
          8328 => x"9c140851",
          8329 => x"eadb3f8b",
          8330 => x"53a01452",
          8331 => x"9c140851",
          8332 => x"eaac3f81",
          8333 => x"0b831734",
          8334 => x"7482b5c8",
          8335 => x"0c873d0d",
          8336 => x"04fd3d0d",
          8337 => x"75700898",
          8338 => x"12085470",
          8339 => x"535553ec",
          8340 => x"9a3f82b5",
          8341 => x"c8088d38",
          8342 => x"9c130853",
          8343 => x"e5733481",
          8344 => x"0b831534",
          8345 => x"853d0d04",
          8346 => x"fa3d0d78",
          8347 => x"7a575780",
          8348 => x"0b891734",
          8349 => x"98170880",
          8350 => x"2e818238",
          8351 => x"80708918",
          8352 => x"5555559c",
          8353 => x"17081470",
          8354 => x"33811656",
          8355 => x"515271a0",
          8356 => x"2ea83871",
          8357 => x"852e0981",
          8358 => x"06843881",
          8359 => x"e5527389",
          8360 => x"2e098106",
          8361 => x"8b38ae73",
          8362 => x"70810555",
          8363 => x"34811555",
          8364 => x"71737081",
          8365 => x"05553481",
          8366 => x"15558a74",
          8367 => x"27c53875",
          8368 => x"15880552",
          8369 => x"800b8113",
          8370 => x"349c1708",
          8371 => x"528b1233",
          8372 => x"8817349c",
          8373 => x"17089c11",
          8374 => x"5252e88a",
          8375 => x"3f82b5c8",
          8376 => x"08760c96",
          8377 => x"1251e7e7",
          8378 => x"3f82b5c8",
          8379 => x"08861723",
          8380 => x"981251e7",
          8381 => x"da3f82b5",
          8382 => x"c8088417",
          8383 => x"23883d0d",
          8384 => x"04f33d0d",
          8385 => x"7f70085e",
          8386 => x"5b806170",
          8387 => x"33515555",
          8388 => x"73af2e83",
          8389 => x"38815573",
          8390 => x"80dc2e91",
          8391 => x"3874802e",
          8392 => x"8c38941d",
          8393 => x"08881c0c",
          8394 => x"aa398115",
          8395 => x"41806170",
          8396 => x"33565656",
          8397 => x"73af2e09",
          8398 => x"81068338",
          8399 => x"81567380",
          8400 => x"dc327030",
          8401 => x"70802578",
          8402 => x"07515154",
          8403 => x"73dc3873",
          8404 => x"881c0c60",
          8405 => x"70335154",
          8406 => x"739f2696",
          8407 => x"38ff800b",
          8408 => x"ab1c3480",
          8409 => x"527a51f6",
          8410 => x"913f82b5",
          8411 => x"c8085585",
          8412 => x"9839913d",
          8413 => x"61a01d5c",
          8414 => x"5a5e8b53",
          8415 => x"a0527951",
          8416 => x"e7ff3f80",
          8417 => x"70595788",
          8418 => x"7933555c",
          8419 => x"73ae2e09",
          8420 => x"810680d4",
          8421 => x"38781870",
          8422 => x"33811a71",
          8423 => x"ae327030",
          8424 => x"709f2a73",
          8425 => x"82260751",
          8426 => x"51535a57",
          8427 => x"54738c38",
          8428 => x"79175475",
          8429 => x"74348117",
          8430 => x"57db3975",
          8431 => x"af327030",
          8432 => x"709f2a51",
          8433 => x"51547580",
          8434 => x"dc2e8c38",
          8435 => x"73802e87",
          8436 => x"3875a026",
          8437 => x"82bd3877",
          8438 => x"197e0ca4",
          8439 => x"54a07627",
          8440 => x"82bd38a0",
          8441 => x"5482b839",
          8442 => x"78187033",
          8443 => x"811a5a57",
          8444 => x"54a07627",
          8445 => x"81fc3875",
          8446 => x"af327030",
          8447 => x"7780dc32",
          8448 => x"70307280",
          8449 => x"25718025",
          8450 => x"07515156",
          8451 => x"51557380",
          8452 => x"2eac3884",
          8453 => x"39811858",
          8454 => x"80781a70",
          8455 => x"33515555",
          8456 => x"73af2e09",
          8457 => x"81068338",
          8458 => x"81557380",
          8459 => x"dc327030",
          8460 => x"70802577",
          8461 => x"07515154",
          8462 => x"73db3881",
          8463 => x"b53975ae",
          8464 => x"2e098106",
          8465 => x"83388154",
          8466 => x"767c2774",
          8467 => x"07547380",
          8468 => x"2ea2387b",
          8469 => x"8b327030",
          8470 => x"77ae3270",
          8471 => x"30728025",
          8472 => x"719f2a07",
          8473 => x"53515651",
          8474 => x"557481a7",
          8475 => x"3888578b",
          8476 => x"5cfef539",
          8477 => x"75982b54",
          8478 => x"7380258c",
          8479 => x"387580ff",
          8480 => x"0682af90",
          8481 => x"11335754",
          8482 => x"7551e6e1",
          8483 => x"3f82b5c8",
          8484 => x"08802eb2",
          8485 => x"38781870",
          8486 => x"33811a71",
          8487 => x"545a5654",
          8488 => x"e6d23f82",
          8489 => x"b5c80880",
          8490 => x"2e80e838",
          8491 => x"ff1c5476",
          8492 => x"742780df",
          8493 => x"38791754",
          8494 => x"75743481",
          8495 => x"177a1155",
          8496 => x"57747434",
          8497 => x"a7397552",
          8498 => x"82aeb051",
          8499 => x"e5fe3f82",
          8500 => x"b5c808bf",
          8501 => x"38ff9f16",
          8502 => x"54739926",
          8503 => x"8938e016",
          8504 => x"7081ff06",
          8505 => x"57547917",
          8506 => x"54757434",
          8507 => x"811757fd",
          8508 => x"f7397719",
          8509 => x"7e0c7680",
          8510 => x"2e993879",
          8511 => x"33547381",
          8512 => x"e52e0981",
          8513 => x"06843885",
          8514 => x"7a348454",
          8515 => x"a076278f",
          8516 => x"388b3986",
          8517 => x"5581f239",
          8518 => x"845680f3",
          8519 => x"39805473",
          8520 => x"8b1b3480",
          8521 => x"7b085852",
          8522 => x"7a51f2ce",
          8523 => x"3f82b5c8",
          8524 => x"085682b5",
          8525 => x"c80880d7",
          8526 => x"38981b08",
          8527 => x"527651e6",
          8528 => x"aa3f82b5",
          8529 => x"c8085682",
          8530 => x"b5c80880",
          8531 => x"c2389c1b",
          8532 => x"08703355",
          8533 => x"5573802e",
          8534 => x"ffbe388b",
          8535 => x"1533bf06",
          8536 => x"5473861c",
          8537 => x"348b1533",
          8538 => x"70832a70",
          8539 => x"81065155",
          8540 => x"58739238",
          8541 => x"8b537952",
          8542 => x"7451e49f",
          8543 => x"3f82b5c8",
          8544 => x"08802e8b",
          8545 => x"3875527a",
          8546 => x"51f3ba3f",
          8547 => x"ff9f3975",
          8548 => x"ab1c3357",
          8549 => x"5574802e",
          8550 => x"bb387484",
          8551 => x"2e098106",
          8552 => x"80e73875",
          8553 => x"852a7081",
          8554 => x"0677822a",
          8555 => x"58515473",
          8556 => x"802e9638",
          8557 => x"75810654",
          8558 => x"73802efb",
          8559 => x"b538ff80",
          8560 => x"0bab1c34",
          8561 => x"805580c1",
          8562 => x"39758106",
          8563 => x"5473ba38",
          8564 => x"8555b639",
          8565 => x"75822a70",
          8566 => x"81065154",
          8567 => x"73ab3886",
          8568 => x"1b337084",
          8569 => x"2a708106",
          8570 => x"51555573",
          8571 => x"802ee138",
          8572 => x"901b0883",
          8573 => x"ff061db4",
          8574 => x"05527c51",
          8575 => x"f5db3f82",
          8576 => x"b5c80888",
          8577 => x"1c0cfaea",
          8578 => x"397482b5",
          8579 => x"c80c8f3d",
          8580 => x"0d04f63d",
          8581 => x"0d7c5bff",
          8582 => x"7b087071",
          8583 => x"7355595c",
          8584 => x"55597380",
          8585 => x"2e81c638",
          8586 => x"75708105",
          8587 => x"573370a0",
          8588 => x"26525271",
          8589 => x"ba2e8d38",
          8590 => x"70ee3871",
          8591 => x"ba2e0981",
          8592 => x"0681a538",
          8593 => x"7333d011",
          8594 => x"7081ff06",
          8595 => x"51525370",
          8596 => x"89269138",
          8597 => x"82147381",
          8598 => x"ff06d005",
          8599 => x"56527176",
          8600 => x"2e80f738",
          8601 => x"800b82af",
          8602 => x"80595577",
          8603 => x"087a5557",
          8604 => x"76708105",
          8605 => x"58337470",
          8606 => x"81055633",
          8607 => x"ff9f1253",
          8608 => x"53537099",
          8609 => x"268938e0",
          8610 => x"137081ff",
          8611 => x"065451ff",
          8612 => x"9f125170",
          8613 => x"99268938",
          8614 => x"e0127081",
          8615 => x"ff065351",
          8616 => x"7230709f",
          8617 => x"2a515172",
          8618 => x"722e0981",
          8619 => x"06853870",
          8620 => x"ffbe3872",
          8621 => x"30747732",
          8622 => x"70307072",
          8623 => x"079f2a73",
          8624 => x"9f2a0753",
          8625 => x"54545170",
          8626 => x"802e8f38",
          8627 => x"81158419",
          8628 => x"59558375",
          8629 => x"25ff9438",
          8630 => x"8b397483",
          8631 => x"24863874",
          8632 => x"767c0c59",
          8633 => x"78518639",
          8634 => x"82cd9433",
          8635 => x"517082b5",
          8636 => x"c80c8c3d",
          8637 => x"0d04fa3d",
          8638 => x"0d785680",
          8639 => x"0b831734",
          8640 => x"ff0bb017",
          8641 => x"0c795275",
          8642 => x"51e2e03f",
          8643 => x"845582b5",
          8644 => x"c8088180",
          8645 => x"3884b216",
          8646 => x"51dfb43f",
          8647 => x"82b5c808",
          8648 => x"83ffff06",
          8649 => x"54835573",
          8650 => x"82d4d52e",
          8651 => x"09810680",
          8652 => x"e338800b",
          8653 => x"b4173356",
          8654 => x"577481e9",
          8655 => x"2e098106",
          8656 => x"83388157",
          8657 => x"7481eb32",
          8658 => x"70307080",
          8659 => x"25790751",
          8660 => x"5154738a",
          8661 => x"387481e8",
          8662 => x"2e098106",
          8663 => x"b5388353",
          8664 => x"82aec052",
          8665 => x"80ea1651",
          8666 => x"e0b13f82",
          8667 => x"b5c80855",
          8668 => x"82b5c808",
          8669 => x"802e9d38",
          8670 => x"855382ae",
          8671 => x"c4528186",
          8672 => x"1651e097",
          8673 => x"3f82b5c8",
          8674 => x"085582b5",
          8675 => x"c808802e",
          8676 => x"83388255",
          8677 => x"7482b5c8",
          8678 => x"0c883d0d",
          8679 => x"04f23d0d",
          8680 => x"61028405",
          8681 => x"80cb0533",
          8682 => x"58558075",
          8683 => x"0c6051fc",
          8684 => x"e13f82b5",
          8685 => x"c808588b",
          8686 => x"56800b82",
          8687 => x"b5c80824",
          8688 => x"86fc3882",
          8689 => x"b5c80884",
          8690 => x"2982cd80",
          8691 => x"05700855",
          8692 => x"538c5673",
          8693 => x"802e86e6",
          8694 => x"3873750c",
          8695 => x"7681fe06",
          8696 => x"74335457",
          8697 => x"72802eae",
          8698 => x"38811433",
          8699 => x"51d7ca3f",
          8700 => x"82b5c808",
          8701 => x"81ff0670",
          8702 => x"81065455",
          8703 => x"72983876",
          8704 => x"802e86b8",
          8705 => x"3874822a",
          8706 => x"70810651",
          8707 => x"538a5672",
          8708 => x"86ac3886",
          8709 => x"a7398074",
          8710 => x"34778115",
          8711 => x"34815281",
          8712 => x"143351d7",
          8713 => x"b23f82b5",
          8714 => x"c80881ff",
          8715 => x"06708106",
          8716 => x"54558356",
          8717 => x"72868738",
          8718 => x"76802e8f",
          8719 => x"3874822a",
          8720 => x"70810651",
          8721 => x"538a5672",
          8722 => x"85f43880",
          8723 => x"70537452",
          8724 => x"5bfda33f",
          8725 => x"82b5c808",
          8726 => x"81ff0657",
          8727 => x"76822e09",
          8728 => x"810680e2",
          8729 => x"388c3d74",
          8730 => x"56588356",
          8731 => x"83f61533",
          8732 => x"70585372",
          8733 => x"802e8d38",
          8734 => x"83fa1551",
          8735 => x"dce83f82",
          8736 => x"b5c80857",
          8737 => x"76787084",
          8738 => x"055a0cff",
          8739 => x"16901656",
          8740 => x"56758025",
          8741 => x"d738800b",
          8742 => x"8d3d5456",
          8743 => x"72708405",
          8744 => x"54085b83",
          8745 => x"577a802e",
          8746 => x"95387a52",
          8747 => x"7351fcc6",
          8748 => x"3f82b5c8",
          8749 => x"0881ff06",
          8750 => x"57817727",
          8751 => x"89388116",
          8752 => x"56837627",
          8753 => x"d7388156",
          8754 => x"76842e84",
          8755 => x"f1388d56",
          8756 => x"76812684",
          8757 => x"e938bf14",
          8758 => x"51dbf43f",
          8759 => x"82b5c808",
          8760 => x"83ffff06",
          8761 => x"53728480",
          8762 => x"2e098106",
          8763 => x"84d03880",
          8764 => x"ca1451db",
          8765 => x"da3f82b5",
          8766 => x"c80883ff",
          8767 => x"ff065877",
          8768 => x"8d3880d8",
          8769 => x"1451dbde",
          8770 => x"3f82b5c8",
          8771 => x"0858779c",
          8772 => x"150c80c4",
          8773 => x"14338215",
          8774 => x"3480c414",
          8775 => x"33ff1170",
          8776 => x"81ff0651",
          8777 => x"54558d56",
          8778 => x"72812684",
          8779 => x"91387481",
          8780 => x"ff067871",
          8781 => x"2980c116",
          8782 => x"33525953",
          8783 => x"728a1523",
          8784 => x"72802e8b",
          8785 => x"38ff1373",
          8786 => x"06537280",
          8787 => x"2e86388d",
          8788 => x"5683eb39",
          8789 => x"80c51451",
          8790 => x"daf53f82",
          8791 => x"b5c80853",
          8792 => x"82b5c808",
          8793 => x"88152372",
          8794 => x"8f06578d",
          8795 => x"567683ce",
          8796 => x"3880c714",
          8797 => x"51dad83f",
          8798 => x"82b5c808",
          8799 => x"83ffff06",
          8800 => x"55748d38",
          8801 => x"80d41451",
          8802 => x"dadc3f82",
          8803 => x"b5c80855",
          8804 => x"80c21451",
          8805 => x"dab93f82",
          8806 => x"b5c80883",
          8807 => x"ffff0653",
          8808 => x"8d567280",
          8809 => x"2e839738",
          8810 => x"88142278",
          8811 => x"1471842a",
          8812 => x"055a5a78",
          8813 => x"75268386",
          8814 => x"388a1422",
          8815 => x"52747931",
          8816 => x"51fef3bf",
          8817 => x"3f82b5c8",
          8818 => x"085582b5",
          8819 => x"c808802e",
          8820 => x"82ec3882",
          8821 => x"b5c80880",
          8822 => x"fffffff5",
          8823 => x"26833883",
          8824 => x"577483ff",
          8825 => x"f5268338",
          8826 => x"8257749f",
          8827 => x"f5268538",
          8828 => x"81578939",
          8829 => x"8d567680",
          8830 => x"2e82c338",
          8831 => x"82157098",
          8832 => x"160c7ba0",
          8833 => x"160c731c",
          8834 => x"70a4170c",
          8835 => x"7a1dac17",
          8836 => x"0c545576",
          8837 => x"832e0981",
          8838 => x"06af3880",
          8839 => x"de1451d9",
          8840 => x"ae3f82b5",
          8841 => x"c80883ff",
          8842 => x"ff06538d",
          8843 => x"5672828e",
          8844 => x"3879828a",
          8845 => x"3880e014",
          8846 => x"51d9ab3f",
          8847 => x"82b5c808",
          8848 => x"a8150c74",
          8849 => x"822b53a2",
          8850 => x"398d5679",
          8851 => x"802e81ee",
          8852 => x"387713a8",
          8853 => x"150c7415",
          8854 => x"5376822e",
          8855 => x"8d387410",
          8856 => x"1570812a",
          8857 => x"76810605",
          8858 => x"515383ff",
          8859 => x"13892a53",
          8860 => x"8d56729c",
          8861 => x"15082681",
          8862 => x"c538ff0b",
          8863 => x"90150cff",
          8864 => x"0b8c150c",
          8865 => x"ff800b84",
          8866 => x"15347683",
          8867 => x"2e098106",
          8868 => x"81923880",
          8869 => x"e41451d8",
          8870 => x"b63f82b5",
          8871 => x"c80883ff",
          8872 => x"ff065372",
          8873 => x"812e0981",
          8874 => x"0680f938",
          8875 => x"811b5273",
          8876 => x"51dbb83f",
          8877 => x"82b5c808",
          8878 => x"80ea3882",
          8879 => x"b5c80884",
          8880 => x"153484b2",
          8881 => x"1451d887",
          8882 => x"3f82b5c8",
          8883 => x"0883ffff",
          8884 => x"06537282",
          8885 => x"d4d52e09",
          8886 => x"810680c8",
          8887 => x"38b41451",
          8888 => x"d8843f82",
          8889 => x"b5c80884",
          8890 => x"8b85a4d2",
          8891 => x"2e098106",
          8892 => x"b3388498",
          8893 => x"1451d7ee",
          8894 => x"3f82b5c8",
          8895 => x"08868a85",
          8896 => x"e4f22e09",
          8897 => x"81069d38",
          8898 => x"849c1451",
          8899 => x"d7d83f82",
          8900 => x"b5c80890",
          8901 => x"150c84a0",
          8902 => x"1451d7ca",
          8903 => x"3f82b5c8",
          8904 => x"088c150c",
          8905 => x"76743482",
          8906 => x"cd902281",
          8907 => x"05537282",
          8908 => x"cd902372",
          8909 => x"86152380",
          8910 => x"0b94150c",
          8911 => x"80567582",
          8912 => x"b5c80c90",
          8913 => x"3d0d04fb",
          8914 => x"3d0d7754",
          8915 => x"89557380",
          8916 => x"2eb93873",
          8917 => x"08537280",
          8918 => x"2eb13872",
          8919 => x"33527180",
          8920 => x"2ea93886",
          8921 => x"13228415",
          8922 => x"22575271",
          8923 => x"762e0981",
          8924 => x"06993881",
          8925 => x"133351d0",
          8926 => x"c03f82b5",
          8927 => x"c8088106",
          8928 => x"52718838",
          8929 => x"71740854",
          8930 => x"55833980",
          8931 => x"53787371",
          8932 => x"0c527482",
          8933 => x"b5c80c87",
          8934 => x"3d0d04fa",
          8935 => x"3d0d02ab",
          8936 => x"05337a58",
          8937 => x"893dfc05",
          8938 => x"5256f4e6",
          8939 => x"3f8b5480",
          8940 => x"0b82b5c8",
          8941 => x"0824bc38",
          8942 => x"82b5c808",
          8943 => x"842982cd",
          8944 => x"80057008",
          8945 => x"55557380",
          8946 => x"2e843880",
          8947 => x"74347854",
          8948 => x"73802e84",
          8949 => x"38807434",
          8950 => x"78750c75",
          8951 => x"5475802e",
          8952 => x"92388053",
          8953 => x"893d7053",
          8954 => x"840551f7",
          8955 => x"b03f82b5",
          8956 => x"c8085473",
          8957 => x"82b5c80c",
          8958 => x"883d0d04",
          8959 => x"eb3d0d67",
          8960 => x"02840580",
          8961 => x"e7053359",
          8962 => x"59895478",
          8963 => x"802e84c8",
          8964 => x"3877bf06",
          8965 => x"7054983d",
          8966 => x"d0055399",
          8967 => x"3d840552",
          8968 => x"58f6fa3f",
          8969 => x"82b5c808",
          8970 => x"5582b5c8",
          8971 => x"0884a438",
          8972 => x"7a5c6852",
          8973 => x"8c3d7052",
          8974 => x"56edc63f",
          8975 => x"82b5c808",
          8976 => x"5582b5c8",
          8977 => x"08923802",
          8978 => x"80d70533",
          8979 => x"70982b55",
          8980 => x"57738025",
          8981 => x"83388655",
          8982 => x"779c0654",
          8983 => x"73802e81",
          8984 => x"ab387480",
          8985 => x"2e953874",
          8986 => x"842e0981",
          8987 => x"06aa3875",
          8988 => x"51eaf83f",
          8989 => x"82b5c808",
          8990 => x"559e3902",
          8991 => x"b2053391",
          8992 => x"06547381",
          8993 => x"b8387782",
          8994 => x"2a708106",
          8995 => x"51547380",
          8996 => x"2e8e3888",
          8997 => x"5583bc39",
          8998 => x"77880758",
          8999 => x"7483b438",
          9000 => x"77832a70",
          9001 => x"81065154",
          9002 => x"73802e81",
          9003 => x"af386252",
          9004 => x"7a51e8a5",
          9005 => x"3f82b5c8",
          9006 => x"08568288",
          9007 => x"b20a5262",
          9008 => x"8e0551d4",
          9009 => x"ea3f6254",
          9010 => x"a00b8b15",
          9011 => x"34805362",
          9012 => x"527a51e8",
          9013 => x"bd3f8052",
          9014 => x"629c0551",
          9015 => x"d4d13f7a",
          9016 => x"54810b83",
          9017 => x"15347580",
          9018 => x"2e80f138",
          9019 => x"7ab01108",
          9020 => x"51548053",
          9021 => x"7552973d",
          9022 => x"d40551dd",
          9023 => x"be3f82b5",
          9024 => x"c8085582",
          9025 => x"b5c80882",
          9026 => x"ca38b739",
          9027 => x"7482c438",
          9028 => x"02b20533",
          9029 => x"70842a70",
          9030 => x"81065155",
          9031 => x"5673802e",
          9032 => x"86388455",
          9033 => x"82ad3977",
          9034 => x"812a7081",
          9035 => x"06515473",
          9036 => x"802ea938",
          9037 => x"75810654",
          9038 => x"73802ea0",
          9039 => x"38875582",
          9040 => x"92397352",
          9041 => x"7a51d6a3",
          9042 => x"3f82b5c8",
          9043 => x"087bff18",
          9044 => x"8c120c55",
          9045 => x"5582b5c8",
          9046 => x"0881f838",
          9047 => x"77832a70",
          9048 => x"81065154",
          9049 => x"73802e86",
          9050 => x"387780c0",
          9051 => x"07587ab0",
          9052 => x"1108a01b",
          9053 => x"0c63a41b",
          9054 => x"0c635370",
          9055 => x"5257e6d9",
          9056 => x"3f82b5c8",
          9057 => x"0882b5c8",
          9058 => x"08881b0c",
          9059 => x"639c0552",
          9060 => x"5ad2d33f",
          9061 => x"82b5c808",
          9062 => x"82b5c808",
          9063 => x"8c1b0c77",
          9064 => x"7a0c5686",
          9065 => x"1722841a",
          9066 => x"2377901a",
          9067 => x"34800b91",
          9068 => x"1a34800b",
          9069 => x"9c1a0c80",
          9070 => x"0b941a0c",
          9071 => x"77852a70",
          9072 => x"81065154",
          9073 => x"73802e81",
          9074 => x"8d3882b5",
          9075 => x"c808802e",
          9076 => x"81843882",
          9077 => x"b5c80894",
          9078 => x"1a0c8a17",
          9079 => x"2270892b",
          9080 => x"7b525957",
          9081 => x"a8397652",
          9082 => x"7851d79f",
          9083 => x"3f82b5c8",
          9084 => x"085782b5",
          9085 => x"c8088126",
          9086 => x"83388255",
          9087 => x"82b5c808",
          9088 => x"ff2e0981",
          9089 => x"06833879",
          9090 => x"55757831",
          9091 => x"56743070",
          9092 => x"76078025",
          9093 => x"51547776",
          9094 => x"278a3881",
          9095 => x"70750655",
          9096 => x"5a73c338",
          9097 => x"76981a0c",
          9098 => x"74a93875",
          9099 => x"83ff0654",
          9100 => x"73802ea2",
          9101 => x"3876527a",
          9102 => x"51d6a63f",
          9103 => x"82b5c808",
          9104 => x"85388255",
          9105 => x"8e397589",
          9106 => x"2a82b5c8",
          9107 => x"08059c1a",
          9108 => x"0c843980",
          9109 => x"790c7454",
          9110 => x"7382b5c8",
          9111 => x"0c973d0d",
          9112 => x"04f23d0d",
          9113 => x"60636564",
          9114 => x"40405d59",
          9115 => x"807e0c90",
          9116 => x"3dfc0552",
          9117 => x"7851f9cf",
          9118 => x"3f82b5c8",
          9119 => x"085582b5",
          9120 => x"c8088a38",
          9121 => x"91193355",
          9122 => x"74802e86",
          9123 => x"38745682",
          9124 => x"c4399019",
          9125 => x"33810655",
          9126 => x"87567480",
          9127 => x"2e82b638",
          9128 => x"9539820b",
          9129 => x"911a3482",
          9130 => x"5682aa39",
          9131 => x"810b911a",
          9132 => x"34815682",
          9133 => x"a0398c19",
          9134 => x"08941a08",
          9135 => x"3155747c",
          9136 => x"27833874",
          9137 => x"5c7b802e",
          9138 => x"82893894",
          9139 => x"19087083",
          9140 => x"ff065656",
          9141 => x"7481b238",
          9142 => x"7e8a1122",
          9143 => x"ff057789",
          9144 => x"2a065b55",
          9145 => x"79a83875",
          9146 => x"87388819",
          9147 => x"08558f39",
          9148 => x"98190852",
          9149 => x"7851d593",
          9150 => x"3f82b5c8",
          9151 => x"08558175",
          9152 => x"27ff9f38",
          9153 => x"74ff2eff",
          9154 => x"a3387498",
          9155 => x"1a0c9819",
          9156 => x"08527e51",
          9157 => x"d4cb3f82",
          9158 => x"b5c80880",
          9159 => x"2eff8338",
          9160 => x"82b5c808",
          9161 => x"1a7c892a",
          9162 => x"59577780",
          9163 => x"2e80d638",
          9164 => x"771a7f8a",
          9165 => x"1122585c",
          9166 => x"55757527",
          9167 => x"8538757a",
          9168 => x"31587754",
          9169 => x"76537c52",
          9170 => x"811b3351",
          9171 => x"ca883f82",
          9172 => x"b5c808fe",
          9173 => x"d7387e83",
          9174 => x"11335656",
          9175 => x"74802e9f",
          9176 => x"38b01608",
          9177 => x"77315574",
          9178 => x"78279438",
          9179 => x"848053b4",
          9180 => x"1652b016",
          9181 => x"08773189",
          9182 => x"2b7d0551",
          9183 => x"cfe03f77",
          9184 => x"892b56b9",
          9185 => x"39769c1a",
          9186 => x"0c941908",
          9187 => x"83ff0684",
          9188 => x"80713157",
          9189 => x"557b7627",
          9190 => x"83387b56",
          9191 => x"9c190852",
          9192 => x"7e51d1c7",
          9193 => x"3f82b5c8",
          9194 => x"08fe8138",
          9195 => x"75539419",
          9196 => x"0883ff06",
          9197 => x"1fb40552",
          9198 => x"7c51cfa2",
          9199 => x"3f7b7631",
          9200 => x"7e08177f",
          9201 => x"0c761e94",
          9202 => x"1b081894",
          9203 => x"1c0c5e5c",
          9204 => x"fdf33980",
          9205 => x"567582b5",
          9206 => x"c80c903d",
          9207 => x"0d04f23d",
          9208 => x"0d606365",
          9209 => x"6440405d",
          9210 => x"58807e0c",
          9211 => x"903dfc05",
          9212 => x"527751f6",
          9213 => x"d23f82b5",
          9214 => x"c8085582",
          9215 => x"b5c8088a",
          9216 => x"38911833",
          9217 => x"5574802e",
          9218 => x"86387456",
          9219 => x"83b83990",
          9220 => x"18337081",
          9221 => x"2a708106",
          9222 => x"51565687",
          9223 => x"5674802e",
          9224 => x"83a43895",
          9225 => x"39820b91",
          9226 => x"19348256",
          9227 => x"83983981",
          9228 => x"0b911934",
          9229 => x"8156838e",
          9230 => x"39941808",
          9231 => x"7c115656",
          9232 => x"74762784",
          9233 => x"3875095c",
          9234 => x"7b802e82",
          9235 => x"ec389418",
          9236 => x"087083ff",
          9237 => x"06565674",
          9238 => x"81fd387e",
          9239 => x"8a1122ff",
          9240 => x"0577892a",
          9241 => x"065c557a",
          9242 => x"bf38758c",
          9243 => x"38881808",
          9244 => x"55749c38",
          9245 => x"7a528539",
          9246 => x"98180852",
          9247 => x"7751d7e7",
          9248 => x"3f82b5c8",
          9249 => x"085582b5",
          9250 => x"c808802e",
          9251 => x"82ab3874",
          9252 => x"812eff91",
          9253 => x"3874ff2e",
          9254 => x"ff953874",
          9255 => x"98190c88",
          9256 => x"18088538",
          9257 => x"7488190c",
          9258 => x"7e55b015",
          9259 => x"089c1908",
          9260 => x"2e098106",
          9261 => x"8d387451",
          9262 => x"cec13f82",
          9263 => x"b5c808fe",
          9264 => x"ee389818",
          9265 => x"08527e51",
          9266 => x"d1973f82",
          9267 => x"b5c80880",
          9268 => x"2efed238",
          9269 => x"82b5c808",
          9270 => x"1b7c892a",
          9271 => x"5a577880",
          9272 => x"2e80d538",
          9273 => x"781b7f8a",
          9274 => x"1122585b",
          9275 => x"55757527",
          9276 => x"8538757b",
          9277 => x"31597854",
          9278 => x"76537c52",
          9279 => x"811a3351",
          9280 => x"c8be3f82",
          9281 => x"b5c808fe",
          9282 => x"a6387eb0",
          9283 => x"11087831",
          9284 => x"56567479",
          9285 => x"279b3884",
          9286 => x"8053b016",
          9287 => x"08773189",
          9288 => x"2b7d0552",
          9289 => x"b41651cc",
          9290 => x"b53f7e55",
          9291 => x"800b8316",
          9292 => x"3478892b",
          9293 => x"5680db39",
          9294 => x"8c180894",
          9295 => x"19082693",
          9296 => x"387e51cd",
          9297 => x"b63f82b5",
          9298 => x"c808fde3",
          9299 => x"387e77b0",
          9300 => x"120c5576",
          9301 => x"9c190c94",
          9302 => x"180883ff",
          9303 => x"06848071",
          9304 => x"3157557b",
          9305 => x"76278338",
          9306 => x"7b569c18",
          9307 => x"08527e51",
          9308 => x"cdf93f82",
          9309 => x"b5c808fd",
          9310 => x"b6387553",
          9311 => x"7c529418",
          9312 => x"0883ff06",
          9313 => x"1fb40551",
          9314 => x"cbd43f7e",
          9315 => x"55810b83",
          9316 => x"16347b76",
          9317 => x"317e0817",
          9318 => x"7f0c761e",
          9319 => x"941a0818",
          9320 => x"70941c0c",
          9321 => x"8c1b0858",
          9322 => x"585e5c74",
          9323 => x"76278338",
          9324 => x"7555748c",
          9325 => x"190cfd90",
          9326 => x"39901833",
          9327 => x"80c00755",
          9328 => x"74901934",
          9329 => x"80567582",
          9330 => x"b5c80c90",
          9331 => x"3d0d04f8",
          9332 => x"3d0d7a8b",
          9333 => x"3dfc0553",
          9334 => x"705256f2",
          9335 => x"ea3f82b5",
          9336 => x"c8085782",
          9337 => x"b5c80880",
          9338 => x"fb389016",
          9339 => x"3370862a",
          9340 => x"70810651",
          9341 => x"55557380",
          9342 => x"2e80e938",
          9343 => x"a0160852",
          9344 => x"7851cce7",
          9345 => x"3f82b5c8",
          9346 => x"085782b5",
          9347 => x"c80880d4",
          9348 => x"38a41608",
          9349 => x"8b1133a0",
          9350 => x"07555573",
          9351 => x"8b163488",
          9352 => x"16085374",
          9353 => x"52750851",
          9354 => x"dde83f8c",
          9355 => x"1608529c",
          9356 => x"1551c9fb",
          9357 => x"3f8288b2",
          9358 => x"0a529615",
          9359 => x"51c9f03f",
          9360 => x"76529215",
          9361 => x"51c9ca3f",
          9362 => x"7854810b",
          9363 => x"83153478",
          9364 => x"51ccdf3f",
          9365 => x"82b5c808",
          9366 => x"90173381",
          9367 => x"bf065557",
          9368 => x"73901734",
          9369 => x"7682b5c8",
          9370 => x"0c8a3d0d",
          9371 => x"04fc3d0d",
          9372 => x"76705254",
          9373 => x"fed93f82",
          9374 => x"b5c80853",
          9375 => x"82b5c808",
          9376 => x"9c38863d",
          9377 => x"fc055273",
          9378 => x"51f1bc3f",
          9379 => x"82b5c808",
          9380 => x"5382b5c8",
          9381 => x"08873882",
          9382 => x"b5c80874",
          9383 => x"0c7282b5",
          9384 => x"c80c863d",
          9385 => x"0d04ff3d",
          9386 => x"0d843d51",
          9387 => x"e6e43f8b",
          9388 => x"52800b82",
          9389 => x"b5c80824",
          9390 => x"8b3882b5",
          9391 => x"c80882cd",
          9392 => x"94348052",
          9393 => x"7182b5c8",
          9394 => x"0c833d0d",
          9395 => x"04ef3d0d",
          9396 => x"8053933d",
          9397 => x"d0055294",
          9398 => x"3d51e9c1",
          9399 => x"3f82b5c8",
          9400 => x"085582b5",
          9401 => x"c80880e0",
          9402 => x"38765863",
          9403 => x"52933dd4",
          9404 => x"0551e08d",
          9405 => x"3f82b5c8",
          9406 => x"085582b5",
          9407 => x"c808bc38",
          9408 => x"0280c705",
          9409 => x"3370982b",
          9410 => x"55567380",
          9411 => x"25893876",
          9412 => x"7a94120c",
          9413 => x"54b23902",
          9414 => x"a2053370",
          9415 => x"842a7081",
          9416 => x"06515556",
          9417 => x"73802e9e",
          9418 => x"38767f53",
          9419 => x"705254db",
          9420 => x"a83f82b5",
          9421 => x"c8089415",
          9422 => x"0c8e3982",
          9423 => x"b5c80884",
          9424 => x"2e098106",
          9425 => x"83388555",
          9426 => x"7482b5c8",
          9427 => x"0c933d0d",
          9428 => x"04e43d0d",
          9429 => x"6f6f5b5b",
          9430 => x"807a3480",
          9431 => x"539e3dff",
          9432 => x"b805529f",
          9433 => x"3d51e8b5",
          9434 => x"3f82b5c8",
          9435 => x"085782b5",
          9436 => x"c80882fc",
          9437 => x"387b437a",
          9438 => x"7c941108",
          9439 => x"47555864",
          9440 => x"5473802e",
          9441 => x"81ed38a0",
          9442 => x"52933d70",
          9443 => x"5255d5ea",
          9444 => x"3f82b5c8",
          9445 => x"085782b5",
          9446 => x"c80882d4",
          9447 => x"3868527b",
          9448 => x"51c9c83f",
          9449 => x"82b5c808",
          9450 => x"5782b5c8",
          9451 => x"0882c138",
          9452 => x"69527b51",
          9453 => x"daa33f82",
          9454 => x"b5c80845",
          9455 => x"76527451",
          9456 => x"d5b83f82",
          9457 => x"b5c80857",
          9458 => x"82b5c808",
          9459 => x"82a23880",
          9460 => x"527451da",
          9461 => x"eb3f82b5",
          9462 => x"c8085782",
          9463 => x"b5c808a4",
          9464 => x"3869527b",
          9465 => x"51d9f23f",
          9466 => x"7382b5c8",
          9467 => x"082ea638",
          9468 => x"76527451",
          9469 => x"d6cf3f82",
          9470 => x"b5c80857",
          9471 => x"82b5c808",
          9472 => x"802ecc38",
          9473 => x"76842e09",
          9474 => x"81068638",
          9475 => x"825781e0",
          9476 => x"397681dc",
          9477 => x"389e3dff",
          9478 => x"bc055274",
          9479 => x"51dcc93f",
          9480 => x"76903d78",
          9481 => x"11811133",
          9482 => x"51565a56",
          9483 => x"73802e91",
          9484 => x"3802b905",
          9485 => x"55811681",
          9486 => x"16703356",
          9487 => x"565673f5",
          9488 => x"38811654",
          9489 => x"73782681",
          9490 => x"90387580",
          9491 => x"2e993878",
          9492 => x"16810555",
          9493 => x"ff186f11",
          9494 => x"ff18ff18",
          9495 => x"58585558",
          9496 => x"74337434",
          9497 => x"75ee38ff",
          9498 => x"186f1155",
          9499 => x"58af7434",
          9500 => x"fe8d3977",
          9501 => x"7b2e0981",
          9502 => x"068a38ff",
          9503 => x"186f1155",
          9504 => x"58af7434",
          9505 => x"800b82cd",
          9506 => x"94337084",
          9507 => x"2982af80",
          9508 => x"05700870",
          9509 => x"33525c56",
          9510 => x"56567376",
          9511 => x"2e8d3881",
          9512 => x"16701a70",
          9513 => x"33515556",
          9514 => x"73f53882",
          9515 => x"16547378",
          9516 => x"26a73880",
          9517 => x"55747627",
          9518 => x"91387419",
          9519 => x"5473337a",
          9520 => x"7081055c",
          9521 => x"34811555",
          9522 => x"ec39ba7a",
          9523 => x"7081055c",
          9524 => x"3474ff2e",
          9525 => x"09810685",
          9526 => x"38915794",
          9527 => x"396e1881",
          9528 => x"19595473",
          9529 => x"337a7081",
          9530 => x"055c347a",
          9531 => x"7826ee38",
          9532 => x"807a3476",
          9533 => x"82b5c80c",
          9534 => x"9e3d0d04",
          9535 => x"f73d0d7b",
          9536 => x"7d8d3dfc",
          9537 => x"05547153",
          9538 => x"5755ecbb",
          9539 => x"3f82b5c8",
          9540 => x"085382b5",
          9541 => x"c80882fa",
          9542 => x"38911533",
          9543 => x"537282f2",
          9544 => x"388c1508",
          9545 => x"54737627",
          9546 => x"92389015",
          9547 => x"3370812a",
          9548 => x"70810651",
          9549 => x"54577283",
          9550 => x"38735694",
          9551 => x"15085480",
          9552 => x"7094170c",
          9553 => x"5875782e",
          9554 => x"82973879",
          9555 => x"8a112270",
          9556 => x"892b5951",
          9557 => x"5373782e",
          9558 => x"b7387652",
          9559 => x"ff1651fe",
          9560 => x"dca13f82",
          9561 => x"b5c808ff",
          9562 => x"15785470",
          9563 => x"535553fe",
          9564 => x"dc913f82",
          9565 => x"b5c80873",
          9566 => x"26963876",
          9567 => x"30707506",
          9568 => x"7094180c",
          9569 => x"77713198",
          9570 => x"18085758",
          9571 => x"5153b139",
          9572 => x"88150854",
          9573 => x"73a63873",
          9574 => x"527451cd",
          9575 => x"ca3f82b5",
          9576 => x"c8085482",
          9577 => x"b5c80881",
          9578 => x"2e819a38",
          9579 => x"82b5c808",
          9580 => x"ff2e819b",
          9581 => x"3882b5c8",
          9582 => x"0888160c",
          9583 => x"7398160c",
          9584 => x"73802e81",
          9585 => x"9c387676",
          9586 => x"2780dc38",
          9587 => x"75773194",
          9588 => x"16081894",
          9589 => x"170c9016",
          9590 => x"3370812a",
          9591 => x"70810651",
          9592 => x"555a5672",
          9593 => x"802e9a38",
          9594 => x"73527451",
          9595 => x"ccf93f82",
          9596 => x"b5c80854",
          9597 => x"82b5c808",
          9598 => x"943882b5",
          9599 => x"c80856a7",
          9600 => x"39735274",
          9601 => x"51c7843f",
          9602 => x"82b5c808",
          9603 => x"5473ff2e",
          9604 => x"be388174",
          9605 => x"27af3879",
          9606 => x"53739814",
          9607 => x"0827a638",
          9608 => x"7398160c",
          9609 => x"ffa03994",
          9610 => x"15081694",
          9611 => x"160c7583",
          9612 => x"ff065372",
          9613 => x"802eaa38",
          9614 => x"73527951",
          9615 => x"c6a33f82",
          9616 => x"b5c80894",
          9617 => x"38820b91",
          9618 => x"16348253",
          9619 => x"80c43981",
          9620 => x"0b911634",
          9621 => x"8153bb39",
          9622 => x"75892a82",
          9623 => x"b5c80805",
          9624 => x"58941508",
          9625 => x"548c1508",
          9626 => x"74279038",
          9627 => x"738c160c",
          9628 => x"90153380",
          9629 => x"c0075372",
          9630 => x"90163473",
          9631 => x"83ff0653",
          9632 => x"72802e8c",
          9633 => x"38779c16",
          9634 => x"082e8538",
          9635 => x"779c160c",
          9636 => x"80537282",
          9637 => x"b5c80c8b",
          9638 => x"3d0d04f9",
          9639 => x"3d0d7956",
          9640 => x"89547580",
          9641 => x"2e818a38",
          9642 => x"8053893d",
          9643 => x"fc05528a",
          9644 => x"3d840551",
          9645 => x"e1e73f82",
          9646 => x"b5c80855",
          9647 => x"82b5c808",
          9648 => x"80ea3877",
          9649 => x"760c7a52",
          9650 => x"7551d8b5",
          9651 => x"3f82b5c8",
          9652 => x"085582b5",
          9653 => x"c80880c3",
          9654 => x"38ab1633",
          9655 => x"70982b55",
          9656 => x"57807424",
          9657 => x"a2388616",
          9658 => x"3370842a",
          9659 => x"70810651",
          9660 => x"55577380",
          9661 => x"2ead389c",
          9662 => x"16085277",
          9663 => x"51d3da3f",
          9664 => x"82b5c808",
          9665 => x"88170c77",
          9666 => x"54861422",
          9667 => x"84172374",
          9668 => x"527551ce",
          9669 => x"e53f82b5",
          9670 => x"c8085574",
          9671 => x"842e0981",
          9672 => x"06853885",
          9673 => x"55863974",
          9674 => x"802e8438",
          9675 => x"80760c74",
          9676 => x"547382b5",
          9677 => x"c80c893d",
          9678 => x"0d04fc3d",
          9679 => x"0d76873d",
          9680 => x"fc055370",
          9681 => x"5253e7ff",
          9682 => x"3f82b5c8",
          9683 => x"08873882",
          9684 => x"b5c80873",
          9685 => x"0c863d0d",
          9686 => x"04fb3d0d",
          9687 => x"7779893d",
          9688 => x"fc055471",
          9689 => x"535654e7",
          9690 => x"de3f82b5",
          9691 => x"c8085382",
          9692 => x"b5c80880",
          9693 => x"df387493",
          9694 => x"3882b5c8",
          9695 => x"08527351",
          9696 => x"cdf83f82",
          9697 => x"b5c80853",
          9698 => x"80ca3982",
          9699 => x"b5c80852",
          9700 => x"7351d3ac",
          9701 => x"3f82b5c8",
          9702 => x"085382b5",
          9703 => x"c808842e",
          9704 => x"09810685",
          9705 => x"38805387",
          9706 => x"3982b5c8",
          9707 => x"08a63874",
          9708 => x"527351d5",
          9709 => x"b33f7252",
          9710 => x"7351cf89",
          9711 => x"3f82b5c8",
          9712 => x"08843270",
          9713 => x"30707207",
          9714 => x"9f2c7082",
          9715 => x"b5c80806",
          9716 => x"51515454",
          9717 => x"7282b5c8",
          9718 => x"0c873d0d",
          9719 => x"04ee3d0d",
          9720 => x"65578053",
          9721 => x"893d7053",
          9722 => x"963d5256",
          9723 => x"dfaf3f82",
          9724 => x"b5c80855",
          9725 => x"82b5c808",
          9726 => x"b2386452",
          9727 => x"7551d681",
          9728 => x"3f82b5c8",
          9729 => x"085582b5",
          9730 => x"c808a038",
          9731 => x"0280cb05",
          9732 => x"3370982b",
          9733 => x"55587380",
          9734 => x"25853886",
          9735 => x"558d3976",
          9736 => x"802e8838",
          9737 => x"76527551",
          9738 => x"d4be3f74",
          9739 => x"82b5c80c",
          9740 => x"943d0d04",
          9741 => x"f03d0d63",
          9742 => x"65555c80",
          9743 => x"53923dec",
          9744 => x"0552933d",
          9745 => x"51ded63f",
          9746 => x"82b5c808",
          9747 => x"5b82b5c8",
          9748 => x"08828038",
          9749 => x"7c740c73",
          9750 => x"08981108",
          9751 => x"fe119013",
          9752 => x"08595658",
          9753 => x"55757426",
          9754 => x"9138757c",
          9755 => x"0c81e439",
          9756 => x"815b81cc",
          9757 => x"39825b81",
          9758 => x"c73982b5",
          9759 => x"c8087533",
          9760 => x"55597381",
          9761 => x"2e098106",
          9762 => x"bf388275",
          9763 => x"5f577652",
          9764 => x"923df005",
          9765 => x"51c1f43f",
          9766 => x"82b5c808",
          9767 => x"ff2ed138",
          9768 => x"82b5c808",
          9769 => x"812ece38",
          9770 => x"82b5c808",
          9771 => x"307082b5",
          9772 => x"c8080780",
          9773 => x"257a0581",
          9774 => x"197f5359",
          9775 => x"5a549814",
          9776 => x"087726ca",
          9777 => x"3880f939",
          9778 => x"a4150882",
          9779 => x"b5c80857",
          9780 => x"58759838",
          9781 => x"77528118",
          9782 => x"7d5258ff",
          9783 => x"bf8d3f82",
          9784 => x"b5c8085b",
          9785 => x"82b5c808",
          9786 => x"80d6387c",
          9787 => x"70337712",
          9788 => x"ff1a5d52",
          9789 => x"56547482",
          9790 => x"2e098106",
          9791 => x"9e38b414",
          9792 => x"51ffbbcb",
          9793 => x"3f82b5c8",
          9794 => x"0883ffff",
          9795 => x"06703070",
          9796 => x"80251b82",
          9797 => x"19595b51",
          9798 => x"549b39b4",
          9799 => x"1451ffbb",
          9800 => x"c53f82b5",
          9801 => x"c808f00a",
          9802 => x"06703070",
          9803 => x"80251b84",
          9804 => x"19595b51",
          9805 => x"547583ff",
          9806 => x"067a5856",
          9807 => x"79ff9238",
          9808 => x"787c0c7c",
          9809 => x"7990120c",
          9810 => x"84113381",
          9811 => x"07565474",
          9812 => x"8415347a",
          9813 => x"82b5c80c",
          9814 => x"923d0d04",
          9815 => x"f93d0d79",
          9816 => x"8a3dfc05",
          9817 => x"53705257",
          9818 => x"e3dd3f82",
          9819 => x"b5c80856",
          9820 => x"82b5c808",
          9821 => x"81a83891",
          9822 => x"17335675",
          9823 => x"81a03890",
          9824 => x"17337081",
          9825 => x"2a708106",
          9826 => x"51555587",
          9827 => x"5573802e",
          9828 => x"818e3894",
          9829 => x"17085473",
          9830 => x"8c180827",
          9831 => x"81803873",
          9832 => x"9b3882b5",
          9833 => x"c8085388",
          9834 => x"17085276",
          9835 => x"51c48c3f",
          9836 => x"82b5c808",
          9837 => x"7488190c",
          9838 => x"5680c939",
          9839 => x"98170852",
          9840 => x"7651ffbf",
          9841 => x"c63f82b5",
          9842 => x"c808ff2e",
          9843 => x"09810683",
          9844 => x"38815682",
          9845 => x"b5c80881",
          9846 => x"2e098106",
          9847 => x"85388256",
          9848 => x"a33975a0",
          9849 => x"38775482",
          9850 => x"b5c80898",
          9851 => x"15082794",
          9852 => x"38981708",
          9853 => x"5382b5c8",
          9854 => x"08527651",
          9855 => x"c3bd3f82",
          9856 => x"b5c80856",
          9857 => x"9417088c",
          9858 => x"180c9017",
          9859 => x"3380c007",
          9860 => x"54739018",
          9861 => x"3475802e",
          9862 => x"85387591",
          9863 => x"18347555",
          9864 => x"7482b5c8",
          9865 => x"0c893d0d",
          9866 => x"04e23d0d",
          9867 => x"8253a03d",
          9868 => x"ffa40552",
          9869 => x"a13d51da",
          9870 => x"e43f82b5",
          9871 => x"c8085582",
          9872 => x"b5c80881",
          9873 => x"f5387845",
          9874 => x"a13d0852",
          9875 => x"953d7052",
          9876 => x"58d1ae3f",
          9877 => x"82b5c808",
          9878 => x"5582b5c8",
          9879 => x"0881db38",
          9880 => x"0280fb05",
          9881 => x"3370852a",
          9882 => x"70810651",
          9883 => x"55568655",
          9884 => x"7381c738",
          9885 => x"75982b54",
          9886 => x"80742481",
          9887 => x"bd380280",
          9888 => x"d6053370",
          9889 => x"81065854",
          9890 => x"87557681",
          9891 => x"ad386b52",
          9892 => x"7851ccc5",
          9893 => x"3f82b5c8",
          9894 => x"0874842a",
          9895 => x"70810651",
          9896 => x"55567380",
          9897 => x"2e80d438",
          9898 => x"785482b5",
          9899 => x"c8089415",
          9900 => x"082e8186",
          9901 => x"38735a82",
          9902 => x"b5c8085c",
          9903 => x"76528a3d",
          9904 => x"705254c7",
          9905 => x"b53f82b5",
          9906 => x"c8085582",
          9907 => x"b5c80880",
          9908 => x"e93882b5",
          9909 => x"c8085273",
          9910 => x"51cce53f",
          9911 => x"82b5c808",
          9912 => x"5582b5c8",
          9913 => x"08863887",
          9914 => x"5580cf39",
          9915 => x"82b5c808",
          9916 => x"842e8838",
          9917 => x"82b5c808",
          9918 => x"80c03877",
          9919 => x"51cec23f",
          9920 => x"82b5c808",
          9921 => x"82b5c808",
          9922 => x"307082b5",
          9923 => x"c8080780",
          9924 => x"25515555",
          9925 => x"75802e94",
          9926 => x"3873802e",
          9927 => x"8f388053",
          9928 => x"75527751",
          9929 => x"c1953f82",
          9930 => x"b5c80855",
          9931 => x"748c3878",
          9932 => x"51ffbafe",
          9933 => x"3f82b5c8",
          9934 => x"08557482",
          9935 => x"b5c80ca0",
          9936 => x"3d0d04e9",
          9937 => x"3d0d8253",
          9938 => x"993dc005",
          9939 => x"529a3d51",
          9940 => x"d8cb3f82",
          9941 => x"b5c80854",
          9942 => x"82b5c808",
          9943 => x"82b03878",
          9944 => x"5e69528e",
          9945 => x"3d705258",
          9946 => x"cf973f82",
          9947 => x"b5c80854",
          9948 => x"82b5c808",
          9949 => x"86388854",
          9950 => x"82943982",
          9951 => x"b5c80884",
          9952 => x"2e098106",
          9953 => x"82883802",
          9954 => x"80df0533",
          9955 => x"70852a81",
          9956 => x"06515586",
          9957 => x"547481f6",
          9958 => x"38785a74",
          9959 => x"528a3d70",
          9960 => x"5257c1c3",
          9961 => x"3f82b5c8",
          9962 => x"08755556",
          9963 => x"82b5c808",
          9964 => x"83388754",
          9965 => x"82b5c808",
          9966 => x"812e0981",
          9967 => x"06833882",
          9968 => x"5482b5c8",
          9969 => x"08ff2e09",
          9970 => x"81068638",
          9971 => x"815481b4",
          9972 => x"397381b0",
          9973 => x"3882b5c8",
          9974 => x"08527851",
          9975 => x"c4a43f82",
          9976 => x"b5c80854",
          9977 => x"82b5c808",
          9978 => x"819a388b",
          9979 => x"53a052b4",
          9980 => x"1951ffb7",
          9981 => x"8c3f7854",
          9982 => x"ae0bb415",
          9983 => x"34785490",
          9984 => x"0bbf1534",
          9985 => x"8288b20a",
          9986 => x"5280ca19",
          9987 => x"51ffb69f",
          9988 => x"3f755378",
          9989 => x"b4115351",
          9990 => x"c9f83fa0",
          9991 => x"5378b411",
          9992 => x"5380d405",
          9993 => x"51ffb6b6",
          9994 => x"3f7854ae",
          9995 => x"0b80d515",
          9996 => x"347f5378",
          9997 => x"80d41153",
          9998 => x"51c9d73f",
          9999 => x"7854810b",
         10000 => x"83153477",
         10001 => x"51cba43f",
         10002 => x"82b5c808",
         10003 => x"5482b5c8",
         10004 => x"08b23882",
         10005 => x"88b20a52",
         10006 => x"64960551",
         10007 => x"ffb5d03f",
         10008 => x"75536452",
         10009 => x"7851c9aa",
         10010 => x"3f645490",
         10011 => x"0b8b1534",
         10012 => x"7854810b",
         10013 => x"83153478",
         10014 => x"51ffb8b6",
         10015 => x"3f82b5c8",
         10016 => x"08548b39",
         10017 => x"80537552",
         10018 => x"7651ffbe",
         10019 => x"ae3f7382",
         10020 => x"b5c80c99",
         10021 => x"3d0d04da",
         10022 => x"3d0da93d",
         10023 => x"840551d2",
         10024 => x"f13f8253",
         10025 => x"a83dff84",
         10026 => x"0552a93d",
         10027 => x"51d5ee3f",
         10028 => x"82b5c808",
         10029 => x"5582b5c8",
         10030 => x"0882d338",
         10031 => x"784da93d",
         10032 => x"08529d3d",
         10033 => x"705258cc",
         10034 => x"b83f82b5",
         10035 => x"c8085582",
         10036 => x"b5c80882",
         10037 => x"b9380281",
         10038 => x"9b053381",
         10039 => x"a0065486",
         10040 => x"557382aa",
         10041 => x"38a053a4",
         10042 => x"3d0852a8",
         10043 => x"3dff8805",
         10044 => x"51ffb4ea",
         10045 => x"3fac5377",
         10046 => x"52923d70",
         10047 => x"5254ffb4",
         10048 => x"dd3faa3d",
         10049 => x"08527351",
         10050 => x"cbf73f82",
         10051 => x"b5c80855",
         10052 => x"82b5c808",
         10053 => x"9538636f",
         10054 => x"2e098106",
         10055 => x"883865a2",
         10056 => x"3d082e92",
         10057 => x"38885581",
         10058 => x"e53982b5",
         10059 => x"c808842e",
         10060 => x"09810681",
         10061 => x"b8387351",
         10062 => x"c9b13f82",
         10063 => x"b5c80855",
         10064 => x"82b5c808",
         10065 => x"81c83868",
         10066 => x"569353a8",
         10067 => x"3dff9505",
         10068 => x"528d1651",
         10069 => x"ffb4873f",
         10070 => x"02af0533",
         10071 => x"8b17348b",
         10072 => x"16337084",
         10073 => x"2a708106",
         10074 => x"51555573",
         10075 => x"893874a0",
         10076 => x"0754738b",
         10077 => x"17347854",
         10078 => x"810b8315",
         10079 => x"348b1633",
         10080 => x"70842a70",
         10081 => x"81065155",
         10082 => x"5573802e",
         10083 => x"80e5386e",
         10084 => x"642e80df",
         10085 => x"38755278",
         10086 => x"51c6be3f",
         10087 => x"82b5c808",
         10088 => x"527851ff",
         10089 => x"b7bb3f82",
         10090 => x"5582b5c8",
         10091 => x"08802e80",
         10092 => x"dd3882b5",
         10093 => x"c8085278",
         10094 => x"51ffb5af",
         10095 => x"3f82b5c8",
         10096 => x"087980d4",
         10097 => x"11585855",
         10098 => x"82b5c808",
         10099 => x"80c03881",
         10100 => x"16335473",
         10101 => x"ae2e0981",
         10102 => x"06993863",
         10103 => x"53755276",
         10104 => x"51c6af3f",
         10105 => x"7854810b",
         10106 => x"83153487",
         10107 => x"3982b5c8",
         10108 => x"089c3877",
         10109 => x"51c8ca3f",
         10110 => x"82b5c808",
         10111 => x"5582b5c8",
         10112 => x"088c3878",
         10113 => x"51ffb5aa",
         10114 => x"3f82b5c8",
         10115 => x"08557482",
         10116 => x"b5c80ca8",
         10117 => x"3d0d04ed",
         10118 => x"3d0d0280",
         10119 => x"db053302",
         10120 => x"840580df",
         10121 => x"05335757",
         10122 => x"8253953d",
         10123 => x"d0055296",
         10124 => x"3d51d2e9",
         10125 => x"3f82b5c8",
         10126 => x"085582b5",
         10127 => x"c80880cf",
         10128 => x"38785a65",
         10129 => x"52953dd4",
         10130 => x"0551c9b5",
         10131 => x"3f82b5c8",
         10132 => x"085582b5",
         10133 => x"c808b838",
         10134 => x"0280cf05",
         10135 => x"3381a006",
         10136 => x"54865573",
         10137 => x"aa3875a7",
         10138 => x"06617109",
         10139 => x"8b123371",
         10140 => x"067a7406",
         10141 => x"07515755",
         10142 => x"56748b15",
         10143 => x"34785481",
         10144 => x"0b831534",
         10145 => x"7851ffb4",
         10146 => x"a93f82b5",
         10147 => x"c8085574",
         10148 => x"82b5c80c",
         10149 => x"953d0d04",
         10150 => x"ef3d0d64",
         10151 => x"56825393",
         10152 => x"3dd00552",
         10153 => x"943d51d1",
         10154 => x"f43f82b5",
         10155 => x"c8085582",
         10156 => x"b5c80880",
         10157 => x"cb387658",
         10158 => x"6352933d",
         10159 => x"d40551c8",
         10160 => x"c03f82b5",
         10161 => x"c8085582",
         10162 => x"b5c808b4",
         10163 => x"380280c7",
         10164 => x"053381a0",
         10165 => x"06548655",
         10166 => x"73a63884",
         10167 => x"16228617",
         10168 => x"2271902b",
         10169 => x"07535496",
         10170 => x"1f51ffb0",
         10171 => x"c23f7654",
         10172 => x"810b8315",
         10173 => x"347651ff",
         10174 => x"b3b83f82",
         10175 => x"b5c80855",
         10176 => x"7482b5c8",
         10177 => x"0c933d0d",
         10178 => x"04ea3d0d",
         10179 => x"696b5c5a",
         10180 => x"8053983d",
         10181 => x"d0055299",
         10182 => x"3d51d181",
         10183 => x"3f82b5c8",
         10184 => x"0882b5c8",
         10185 => x"08307082",
         10186 => x"b5c80807",
         10187 => x"80255155",
         10188 => x"5779802e",
         10189 => x"81853881",
         10190 => x"70750655",
         10191 => x"5573802e",
         10192 => x"80f9387b",
         10193 => x"5d805f80",
         10194 => x"528d3d70",
         10195 => x"5254ffbe",
         10196 => x"a93f82b5",
         10197 => x"c8085782",
         10198 => x"b5c80880",
         10199 => x"d1387452",
         10200 => x"7351c3dc",
         10201 => x"3f82b5c8",
         10202 => x"085782b5",
         10203 => x"c808bf38",
         10204 => x"82b5c808",
         10205 => x"82b5c808",
         10206 => x"655b5956",
         10207 => x"78188119",
         10208 => x"7b185659",
         10209 => x"55743374",
         10210 => x"34811656",
         10211 => x"8a7827ec",
         10212 => x"388b5675",
         10213 => x"1a548074",
         10214 => x"3475802e",
         10215 => x"9e38ff16",
         10216 => x"701b7033",
         10217 => x"51555673",
         10218 => x"a02ee838",
         10219 => x"8e397684",
         10220 => x"2e098106",
         10221 => x"8638807a",
         10222 => x"34805776",
         10223 => x"30707807",
         10224 => x"80255154",
         10225 => x"7a802e80",
         10226 => x"c1387380",
         10227 => x"2ebc387b",
         10228 => x"a0110853",
         10229 => x"51ffb193",
         10230 => x"3f82b5c8",
         10231 => x"085782b5",
         10232 => x"c808a738",
         10233 => x"7b703355",
         10234 => x"5580c356",
         10235 => x"73832e8b",
         10236 => x"3880e456",
         10237 => x"73842e83",
         10238 => x"38a75675",
         10239 => x"15b40551",
         10240 => x"ffade33f",
         10241 => x"82b5c808",
         10242 => x"7b0c7682",
         10243 => x"b5c80c98",
         10244 => x"3d0d04e6",
         10245 => x"3d0d8253",
         10246 => x"9c3dffb8",
         10247 => x"05529d3d",
         10248 => x"51cefa3f",
         10249 => x"82b5c808",
         10250 => x"82b5c808",
         10251 => x"565482b5",
         10252 => x"c8088398",
         10253 => x"388b53a0",
         10254 => x"528b3d70",
         10255 => x"5259ffae",
         10256 => x"c03f736d",
         10257 => x"70337081",
         10258 => x"ff065257",
         10259 => x"55579f74",
         10260 => x"2781bc38",
         10261 => x"78587481",
         10262 => x"ff066d81",
         10263 => x"054e7052",
         10264 => x"55ffaf89",
         10265 => x"3f82b5c8",
         10266 => x"08802ea5",
         10267 => x"386c7033",
         10268 => x"70535754",
         10269 => x"ffaefd3f",
         10270 => x"82b5c808",
         10271 => x"802e8d38",
         10272 => x"74882b76",
         10273 => x"076d8105",
         10274 => x"4e558639",
         10275 => x"82b5c808",
         10276 => x"55ff9f15",
         10277 => x"7083ffff",
         10278 => x"06515473",
         10279 => x"99268a38",
         10280 => x"e0157083",
         10281 => x"ffff0656",
         10282 => x"5480ff75",
         10283 => x"27873882",
         10284 => x"ae901533",
         10285 => x"5574802e",
         10286 => x"a3387452",
         10287 => x"82b09051",
         10288 => x"ffae893f",
         10289 => x"82b5c808",
         10290 => x"933881ff",
         10291 => x"75278838",
         10292 => x"76892688",
         10293 => x"388b398a",
         10294 => x"77278638",
         10295 => x"865581ec",
         10296 => x"3981ff75",
         10297 => x"278f3874",
         10298 => x"882a5473",
         10299 => x"78708105",
         10300 => x"5a348117",
         10301 => x"57747870",
         10302 => x"81055a34",
         10303 => x"81176d70",
         10304 => x"337081ff",
         10305 => x"06525755",
         10306 => x"57739f26",
         10307 => x"fec8388b",
         10308 => x"3d335486",
         10309 => x"557381e5",
         10310 => x"2e81b138",
         10311 => x"76802e99",
         10312 => x"3802a705",
         10313 => x"55761570",
         10314 => x"33515473",
         10315 => x"a02e0981",
         10316 => x"068738ff",
         10317 => x"175776ed",
         10318 => x"38794180",
         10319 => x"43805291",
         10320 => x"3d705255",
         10321 => x"ffbab33f",
         10322 => x"82b5c808",
         10323 => x"5482b5c8",
         10324 => x"0880f738",
         10325 => x"81527451",
         10326 => x"ffbfe53f",
         10327 => x"82b5c808",
         10328 => x"5482b5c8",
         10329 => x"088d3876",
         10330 => x"80c43867",
         10331 => x"54e57434",
         10332 => x"80c63982",
         10333 => x"b5c80884",
         10334 => x"2e098106",
         10335 => x"80cc3880",
         10336 => x"5476742e",
         10337 => x"80c43881",
         10338 => x"527451ff",
         10339 => x"bdb03f82",
         10340 => x"b5c80854",
         10341 => x"82b5c808",
         10342 => x"b138a053",
         10343 => x"82b5c808",
         10344 => x"526751ff",
         10345 => x"abdb3f67",
         10346 => x"54880b8b",
         10347 => x"15348b53",
         10348 => x"78526751",
         10349 => x"ffaba73f",
         10350 => x"7954810b",
         10351 => x"83153479",
         10352 => x"51ffadee",
         10353 => x"3f82b5c8",
         10354 => x"08547355",
         10355 => x"7482b5c8",
         10356 => x"0c9c3d0d",
         10357 => x"04f23d0d",
         10358 => x"60620288",
         10359 => x"0580cb05",
         10360 => x"33933dfc",
         10361 => x"05557254",
         10362 => x"405e5ad2",
         10363 => x"da3f82b5",
         10364 => x"c8085882",
         10365 => x"b5c80882",
         10366 => x"bd38911a",
         10367 => x"33587782",
         10368 => x"b5387c80",
         10369 => x"2e97388c",
         10370 => x"1a085978",
         10371 => x"9038901a",
         10372 => x"3370812a",
         10373 => x"70810651",
         10374 => x"55557390",
         10375 => x"38875482",
         10376 => x"97398258",
         10377 => x"82903981",
         10378 => x"58828b39",
         10379 => x"7e8a1122",
         10380 => x"70892b70",
         10381 => x"557f5456",
         10382 => x"5656fec2",
         10383 => x"c63fff14",
         10384 => x"7d067030",
         10385 => x"7072079f",
         10386 => x"2a82b5c8",
         10387 => x"08058c19",
         10388 => x"087c405a",
         10389 => x"5d555581",
         10390 => x"77278838",
         10391 => x"98160877",
         10392 => x"26833882",
         10393 => x"57767756",
         10394 => x"59805674",
         10395 => x"527951ff",
         10396 => x"ae993f81",
         10397 => x"157f5555",
         10398 => x"98140875",
         10399 => x"26833882",
         10400 => x"5582b5c8",
         10401 => x"08812eff",
         10402 => x"993882b5",
         10403 => x"c808ff2e",
         10404 => x"ff953882",
         10405 => x"b5c8088e",
         10406 => x"38811656",
         10407 => x"757b2e09",
         10408 => x"81068738",
         10409 => x"93397459",
         10410 => x"80567477",
         10411 => x"2e098106",
         10412 => x"ffb93887",
         10413 => x"5880ff39",
         10414 => x"7d802eba",
         10415 => x"38787b55",
         10416 => x"557a802e",
         10417 => x"b4388115",
         10418 => x"5673812e",
         10419 => x"09810683",
         10420 => x"38ff5675",
         10421 => x"5374527e",
         10422 => x"51ffafa8",
         10423 => x"3f82b5c8",
         10424 => x"085882b5",
         10425 => x"c80880ce",
         10426 => x"38748116",
         10427 => x"ff165656",
         10428 => x"5c73d338",
         10429 => x"8439ff19",
         10430 => x"5c7e7c8c",
         10431 => x"120c557d",
         10432 => x"802eb338",
         10433 => x"78881b0c",
         10434 => x"7c8c1b0c",
         10435 => x"901a3380",
         10436 => x"c0075473",
         10437 => x"901b3498",
         10438 => x"1508fe05",
         10439 => x"90160857",
         10440 => x"54757426",
         10441 => x"9138757b",
         10442 => x"3190160c",
         10443 => x"84153381",
         10444 => x"07547384",
         10445 => x"16347754",
         10446 => x"7382b5c8",
         10447 => x"0c903d0d",
         10448 => x"04e93d0d",
         10449 => x"6b6d0288",
         10450 => x"0580eb05",
         10451 => x"339d3d54",
         10452 => x"5a5c59c5",
         10453 => x"bd3f8b56",
         10454 => x"800b82b5",
         10455 => x"c808248b",
         10456 => x"f83882b5",
         10457 => x"c8088429",
         10458 => x"82cd8005",
         10459 => x"70085155",
         10460 => x"74802e84",
         10461 => x"38807534",
         10462 => x"82b5c808",
         10463 => x"81ff065f",
         10464 => x"81527e51",
         10465 => x"ffa0d03f",
         10466 => x"82b5c808",
         10467 => x"81ff0670",
         10468 => x"81065657",
         10469 => x"8356748b",
         10470 => x"c0387682",
         10471 => x"2a708106",
         10472 => x"51558a56",
         10473 => x"748bb238",
         10474 => x"993dfc05",
         10475 => x"5383527e",
         10476 => x"51ffa4f0",
         10477 => x"3f82b5c8",
         10478 => x"08993867",
         10479 => x"5574802e",
         10480 => x"92387482",
         10481 => x"8080268b",
         10482 => x"38ff1575",
         10483 => x"06557480",
         10484 => x"2e833881",
         10485 => x"4878802e",
         10486 => x"87388480",
         10487 => x"79269238",
         10488 => x"7881800a",
         10489 => x"268b38ff",
         10490 => x"19790655",
         10491 => x"74802e86",
         10492 => x"3893568a",
         10493 => x"e4397889",
         10494 => x"2a6e892a",
         10495 => x"70892b77",
         10496 => x"59484359",
         10497 => x"7a833881",
         10498 => x"56613070",
         10499 => x"80257707",
         10500 => x"51559156",
         10501 => x"748ac238",
         10502 => x"993df805",
         10503 => x"5381527e",
         10504 => x"51ffa480",
         10505 => x"3f815682",
         10506 => x"b5c8088a",
         10507 => x"ac387783",
         10508 => x"2a707706",
         10509 => x"82b5c808",
         10510 => x"43564574",
         10511 => x"8338bf41",
         10512 => x"66558e56",
         10513 => x"6075268a",
         10514 => x"90387461",
         10515 => x"31704855",
         10516 => x"80ff7527",
         10517 => x"8a833893",
         10518 => x"56788180",
         10519 => x"2689fa38",
         10520 => x"77812a70",
         10521 => x"81065643",
         10522 => x"74802e95",
         10523 => x"38778706",
         10524 => x"5574822e",
         10525 => x"838d3877",
         10526 => x"81065574",
         10527 => x"802e8383",
         10528 => x"38778106",
         10529 => x"55935682",
         10530 => x"5e74802e",
         10531 => x"89cb3878",
         10532 => x"5a7d832e",
         10533 => x"09810680",
         10534 => x"e13878ae",
         10535 => x"3866912a",
         10536 => x"57810b82",
         10537 => x"b0b42256",
         10538 => x"5a74802e",
         10539 => x"9d387477",
         10540 => x"26983882",
         10541 => x"b0b45679",
         10542 => x"10821770",
         10543 => x"2257575a",
         10544 => x"74802e86",
         10545 => x"38767527",
         10546 => x"ee387952",
         10547 => x"6651febd",
         10548 => x"b23f82b5",
         10549 => x"c8088429",
         10550 => x"84870570",
         10551 => x"892a5e55",
         10552 => x"a05c800b",
         10553 => x"82b5c808",
         10554 => x"fc808a05",
         10555 => x"5644fdff",
         10556 => x"f00a7527",
         10557 => x"80ec3888",
         10558 => x"d33978ae",
         10559 => x"38668c2a",
         10560 => x"57810b82",
         10561 => x"b0a42256",
         10562 => x"5a74802e",
         10563 => x"9d387477",
         10564 => x"26983882",
         10565 => x"b0a45679",
         10566 => x"10821770",
         10567 => x"2257575a",
         10568 => x"74802e86",
         10569 => x"38767527",
         10570 => x"ee387952",
         10571 => x"6651febc",
         10572 => x"d23f82b5",
         10573 => x"c8081084",
         10574 => x"055782b5",
         10575 => x"c8089ff5",
         10576 => x"26963881",
         10577 => x"0b82b5c8",
         10578 => x"081082b5",
         10579 => x"c8080571",
         10580 => x"11722a83",
         10581 => x"0559565e",
         10582 => x"83ff1789",
         10583 => x"2a5d815c",
         10584 => x"a044601c",
         10585 => x"7d116505",
         10586 => x"697012ff",
         10587 => x"05713070",
         10588 => x"72067431",
         10589 => x"5c525957",
         10590 => x"59407d83",
         10591 => x"2e098106",
         10592 => x"8938761c",
         10593 => x"6018415c",
         10594 => x"8439761d",
         10595 => x"5d799029",
         10596 => x"18706231",
         10597 => x"68585155",
         10598 => x"74762687",
         10599 => x"af38757c",
         10600 => x"317d317a",
         10601 => x"53706531",
         10602 => x"5255febb",
         10603 => x"d63f82b5",
         10604 => x"c808587d",
         10605 => x"832e0981",
         10606 => x"069b3882",
         10607 => x"b5c80883",
         10608 => x"fff52680",
         10609 => x"dd387887",
         10610 => x"83387981",
         10611 => x"2a5978fd",
         10612 => x"be3886f8",
         10613 => x"397d822e",
         10614 => x"09810680",
         10615 => x"c53883ff",
         10616 => x"f50b82b5",
         10617 => x"c80827a0",
         10618 => x"38788f38",
         10619 => x"791a5574",
         10620 => x"80c02686",
         10621 => x"387459fd",
         10622 => x"96396281",
         10623 => x"06557480",
         10624 => x"2e8f3883",
         10625 => x"5efd8839",
         10626 => x"82b5c808",
         10627 => x"9ff52692",
         10628 => x"387886b8",
         10629 => x"38791a59",
         10630 => x"81807927",
         10631 => x"fcf13886",
         10632 => x"ab398055",
         10633 => x"7d812e09",
         10634 => x"81068338",
         10635 => x"7d559ff5",
         10636 => x"78278b38",
         10637 => x"74810655",
         10638 => x"8e567486",
         10639 => x"9c388480",
         10640 => x"5380527a",
         10641 => x"51ffa2b9",
         10642 => x"3f8b5382",
         10643 => x"aecc527a",
         10644 => x"51ffa28a",
         10645 => x"3f848052",
         10646 => x"8b1b51ff",
         10647 => x"a1b33f79",
         10648 => x"8d1c347b",
         10649 => x"83ffff06",
         10650 => x"528e1b51",
         10651 => x"ffa1a23f",
         10652 => x"810b901c",
         10653 => x"347d8332",
         10654 => x"70307096",
         10655 => x"2a848006",
         10656 => x"54515591",
         10657 => x"1b51ffa1",
         10658 => x"883f6655",
         10659 => x"7483ffff",
         10660 => x"26903874",
         10661 => x"83ffff06",
         10662 => x"52931b51",
         10663 => x"ffa0f23f",
         10664 => x"8a397452",
         10665 => x"a01b51ff",
         10666 => x"a1853ff8",
         10667 => x"0b951c34",
         10668 => x"bf52981b",
         10669 => x"51ffa0d9",
         10670 => x"3f81ff52",
         10671 => x"9a1b51ff",
         10672 => x"a0cf3f60",
         10673 => x"529c1b51",
         10674 => x"ffa0e43f",
         10675 => x"7d832e09",
         10676 => x"810680cb",
         10677 => x"388288b2",
         10678 => x"0a5280c3",
         10679 => x"1b51ffa0",
         10680 => x"ce3f7c52",
         10681 => x"a41b51ff",
         10682 => x"a0c53f82",
         10683 => x"52ac1b51",
         10684 => x"ffa0bc3f",
         10685 => x"8152b01b",
         10686 => x"51ffa095",
         10687 => x"3f8652b2",
         10688 => x"1b51ffa0",
         10689 => x"8c3fff80",
         10690 => x"0b80c01c",
         10691 => x"34a90b80",
         10692 => x"c21c3493",
         10693 => x"5382aed8",
         10694 => x"5280c71b",
         10695 => x"51ae3982",
         10696 => x"88b20a52",
         10697 => x"a71b51ff",
         10698 => x"a0853f7c",
         10699 => x"83ffff06",
         10700 => x"52961b51",
         10701 => x"ff9fda3f",
         10702 => x"ff800ba4",
         10703 => x"1c34a90b",
         10704 => x"a61c3493",
         10705 => x"5382aeec",
         10706 => x"52ab1b51",
         10707 => x"ffa08f3f",
         10708 => x"82d4d552",
         10709 => x"83fe1b70",
         10710 => x"5259ff9f",
         10711 => x"b43f8154",
         10712 => x"60537a52",
         10713 => x"7e51ff9b",
         10714 => x"d73f8156",
         10715 => x"82b5c808",
         10716 => x"83e7387d",
         10717 => x"832e0981",
         10718 => x"0680ee38",
         10719 => x"75546086",
         10720 => x"05537a52",
         10721 => x"7e51ff9b",
         10722 => x"b73f8480",
         10723 => x"5380527a",
         10724 => x"51ff9fed",
         10725 => x"3f848b85",
         10726 => x"a4d2527a",
         10727 => x"51ff9f8f",
         10728 => x"3f868a85",
         10729 => x"e4f25283",
         10730 => x"e41b51ff",
         10731 => x"9f813fff",
         10732 => x"185283e8",
         10733 => x"1b51ff9e",
         10734 => x"f63f8252",
         10735 => x"83ec1b51",
         10736 => x"ff9eec3f",
         10737 => x"82d4d552",
         10738 => x"7851ff9e",
         10739 => x"c43f7554",
         10740 => x"60870553",
         10741 => x"7a527e51",
         10742 => x"ff9ae53f",
         10743 => x"75546016",
         10744 => x"537a527e",
         10745 => x"51ff9ad8",
         10746 => x"3f655380",
         10747 => x"527a51ff",
         10748 => x"9f8f3f7f",
         10749 => x"5680587d",
         10750 => x"832e0981",
         10751 => x"069a38f8",
         10752 => x"527a51ff",
         10753 => x"9ea93fff",
         10754 => x"52841b51",
         10755 => x"ff9ea03f",
         10756 => x"f00a5288",
         10757 => x"1b519139",
         10758 => x"87fffff8",
         10759 => x"557d812e",
         10760 => x"8338f855",
         10761 => x"74527a51",
         10762 => x"ff9e843f",
         10763 => x"7c556157",
         10764 => x"74622683",
         10765 => x"38745776",
         10766 => x"5475537a",
         10767 => x"527e51ff",
         10768 => x"99fe3f82",
         10769 => x"b5c80882",
         10770 => x"87388480",
         10771 => x"5382b5c8",
         10772 => x"08527a51",
         10773 => x"ff9eaa3f",
         10774 => x"76167578",
         10775 => x"31565674",
         10776 => x"cd388118",
         10777 => x"5877802e",
         10778 => x"ff8d3879",
         10779 => x"557d832e",
         10780 => x"83386355",
         10781 => x"61577462",
         10782 => x"26833874",
         10783 => x"57765475",
         10784 => x"537a527e",
         10785 => x"51ff99b8",
         10786 => x"3f82b5c8",
         10787 => x"0881c138",
         10788 => x"76167578",
         10789 => x"31565674",
         10790 => x"db388c56",
         10791 => x"7d832e93",
         10792 => x"38865666",
         10793 => x"83ffff26",
         10794 => x"8a388456",
         10795 => x"7d822e83",
         10796 => x"38815664",
         10797 => x"81065877",
         10798 => x"80fe3884",
         10799 => x"80537752",
         10800 => x"7a51ff9d",
         10801 => x"bc3f82d4",
         10802 => x"d5527851",
         10803 => x"ff9cc23f",
         10804 => x"83be1b55",
         10805 => x"77753481",
         10806 => x"0b811634",
         10807 => x"810b8216",
         10808 => x"34778316",
         10809 => x"34758416",
         10810 => x"34606705",
         10811 => x"5680fdc1",
         10812 => x"527551fe",
         10813 => x"b58d3ffe",
         10814 => x"0b851634",
         10815 => x"82b5c808",
         10816 => x"822abf07",
         10817 => x"56758616",
         10818 => x"3482b5c8",
         10819 => x"08871634",
         10820 => x"605283c6",
         10821 => x"1b51ff9c",
         10822 => x"963f6652",
         10823 => x"83ca1b51",
         10824 => x"ff9c8c3f",
         10825 => x"81547753",
         10826 => x"7a527e51",
         10827 => x"ff98913f",
         10828 => x"815682b5",
         10829 => x"c808a238",
         10830 => x"80538052",
         10831 => x"7e51ff99",
         10832 => x"e33f8156",
         10833 => x"82b5c808",
         10834 => x"90388939",
         10835 => x"8e568a39",
         10836 => x"81568639",
         10837 => x"82b5c808",
         10838 => x"567582b5",
         10839 => x"c80c993d",
         10840 => x"0d04f53d",
         10841 => x"0d7d605b",
         10842 => x"59807960",
         10843 => x"ff055a57",
         10844 => x"57767825",
         10845 => x"b4388d3d",
         10846 => x"f8115555",
         10847 => x"8153fc15",
         10848 => x"527951c9",
         10849 => x"dc3f7a81",
         10850 => x"2e098106",
         10851 => x"9c388c3d",
         10852 => x"3355748d",
         10853 => x"2edb3874",
         10854 => x"76708105",
         10855 => x"58348117",
         10856 => x"57748a2e",
         10857 => x"098106c9",
         10858 => x"38807634",
         10859 => x"78557683",
         10860 => x"38765574",
         10861 => x"82b5c80c",
         10862 => x"8d3d0d04",
         10863 => x"f73d0d7b",
         10864 => x"028405b3",
         10865 => x"05335957",
         10866 => x"778a2e09",
         10867 => x"81068738",
         10868 => x"8d527651",
         10869 => x"e73f8417",
         10870 => x"08568076",
         10871 => x"24be3888",
         10872 => x"17087717",
         10873 => x"8c055659",
         10874 => x"77753481",
         10875 => x"1656bb76",
         10876 => x"25a1388b",
         10877 => x"3dfc0554",
         10878 => x"75538c17",
         10879 => x"52760851",
         10880 => x"cbdc3f79",
         10881 => x"76327030",
         10882 => x"7072079f",
         10883 => x"2a703053",
         10884 => x"51565675",
         10885 => x"84180c81",
         10886 => x"1988180c",
         10887 => x"8b3d0d04",
         10888 => x"f93d0d79",
         10889 => x"84110856",
         10890 => x"56807524",
         10891 => x"a738893d",
         10892 => x"fc055474",
         10893 => x"538c1652",
         10894 => x"750851cb",
         10895 => x"a13f82b5",
         10896 => x"c8089138",
         10897 => x"84160878",
         10898 => x"2e098106",
         10899 => x"87388816",
         10900 => x"08558339",
         10901 => x"ff557482",
         10902 => x"b5c80c89",
         10903 => x"3d0d04fd",
         10904 => x"3d0d7554",
         10905 => x"80cc5380",
         10906 => x"527351ff",
         10907 => x"9a933f76",
         10908 => x"740c853d",
         10909 => x"0d04ea3d",
         10910 => x"0d0280e3",
         10911 => x"05336a53",
         10912 => x"863d7053",
         10913 => x"5454d83f",
         10914 => x"73527251",
         10915 => x"feae3f72",
         10916 => x"51ff8d3f",
         10917 => x"983d0d04",
         10918 => x"00ffffff",
         10919 => x"ff00ffff",
         10920 => x"ffff00ff",
         10921 => x"ffffff00",
         10922 => x"00002baa",
         10923 => x"00002b2e",
         10924 => x"00002b35",
         10925 => x"00002b3c",
         10926 => x"00002b43",
         10927 => x"00002b4a",
         10928 => x"00002b51",
         10929 => x"00002b58",
         10930 => x"00002b5f",
         10931 => x"00002b66",
         10932 => x"00002b6d",
         10933 => x"00002b74",
         10934 => x"00002b7a",
         10935 => x"00002b80",
         10936 => x"00002b86",
         10937 => x"00002b8c",
         10938 => x"00002b92",
         10939 => x"00002b98",
         10940 => x"00002b9e",
         10941 => x"00002ba4",
         10942 => x"0000414f",
         10943 => x"00004155",
         10944 => x"0000415b",
         10945 => x"00004161",
         10946 => x"00004167",
         10947 => x"00004745",
         10948 => x"00004845",
         10949 => x"00004956",
         10950 => x"00004bae",
         10951 => x"0000482d",
         10952 => x"0000461a",
         10953 => x"00004a1e",
         10954 => x"00004b7f",
         10955 => x"00004a61",
         10956 => x"00004af7",
         10957 => x"00004a7d",
         10958 => x"00004900",
         10959 => x"0000461a",
         10960 => x"00004956",
         10961 => x"0000497f",
         10962 => x"00004a1e",
         10963 => x"0000461a",
         10964 => x"0000461a",
         10965 => x"00004a7d",
         10966 => x"00004af7",
         10967 => x"00004b7f",
         10968 => x"00004bae",
         10969 => x"00000e31",
         10970 => x"0000171a",
         10971 => x"0000171a",
         10972 => x"00000e60",
         10973 => x"0000171a",
         10974 => x"0000171a",
         10975 => x"0000171a",
         10976 => x"0000171a",
         10977 => x"0000171a",
         10978 => x"0000171a",
         10979 => x"0000171a",
         10980 => x"00000e1d",
         10981 => x"0000171a",
         10982 => x"00000e48",
         10983 => x"00000e78",
         10984 => x"0000171a",
         10985 => x"0000171a",
         10986 => x"0000171a",
         10987 => x"0000171a",
         10988 => x"0000171a",
         10989 => x"0000171a",
         10990 => x"0000171a",
         10991 => x"0000171a",
         10992 => x"0000171a",
         10993 => x"0000171a",
         10994 => x"0000171a",
         10995 => x"0000171a",
         10996 => x"0000171a",
         10997 => x"0000171a",
         10998 => x"0000171a",
         10999 => x"0000171a",
         11000 => x"0000171a",
         11001 => x"0000171a",
         11002 => x"0000171a",
         11003 => x"0000171a",
         11004 => x"0000171a",
         11005 => x"0000171a",
         11006 => x"0000171a",
         11007 => x"0000171a",
         11008 => x"0000171a",
         11009 => x"0000171a",
         11010 => x"0000171a",
         11011 => x"0000171a",
         11012 => x"0000171a",
         11013 => x"0000171a",
         11014 => x"0000171a",
         11015 => x"0000171a",
         11016 => x"0000171a",
         11017 => x"0000171a",
         11018 => x"0000171a",
         11019 => x"0000171a",
         11020 => x"00000fa8",
         11021 => x"0000171a",
         11022 => x"0000171a",
         11023 => x"0000171a",
         11024 => x"0000171a",
         11025 => x"00001116",
         11026 => x"0000171a",
         11027 => x"0000171a",
         11028 => x"0000171a",
         11029 => x"0000171a",
         11030 => x"0000171a",
         11031 => x"0000171a",
         11032 => x"0000171a",
         11033 => x"0000171a",
         11034 => x"0000171a",
         11035 => x"0000171a",
         11036 => x"00000ed8",
         11037 => x"0000103f",
         11038 => x"00000eaf",
         11039 => x"00000eaf",
         11040 => x"00000eaf",
         11041 => x"0000171a",
         11042 => x"0000103f",
         11043 => x"0000171a",
         11044 => x"0000171a",
         11045 => x"00000e98",
         11046 => x"0000171a",
         11047 => x"0000171a",
         11048 => x"000010ec",
         11049 => x"000010f7",
         11050 => x"0000171a",
         11051 => x"0000171a",
         11052 => x"00000f11",
         11053 => x"0000171a",
         11054 => x"0000111f",
         11055 => x"0000171a",
         11056 => x"0000171a",
         11057 => x"00001116",
         11058 => x"64696e69",
         11059 => x"74000000",
         11060 => x"64696f63",
         11061 => x"746c0000",
         11062 => x"66696e69",
         11063 => x"74000000",
         11064 => x"666c6f61",
         11065 => x"64000000",
         11066 => x"66657865",
         11067 => x"63000000",
         11068 => x"6d636c65",
         11069 => x"61720000",
         11070 => x"6d636f70",
         11071 => x"79000000",
         11072 => x"6d646966",
         11073 => x"66000000",
         11074 => x"6d64756d",
         11075 => x"70000000",
         11076 => x"6d656200",
         11077 => x"6d656800",
         11078 => x"6d657700",
         11079 => x"68696400",
         11080 => x"68696500",
         11081 => x"68666400",
         11082 => x"68666500",
         11083 => x"63616c6c",
         11084 => x"00000000",
         11085 => x"6a6d7000",
         11086 => x"72657374",
         11087 => x"61727400",
         11088 => x"72657365",
         11089 => x"74000000",
         11090 => x"696e666f",
         11091 => x"00000000",
         11092 => x"74657374",
         11093 => x"00000000",
         11094 => x"74626173",
         11095 => x"69630000",
         11096 => x"6d626173",
         11097 => x"69630000",
         11098 => x"6b696c6f",
         11099 => x"00000000",
         11100 => x"65640000",
         11101 => x"4469736b",
         11102 => x"20457272",
         11103 => x"6f720000",
         11104 => x"496e7465",
         11105 => x"726e616c",
         11106 => x"20657272",
         11107 => x"6f722e00",
         11108 => x"4469736b",
         11109 => x"206e6f74",
         11110 => x"20726561",
         11111 => x"64792e00",
         11112 => x"4e6f2066",
         11113 => x"696c6520",
         11114 => x"666f756e",
         11115 => x"642e0000",
         11116 => x"4e6f2070",
         11117 => x"61746820",
         11118 => x"666f756e",
         11119 => x"642e0000",
         11120 => x"496e7661",
         11121 => x"6c696420",
         11122 => x"66696c65",
         11123 => x"6e616d65",
         11124 => x"2e000000",
         11125 => x"41636365",
         11126 => x"73732064",
         11127 => x"656e6965",
         11128 => x"642e0000",
         11129 => x"46696c65",
         11130 => x"20616c72",
         11131 => x"65616479",
         11132 => x"20657869",
         11133 => x"7374732e",
         11134 => x"00000000",
         11135 => x"46696c65",
         11136 => x"2068616e",
         11137 => x"646c6520",
         11138 => x"696e7661",
         11139 => x"6c69642e",
         11140 => x"00000000",
         11141 => x"53442069",
         11142 => x"73207772",
         11143 => x"69746520",
         11144 => x"70726f74",
         11145 => x"65637465",
         11146 => x"642e0000",
         11147 => x"44726976",
         11148 => x"65206e75",
         11149 => x"6d626572",
         11150 => x"20697320",
         11151 => x"696e7661",
         11152 => x"6c69642e",
         11153 => x"00000000",
         11154 => x"4469736b",
         11155 => x"206e6f74",
         11156 => x"20656e61",
         11157 => x"626c6564",
         11158 => x"2e000000",
         11159 => x"4e6f2063",
         11160 => x"6f6d7061",
         11161 => x"7469626c",
         11162 => x"65206669",
         11163 => x"6c657379",
         11164 => x"7374656d",
         11165 => x"20666f75",
         11166 => x"6e64206f",
         11167 => x"6e206469",
         11168 => x"736b2e00",
         11169 => x"466f726d",
         11170 => x"61742061",
         11171 => x"626f7274",
         11172 => x"65642e00",
         11173 => x"54696d65",
         11174 => x"6f75742c",
         11175 => x"206f7065",
         11176 => x"72617469",
         11177 => x"6f6e2063",
         11178 => x"616e6365",
         11179 => x"6c6c6564",
         11180 => x"2e000000",
         11181 => x"46696c65",
         11182 => x"20697320",
         11183 => x"6c6f636b",
         11184 => x"65642e00",
         11185 => x"496e7375",
         11186 => x"66666963",
         11187 => x"69656e74",
         11188 => x"206d656d",
         11189 => x"6f72792e",
         11190 => x"00000000",
         11191 => x"546f6f20",
         11192 => x"6d616e79",
         11193 => x"206f7065",
         11194 => x"6e206669",
         11195 => x"6c65732e",
         11196 => x"00000000",
         11197 => x"50617261",
         11198 => x"6d657465",
         11199 => x"72732069",
         11200 => x"6e636f72",
         11201 => x"72656374",
         11202 => x"2e000000",
         11203 => x"53756363",
         11204 => x"6573732e",
         11205 => x"00000000",
         11206 => x"556e6b6e",
         11207 => x"6f776e20",
         11208 => x"6572726f",
         11209 => x"722e0000",
         11210 => x"0a256c75",
         11211 => x"20627974",
         11212 => x"65732025",
         11213 => x"73206174",
         11214 => x"20256c75",
         11215 => x"20627974",
         11216 => x"65732f73",
         11217 => x"65632e0a",
         11218 => x"00000000",
         11219 => x"72656164",
         11220 => x"00000000",
         11221 => x"2530386c",
         11222 => x"58000000",
         11223 => x"3a202000",
         11224 => x"25303458",
         11225 => x"00000000",
         11226 => x"20202020",
         11227 => x"20202020",
         11228 => x"00000000",
         11229 => x"25303258",
         11230 => x"00000000",
         11231 => x"20200000",
         11232 => x"207c0000",
         11233 => x"7c000000",
         11234 => x"7a4f5300",
         11235 => x"0a2a2a20",
         11236 => x"25732028",
         11237 => x"00000000",
         11238 => x"30322f30",
         11239 => x"352f3230",
         11240 => x"32300000",
         11241 => x"76312e30",
         11242 => x"32000000",
         11243 => x"205a5055",
         11244 => x"2c207265",
         11245 => x"76202530",
         11246 => x"32782920",
         11247 => x"25732025",
         11248 => x"73202a2a",
         11249 => x"0a0a0000",
         11250 => x"5a505520",
         11251 => x"496e7465",
         11252 => x"72727570",
         11253 => x"74204861",
         11254 => x"6e646c65",
         11255 => x"72000000",
         11256 => x"54696d65",
         11257 => x"7220696e",
         11258 => x"74657272",
         11259 => x"75707400",
         11260 => x"50533220",
         11261 => x"696e7465",
         11262 => x"72727570",
         11263 => x"74000000",
         11264 => x"494f4354",
         11265 => x"4c205244",
         11266 => x"20696e74",
         11267 => x"65727275",
         11268 => x"70740000",
         11269 => x"494f4354",
         11270 => x"4c205752",
         11271 => x"20696e74",
         11272 => x"65727275",
         11273 => x"70740000",
         11274 => x"55415254",
         11275 => x"30205258",
         11276 => x"20696e74",
         11277 => x"65727275",
         11278 => x"70740000",
         11279 => x"55415254",
         11280 => x"30205458",
         11281 => x"20696e74",
         11282 => x"65727275",
         11283 => x"70740000",
         11284 => x"55415254",
         11285 => x"31205258",
         11286 => x"20696e74",
         11287 => x"65727275",
         11288 => x"70740000",
         11289 => x"55415254",
         11290 => x"31205458",
         11291 => x"20696e74",
         11292 => x"65727275",
         11293 => x"70740000",
         11294 => x"53657474",
         11295 => x"696e6720",
         11296 => x"75702074",
         11297 => x"696d6572",
         11298 => x"2e2e2e00",
         11299 => x"456e6162",
         11300 => x"6c696e67",
         11301 => x"2074696d",
         11302 => x"65722e2e",
         11303 => x"2e000000",
         11304 => x"6175746f",
         11305 => x"65786563",
         11306 => x"2e626174",
         11307 => x"00000000",
         11308 => x"7a4f532e",
         11309 => x"68737400",
         11310 => x"303a0000",
         11311 => x"4661696c",
         11312 => x"65642074",
         11313 => x"6f20696e",
         11314 => x"69746961",
         11315 => x"6c697365",
         11316 => x"20736420",
         11317 => x"63617264",
         11318 => x"20302c20",
         11319 => x"706c6561",
         11320 => x"73652069",
         11321 => x"6e697420",
         11322 => x"6d616e75",
         11323 => x"616c6c79",
         11324 => x"2e000000",
         11325 => x"2a200000",
         11326 => x"436c6561",
         11327 => x"72696e67",
         11328 => x"2e2e2e2e",
         11329 => x"00000000",
         11330 => x"436f7079",
         11331 => x"696e672e",
         11332 => x"2e2e0000",
         11333 => x"436f6d70",
         11334 => x"6172696e",
         11335 => x"672e2e2e",
         11336 => x"00000000",
         11337 => x"2530386c",
         11338 => x"78282530",
         11339 => x"3878292d",
         11340 => x"3e253038",
         11341 => x"6c782825",
         11342 => x"30387829",
         11343 => x"0a000000",
         11344 => x"44756d70",
         11345 => x"204d656d",
         11346 => x"6f727900",
         11347 => x"0a436f6d",
         11348 => x"706c6574",
         11349 => x"652e0000",
         11350 => x"2530386c",
         11351 => x"58202530",
         11352 => x"32582d00",
         11353 => x"3f3f3f00",
         11354 => x"2530386c",
         11355 => x"58202530",
         11356 => x"34582d00",
         11357 => x"2530386c",
         11358 => x"58202530",
         11359 => x"386c582d",
         11360 => x"00000000",
         11361 => x"45786563",
         11362 => x"7574696e",
         11363 => x"6720636f",
         11364 => x"64652040",
         11365 => x"20253038",
         11366 => x"6c78202e",
         11367 => x"2e2e0a00",
         11368 => x"43616c6c",
         11369 => x"696e6720",
         11370 => x"636f6465",
         11371 => x"20402025",
         11372 => x"30386c78",
         11373 => x"202e2e2e",
         11374 => x"0a000000",
         11375 => x"43616c6c",
         11376 => x"20726574",
         11377 => x"75726e65",
         11378 => x"6420636f",
         11379 => x"64652028",
         11380 => x"2564292e",
         11381 => x"0a000000",
         11382 => x"52657374",
         11383 => x"61727469",
         11384 => x"6e672061",
         11385 => x"70706c69",
         11386 => x"63617469",
         11387 => x"6f6e2e2e",
         11388 => x"2e000000",
         11389 => x"436f6c64",
         11390 => x"20726562",
         11391 => x"6f6f7469",
         11392 => x"6e672e2e",
         11393 => x"2e000000",
         11394 => x"5a505500",
         11395 => x"62696e00",
         11396 => x"25643a5c",
         11397 => x"25735c25",
         11398 => x"732e2573",
         11399 => x"00000000",
         11400 => x"25643a5c",
         11401 => x"25735c25",
         11402 => x"73000000",
         11403 => x"25643a5c",
         11404 => x"25730000",
         11405 => x"42616420",
         11406 => x"636f6d6d",
         11407 => x"616e642e",
         11408 => x"00000000",
         11409 => x"52756e6e",
         11410 => x"696e672e",
         11411 => x"2e2e0000",
         11412 => x"456e6162",
         11413 => x"6c696e67",
         11414 => x"20696e74",
         11415 => x"65727275",
         11416 => x"7074732e",
         11417 => x"2e2e0000",
         11418 => x"25642f25",
         11419 => x"642f2564",
         11420 => x"2025643a",
         11421 => x"25643a25",
         11422 => x"642e2564",
         11423 => x"25640a00",
         11424 => x"536f4320",
         11425 => x"436f6e66",
         11426 => x"69677572",
         11427 => x"6174696f",
         11428 => x"6e000000",
         11429 => x"20286672",
         11430 => x"6f6d2053",
         11431 => x"6f432063",
         11432 => x"6f6e6669",
         11433 => x"67290000",
         11434 => x"3a0a4465",
         11435 => x"76696365",
         11436 => x"7320696d",
         11437 => x"706c656d",
         11438 => x"656e7465",
         11439 => x"643a0a00",
         11440 => x"20202020",
         11441 => x"57422053",
         11442 => x"4452414d",
         11443 => x"20202825",
         11444 => x"3038583a",
         11445 => x"25303858",
         11446 => x"292e0a00",
         11447 => x"20202020",
         11448 => x"53445241",
         11449 => x"4d202020",
         11450 => x"20202825",
         11451 => x"3038583a",
         11452 => x"25303858",
         11453 => x"292e0a00",
         11454 => x"20202020",
         11455 => x"494e534e",
         11456 => x"20425241",
         11457 => x"4d202825",
         11458 => x"3038583a",
         11459 => x"25303858",
         11460 => x"292e0a00",
         11461 => x"20202020",
         11462 => x"4252414d",
         11463 => x"20202020",
         11464 => x"20202825",
         11465 => x"3038583a",
         11466 => x"25303858",
         11467 => x"292e0a00",
         11468 => x"20202020",
         11469 => x"52414d20",
         11470 => x"20202020",
         11471 => x"20202825",
         11472 => x"3038583a",
         11473 => x"25303858",
         11474 => x"292e0a00",
         11475 => x"20202020",
         11476 => x"53442043",
         11477 => x"41524420",
         11478 => x"20202844",
         11479 => x"65766963",
         11480 => x"6573203d",
         11481 => x"25303264",
         11482 => x"292e0a00",
         11483 => x"20202020",
         11484 => x"54494d45",
         11485 => x"52312020",
         11486 => x"20202854",
         11487 => x"696d6572",
         11488 => x"7320203d",
         11489 => x"25303264",
         11490 => x"292e0a00",
         11491 => x"20202020",
         11492 => x"494e5452",
         11493 => x"20435452",
         11494 => x"4c202843",
         11495 => x"68616e6e",
         11496 => x"656c733d",
         11497 => x"25303264",
         11498 => x"292e0a00",
         11499 => x"20202020",
         11500 => x"57495348",
         11501 => x"424f4e45",
         11502 => x"20425553",
         11503 => x"0a000000",
         11504 => x"20202020",
         11505 => x"57422049",
         11506 => x"32430a00",
         11507 => x"20202020",
         11508 => x"494f4354",
         11509 => x"4c0a0000",
         11510 => x"20202020",
         11511 => x"5053320a",
         11512 => x"00000000",
         11513 => x"20202020",
         11514 => x"5350490a",
         11515 => x"00000000",
         11516 => x"41646472",
         11517 => x"65737365",
         11518 => x"733a0a00",
         11519 => x"20202020",
         11520 => x"43505520",
         11521 => x"52657365",
         11522 => x"74205665",
         11523 => x"63746f72",
         11524 => x"20416464",
         11525 => x"72657373",
         11526 => x"203d2025",
         11527 => x"3038580a",
         11528 => x"00000000",
         11529 => x"20202020",
         11530 => x"43505520",
         11531 => x"4d656d6f",
         11532 => x"72792053",
         11533 => x"74617274",
         11534 => x"20416464",
         11535 => x"72657373",
         11536 => x"203d2025",
         11537 => x"3038580a",
         11538 => x"00000000",
         11539 => x"20202020",
         11540 => x"53746163",
         11541 => x"6b205374",
         11542 => x"61727420",
         11543 => x"41646472",
         11544 => x"65737320",
         11545 => x"20202020",
         11546 => x"203d2025",
         11547 => x"3038580a",
         11548 => x"00000000",
         11549 => x"4d697363",
         11550 => x"3a0a0000",
         11551 => x"20202020",
         11552 => x"5a505520",
         11553 => x"49642020",
         11554 => x"20202020",
         11555 => x"20202020",
         11556 => x"20202020",
         11557 => x"20202020",
         11558 => x"203d2025",
         11559 => x"3034580a",
         11560 => x"00000000",
         11561 => x"20202020",
         11562 => x"53797374",
         11563 => x"656d2043",
         11564 => x"6c6f636b",
         11565 => x"20467265",
         11566 => x"71202020",
         11567 => x"20202020",
         11568 => x"203d2025",
         11569 => x"642e2530",
         11570 => x"34644d48",
         11571 => x"7a0a0000",
         11572 => x"20202020",
         11573 => x"53445241",
         11574 => x"4d20436c",
         11575 => x"6f636b20",
         11576 => x"46726571",
         11577 => x"20202020",
         11578 => x"20202020",
         11579 => x"203d2025",
         11580 => x"642e2530",
         11581 => x"34644d48",
         11582 => x"7a0a0000",
         11583 => x"20202020",
         11584 => x"57697368",
         11585 => x"626f6e65",
         11586 => x"20534452",
         11587 => x"414d2043",
         11588 => x"6c6f636b",
         11589 => x"20467265",
         11590 => x"713d2025",
         11591 => x"642e2530",
         11592 => x"34644d48",
         11593 => x"7a0a0000",
         11594 => x"536d616c",
         11595 => x"6c000000",
         11596 => x"4d656469",
         11597 => x"756d0000",
         11598 => x"466c6578",
         11599 => x"00000000",
         11600 => x"45564f00",
         11601 => x"45564f6d",
         11602 => x"696e0000",
         11603 => x"556e6b6e",
         11604 => x"6f776e00",
         11605 => x"000096b0",
         11606 => x"01000000",
         11607 => x"00000002",
         11608 => x"000096ac",
         11609 => x"01000000",
         11610 => x"00000003",
         11611 => x"000096a8",
         11612 => x"01000000",
         11613 => x"00000004",
         11614 => x"000096a4",
         11615 => x"01000000",
         11616 => x"00000005",
         11617 => x"000096a0",
         11618 => x"01000000",
         11619 => x"00000006",
         11620 => x"0000969c",
         11621 => x"01000000",
         11622 => x"00000007",
         11623 => x"00009698",
         11624 => x"01000000",
         11625 => x"00000001",
         11626 => x"00009694",
         11627 => x"01000000",
         11628 => x"00000008",
         11629 => x"00009690",
         11630 => x"01000000",
         11631 => x"0000000b",
         11632 => x"0000968c",
         11633 => x"01000000",
         11634 => x"00000009",
         11635 => x"00009688",
         11636 => x"01000000",
         11637 => x"0000000a",
         11638 => x"00009684",
         11639 => x"04000000",
         11640 => x"0000000d",
         11641 => x"00009680",
         11642 => x"04000000",
         11643 => x"0000000c",
         11644 => x"0000967c",
         11645 => x"04000000",
         11646 => x"0000000e",
         11647 => x"00009678",
         11648 => x"03000000",
         11649 => x"0000000f",
         11650 => x"00009674",
         11651 => x"04000000",
         11652 => x"0000000f",
         11653 => x"00009670",
         11654 => x"04000000",
         11655 => x"00000010",
         11656 => x"0000966c",
         11657 => x"04000000",
         11658 => x"00000011",
         11659 => x"00009668",
         11660 => x"03000000",
         11661 => x"00000012",
         11662 => x"00009664",
         11663 => x"03000000",
         11664 => x"00000013",
         11665 => x"00009660",
         11666 => x"03000000",
         11667 => x"00000014",
         11668 => x"0000965c",
         11669 => x"03000000",
         11670 => x"00000015",
         11671 => x"1b5b4400",
         11672 => x"1b5b4300",
         11673 => x"1b5b4200",
         11674 => x"1b5b4100",
         11675 => x"1b5b367e",
         11676 => x"1b5b357e",
         11677 => x"1b5b347e",
         11678 => x"1b304600",
         11679 => x"1b5b337e",
         11680 => x"1b5b327e",
         11681 => x"1b5b317e",
         11682 => x"10000000",
         11683 => x"0e000000",
         11684 => x"0d000000",
         11685 => x"0b000000",
         11686 => x"08000000",
         11687 => x"06000000",
         11688 => x"05000000",
         11689 => x"04000000",
         11690 => x"03000000",
         11691 => x"02000000",
         11692 => x"01000000",
         11693 => x"68697374",
         11694 => x"6f727900",
         11695 => x"68697374",
         11696 => x"00000000",
         11697 => x"21000000",
         11698 => x"2530346c",
         11699 => x"75202025",
         11700 => x"730a0000",
         11701 => x"4661696c",
         11702 => x"65642074",
         11703 => x"6f207265",
         11704 => x"73657420",
         11705 => x"74686520",
         11706 => x"68697374",
         11707 => x"6f727920",
         11708 => x"66696c65",
         11709 => x"20746f20",
         11710 => x"454f462e",
         11711 => x"00000000",
         11712 => x"43616e6e",
         11713 => x"6f74206f",
         11714 => x"70656e2f",
         11715 => x"63726561",
         11716 => x"74652068",
         11717 => x"6973746f",
         11718 => x"72792066",
         11719 => x"696c652c",
         11720 => x"20646973",
         11721 => x"61626c69",
         11722 => x"6e672e00",
         11723 => x"53440000",
         11724 => x"222a2b2c",
         11725 => x"3a3b3c3d",
         11726 => x"3e3f5b5d",
         11727 => x"7c7f0000",
         11728 => x"46415400",
         11729 => x"46415433",
         11730 => x"32000000",
         11731 => x"ebfe904d",
         11732 => x"53444f53",
         11733 => x"352e3000",
         11734 => x"4e4f204e",
         11735 => x"414d4520",
         11736 => x"20202046",
         11737 => x"41543332",
         11738 => x"20202000",
         11739 => x"4e4f204e",
         11740 => x"414d4520",
         11741 => x"20202046",
         11742 => x"41542020",
         11743 => x"20202000",
         11744 => x"0000972c",
         11745 => x"00000000",
         11746 => x"00000000",
         11747 => x"00000000",
         11748 => x"809a4541",
         11749 => x"8e418f80",
         11750 => x"45454549",
         11751 => x"49498e8f",
         11752 => x"9092924f",
         11753 => x"994f5555",
         11754 => x"59999a9b",
         11755 => x"9c9d9e9f",
         11756 => x"41494f55",
         11757 => x"a5a5a6a7",
         11758 => x"a8a9aaab",
         11759 => x"acadaeaf",
         11760 => x"b0b1b2b3",
         11761 => x"b4b5b6b7",
         11762 => x"b8b9babb",
         11763 => x"bcbdbebf",
         11764 => x"c0c1c2c3",
         11765 => x"c4c5c6c7",
         11766 => x"c8c9cacb",
         11767 => x"cccdcecf",
         11768 => x"d0d1d2d3",
         11769 => x"d4d5d6d7",
         11770 => x"d8d9dadb",
         11771 => x"dcdddedf",
         11772 => x"e0e1e2e3",
         11773 => x"e4e5e6e7",
         11774 => x"e8e9eaeb",
         11775 => x"ecedeeef",
         11776 => x"f0f1f2f3",
         11777 => x"f4f5f6f7",
         11778 => x"f8f9fafb",
         11779 => x"fcfdfeff",
         11780 => x"2b2e2c3b",
         11781 => x"3d5b5d2f",
         11782 => x"5c222a3a",
         11783 => x"3c3e3f7c",
         11784 => x"7f000000",
         11785 => x"00010004",
         11786 => x"00100040",
         11787 => x"01000200",
         11788 => x"00000000",
         11789 => x"00010002",
         11790 => x"00040008",
         11791 => x"00100020",
         11792 => x"00000000",
         11793 => x"00000000",
         11794 => x"00008cc8",
         11795 => x"01020100",
         11796 => x"00000000",
         11797 => x"00000000",
         11798 => x"00008cd0",
         11799 => x"01040100",
         11800 => x"00000000",
         11801 => x"00000000",
         11802 => x"00008cd8",
         11803 => x"01140300",
         11804 => x"00000000",
         11805 => x"00000000",
         11806 => x"00008ce0",
         11807 => x"012b0300",
         11808 => x"00000000",
         11809 => x"00000000",
         11810 => x"00008ce8",
         11811 => x"01300300",
         11812 => x"00000000",
         11813 => x"00000000",
         11814 => x"00008cf0",
         11815 => x"013c0400",
         11816 => x"00000000",
         11817 => x"00000000",
         11818 => x"00008cf8",
         11819 => x"013d0400",
         11820 => x"00000000",
         11821 => x"00000000",
         11822 => x"00008d00",
         11823 => x"013f0400",
         11824 => x"00000000",
         11825 => x"00000000",
         11826 => x"00008d08",
         11827 => x"01400400",
         11828 => x"00000000",
         11829 => x"00000000",
         11830 => x"00008d10",
         11831 => x"01410400",
         11832 => x"00000000",
         11833 => x"00000000",
         11834 => x"00008d14",
         11835 => x"01420400",
         11836 => x"00000000",
         11837 => x"00000000",
         11838 => x"00008d18",
         11839 => x"01430400",
         11840 => x"00000000",
         11841 => x"00000000",
         11842 => x"00008d1c",
         11843 => x"01500500",
         11844 => x"00000000",
         11845 => x"00000000",
         11846 => x"00008d20",
         11847 => x"01510500",
         11848 => x"00000000",
         11849 => x"00000000",
         11850 => x"00008d24",
         11851 => x"01540500",
         11852 => x"00000000",
         11853 => x"00000000",
         11854 => x"00008d28",
         11855 => x"01550500",
         11856 => x"00000000",
         11857 => x"00000000",
         11858 => x"00008d2c",
         11859 => x"01790700",
         11860 => x"00000000",
         11861 => x"00000000",
         11862 => x"00008d34",
         11863 => x"01780700",
         11864 => x"00000000",
         11865 => x"00000000",
         11866 => x"00008d38",
         11867 => x"01820800",
         11868 => x"00000000",
         11869 => x"00000000",
         11870 => x"00008d40",
         11871 => x"01830800",
         11872 => x"00000000",
         11873 => x"00000000",
         11874 => x"00008d48",
         11875 => x"01850800",
         11876 => x"00000000",
         11877 => x"00000000",
         11878 => x"00008d50",
         11879 => x"01870800",
         11880 => x"00000000",
         11881 => x"00000000",
         11882 => x"00008d58",
         11883 => x"018c0900",
         11884 => x"00000000",
         11885 => x"00000000",
         11886 => x"00008d60",
         11887 => x"018d0900",
         11888 => x"00000000",
         11889 => x"00000000",
         11890 => x"00008d68",
         11891 => x"018e0900",
         11892 => x"00000000",
         11893 => x"00000000",
         11894 => x"00008d70",
         11895 => x"018f0900",
         11896 => x"00000000",
         11897 => x"00000000",
         11898 => x"00000000",
         11899 => x"00000000",
         11900 => x"00007fff",
         11901 => x"00000000",
         11902 => x"00007fff",
         11903 => x"00010000",
         11904 => x"00007fff",
         11905 => x"00010000",
         11906 => x"00810000",
         11907 => x"01000000",
         11908 => x"017fffff",
         11909 => x"00000000",
         11910 => x"00000000",
         11911 => x"00007800",
         11912 => x"00000000",
         11913 => x"05f5e100",
         11914 => x"05f5e100",
         11915 => x"05f5e100",
         11916 => x"00000000",
         11917 => x"01010101",
         11918 => x"01010101",
         11919 => x"01011001",
         11920 => x"01000000",
         11921 => x"00000000",
         11922 => x"00000000",
         11923 => x"00000000",
         11924 => x"00000000",
         11925 => x"00000000",
         11926 => x"00000000",
         11927 => x"00000000",
         11928 => x"00000000",
         11929 => x"00000000",
         11930 => x"00000000",
         11931 => x"00000000",
         11932 => x"00000000",
         11933 => x"00000000",
         11934 => x"00000000",
         11935 => x"00000000",
         11936 => x"00000000",
         11937 => x"00000000",
         11938 => x"00000000",
         11939 => x"00000000",
         11940 => x"00000000",
         11941 => x"00000000",
         11942 => x"00000000",
         11943 => x"00000000",
         11944 => x"00000000",
         11945 => x"000096b4",
         11946 => x"01000000",
         11947 => x"000096bc",
         11948 => x"01000000",
         11949 => x"000096c4",
         11950 => x"02000000",
         11951 => x"00000000",
         11952 => x"00000000",
         11953 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

