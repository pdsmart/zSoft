-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b83ff",
             1 => x"f80d0b0b",
             2 => x"0b93b904",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"9d040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b9380",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b8295",
           162 => x"98738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93850400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b80c3",
           171 => x"f42d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b80c5",
           179 => x"e02d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"95040b0b",
           269 => x"0b8ca404",
           270 => x"0b0b0b8c",
           271 => x"b3040b0b",
           272 => x"0b8cc204",
           273 => x"0b0b0b8c",
           274 => x"d1040b0b",
           275 => x"0b8ce004",
           276 => x"0b0b0b8c",
           277 => x"f0040b0b",
           278 => x"0b8d8004",
           279 => x"0b0b0b8d",
           280 => x"8f040b0b",
           281 => x"0b8d9e04",
           282 => x"0b0b0b8d",
           283 => x"ad040b0b",
           284 => x"0b8dbd04",
           285 => x"0b0b0b8d",
           286 => x"cd040b0b",
           287 => x"0b8ddd04",
           288 => x"0b0b0b8d",
           289 => x"ed040b0b",
           290 => x"0b8dfd04",
           291 => x"0b0b0b8e",
           292 => x"8d040b0b",
           293 => x"0b8e9d04",
           294 => x"0b0b0b8e",
           295 => x"ad040b0b",
           296 => x"0b8ebd04",
           297 => x"0b0b0b8e",
           298 => x"cd040b0b",
           299 => x"0b8edd04",
           300 => x"0b0b0b8e",
           301 => x"ed040b0b",
           302 => x"0b8efd04",
           303 => x"0b0b0b8f",
           304 => x"8d040b0b",
           305 => x"0b8f9d04",
           306 => x"0b0b0b8f",
           307 => x"ad040b0b",
           308 => x"0b8fbd04",
           309 => x"0b0b0b8f",
           310 => x"cd040b0b",
           311 => x"0b8fdd04",
           312 => x"0b0b0b8f",
           313 => x"ed040b0b",
           314 => x"0b8ffd04",
           315 => x"0b0b0b90",
           316 => x"8d040b0b",
           317 => x"0b909d04",
           318 => x"0b0b0b90",
           319 => x"ad040b0b",
           320 => x"0b90bd04",
           321 => x"0b0b0b90",
           322 => x"cd040b0b",
           323 => x"0b90dd04",
           324 => x"0b0b0b90",
           325 => x"ed040b0b",
           326 => x"0b90fd04",
           327 => x"0b0b0b91",
           328 => x"8d040b0b",
           329 => x"0b919d04",
           330 => x"0b0b0b91",
           331 => x"ad040b0b",
           332 => x"0b91bd04",
           333 => x"0b0b0b91",
           334 => x"cd040b0b",
           335 => x"0b91dd04",
           336 => x"0b0b0b91",
           337 => x"ed040b0b",
           338 => x"0b91fd04",
           339 => x"0b0b0b92",
           340 => x"8d040b0b",
           341 => x"0b929d04",
           342 => x"0b0b0b92",
           343 => x"ad040b0b",
           344 => x"0b92bd04",
           345 => x"0b0b0b92",
           346 => x"cd04ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0482b5d4",
           386 => x"0c80f4da",
           387 => x"2d82b5d4",
           388 => x"0882d090",
           389 => x"0482b5d4",
           390 => x"0cb3b22d",
           391 => x"82b5d408",
           392 => x"82d09004",
           393 => x"82b5d40c",
           394 => x"afe32d82",
           395 => x"b5d40882",
           396 => x"d0900482",
           397 => x"b5d40caf",
           398 => x"ad2d82b5",
           399 => x"d40882d0",
           400 => x"900482b5",
           401 => x"d40c94ad",
           402 => x"2d82b5d4",
           403 => x"0882d090",
           404 => x"0482b5d4",
           405 => x"0cb1c22d",
           406 => x"82b5d408",
           407 => x"82d09004",
           408 => x"82b5d40c",
           409 => x"80cfcc2d",
           410 => x"82b5d408",
           411 => x"82d09004",
           412 => x"82b5d40c",
           413 => x"80c9fb2d",
           414 => x"82b5d408",
           415 => x"82d09004",
           416 => x"82b5d40c",
           417 => x"93d82d82",
           418 => x"b5d40882",
           419 => x"d0900482",
           420 => x"b5d40c96",
           421 => x"c02d82b5",
           422 => x"d40882d0",
           423 => x"900482b5",
           424 => x"d40c97cd",
           425 => x"2d82b5d4",
           426 => x"0882d090",
           427 => x"0482b5d4",
           428 => x"0c80f884",
           429 => x"2d82b5d4",
           430 => x"0882d090",
           431 => x"0482b5d4",
           432 => x"0c80f8e2",
           433 => x"2d82b5d4",
           434 => x"0882d090",
           435 => x"0482b5d4",
           436 => x"0c80f09f",
           437 => x"2d82b5d4",
           438 => x"0882d090",
           439 => x"0482b5d4",
           440 => x"0c80f296",
           441 => x"2d82b5d4",
           442 => x"0882d090",
           443 => x"0482b5d4",
           444 => x"0c80f3c9",
           445 => x"2d82b5d4",
           446 => x"0882d090",
           447 => x"0482b5d4",
           448 => x"0c81d7fc",
           449 => x"2d82b5d4",
           450 => x"0882d090",
           451 => x"0482b5d4",
           452 => x"0c81e4ed",
           453 => x"2d82b5d4",
           454 => x"0882d090",
           455 => x"0482b5d4",
           456 => x"0c81dce1",
           457 => x"2d82b5d4",
           458 => x"0882d090",
           459 => x"0482b5d4",
           460 => x"0c81dfde",
           461 => x"2d82b5d4",
           462 => x"0882d090",
           463 => x"0482b5d4",
           464 => x"0c81e9fc",
           465 => x"2d82b5d4",
           466 => x"0882d090",
           467 => x"0482b5d4",
           468 => x"0c81f2dc",
           469 => x"2d82b5d4",
           470 => x"0882d090",
           471 => x"0482b5d4",
           472 => x"0c81e3cf",
           473 => x"2d82b5d4",
           474 => x"0882d090",
           475 => x"0482b5d4",
           476 => x"0c81ed9b",
           477 => x"2d82b5d4",
           478 => x"0882d090",
           479 => x"0482b5d4",
           480 => x"0c81eeba",
           481 => x"2d82b5d4",
           482 => x"0882d090",
           483 => x"0482b5d4",
           484 => x"0c81eed9",
           485 => x"2d82b5d4",
           486 => x"0882d090",
           487 => x"0482b5d4",
           488 => x"0c81f6c3",
           489 => x"2d82b5d4",
           490 => x"0882d090",
           491 => x"0482b5d4",
           492 => x"0c81f4a9",
           493 => x"2d82b5d4",
           494 => x"0882d090",
           495 => x"0482b5d4",
           496 => x"0c81f997",
           497 => x"2d82b5d4",
           498 => x"0882d090",
           499 => x"0482b5d4",
           500 => x"0c81efdd",
           501 => x"2d82b5d4",
           502 => x"0882d090",
           503 => x"0482b5d4",
           504 => x"0c81fc97",
           505 => x"2d82b5d4",
           506 => x"0882d090",
           507 => x"0482b5d4",
           508 => x"0c81fd98",
           509 => x"2d82b5d4",
           510 => x"0882d090",
           511 => x"0482b5d4",
           512 => x"0c81e5cd",
           513 => x"2d82b5d4",
           514 => x"0882d090",
           515 => x"0482b5d4",
           516 => x"0c81e5a6",
           517 => x"2d82b5d4",
           518 => x"0882d090",
           519 => x"0482b5d4",
           520 => x"0c81e6d1",
           521 => x"2d82b5d4",
           522 => x"0882d090",
           523 => x"0482b5d4",
           524 => x"0c81f0b4",
           525 => x"2d82b5d4",
           526 => x"0882d090",
           527 => x"0482b5d4",
           528 => x"0c81fe89",
           529 => x"2d82b5d4",
           530 => x"0882d090",
           531 => x"0482b5d4",
           532 => x"0c828093",
           533 => x"2d82b5d4",
           534 => x"0882d090",
           535 => x"0482b5d4",
           536 => x"0c8283d5",
           537 => x"2d82b5d4",
           538 => x"0882d090",
           539 => x"0482b5d4",
           540 => x"0c81d79b",
           541 => x"2d82b5d4",
           542 => x"0882d090",
           543 => x"0482b5d4",
           544 => x"0c8286c1",
           545 => x"2d82b5d4",
           546 => x"0882d090",
           547 => x"0482b5d4",
           548 => x"0c8294f6",
           549 => x"2d82b5d4",
           550 => x"0882d090",
           551 => x"0482b5d4",
           552 => x"0c8292e2",
           553 => x"2d82b5d4",
           554 => x"0882d090",
           555 => x"0482b5d4",
           556 => x"0c81a8d6",
           557 => x"2d82b5d4",
           558 => x"0882d090",
           559 => x"0482b5d4",
           560 => x"0c81aac0",
           561 => x"2d82b5d4",
           562 => x"0882d090",
           563 => x"0482b5d4",
           564 => x"0c81aca4",
           565 => x"2d82b5d4",
           566 => x"0882d090",
           567 => x"0482b5d4",
           568 => x"0c80f0c8",
           569 => x"2d82b5d4",
           570 => x"0882d090",
           571 => x"0482b5d4",
           572 => x"0c80f1ec",
           573 => x"2d82b5d4",
           574 => x"0882d090",
           575 => x"0482b5d4",
           576 => x"0c80f5cf",
           577 => x"2d82b5d4",
           578 => x"0882d090",
           579 => x"0482b5d4",
           580 => x"0c80d698",
           581 => x"2d82b5d4",
           582 => x"0882d090",
           583 => x"0482b5d4",
           584 => x"0c81a2ea",
           585 => x"2d82b5d4",
           586 => x"0882d090",
           587 => x"0482b5d4",
           588 => x"0c81a392",
           589 => x"2d82b5d4",
           590 => x"0882d090",
           591 => x"0482b5d4",
           592 => x"0c81a78a",
           593 => x"2d82b5d4",
           594 => x"0882d090",
           595 => x"0482b5d4",
           596 => x"0c819fd4",
           597 => x"2d82b5d4",
           598 => x"0882d090",
           599 => x"043c0400",
           600 => x"00101010",
           601 => x"10101010",
           602 => x"10101010",
           603 => x"10101010",
           604 => x"10101010",
           605 => x"10101010",
           606 => x"10101010",
           607 => x"10101010",
           608 => x"53510400",
           609 => x"007381ff",
           610 => x"06738306",
           611 => x"09810583",
           612 => x"05101010",
           613 => x"2b0772fc",
           614 => x"060c5151",
           615 => x"04727280",
           616 => x"728106ff",
           617 => x"05097206",
           618 => x"05711052",
           619 => x"720a100a",
           620 => x"5372ed38",
           621 => x"51515351",
           622 => x"0482b5c8",
           623 => x"7082cda4",
           624 => x"278e3880",
           625 => x"71708405",
           626 => x"530c0b0b",
           627 => x"0b93bc04",
           628 => x"8c815180",
           629 => x"eee20400",
           630 => x"82b5d408",
           631 => x"0282b5d4",
           632 => x"0cfb3d0d",
           633 => x"82b5d408",
           634 => x"8c057082",
           635 => x"b5d408fc",
           636 => x"050c82b5",
           637 => x"d408fc05",
           638 => x"085482b5",
           639 => x"d4088805",
           640 => x"085382cd",
           641 => x"9c085254",
           642 => x"849a3f82",
           643 => x"b5c80870",
           644 => x"82b5d408",
           645 => x"f8050c82",
           646 => x"b5d408f8",
           647 => x"05087082",
           648 => x"b5c80c51",
           649 => x"54873d0d",
           650 => x"82b5d40c",
           651 => x"0482b5d4",
           652 => x"080282b5",
           653 => x"d40cfb3d",
           654 => x"0d82b5d4",
           655 => x"08900508",
           656 => x"85113370",
           657 => x"81327081",
           658 => x"06515151",
           659 => x"52718f38",
           660 => x"800b82b5",
           661 => x"d4088c05",
           662 => x"08258338",
           663 => x"8d39800b",
           664 => x"82b5d408",
           665 => x"f4050c81",
           666 => x"c43982b5",
           667 => x"d4088c05",
           668 => x"08ff0582",
           669 => x"b5d4088c",
           670 => x"050c800b",
           671 => x"82b5d408",
           672 => x"f8050c82",
           673 => x"b5d40888",
           674 => x"050882b5",
           675 => x"d408fc05",
           676 => x"0c82b5d4",
           677 => x"08f80508",
           678 => x"8a2e80f6",
           679 => x"38800b82",
           680 => x"b5d4088c",
           681 => x"05082580",
           682 => x"e93882b5",
           683 => x"d4089005",
           684 => x"0851a090",
           685 => x"3f82b5c8",
           686 => x"087082b5",
           687 => x"d408f805",
           688 => x"0c5282b5",
           689 => x"d408f805",
           690 => x"08ff2e09",
           691 => x"81068d38",
           692 => x"800b82b5",
           693 => x"d408f405",
           694 => x"0c80d239",
           695 => x"82b5d408",
           696 => x"fc050882",
           697 => x"b5d408f8",
           698 => x"05085353",
           699 => x"71733482",
           700 => x"b5d4088c",
           701 => x"0508ff05",
           702 => x"82b5d408",
           703 => x"8c050c82",
           704 => x"b5d408fc",
           705 => x"05088105",
           706 => x"82b5d408",
           707 => x"fc050cff",
           708 => x"803982b5",
           709 => x"d408fc05",
           710 => x"08528072",
           711 => x"3482b5d4",
           712 => x"08880508",
           713 => x"7082b5d4",
           714 => x"08f4050c",
           715 => x"5282b5d4",
           716 => x"08f40508",
           717 => x"82b5c80c",
           718 => x"873d0d82",
           719 => x"b5d40c04",
           720 => x"82b5d408",
           721 => x"0282b5d4",
           722 => x"0cf43d0d",
           723 => x"860b82b5",
           724 => x"d408e505",
           725 => x"3482b5d4",
           726 => x"08880508",
           727 => x"82b5d408",
           728 => x"e0050cfe",
           729 => x"0a0b82b5",
           730 => x"d408e805",
           731 => x"0c82b5d4",
           732 => x"08900570",
           733 => x"82b5d408",
           734 => x"fc050c82",
           735 => x"b5d408fc",
           736 => x"05085482",
           737 => x"b5d4088c",
           738 => x"05085382",
           739 => x"b5d408e0",
           740 => x"05705351",
           741 => x"54818d3f",
           742 => x"82b5c808",
           743 => x"7082b5d4",
           744 => x"08dc050c",
           745 => x"82b5d408",
           746 => x"ec050882",
           747 => x"b5d40888",
           748 => x"05080551",
           749 => x"54807434",
           750 => x"82b5d408",
           751 => x"dc050870",
           752 => x"82b5c80c",
           753 => x"548e3d0d",
           754 => x"82b5d40c",
           755 => x"0482b5d4",
           756 => x"080282b5",
           757 => x"d40cfb3d",
           758 => x"0d82b5d4",
           759 => x"08900570",
           760 => x"82b5d408",
           761 => x"fc050c82",
           762 => x"b5d408fc",
           763 => x"05085482",
           764 => x"b5d4088c",
           765 => x"05085382",
           766 => x"b5d40888",
           767 => x"05085254",
           768 => x"a33f82b5",
           769 => x"c8087082",
           770 => x"b5d408f8",
           771 => x"050c82b5",
           772 => x"d408f805",
           773 => x"087082b5",
           774 => x"c80c5154",
           775 => x"873d0d82",
           776 => x"b5d40c04",
           777 => x"82b5d408",
           778 => x"0282b5d4",
           779 => x"0ced3d0d",
           780 => x"800b82b5",
           781 => x"d408e405",
           782 => x"2382b5d4",
           783 => x"08880508",
           784 => x"53800b8c",
           785 => x"140c82b5",
           786 => x"d4088805",
           787 => x"08851133",
           788 => x"70812a70",
           789 => x"81327081",
           790 => x"06515151",
           791 => x"51537280",
           792 => x"2e8d38ff",
           793 => x"0b82b5d4",
           794 => x"08e0050c",
           795 => x"96ac3982",
           796 => x"b5d4088c",
           797 => x"05085372",
           798 => x"33537282",
           799 => x"b5d408f8",
           800 => x"05347281",
           801 => x"ff065372",
           802 => x"802e95fa",
           803 => x"3882b5d4",
           804 => x"088c0508",
           805 => x"810582b5",
           806 => x"d4088c05",
           807 => x"0c82b5d4",
           808 => x"08e40522",
           809 => x"70810651",
           810 => x"5372802e",
           811 => x"958b3882",
           812 => x"b5d408f8",
           813 => x"053353af",
           814 => x"732781fc",
           815 => x"3882b5d4",
           816 => x"08f80533",
           817 => x"5372b926",
           818 => x"81ee3882",
           819 => x"b5d408f8",
           820 => x"05335372",
           821 => x"b02e0981",
           822 => x"0680c538",
           823 => x"82b5d408",
           824 => x"e8053370",
           825 => x"982b7098",
           826 => x"2c515153",
           827 => x"72b23882",
           828 => x"b5d408e4",
           829 => x"05227083",
           830 => x"2a708132",
           831 => x"70810651",
           832 => x"51515372",
           833 => x"802e9938",
           834 => x"82b5d408",
           835 => x"e4052270",
           836 => x"82800751",
           837 => x"537282b5",
           838 => x"d408e405",
           839 => x"23fed039",
           840 => x"82b5d408",
           841 => x"e8053370",
           842 => x"982b7098",
           843 => x"2c707083",
           844 => x"2b721173",
           845 => x"11515151",
           846 => x"53515553",
           847 => x"7282b5d4",
           848 => x"08e80534",
           849 => x"82b5d408",
           850 => x"e8053354",
           851 => x"82b5d408",
           852 => x"f8053370",
           853 => x"15d01151",
           854 => x"51537282",
           855 => x"b5d408e8",
           856 => x"053482b5",
           857 => x"d408e805",
           858 => x"3370982b",
           859 => x"70982c51",
           860 => x"51537280",
           861 => x"258b3880",
           862 => x"ff0b82b5",
           863 => x"d408e805",
           864 => x"3482b5d4",
           865 => x"08e40522",
           866 => x"70832a70",
           867 => x"81065151",
           868 => x"5372fddb",
           869 => x"3882b5d4",
           870 => x"08e80533",
           871 => x"70882b70",
           872 => x"902b7090",
           873 => x"2c70882c",
           874 => x"51515151",
           875 => x"537282b5",
           876 => x"d408ec05",
           877 => x"23fdb839",
           878 => x"82b5d408",
           879 => x"e4052270",
           880 => x"832a7081",
           881 => x"06515153",
           882 => x"72802e9d",
           883 => x"3882b5d4",
           884 => x"08e80533",
           885 => x"70982b70",
           886 => x"982c5151",
           887 => x"53728a38",
           888 => x"810b82b5",
           889 => x"d408e805",
           890 => x"3482b5d4",
           891 => x"08f80533",
           892 => x"e01182b5",
           893 => x"d408c405",
           894 => x"0c5382b5",
           895 => x"d408c405",
           896 => x"0880d826",
           897 => x"92943882",
           898 => x"b5d408c4",
           899 => x"05087082",
           900 => x"2b8296e4",
           901 => x"11700851",
           902 => x"51515372",
           903 => x"0482b5d4",
           904 => x"08e40522",
           905 => x"70900751",
           906 => x"537282b5",
           907 => x"d408e405",
           908 => x"2382b5d4",
           909 => x"08e40522",
           910 => x"70a00751",
           911 => x"537282b5",
           912 => x"d408e405",
           913 => x"23fca839",
           914 => x"82b5d408",
           915 => x"e4052270",
           916 => x"81800751",
           917 => x"537282b5",
           918 => x"d408e405",
           919 => x"23fc9039",
           920 => x"82b5d408",
           921 => x"e4052270",
           922 => x"80c00751",
           923 => x"537282b5",
           924 => x"d408e405",
           925 => x"23fbf839",
           926 => x"82b5d408",
           927 => x"e4052270",
           928 => x"88075153",
           929 => x"7282b5d4",
           930 => x"08e40523",
           931 => x"800b82b5",
           932 => x"d408e805",
           933 => x"34fbd839",
           934 => x"82b5d408",
           935 => x"e4052270",
           936 => x"84075153",
           937 => x"7282b5d4",
           938 => x"08e40523",
           939 => x"fbc139bf",
           940 => x"0b82b5d4",
           941 => x"08fc0534",
           942 => x"82b5d408",
           943 => x"ec0522ff",
           944 => x"11515372",
           945 => x"82b5d408",
           946 => x"ec052380",
           947 => x"e30b82b5",
           948 => x"d408f805",
           949 => x"348da839",
           950 => x"82b5d408",
           951 => x"90050882",
           952 => x"b5d40890",
           953 => x"05088405",
           954 => x"82b5d408",
           955 => x"90050c70",
           956 => x"08515372",
           957 => x"82b5d408",
           958 => x"fc053482",
           959 => x"b5d408ec",
           960 => x"0522ff11",
           961 => x"51537282",
           962 => x"b5d408ec",
           963 => x"05238cef",
           964 => x"3982b5d4",
           965 => x"08900508",
           966 => x"82b5d408",
           967 => x"90050884",
           968 => x"0582b5d4",
           969 => x"0890050c",
           970 => x"700882b5",
           971 => x"d408fc05",
           972 => x"0c82b5d4",
           973 => x"08e40522",
           974 => x"70832a70",
           975 => x"81065151",
           976 => x"51537280",
           977 => x"2eab3882",
           978 => x"b5d408e8",
           979 => x"05337098",
           980 => x"2b537298",
           981 => x"2c5382b5",
           982 => x"d408fc05",
           983 => x"085253a2",
           984 => x"d83f82b5",
           985 => x"c8085372",
           986 => x"82b5d408",
           987 => x"f4052399",
           988 => x"3982b5d4",
           989 => x"08fc0508",
           990 => x"519d8a3f",
           991 => x"82b5c808",
           992 => x"537282b5",
           993 => x"d408f405",
           994 => x"2382b5d4",
           995 => x"08ec0522",
           996 => x"5382b5d4",
           997 => x"08f40522",
           998 => x"73713154",
           999 => x"547282b5",
          1000 => x"d408ec05",
          1001 => x"238bd839",
          1002 => x"82b5d408",
          1003 => x"90050882",
          1004 => x"b5d40890",
          1005 => x"05088405",
          1006 => x"82b5d408",
          1007 => x"90050c70",
          1008 => x"0882b5d4",
          1009 => x"08fc050c",
          1010 => x"82b5d408",
          1011 => x"e4052270",
          1012 => x"832a7081",
          1013 => x"06515151",
          1014 => x"5372802e",
          1015 => x"ab3882b5",
          1016 => x"d408e805",
          1017 => x"3370982b",
          1018 => x"5372982c",
          1019 => x"5382b5d4",
          1020 => x"08fc0508",
          1021 => x"5253a1c1",
          1022 => x"3f82b5c8",
          1023 => x"08537282",
          1024 => x"b5d408f4",
          1025 => x"05239939",
          1026 => x"82b5d408",
          1027 => x"fc050851",
          1028 => x"9bf33f82",
          1029 => x"b5c80853",
          1030 => x"7282b5d4",
          1031 => x"08f40523",
          1032 => x"82b5d408",
          1033 => x"ec052253",
          1034 => x"82b5d408",
          1035 => x"f4052273",
          1036 => x"71315454",
          1037 => x"7282b5d4",
          1038 => x"08ec0523",
          1039 => x"8ac13982",
          1040 => x"b5d408e4",
          1041 => x"05227082",
          1042 => x"2a708106",
          1043 => x"51515372",
          1044 => x"802ea438",
          1045 => x"82b5d408",
          1046 => x"90050882",
          1047 => x"b5d40890",
          1048 => x"05088405",
          1049 => x"82b5d408",
          1050 => x"90050c70",
          1051 => x"0882b5d4",
          1052 => x"08dc050c",
          1053 => x"53a23982",
          1054 => x"b5d40890",
          1055 => x"050882b5",
          1056 => x"d4089005",
          1057 => x"08840582",
          1058 => x"b5d40890",
          1059 => x"050c7008",
          1060 => x"82b5d408",
          1061 => x"dc050c53",
          1062 => x"82b5d408",
          1063 => x"dc050882",
          1064 => x"b5d408fc",
          1065 => x"050c82b5",
          1066 => x"d408fc05",
          1067 => x"088025a4",
          1068 => x"3882b5d4",
          1069 => x"08e40522",
          1070 => x"70820751",
          1071 => x"537282b5",
          1072 => x"d408e405",
          1073 => x"2382b5d4",
          1074 => x"08fc0508",
          1075 => x"3082b5d4",
          1076 => x"08fc050c",
          1077 => x"82b5d408",
          1078 => x"e4052270",
          1079 => x"ffbf0651",
          1080 => x"537282b5",
          1081 => x"d408e405",
          1082 => x"2381af39",
          1083 => x"880b82b5",
          1084 => x"d408f405",
          1085 => x"23a93982",
          1086 => x"b5d408e4",
          1087 => x"05227080",
          1088 => x"c0075153",
          1089 => x"7282b5d4",
          1090 => x"08e40523",
          1091 => x"80f80b82",
          1092 => x"b5d408f8",
          1093 => x"0534900b",
          1094 => x"82b5d408",
          1095 => x"f4052382",
          1096 => x"b5d408e4",
          1097 => x"05227082",
          1098 => x"2a708106",
          1099 => x"51515372",
          1100 => x"802ea438",
          1101 => x"82b5d408",
          1102 => x"90050882",
          1103 => x"b5d40890",
          1104 => x"05088405",
          1105 => x"82b5d408",
          1106 => x"90050c70",
          1107 => x"0882b5d4",
          1108 => x"08d8050c",
          1109 => x"53a23982",
          1110 => x"b5d40890",
          1111 => x"050882b5",
          1112 => x"d4089005",
          1113 => x"08840582",
          1114 => x"b5d40890",
          1115 => x"050c7008",
          1116 => x"82b5d408",
          1117 => x"d8050c53",
          1118 => x"82b5d408",
          1119 => x"d8050882",
          1120 => x"b5d408fc",
          1121 => x"050c82b5",
          1122 => x"d408e405",
          1123 => x"2270cf06",
          1124 => x"51537282",
          1125 => x"b5d408e4",
          1126 => x"052382b5",
          1127 => x"d80b82b5",
          1128 => x"d408f005",
          1129 => x"0c82b5d4",
          1130 => x"08f00508",
          1131 => x"82b5d408",
          1132 => x"f4052282",
          1133 => x"b5d408fc",
          1134 => x"05087155",
          1135 => x"70545654",
          1136 => x"55a3f33f",
          1137 => x"82b5c808",
          1138 => x"53727534",
          1139 => x"82b5d408",
          1140 => x"f0050882",
          1141 => x"b5d408d4",
          1142 => x"050c82b5",
          1143 => x"d408f005",
          1144 => x"08703351",
          1145 => x"53897327",
          1146 => x"a43882b5",
          1147 => x"d408f005",
          1148 => x"08537233",
          1149 => x"5482b5d4",
          1150 => x"08f80533",
          1151 => x"7015df11",
          1152 => x"51515372",
          1153 => x"82b5d408",
          1154 => x"d0053497",
          1155 => x"3982b5d4",
          1156 => x"08f00508",
          1157 => x"537233b0",
          1158 => x"11515372",
          1159 => x"82b5d408",
          1160 => x"d0053482",
          1161 => x"b5d408d4",
          1162 => x"05085382",
          1163 => x"b5d408d0",
          1164 => x"05337334",
          1165 => x"82b5d408",
          1166 => x"f0050881",
          1167 => x"0582b5d4",
          1168 => x"08f0050c",
          1169 => x"82b5d408",
          1170 => x"f4052270",
          1171 => x"5382b5d4",
          1172 => x"08fc0508",
          1173 => x"5253a2ab",
          1174 => x"3f82b5c8",
          1175 => x"087082b5",
          1176 => x"d408fc05",
          1177 => x"0c5382b5",
          1178 => x"d408fc05",
          1179 => x"08802e84",
          1180 => x"38feb239",
          1181 => x"82b5d408",
          1182 => x"f0050882",
          1183 => x"b5d85455",
          1184 => x"72547470",
          1185 => x"75315153",
          1186 => x"7282b5d4",
          1187 => x"08fc0534",
          1188 => x"82b5d408",
          1189 => x"e4052270",
          1190 => x"b2065153",
          1191 => x"72802e94",
          1192 => x"3882b5d4",
          1193 => x"08ec0522",
          1194 => x"ff115153",
          1195 => x"7282b5d4",
          1196 => x"08ec0523",
          1197 => x"82b5d408",
          1198 => x"e4052270",
          1199 => x"862a7081",
          1200 => x"06515153",
          1201 => x"72802e80",
          1202 => x"e73882b5",
          1203 => x"d408ec05",
          1204 => x"2270902b",
          1205 => x"82b5d408",
          1206 => x"cc050c82",
          1207 => x"b5d408cc",
          1208 => x"0508902c",
          1209 => x"82b5d408",
          1210 => x"cc050c82",
          1211 => x"b5d408f4",
          1212 => x"05225153",
          1213 => x"72902e09",
          1214 => x"81069538",
          1215 => x"82b5d408",
          1216 => x"cc0508fe",
          1217 => x"05537282",
          1218 => x"b5d408c8",
          1219 => x"05239339",
          1220 => x"82b5d408",
          1221 => x"cc0508ff",
          1222 => x"05537282",
          1223 => x"b5d408c8",
          1224 => x"052382b5",
          1225 => x"d408c805",
          1226 => x"2282b5d4",
          1227 => x"08ec0523",
          1228 => x"82b5d408",
          1229 => x"e4052270",
          1230 => x"832a7081",
          1231 => x"06515153",
          1232 => x"72802e80",
          1233 => x"d03882b5",
          1234 => x"d408e805",
          1235 => x"3370982b",
          1236 => x"70982c82",
          1237 => x"b5d408fc",
          1238 => x"05335751",
          1239 => x"51537274",
          1240 => x"24973882",
          1241 => x"b5d408e4",
          1242 => x"052270f7",
          1243 => x"06515372",
          1244 => x"82b5d408",
          1245 => x"e405239d",
          1246 => x"3982b5d4",
          1247 => x"08e80533",
          1248 => x"5382b5d4",
          1249 => x"08fc0533",
          1250 => x"73713154",
          1251 => x"547282b5",
          1252 => x"d408e805",
          1253 => x"3482b5d4",
          1254 => x"08e40522",
          1255 => x"70832a70",
          1256 => x"81065151",
          1257 => x"5372802e",
          1258 => x"b13882b5",
          1259 => x"d408e805",
          1260 => x"3370882b",
          1261 => x"70902b70",
          1262 => x"902c7088",
          1263 => x"2c515151",
          1264 => x"51537254",
          1265 => x"82b5d408",
          1266 => x"ec052270",
          1267 => x"75315153",
          1268 => x"7282b5d4",
          1269 => x"08ec0523",
          1270 => x"af3982b5",
          1271 => x"d408fc05",
          1272 => x"3370882b",
          1273 => x"70902b70",
          1274 => x"902c7088",
          1275 => x"2c515151",
          1276 => x"51537254",
          1277 => x"82b5d408",
          1278 => x"ec052270",
          1279 => x"75315153",
          1280 => x"7282b5d4",
          1281 => x"08ec0523",
          1282 => x"82b5d408",
          1283 => x"e4052270",
          1284 => x"83800651",
          1285 => x"5372b038",
          1286 => x"82b5d408",
          1287 => x"ec0522ff",
          1288 => x"11545472",
          1289 => x"82b5d408",
          1290 => x"ec052373",
          1291 => x"902b7090",
          1292 => x"2c515380",
          1293 => x"73259038",
          1294 => x"82b5d408",
          1295 => x"88050852",
          1296 => x"a0518aee",
          1297 => x"3fd23982",
          1298 => x"b5d408e4",
          1299 => x"05227081",
          1300 => x"2a708106",
          1301 => x"51515372",
          1302 => x"802e9138",
          1303 => x"82b5d408",
          1304 => x"88050852",
          1305 => x"ad518aca",
          1306 => x"3f80c739",
          1307 => x"82b5d408",
          1308 => x"e4052270",
          1309 => x"842a7081",
          1310 => x"06515153",
          1311 => x"72802e90",
          1312 => x"3882b5d4",
          1313 => x"08880508",
          1314 => x"52ab518a",
          1315 => x"a53fa339",
          1316 => x"82b5d408",
          1317 => x"e4052270",
          1318 => x"852a7081",
          1319 => x"06515153",
          1320 => x"72802e8e",
          1321 => x"3882b5d4",
          1322 => x"08880508",
          1323 => x"52a0518a",
          1324 => x"813f82b5",
          1325 => x"d408e405",
          1326 => x"2270862a",
          1327 => x"70810651",
          1328 => x"51537280",
          1329 => x"2eb13882",
          1330 => x"b5d40888",
          1331 => x"050852b0",
          1332 => x"5189df3f",
          1333 => x"82b5d408",
          1334 => x"f4052253",
          1335 => x"72902e09",
          1336 => x"81069438",
          1337 => x"82b5d408",
          1338 => x"88050852",
          1339 => x"82b5d408",
          1340 => x"f8053351",
          1341 => x"89bc3f82",
          1342 => x"b5d408e4",
          1343 => x"05227088",
          1344 => x"2a708106",
          1345 => x"51515372",
          1346 => x"802eb038",
          1347 => x"82b5d408",
          1348 => x"ec0522ff",
          1349 => x"11545472",
          1350 => x"82b5d408",
          1351 => x"ec052373",
          1352 => x"902b7090",
          1353 => x"2c515380",
          1354 => x"73259038",
          1355 => x"82b5d408",
          1356 => x"88050852",
          1357 => x"b05188fa",
          1358 => x"3fd23982",
          1359 => x"b5d408e4",
          1360 => x"05227083",
          1361 => x"2a708106",
          1362 => x"51515372",
          1363 => x"802eb038",
          1364 => x"82b5d408",
          1365 => x"e80533ff",
          1366 => x"11545472",
          1367 => x"82b5d408",
          1368 => x"e8053473",
          1369 => x"982b7098",
          1370 => x"2c515380",
          1371 => x"73259038",
          1372 => x"82b5d408",
          1373 => x"88050852",
          1374 => x"b05188b6",
          1375 => x"3fd23982",
          1376 => x"b5d408e4",
          1377 => x"05227087",
          1378 => x"2a708106",
          1379 => x"51515372",
          1380 => x"b03882b5",
          1381 => x"d408ec05",
          1382 => x"22ff1154",
          1383 => x"547282b5",
          1384 => x"d408ec05",
          1385 => x"2373902b",
          1386 => x"70902c51",
          1387 => x"53807325",
          1388 => x"903882b5",
          1389 => x"d4088805",
          1390 => x"0852a051",
          1391 => x"87f43fd2",
          1392 => x"3982b5d4",
          1393 => x"08f80533",
          1394 => x"537280e3",
          1395 => x"2e098106",
          1396 => x"973882b5",
          1397 => x"d4088805",
          1398 => x"085282b5",
          1399 => x"d408fc05",
          1400 => x"335187ce",
          1401 => x"3f81ee39",
          1402 => x"82b5d408",
          1403 => x"f8053353",
          1404 => x"7280f32e",
          1405 => x"09810680",
          1406 => x"cb3882b5",
          1407 => x"d408f405",
          1408 => x"22ff1151",
          1409 => x"537282b5",
          1410 => x"d408f405",
          1411 => x"237283ff",
          1412 => x"ff065372",
          1413 => x"83ffff2e",
          1414 => x"81bb3882",
          1415 => x"b5d40888",
          1416 => x"05085282",
          1417 => x"b5d408fc",
          1418 => x"05087033",
          1419 => x"5282b5d4",
          1420 => x"08fc0508",
          1421 => x"810582b5",
          1422 => x"d408fc05",
          1423 => x"0c5386f2",
          1424 => x"3fffb739",
          1425 => x"82b5d408",
          1426 => x"f8053353",
          1427 => x"7280d32e",
          1428 => x"09810680",
          1429 => x"cb3882b5",
          1430 => x"d408f405",
          1431 => x"22ff1151",
          1432 => x"537282b5",
          1433 => x"d408f405",
          1434 => x"237283ff",
          1435 => x"ff065372",
          1436 => x"83ffff2e",
          1437 => x"80df3882",
          1438 => x"b5d40888",
          1439 => x"05085282",
          1440 => x"b5d408fc",
          1441 => x"05087033",
          1442 => x"525386a6",
          1443 => x"3f82b5d4",
          1444 => x"08fc0508",
          1445 => x"810582b5",
          1446 => x"d408fc05",
          1447 => x"0cffb739",
          1448 => x"82b5d408",
          1449 => x"f0050882",
          1450 => x"b5d82ea9",
          1451 => x"3882b5d4",
          1452 => x"08880508",
          1453 => x"5282b5d4",
          1454 => x"08f00508",
          1455 => x"ff0582b5",
          1456 => x"d408f005",
          1457 => x"0c82b5d4",
          1458 => x"08f00508",
          1459 => x"70335253",
          1460 => x"85e03fcc",
          1461 => x"3982b5d4",
          1462 => x"08e40522",
          1463 => x"70872a70",
          1464 => x"81065151",
          1465 => x"5372802e",
          1466 => x"80c33882",
          1467 => x"b5d408ec",
          1468 => x"0522ff11",
          1469 => x"54547282",
          1470 => x"b5d408ec",
          1471 => x"05237390",
          1472 => x"2b70902c",
          1473 => x"51538073",
          1474 => x"25a33882",
          1475 => x"b5d40888",
          1476 => x"050852a0",
          1477 => x"51859b3f",
          1478 => x"d23982b5",
          1479 => x"d4088805",
          1480 => x"085282b5",
          1481 => x"d408f805",
          1482 => x"33518586",
          1483 => x"3f800b82",
          1484 => x"b5d408e4",
          1485 => x"0523eab7",
          1486 => x"3982b5d4",
          1487 => x"08f80533",
          1488 => x"5372a52e",
          1489 => x"098106a8",
          1490 => x"38810b82",
          1491 => x"b5d408e4",
          1492 => x"0523800b",
          1493 => x"82b5d408",
          1494 => x"ec052380",
          1495 => x"0b82b5d4",
          1496 => x"08e80534",
          1497 => x"8a0b82b5",
          1498 => x"d408f405",
          1499 => x"23ea8039",
          1500 => x"82b5d408",
          1501 => x"88050852",
          1502 => x"82b5d408",
          1503 => x"f8053351",
          1504 => x"84b03fe9",
          1505 => x"ea3982b5",
          1506 => x"d4088805",
          1507 => x"088c1108",
          1508 => x"7082b5d4",
          1509 => x"08e0050c",
          1510 => x"515382b5",
          1511 => x"d408e005",
          1512 => x"0882b5c8",
          1513 => x"0c953d0d",
          1514 => x"82b5d40c",
          1515 => x"0482b5d4",
          1516 => x"080282b5",
          1517 => x"d40cfd3d",
          1518 => x"0d82cd98",
          1519 => x"085382b5",
          1520 => x"d4088c05",
          1521 => x"085282b5",
          1522 => x"d4088805",
          1523 => x"0851e4dd",
          1524 => x"3f82b5c8",
          1525 => x"087082b5",
          1526 => x"c80c5485",
          1527 => x"3d0d82b5",
          1528 => x"d40c0482",
          1529 => x"b5d40802",
          1530 => x"82b5d40c",
          1531 => x"fb3d0d80",
          1532 => x"0b82b5d4",
          1533 => x"08f8050c",
          1534 => x"82cd9c08",
          1535 => x"85113370",
          1536 => x"812a7081",
          1537 => x"32708106",
          1538 => x"51515151",
          1539 => x"5372802e",
          1540 => x"8d38ff0b",
          1541 => x"82b5d408",
          1542 => x"f4050c81",
          1543 => x"923982b5",
          1544 => x"d4088805",
          1545 => x"08537233",
          1546 => x"82b5d408",
          1547 => x"88050881",
          1548 => x"0582b5d4",
          1549 => x"0888050c",
          1550 => x"537282b5",
          1551 => x"d408fc05",
          1552 => x"347281ff",
          1553 => x"06537280",
          1554 => x"2eb03882",
          1555 => x"cd9c0882",
          1556 => x"cd9c0853",
          1557 => x"82b5d408",
          1558 => x"fc053352",
          1559 => x"90110851",
          1560 => x"53722d82",
          1561 => x"b5c80853",
          1562 => x"72802eff",
          1563 => x"b138ff0b",
          1564 => x"82b5d408",
          1565 => x"f8050cff",
          1566 => x"a53982cd",
          1567 => x"9c0882cd",
          1568 => x"9c085353",
          1569 => x"8a519013",
          1570 => x"0853722d",
          1571 => x"82b5c808",
          1572 => x"5372802e",
          1573 => x"8a38ff0b",
          1574 => x"82b5d408",
          1575 => x"f8050c82",
          1576 => x"b5d408f8",
          1577 => x"05087082",
          1578 => x"b5d408f4",
          1579 => x"050c5382",
          1580 => x"b5d408f4",
          1581 => x"050882b5",
          1582 => x"c80c873d",
          1583 => x"0d82b5d4",
          1584 => x"0c0482b5",
          1585 => x"d4080282",
          1586 => x"b5d40cfb",
          1587 => x"3d0d800b",
          1588 => x"82b5d408",
          1589 => x"f8050c82",
          1590 => x"b5d4088c",
          1591 => x"05088511",
          1592 => x"3370812a",
          1593 => x"70813270",
          1594 => x"81065151",
          1595 => x"51515372",
          1596 => x"802e8d38",
          1597 => x"ff0b82b5",
          1598 => x"d408f405",
          1599 => x"0c80f339",
          1600 => x"82b5d408",
          1601 => x"88050853",
          1602 => x"723382b5",
          1603 => x"d4088805",
          1604 => x"08810582",
          1605 => x"b5d40888",
          1606 => x"050c5372",
          1607 => x"82b5d408",
          1608 => x"fc053472",
          1609 => x"81ff0653",
          1610 => x"72802eb6",
          1611 => x"3882b5d4",
          1612 => x"088c0508",
          1613 => x"82b5d408",
          1614 => x"8c050853",
          1615 => x"82b5d408",
          1616 => x"fc053352",
          1617 => x"90110851",
          1618 => x"53722d82",
          1619 => x"b5c80853",
          1620 => x"72802eff",
          1621 => x"ab38ff0b",
          1622 => x"82b5d408",
          1623 => x"f8050cff",
          1624 => x"9f3982b5",
          1625 => x"d408f805",
          1626 => x"087082b5",
          1627 => x"d408f405",
          1628 => x"0c5382b5",
          1629 => x"d408f405",
          1630 => x"0882b5c8",
          1631 => x"0c873d0d",
          1632 => x"82b5d40c",
          1633 => x"0482b5d4",
          1634 => x"080282b5",
          1635 => x"d40cfe3d",
          1636 => x"0d82cd9c",
          1637 => x"085282b5",
          1638 => x"d4088805",
          1639 => x"0851933f",
          1640 => x"82b5c808",
          1641 => x"7082b5c8",
          1642 => x"0c53843d",
          1643 => x"0d82b5d4",
          1644 => x"0c0482b5",
          1645 => x"d4080282",
          1646 => x"b5d40cfb",
          1647 => x"3d0d82b5",
          1648 => x"d4088c05",
          1649 => x"08851133",
          1650 => x"70812a70",
          1651 => x"81327081",
          1652 => x"06515151",
          1653 => x"51537280",
          1654 => x"2e8d38ff",
          1655 => x"0b82b5d4",
          1656 => x"08fc050c",
          1657 => x"81cb3982",
          1658 => x"b5d4088c",
          1659 => x"05088511",
          1660 => x"3370822a",
          1661 => x"70810651",
          1662 => x"51515372",
          1663 => x"802e80db",
          1664 => x"3882b5d4",
          1665 => x"088c0508",
          1666 => x"82b5d408",
          1667 => x"8c050854",
          1668 => x"548c1408",
          1669 => x"88140825",
          1670 => x"9f3882b5",
          1671 => x"d4088c05",
          1672 => x"08700870",
          1673 => x"82b5d408",
          1674 => x"88050852",
          1675 => x"57545472",
          1676 => x"75347308",
          1677 => x"8105740c",
          1678 => x"82b5d408",
          1679 => x"8c05088c",
          1680 => x"11088105",
          1681 => x"8c120c82",
          1682 => x"b5d40888",
          1683 => x"05087082",
          1684 => x"b5d408fc",
          1685 => x"050c5153",
          1686 => x"80d73982",
          1687 => x"b5d4088c",
          1688 => x"050882b5",
          1689 => x"d4088c05",
          1690 => x"085382b5",
          1691 => x"d4088805",
          1692 => x"087081ff",
          1693 => x"06539012",
          1694 => x"08515454",
          1695 => x"722d82b5",
          1696 => x"c8085372",
          1697 => x"a33882b5",
          1698 => x"d4088c05",
          1699 => x"088c1108",
          1700 => x"81058c12",
          1701 => x"0c82b5d4",
          1702 => x"08880508",
          1703 => x"7082b5d4",
          1704 => x"08fc050c",
          1705 => x"51538a39",
          1706 => x"ff0b82b5",
          1707 => x"d408fc05",
          1708 => x"0c82b5d4",
          1709 => x"08fc0508",
          1710 => x"82b5c80c",
          1711 => x"873d0d82",
          1712 => x"b5d40c04",
          1713 => x"82b5d408",
          1714 => x"0282b5d4",
          1715 => x"0cf93d0d",
          1716 => x"82b5d408",
          1717 => x"88050885",
          1718 => x"11337081",
          1719 => x"32708106",
          1720 => x"51515152",
          1721 => x"71802e8d",
          1722 => x"38ff0b82",
          1723 => x"b5d408f8",
          1724 => x"050c8394",
          1725 => x"3982b5d4",
          1726 => x"08880508",
          1727 => x"85113370",
          1728 => x"862a7081",
          1729 => x"06515151",
          1730 => x"5271802e",
          1731 => x"80c53882",
          1732 => x"b5d40888",
          1733 => x"050882b5",
          1734 => x"d4088805",
          1735 => x"08535385",
          1736 => x"123370ff",
          1737 => x"bf065152",
          1738 => x"71851434",
          1739 => x"82b5d408",
          1740 => x"8805088c",
          1741 => x"11088105",
          1742 => x"8c120c82",
          1743 => x"b5d40888",
          1744 => x"05088411",
          1745 => x"337082b5",
          1746 => x"d408f805",
          1747 => x"0c515152",
          1748 => x"82b63982",
          1749 => x"b5d40888",
          1750 => x"05088511",
          1751 => x"3370822a",
          1752 => x"70810651",
          1753 => x"51515271",
          1754 => x"802e80d7",
          1755 => x"3882b5d4",
          1756 => x"08880508",
          1757 => x"70087033",
          1758 => x"82b5d408",
          1759 => x"fc050c51",
          1760 => x"5282b5d4",
          1761 => x"08fc0508",
          1762 => x"a93882b5",
          1763 => x"d4088805",
          1764 => x"0882b5d4",
          1765 => x"08880508",
          1766 => x"53538512",
          1767 => x"3370a007",
          1768 => x"51527185",
          1769 => x"1434ff0b",
          1770 => x"82b5d408",
          1771 => x"f8050c81",
          1772 => x"d73982b5",
          1773 => x"d4088805",
          1774 => x"08700881",
          1775 => x"05710c52",
          1776 => x"81a13982",
          1777 => x"b5d40888",
          1778 => x"050882b5",
          1779 => x"d4088805",
          1780 => x"08529411",
          1781 => x"08515271",
          1782 => x"2d82b5c8",
          1783 => x"087082b5",
          1784 => x"d408fc05",
          1785 => x"0c5282b5",
          1786 => x"d408fc05",
          1787 => x"08802580",
          1788 => x"f23882b5",
          1789 => x"d4088805",
          1790 => x"0882b5d4",
          1791 => x"08f4050c",
          1792 => x"82b5d408",
          1793 => x"88050885",
          1794 => x"113382b5",
          1795 => x"d408f005",
          1796 => x"0c5282b5",
          1797 => x"d408fc05",
          1798 => x"08ff2e09",
          1799 => x"81069538",
          1800 => x"82b5d408",
          1801 => x"f0050890",
          1802 => x"07527182",
          1803 => x"b5d408ec",
          1804 => x"05349339",
          1805 => x"82b5d408",
          1806 => x"f00508a0",
          1807 => x"07527182",
          1808 => x"b5d408ec",
          1809 => x"053482b5",
          1810 => x"d408f405",
          1811 => x"085282b5",
          1812 => x"d408ec05",
          1813 => x"33851334",
          1814 => x"ff0b82b5",
          1815 => x"d408f805",
          1816 => x"0ca63982",
          1817 => x"b5d40888",
          1818 => x"05088c11",
          1819 => x"0881058c",
          1820 => x"120c82b5",
          1821 => x"d408fc05",
          1822 => x"087081ff",
          1823 => x"067082b5",
          1824 => x"d408f805",
          1825 => x"0c515152",
          1826 => x"82b5d408",
          1827 => x"f8050882",
          1828 => x"b5c80c89",
          1829 => x"3d0d82b5",
          1830 => x"d40c0482",
          1831 => x"b5d40802",
          1832 => x"82b5d40c",
          1833 => x"fd3d0d82",
          1834 => x"b5d40888",
          1835 => x"050882b5",
          1836 => x"d408fc05",
          1837 => x"0c82b5d4",
          1838 => x"088c0508",
          1839 => x"82b5d408",
          1840 => x"f8050c82",
          1841 => x"b5d40890",
          1842 => x"0508802e",
          1843 => x"82a23882",
          1844 => x"b5d408f8",
          1845 => x"050882b5",
          1846 => x"d408fc05",
          1847 => x"082681ac",
          1848 => x"3882b5d4",
          1849 => x"08f80508",
          1850 => x"82b5d408",
          1851 => x"90050805",
          1852 => x"5182b5d4",
          1853 => x"08fc0508",
          1854 => x"71278190",
          1855 => x"3882b5d4",
          1856 => x"08fc0508",
          1857 => x"82b5d408",
          1858 => x"90050805",
          1859 => x"82b5d408",
          1860 => x"fc050c82",
          1861 => x"b5d408f8",
          1862 => x"050882b5",
          1863 => x"d4089005",
          1864 => x"080582b5",
          1865 => x"d408f805",
          1866 => x"0c82b5d4",
          1867 => x"08900508",
          1868 => x"810582b5",
          1869 => x"d4089005",
          1870 => x"0c82b5d4",
          1871 => x"08900508",
          1872 => x"ff0582b5",
          1873 => x"d4089005",
          1874 => x"0c82b5d4",
          1875 => x"08900508",
          1876 => x"802e819c",
          1877 => x"3882b5d4",
          1878 => x"08fc0508",
          1879 => x"ff0582b5",
          1880 => x"d408fc05",
          1881 => x"0c82b5d4",
          1882 => x"08f80508",
          1883 => x"ff0582b5",
          1884 => x"d408f805",
          1885 => x"0c82b5d4",
          1886 => x"08fc0508",
          1887 => x"82b5d408",
          1888 => x"f8050853",
          1889 => x"51713371",
          1890 => x"34ffae39",
          1891 => x"82b5d408",
          1892 => x"90050881",
          1893 => x"0582b5d4",
          1894 => x"0890050c",
          1895 => x"82b5d408",
          1896 => x"900508ff",
          1897 => x"0582b5d4",
          1898 => x"0890050c",
          1899 => x"82b5d408",
          1900 => x"90050880",
          1901 => x"2eba3882",
          1902 => x"b5d408f8",
          1903 => x"05085170",
          1904 => x"3382b5d4",
          1905 => x"08f80508",
          1906 => x"810582b5",
          1907 => x"d408f805",
          1908 => x"0c82b5d4",
          1909 => x"08fc0508",
          1910 => x"52527171",
          1911 => x"3482b5d4",
          1912 => x"08fc0508",
          1913 => x"810582b5",
          1914 => x"d408fc05",
          1915 => x"0cffad39",
          1916 => x"82b5d408",
          1917 => x"88050870",
          1918 => x"82b5c80c",
          1919 => x"51853d0d",
          1920 => x"82b5d40c",
          1921 => x"0482b5d4",
          1922 => x"080282b5",
          1923 => x"d40cfe3d",
          1924 => x"0d82b5d4",
          1925 => x"08880508",
          1926 => x"82b5d408",
          1927 => x"fc050c82",
          1928 => x"b5d408fc",
          1929 => x"05085271",
          1930 => x"3382b5d4",
          1931 => x"08fc0508",
          1932 => x"810582b5",
          1933 => x"d408fc05",
          1934 => x"0c7081ff",
          1935 => x"06515170",
          1936 => x"802e8338",
          1937 => x"da3982b5",
          1938 => x"d408fc05",
          1939 => x"08ff0582",
          1940 => x"b5d408fc",
          1941 => x"050c82b5",
          1942 => x"d408fc05",
          1943 => x"0882b5d4",
          1944 => x"08880508",
          1945 => x"317082b5",
          1946 => x"c80c5184",
          1947 => x"3d0d82b5",
          1948 => x"d40c0482",
          1949 => x"b5d40802",
          1950 => x"82b5d40c",
          1951 => x"fe3d0d82",
          1952 => x"b5d40888",
          1953 => x"050882b5",
          1954 => x"d408fc05",
          1955 => x"0c82b5d4",
          1956 => x"088c0508",
          1957 => x"52713382",
          1958 => x"b5d4088c",
          1959 => x"05088105",
          1960 => x"82b5d408",
          1961 => x"8c050c82",
          1962 => x"b5d408fc",
          1963 => x"05085351",
          1964 => x"70723482",
          1965 => x"b5d408fc",
          1966 => x"05088105",
          1967 => x"82b5d408",
          1968 => x"fc050c70",
          1969 => x"81ff0651",
          1970 => x"70802e84",
          1971 => x"38ffbe39",
          1972 => x"82b5d408",
          1973 => x"88050870",
          1974 => x"82b5c80c",
          1975 => x"51843d0d",
          1976 => x"82b5d40c",
          1977 => x"0482b5d4",
          1978 => x"080282b5",
          1979 => x"d40cfd3d",
          1980 => x"0d82b5d4",
          1981 => x"08880508",
          1982 => x"82b5d408",
          1983 => x"fc050c82",
          1984 => x"b5d4088c",
          1985 => x"050882b5",
          1986 => x"d408f805",
          1987 => x"0c82b5d4",
          1988 => x"08900508",
          1989 => x"802e80e5",
          1990 => x"3882b5d4",
          1991 => x"08900508",
          1992 => x"810582b5",
          1993 => x"d4089005",
          1994 => x"0c82b5d4",
          1995 => x"08900508",
          1996 => x"ff0582b5",
          1997 => x"d4089005",
          1998 => x"0c82b5d4",
          1999 => x"08900508",
          2000 => x"802eba38",
          2001 => x"82b5d408",
          2002 => x"f8050851",
          2003 => x"703382b5",
          2004 => x"d408f805",
          2005 => x"08810582",
          2006 => x"b5d408f8",
          2007 => x"050c82b5",
          2008 => x"d408fc05",
          2009 => x"08525271",
          2010 => x"713482b5",
          2011 => x"d408fc05",
          2012 => x"08810582",
          2013 => x"b5d408fc",
          2014 => x"050cffad",
          2015 => x"3982b5d4",
          2016 => x"08880508",
          2017 => x"7082b5c8",
          2018 => x"0c51853d",
          2019 => x"0d82b5d4",
          2020 => x"0c0482b5",
          2021 => x"d4080282",
          2022 => x"b5d40cfd",
          2023 => x"3d0d82b5",
          2024 => x"d4089005",
          2025 => x"08802e81",
          2026 => x"f43882b5",
          2027 => x"d4088c05",
          2028 => x"08527133",
          2029 => x"82b5d408",
          2030 => x"8c050881",
          2031 => x"0582b5d4",
          2032 => x"088c050c",
          2033 => x"82b5d408",
          2034 => x"88050870",
          2035 => x"337281ff",
          2036 => x"06535454",
          2037 => x"5171712e",
          2038 => x"843880ce",
          2039 => x"3982b5d4",
          2040 => x"08880508",
          2041 => x"52713382",
          2042 => x"b5d40888",
          2043 => x"05088105",
          2044 => x"82b5d408",
          2045 => x"88050c70",
          2046 => x"81ff0651",
          2047 => x"51708d38",
          2048 => x"800b82b5",
          2049 => x"d408fc05",
          2050 => x"0c819b39",
          2051 => x"82b5d408",
          2052 => x"900508ff",
          2053 => x"0582b5d4",
          2054 => x"0890050c",
          2055 => x"82b5d408",
          2056 => x"90050880",
          2057 => x"2e8438ff",
          2058 => x"813982b5",
          2059 => x"d4089005",
          2060 => x"08802e80",
          2061 => x"e83882b5",
          2062 => x"d4088805",
          2063 => x"08703352",
          2064 => x"53708d38",
          2065 => x"ff0b82b5",
          2066 => x"d408fc05",
          2067 => x"0c80d739",
          2068 => x"82b5d408",
          2069 => x"8c0508ff",
          2070 => x"0582b5d4",
          2071 => x"088c050c",
          2072 => x"82b5d408",
          2073 => x"8c050870",
          2074 => x"33525270",
          2075 => x"8c38810b",
          2076 => x"82b5d408",
          2077 => x"fc050cae",
          2078 => x"3982b5d4",
          2079 => x"08880508",
          2080 => x"703382b5",
          2081 => x"d4088c05",
          2082 => x"08703372",
          2083 => x"71317082",
          2084 => x"b5d408fc",
          2085 => x"050c5355",
          2086 => x"5252538a",
          2087 => x"39800b82",
          2088 => x"b5d408fc",
          2089 => x"050c82b5",
          2090 => x"d408fc05",
          2091 => x"0882b5c8",
          2092 => x"0c853d0d",
          2093 => x"82b5d40c",
          2094 => x"0482b5d4",
          2095 => x"080282b5",
          2096 => x"d40cfd3d",
          2097 => x"0d82b5d4",
          2098 => x"08880508",
          2099 => x"82b5d408",
          2100 => x"f8050c82",
          2101 => x"b5d4088c",
          2102 => x"05088d38",
          2103 => x"800b82b5",
          2104 => x"d408fc05",
          2105 => x"0c80ec39",
          2106 => x"82b5d408",
          2107 => x"f8050852",
          2108 => x"713382b5",
          2109 => x"d408f805",
          2110 => x"08810582",
          2111 => x"b5d408f8",
          2112 => x"050c7081",
          2113 => x"ff065151",
          2114 => x"70802e9f",
          2115 => x"3882b5d4",
          2116 => x"088c0508",
          2117 => x"ff0582b5",
          2118 => x"d4088c05",
          2119 => x"0c82b5d4",
          2120 => x"088c0508",
          2121 => x"ff2e8438",
          2122 => x"ffbe3982",
          2123 => x"b5d408f8",
          2124 => x"0508ff05",
          2125 => x"82b5d408",
          2126 => x"f8050c82",
          2127 => x"b5d408f8",
          2128 => x"050882b5",
          2129 => x"d4088805",
          2130 => x"08317082",
          2131 => x"b5d408fc",
          2132 => x"050c5182",
          2133 => x"b5d408fc",
          2134 => x"050882b5",
          2135 => x"c80c853d",
          2136 => x"0d82b5d4",
          2137 => x"0c0482b5",
          2138 => x"d4080282",
          2139 => x"b5d40cfe",
          2140 => x"3d0d82b5",
          2141 => x"d4088805",
          2142 => x"0882b5d4",
          2143 => x"08fc050c",
          2144 => x"82b5d408",
          2145 => x"90050880",
          2146 => x"2e80d438",
          2147 => x"82b5d408",
          2148 => x"90050881",
          2149 => x"0582b5d4",
          2150 => x"0890050c",
          2151 => x"82b5d408",
          2152 => x"900508ff",
          2153 => x"0582b5d4",
          2154 => x"0890050c",
          2155 => x"82b5d408",
          2156 => x"90050880",
          2157 => x"2ea93882",
          2158 => x"b5d4088c",
          2159 => x"05085170",
          2160 => x"82b5d408",
          2161 => x"fc050852",
          2162 => x"52717134",
          2163 => x"82b5d408",
          2164 => x"fc050881",
          2165 => x"0582b5d4",
          2166 => x"08fc050c",
          2167 => x"ffbe3982",
          2168 => x"b5d40888",
          2169 => x"05087082",
          2170 => x"b5c80c51",
          2171 => x"843d0d82",
          2172 => x"b5d40c04",
          2173 => x"82b5d408",
          2174 => x"0282b5d4",
          2175 => x"0cf93d0d",
          2176 => x"800b82b5",
          2177 => x"d408fc05",
          2178 => x"0c82b5d4",
          2179 => x"08880508",
          2180 => x"8025b938",
          2181 => x"82b5d408",
          2182 => x"88050830",
          2183 => x"82b5d408",
          2184 => x"88050c80",
          2185 => x"0b82b5d4",
          2186 => x"08f4050c",
          2187 => x"82b5d408",
          2188 => x"fc05088a",
          2189 => x"38810b82",
          2190 => x"b5d408f4",
          2191 => x"050c82b5",
          2192 => x"d408f405",
          2193 => x"0882b5d4",
          2194 => x"08fc050c",
          2195 => x"82b5d408",
          2196 => x"8c050880",
          2197 => x"25b93882",
          2198 => x"b5d4088c",
          2199 => x"05083082",
          2200 => x"b5d4088c",
          2201 => x"050c800b",
          2202 => x"82b5d408",
          2203 => x"f0050c82",
          2204 => x"b5d408fc",
          2205 => x"05088a38",
          2206 => x"810b82b5",
          2207 => x"d408f005",
          2208 => x"0c82b5d4",
          2209 => x"08f00508",
          2210 => x"82b5d408",
          2211 => x"fc050c80",
          2212 => x"5382b5d4",
          2213 => x"088c0508",
          2214 => x"5282b5d4",
          2215 => x"08880508",
          2216 => x"5182c53f",
          2217 => x"82b5c808",
          2218 => x"7082b5d4",
          2219 => x"08f8050c",
          2220 => x"5482b5d4",
          2221 => x"08fc0508",
          2222 => x"802e9038",
          2223 => x"82b5d408",
          2224 => x"f8050830",
          2225 => x"82b5d408",
          2226 => x"f8050c82",
          2227 => x"b5d408f8",
          2228 => x"05087082",
          2229 => x"b5c80c54",
          2230 => x"893d0d82",
          2231 => x"b5d40c04",
          2232 => x"82b5d408",
          2233 => x"0282b5d4",
          2234 => x"0cfb3d0d",
          2235 => x"800b82b5",
          2236 => x"d408fc05",
          2237 => x"0c82b5d4",
          2238 => x"08880508",
          2239 => x"80259938",
          2240 => x"82b5d408",
          2241 => x"88050830",
          2242 => x"82b5d408",
          2243 => x"88050c81",
          2244 => x"0b82b5d4",
          2245 => x"08fc050c",
          2246 => x"82b5d408",
          2247 => x"8c050880",
          2248 => x"25903882",
          2249 => x"b5d4088c",
          2250 => x"05083082",
          2251 => x"b5d4088c",
          2252 => x"050c8153",
          2253 => x"82b5d408",
          2254 => x"8c050852",
          2255 => x"82b5d408",
          2256 => x"88050851",
          2257 => x"81a23f82",
          2258 => x"b5c80870",
          2259 => x"82b5d408",
          2260 => x"f8050c54",
          2261 => x"82b5d408",
          2262 => x"fc050880",
          2263 => x"2e903882",
          2264 => x"b5d408f8",
          2265 => x"05083082",
          2266 => x"b5d408f8",
          2267 => x"050c82b5",
          2268 => x"d408f805",
          2269 => x"087082b5",
          2270 => x"c80c5487",
          2271 => x"3d0d82b5",
          2272 => x"d40c0482",
          2273 => x"b5d40802",
          2274 => x"82b5d40c",
          2275 => x"fd3d0d80",
          2276 => x"5382b5d4",
          2277 => x"088c0508",
          2278 => x"5282b5d4",
          2279 => x"08880508",
          2280 => x"5180c53f",
          2281 => x"82b5c808",
          2282 => x"7082b5c8",
          2283 => x"0c54853d",
          2284 => x"0d82b5d4",
          2285 => x"0c0482b5",
          2286 => x"d4080282",
          2287 => x"b5d40cfd",
          2288 => x"3d0d8153",
          2289 => x"82b5d408",
          2290 => x"8c050852",
          2291 => x"82b5d408",
          2292 => x"88050851",
          2293 => x"933f82b5",
          2294 => x"c8087082",
          2295 => x"b5c80c54",
          2296 => x"853d0d82",
          2297 => x"b5d40c04",
          2298 => x"82b5d408",
          2299 => x"0282b5d4",
          2300 => x"0cfd3d0d",
          2301 => x"810b82b5",
          2302 => x"d408fc05",
          2303 => x"0c800b82",
          2304 => x"b5d408f8",
          2305 => x"050c82b5",
          2306 => x"d4088c05",
          2307 => x"0882b5d4",
          2308 => x"08880508",
          2309 => x"27b93882",
          2310 => x"b5d408fc",
          2311 => x"0508802e",
          2312 => x"ae38800b",
          2313 => x"82b5d408",
          2314 => x"8c050824",
          2315 => x"a23882b5",
          2316 => x"d4088c05",
          2317 => x"081082b5",
          2318 => x"d4088c05",
          2319 => x"0c82b5d4",
          2320 => x"08fc0508",
          2321 => x"1082b5d4",
          2322 => x"08fc050c",
          2323 => x"ffb83982",
          2324 => x"b5d408fc",
          2325 => x"0508802e",
          2326 => x"80e13882",
          2327 => x"b5d4088c",
          2328 => x"050882b5",
          2329 => x"d4088805",
          2330 => x"0826ad38",
          2331 => x"82b5d408",
          2332 => x"88050882",
          2333 => x"b5d4088c",
          2334 => x"05083182",
          2335 => x"b5d40888",
          2336 => x"050c82b5",
          2337 => x"d408f805",
          2338 => x"0882b5d4",
          2339 => x"08fc0508",
          2340 => x"0782b5d4",
          2341 => x"08f8050c",
          2342 => x"82b5d408",
          2343 => x"fc050881",
          2344 => x"2a82b5d4",
          2345 => x"08fc050c",
          2346 => x"82b5d408",
          2347 => x"8c050881",
          2348 => x"2a82b5d4",
          2349 => x"088c050c",
          2350 => x"ff953982",
          2351 => x"b5d40890",
          2352 => x"0508802e",
          2353 => x"933882b5",
          2354 => x"d4088805",
          2355 => x"087082b5",
          2356 => x"d408f405",
          2357 => x"0c519139",
          2358 => x"82b5d408",
          2359 => x"f8050870",
          2360 => x"82b5d408",
          2361 => x"f4050c51",
          2362 => x"82b5d408",
          2363 => x"f4050882",
          2364 => x"b5c80c85",
          2365 => x"3d0d82b5",
          2366 => x"d40c0482",
          2367 => x"b5d40802",
          2368 => x"82b5d40c",
          2369 => x"f73d0d80",
          2370 => x"0b82b5d4",
          2371 => x"08f00534",
          2372 => x"82b5d408",
          2373 => x"8c050853",
          2374 => x"80730c82",
          2375 => x"b5d40888",
          2376 => x"05087008",
          2377 => x"51537233",
          2378 => x"537282b5",
          2379 => x"d408f805",
          2380 => x"347281ff",
          2381 => x"065372a0",
          2382 => x"2e098106",
          2383 => x"913882b5",
          2384 => x"d4088805",
          2385 => x"08700881",
          2386 => x"05710c53",
          2387 => x"ce3982b5",
          2388 => x"d408f805",
          2389 => x"335372ad",
          2390 => x"2e098106",
          2391 => x"a438810b",
          2392 => x"82b5d408",
          2393 => x"f0053482",
          2394 => x"b5d40888",
          2395 => x"05087008",
          2396 => x"8105710c",
          2397 => x"70085153",
          2398 => x"723382b5",
          2399 => x"d408f805",
          2400 => x"3482b5d4",
          2401 => x"08f80533",
          2402 => x"5372b02e",
          2403 => x"09810681",
          2404 => x"dc3882b5",
          2405 => x"d4088805",
          2406 => x"08700881",
          2407 => x"05710c70",
          2408 => x"08515372",
          2409 => x"3382b5d4",
          2410 => x"08f80534",
          2411 => x"82b5d408",
          2412 => x"f8053382",
          2413 => x"b5d408e8",
          2414 => x"050c82b5",
          2415 => x"d408e805",
          2416 => x"0880e22e",
          2417 => x"b63882b5",
          2418 => x"d408e805",
          2419 => x"0880f82e",
          2420 => x"843880cd",
          2421 => x"39900b82",
          2422 => x"b5d408f4",
          2423 => x"053482b5",
          2424 => x"d4088805",
          2425 => x"08700881",
          2426 => x"05710c70",
          2427 => x"08515372",
          2428 => x"3382b5d4",
          2429 => x"08f80534",
          2430 => x"81a43982",
          2431 => x"0b82b5d4",
          2432 => x"08f40534",
          2433 => x"82b5d408",
          2434 => x"88050870",
          2435 => x"08810571",
          2436 => x"0c700851",
          2437 => x"53723382",
          2438 => x"b5d408f8",
          2439 => x"053480fe",
          2440 => x"3982b5d4",
          2441 => x"08f80533",
          2442 => x"5372a026",
          2443 => x"8d38810b",
          2444 => x"82b5d408",
          2445 => x"ec050c83",
          2446 => x"803982b5",
          2447 => x"d408f805",
          2448 => x"3353af73",
          2449 => x"27903882",
          2450 => x"b5d408f8",
          2451 => x"05335372",
          2452 => x"b9268338",
          2453 => x"8d39800b",
          2454 => x"82b5d408",
          2455 => x"ec050c82",
          2456 => x"d839880b",
          2457 => x"82b5d408",
          2458 => x"f40534b2",
          2459 => x"3982b5d4",
          2460 => x"08f80533",
          2461 => x"53af7327",
          2462 => x"903882b5",
          2463 => x"d408f805",
          2464 => x"335372b9",
          2465 => x"2683388d",
          2466 => x"39800b82",
          2467 => x"b5d408ec",
          2468 => x"050c82a5",
          2469 => x"398a0b82",
          2470 => x"b5d408f4",
          2471 => x"0534800b",
          2472 => x"82b5d408",
          2473 => x"fc050c82",
          2474 => x"b5d408f8",
          2475 => x"053353a0",
          2476 => x"732781cf",
          2477 => x"3882b5d4",
          2478 => x"08f80533",
          2479 => x"5380e073",
          2480 => x"27943882",
          2481 => x"b5d408f8",
          2482 => x"0533e011",
          2483 => x"51537282",
          2484 => x"b5d408f8",
          2485 => x"053482b5",
          2486 => x"d408f805",
          2487 => x"33d01151",
          2488 => x"537282b5",
          2489 => x"d408f805",
          2490 => x"3482b5d4",
          2491 => x"08f80533",
          2492 => x"53907327",
          2493 => x"ad3882b5",
          2494 => x"d408f805",
          2495 => x"33f91151",
          2496 => x"537282b5",
          2497 => x"d408f805",
          2498 => x"3482b5d4",
          2499 => x"08f80533",
          2500 => x"53728926",
          2501 => x"8d38800b",
          2502 => x"82b5d408",
          2503 => x"ec050c81",
          2504 => x"983982b5",
          2505 => x"d408f805",
          2506 => x"3382b5d4",
          2507 => x"08f40533",
          2508 => x"54547274",
          2509 => x"268d3880",
          2510 => x"0b82b5d4",
          2511 => x"08ec050c",
          2512 => x"80f73982",
          2513 => x"b5d408f4",
          2514 => x"05337082",
          2515 => x"b5d408fc",
          2516 => x"05082982",
          2517 => x"b5d408f8",
          2518 => x"05337012",
          2519 => x"82b5d408",
          2520 => x"fc050c82",
          2521 => x"b5d40888",
          2522 => x"05087008",
          2523 => x"8105710c",
          2524 => x"70085151",
          2525 => x"52555372",
          2526 => x"3382b5d4",
          2527 => x"08f80534",
          2528 => x"fea53982",
          2529 => x"b5d408f0",
          2530 => x"05335372",
          2531 => x"802e9038",
          2532 => x"82b5d408",
          2533 => x"fc050830",
          2534 => x"82b5d408",
          2535 => x"fc050c82",
          2536 => x"b5d4088c",
          2537 => x"050882b5",
          2538 => x"d408fc05",
          2539 => x"08710c53",
          2540 => x"810b82b5",
          2541 => x"d408ec05",
          2542 => x"0c82b5d4",
          2543 => x"08ec0508",
          2544 => x"82b5c80c",
          2545 => x"8b3d0d82",
          2546 => x"b5d40c04",
          2547 => x"82b5d408",
          2548 => x"0282b5d4",
          2549 => x"0cf73d0d",
          2550 => x"800b82b5",
          2551 => x"d408f005",
          2552 => x"3482b5d4",
          2553 => x"088c0508",
          2554 => x"5380730c",
          2555 => x"82b5d408",
          2556 => x"88050870",
          2557 => x"08515372",
          2558 => x"33537282",
          2559 => x"b5d408f8",
          2560 => x"05347281",
          2561 => x"ff065372",
          2562 => x"a02e0981",
          2563 => x"06913882",
          2564 => x"b5d40888",
          2565 => x"05087008",
          2566 => x"8105710c",
          2567 => x"53ce3982",
          2568 => x"b5d408f8",
          2569 => x"05335372",
          2570 => x"ad2e0981",
          2571 => x"06a43881",
          2572 => x"0b82b5d4",
          2573 => x"08f00534",
          2574 => x"82b5d408",
          2575 => x"88050870",
          2576 => x"08810571",
          2577 => x"0c700851",
          2578 => x"53723382",
          2579 => x"b5d408f8",
          2580 => x"053482b5",
          2581 => x"d408f805",
          2582 => x"335372b0",
          2583 => x"2e098106",
          2584 => x"81dc3882",
          2585 => x"b5d40888",
          2586 => x"05087008",
          2587 => x"8105710c",
          2588 => x"70085153",
          2589 => x"723382b5",
          2590 => x"d408f805",
          2591 => x"3482b5d4",
          2592 => x"08f80533",
          2593 => x"82b5d408",
          2594 => x"e8050c82",
          2595 => x"b5d408e8",
          2596 => x"050880e2",
          2597 => x"2eb63882",
          2598 => x"b5d408e8",
          2599 => x"050880f8",
          2600 => x"2e843880",
          2601 => x"cd39900b",
          2602 => x"82b5d408",
          2603 => x"f4053482",
          2604 => x"b5d40888",
          2605 => x"05087008",
          2606 => x"8105710c",
          2607 => x"70085153",
          2608 => x"723382b5",
          2609 => x"d408f805",
          2610 => x"3481a439",
          2611 => x"820b82b5",
          2612 => x"d408f405",
          2613 => x"3482b5d4",
          2614 => x"08880508",
          2615 => x"70088105",
          2616 => x"710c7008",
          2617 => x"51537233",
          2618 => x"82b5d408",
          2619 => x"f8053480",
          2620 => x"fe3982b5",
          2621 => x"d408f805",
          2622 => x"335372a0",
          2623 => x"268d3881",
          2624 => x"0b82b5d4",
          2625 => x"08ec050c",
          2626 => x"83803982",
          2627 => x"b5d408f8",
          2628 => x"053353af",
          2629 => x"73279038",
          2630 => x"82b5d408",
          2631 => x"f8053353",
          2632 => x"72b92683",
          2633 => x"388d3980",
          2634 => x"0b82b5d4",
          2635 => x"08ec050c",
          2636 => x"82d83988",
          2637 => x"0b82b5d4",
          2638 => x"08f40534",
          2639 => x"b23982b5",
          2640 => x"d408f805",
          2641 => x"3353af73",
          2642 => x"27903882",
          2643 => x"b5d408f8",
          2644 => x"05335372",
          2645 => x"b9268338",
          2646 => x"8d39800b",
          2647 => x"82b5d408",
          2648 => x"ec050c82",
          2649 => x"a5398a0b",
          2650 => x"82b5d408",
          2651 => x"f4053480",
          2652 => x"0b82b5d4",
          2653 => x"08fc050c",
          2654 => x"82b5d408",
          2655 => x"f8053353",
          2656 => x"a0732781",
          2657 => x"cf3882b5",
          2658 => x"d408f805",
          2659 => x"335380e0",
          2660 => x"73279438",
          2661 => x"82b5d408",
          2662 => x"f80533e0",
          2663 => x"11515372",
          2664 => x"82b5d408",
          2665 => x"f8053482",
          2666 => x"b5d408f8",
          2667 => x"0533d011",
          2668 => x"51537282",
          2669 => x"b5d408f8",
          2670 => x"053482b5",
          2671 => x"d408f805",
          2672 => x"33539073",
          2673 => x"27ad3882",
          2674 => x"b5d408f8",
          2675 => x"0533f911",
          2676 => x"51537282",
          2677 => x"b5d408f8",
          2678 => x"053482b5",
          2679 => x"d408f805",
          2680 => x"33537289",
          2681 => x"268d3880",
          2682 => x"0b82b5d4",
          2683 => x"08ec050c",
          2684 => x"81983982",
          2685 => x"b5d408f8",
          2686 => x"053382b5",
          2687 => x"d408f405",
          2688 => x"33545472",
          2689 => x"74268d38",
          2690 => x"800b82b5",
          2691 => x"d408ec05",
          2692 => x"0c80f739",
          2693 => x"82b5d408",
          2694 => x"f4053370",
          2695 => x"82b5d408",
          2696 => x"fc050829",
          2697 => x"82b5d408",
          2698 => x"f8053370",
          2699 => x"1282b5d4",
          2700 => x"08fc050c",
          2701 => x"82b5d408",
          2702 => x"88050870",
          2703 => x"08810571",
          2704 => x"0c700851",
          2705 => x"51525553",
          2706 => x"723382b5",
          2707 => x"d408f805",
          2708 => x"34fea539",
          2709 => x"82b5d408",
          2710 => x"f0053353",
          2711 => x"72802e90",
          2712 => x"3882b5d4",
          2713 => x"08fc0508",
          2714 => x"3082b5d4",
          2715 => x"08fc050c",
          2716 => x"82b5d408",
          2717 => x"8c050882",
          2718 => x"b5d408fc",
          2719 => x"0508710c",
          2720 => x"53810b82",
          2721 => x"b5d408ec",
          2722 => x"050c82b5",
          2723 => x"d408ec05",
          2724 => x"0882b5c8",
          2725 => x"0c8b3d0d",
          2726 => x"82b5d40c",
          2727 => x"04f93d0d",
          2728 => x"79700870",
          2729 => x"56565874",
          2730 => x"802e80e3",
          2731 => x"38953975",
          2732 => x"0851e6d1",
          2733 => x"3f82b5c8",
          2734 => x"0815780c",
          2735 => x"85163354",
          2736 => x"80cd3974",
          2737 => x"335473a0",
          2738 => x"2e098106",
          2739 => x"86388115",
          2740 => x"55f13980",
          2741 => x"57769029",
          2742 => x"82b0c805",
          2743 => x"70085256",
          2744 => x"e6a33f82",
          2745 => x"b5c80853",
          2746 => x"74527508",
          2747 => x"51e9a33f",
          2748 => x"82b5c808",
          2749 => x"8b388416",
          2750 => x"33547381",
          2751 => x"2effb038",
          2752 => x"81177081",
          2753 => x"ff065854",
          2754 => x"997727c9",
          2755 => x"38ff5473",
          2756 => x"82b5c80c",
          2757 => x"893d0d04",
          2758 => x"ff3d0d73",
          2759 => x"52719326",
          2760 => x"818e3871",
          2761 => x"84298295",
          2762 => x"a8055271",
          2763 => x"0804829a",
          2764 => x"f4518180",
          2765 => x"39829b80",
          2766 => x"5180f939",
          2767 => x"829b9051",
          2768 => x"80f23982",
          2769 => x"9ba05180",
          2770 => x"eb39829b",
          2771 => x"b05180e4",
          2772 => x"39829bc0",
          2773 => x"5180dd39",
          2774 => x"829bd451",
          2775 => x"80d63982",
          2776 => x"9be45180",
          2777 => x"cf39829b",
          2778 => x"fc5180c8",
          2779 => x"39829c94",
          2780 => x"5180c139",
          2781 => x"829cac51",
          2782 => x"bb39829c",
          2783 => x"c851b539",
          2784 => x"829cdc51",
          2785 => x"af39829d",
          2786 => x"8451a939",
          2787 => x"829d9451",
          2788 => x"a339829d",
          2789 => x"b4519d39",
          2790 => x"829dc451",
          2791 => x"9739829d",
          2792 => x"dc519139",
          2793 => x"829df451",
          2794 => x"8b39829e",
          2795 => x"8c518539",
          2796 => x"829e9851",
          2797 => x"d8ad3f83",
          2798 => x"3d0d04fb",
          2799 => x"3d0d7779",
          2800 => x"56567487",
          2801 => x"e7268a38",
          2802 => x"74527587",
          2803 => x"e8295190",
          2804 => x"3987e852",
          2805 => x"7451efab",
          2806 => x"3f82b5c8",
          2807 => x"08527551",
          2808 => x"efa13f82",
          2809 => x"b5c80854",
          2810 => x"79537552",
          2811 => x"829ea851",
          2812 => x"ffbbe53f",
          2813 => x"873d0d04",
          2814 => x"ec3d0d66",
          2815 => x"02840580",
          2816 => x"e305335b",
          2817 => x"57806878",
          2818 => x"30707a07",
          2819 => x"73255157",
          2820 => x"59597856",
          2821 => x"7787ff26",
          2822 => x"83388156",
          2823 => x"74760770",
          2824 => x"81ff0651",
          2825 => x"55935674",
          2826 => x"81823881",
          2827 => x"5376528c",
          2828 => x"3d705256",
          2829 => x"80ffc53f",
          2830 => x"82b5c808",
          2831 => x"5782b5c8",
          2832 => x"08b93882",
          2833 => x"b5c80887",
          2834 => x"c098880c",
          2835 => x"82b5c808",
          2836 => x"59963dd4",
          2837 => x"05548480",
          2838 => x"53775275",
          2839 => x"51818481",
          2840 => x"3f82b5c8",
          2841 => x"085782b5",
          2842 => x"c8089038",
          2843 => x"7a557480",
          2844 => x"2e893874",
          2845 => x"19751959",
          2846 => x"59d73996",
          2847 => x"3dd80551",
          2848 => x"818bea3f",
          2849 => x"76307078",
          2850 => x"0780257b",
          2851 => x"30709f2a",
          2852 => x"72065157",
          2853 => x"51567480",
          2854 => x"2e903882",
          2855 => x"9ecc5387",
          2856 => x"c0988808",
          2857 => x"527851fe",
          2858 => x"923f7656",
          2859 => x"7582b5c8",
          2860 => x"0c963d0d",
          2861 => x"04f83d0d",
          2862 => x"7c028405",
          2863 => x"b7053358",
          2864 => x"59ff5880",
          2865 => x"537b527a",
          2866 => x"51fead3f",
          2867 => x"82b5c808",
          2868 => x"a8387680",
          2869 => x"2e883876",
          2870 => x"812e9c38",
          2871 => x"9c3982cd",
          2872 => x"98566155",
          2873 => x"605482b5",
          2874 => x"c8537f52",
          2875 => x"7e51782d",
          2876 => x"82b5c808",
          2877 => x"58833978",
          2878 => x"047782b5",
          2879 => x"c80c8a3d",
          2880 => x"0d04f33d",
          2881 => x"0d7f6163",
          2882 => x"028c0580",
          2883 => x"cf053373",
          2884 => x"73156841",
          2885 => x"5f5c5c5e",
          2886 => x"5e5e7a52",
          2887 => x"829ed451",
          2888 => x"ffb9b53f",
          2889 => x"829edc51",
          2890 => x"ffb9ad3f",
          2891 => x"80557479",
          2892 => x"27818038",
          2893 => x"7b902e89",
          2894 => x"387ba02e",
          2895 => x"a73880c6",
          2896 => x"39741853",
          2897 => x"727a278e",
          2898 => x"38722252",
          2899 => x"829ee051",
          2900 => x"ffb9853f",
          2901 => x"8939829e",
          2902 => x"ec51ffb8",
          2903 => x"fb3f8215",
          2904 => x"5580c339",
          2905 => x"74185372",
          2906 => x"7a278e38",
          2907 => x"72085282",
          2908 => x"9ed451ff",
          2909 => x"b8e23f89",
          2910 => x"39829ee8",
          2911 => x"51ffb8d8",
          2912 => x"3f841555",
          2913 => x"a1397418",
          2914 => x"53727a27",
          2915 => x"8e387233",
          2916 => x"52829ef4",
          2917 => x"51ffb8c0",
          2918 => x"3f893982",
          2919 => x"9efc51ff",
          2920 => x"b8b63f81",
          2921 => x"155582cd",
          2922 => x"9c0852a0",
          2923 => x"51d8833f",
          2924 => x"fefc3982",
          2925 => x"9f8051ff",
          2926 => x"b89e3f80",
          2927 => x"55747927",
          2928 => x"80c63874",
          2929 => x"18703355",
          2930 => x"53805672",
          2931 => x"7a278338",
          2932 => x"81568053",
          2933 => x"9f742783",
          2934 => x"38815375",
          2935 => x"73067081",
          2936 => x"ff065153",
          2937 => x"72802e90",
          2938 => x"387380fe",
          2939 => x"268a3882",
          2940 => x"cd9c0852",
          2941 => x"73518839",
          2942 => x"82cd9c08",
          2943 => x"52a051d7",
          2944 => x"b13f8115",
          2945 => x"55ffb639",
          2946 => x"829f8451",
          2947 => x"d3d53f78",
          2948 => x"18791c5c",
          2949 => x"589ccb3f",
          2950 => x"82b5c808",
          2951 => x"982b7098",
          2952 => x"2c515776",
          2953 => x"a02e0981",
          2954 => x"06aa389c",
          2955 => x"b53f82b5",
          2956 => x"c808982b",
          2957 => x"70982c70",
          2958 => x"a0327030",
          2959 => x"729b3270",
          2960 => x"30707207",
          2961 => x"73750706",
          2962 => x"51585859",
          2963 => x"57515780",
          2964 => x"7324d838",
          2965 => x"769b2e09",
          2966 => x"81068538",
          2967 => x"80538c39",
          2968 => x"7c1e5372",
          2969 => x"7826fdb2",
          2970 => x"38ff5372",
          2971 => x"82b5c80c",
          2972 => x"8f3d0d04",
          2973 => x"fc3d0d02",
          2974 => x"9b053382",
          2975 => x"9f885382",
          2976 => x"9f8c5255",
          2977 => x"ffb6d13f",
          2978 => x"82b4a022",
          2979 => x"51a5a63f",
          2980 => x"829f9854",
          2981 => x"829fa453",
          2982 => x"82b4a133",
          2983 => x"52829fac",
          2984 => x"51ffb6b4",
          2985 => x"3f74802e",
          2986 => x"8438a0d8",
          2987 => x"3f863d0d",
          2988 => x"04fe3d0d",
          2989 => x"87c09680",
          2990 => x"0853a5c2",
          2991 => x"3f815198",
          2992 => x"8e3f829f",
          2993 => x"c85199a3",
          2994 => x"3f805198",
          2995 => x"823f7281",
          2996 => x"2a708106",
          2997 => x"51527180",
          2998 => x"2e923881",
          2999 => x"5197f03f",
          3000 => x"829fe051",
          3001 => x"99853f80",
          3002 => x"5197e43f",
          3003 => x"72822a70",
          3004 => x"81065152",
          3005 => x"71802e92",
          3006 => x"38815197",
          3007 => x"d23f829f",
          3008 => x"f05198e7",
          3009 => x"3f805197",
          3010 => x"c63f7283",
          3011 => x"2a708106",
          3012 => x"51527180",
          3013 => x"2e923881",
          3014 => x"5197b43f",
          3015 => x"82a08051",
          3016 => x"98c93f80",
          3017 => x"5197a83f",
          3018 => x"72842a70",
          3019 => x"81065152",
          3020 => x"71802e92",
          3021 => x"38815197",
          3022 => x"963f82a0",
          3023 => x"945198ab",
          3024 => x"3f805197",
          3025 => x"8a3f7285",
          3026 => x"2a708106",
          3027 => x"51527180",
          3028 => x"2e923881",
          3029 => x"5196f83f",
          3030 => x"82a0a851",
          3031 => x"988d3f80",
          3032 => x"5196ec3f",
          3033 => x"72862a70",
          3034 => x"81065152",
          3035 => x"71802e92",
          3036 => x"38815196",
          3037 => x"da3f82a0",
          3038 => x"bc5197ef",
          3039 => x"3f805196",
          3040 => x"ce3f7287",
          3041 => x"2a708106",
          3042 => x"51527180",
          3043 => x"2e923881",
          3044 => x"5196bc3f",
          3045 => x"82a0d051",
          3046 => x"97d13f80",
          3047 => x"5196b03f",
          3048 => x"72882a70",
          3049 => x"81065152",
          3050 => x"71802e92",
          3051 => x"38815196",
          3052 => x"9e3f82a0",
          3053 => x"e45197b3",
          3054 => x"3f805196",
          3055 => x"923fa3c6",
          3056 => x"3f843d0d",
          3057 => x"04fb3d0d",
          3058 => x"77028405",
          3059 => x"a3053370",
          3060 => x"55565680",
          3061 => x"527551e3",
          3062 => x"8d3f0b0b",
          3063 => x"82b0c433",
          3064 => x"5473a938",
          3065 => x"815382a1",
          3066 => x"a05282cc",
          3067 => x"c85180f8",
          3068 => x"8b3f82b5",
          3069 => x"c8083070",
          3070 => x"82b5c808",
          3071 => x"07802582",
          3072 => x"71315151",
          3073 => x"54730b0b",
          3074 => x"82b0c434",
          3075 => x"0b0b82b0",
          3076 => x"c4335473",
          3077 => x"812e0981",
          3078 => x"06af3882",
          3079 => x"ccc85374",
          3080 => x"52755181",
          3081 => x"b2bc3f82",
          3082 => x"b5c80880",
          3083 => x"2e8b3882",
          3084 => x"b5c80851",
          3085 => x"cfad3f91",
          3086 => x"3982ccc8",
          3087 => x"518184ad",
          3088 => x"3f820b0b",
          3089 => x"0b82b0c4",
          3090 => x"340b0b82",
          3091 => x"b0c43354",
          3092 => x"73822e09",
          3093 => x"81068c38",
          3094 => x"82a1b053",
          3095 => x"74527551",
          3096 => x"a9be3f80",
          3097 => x"0b82b5c8",
          3098 => x"0c873d0d",
          3099 => x"04ce3d0d",
          3100 => x"80707182",
          3101 => x"ccc40c5f",
          3102 => x"5d81527c",
          3103 => x"5180c6d7",
          3104 => x"3f82b5c8",
          3105 => x"0881ff06",
          3106 => x"59787d2e",
          3107 => x"098106a3",
          3108 => x"38963d59",
          3109 => x"835382a1",
          3110 => x"b8527851",
          3111 => x"dcc73f7c",
          3112 => x"53785282",
          3113 => x"b6f45180",
          3114 => x"f5f13f82",
          3115 => x"b5c8087d",
          3116 => x"2e883882",
          3117 => x"a1bc518d",
          3118 => x"a3398170",
          3119 => x"5f5d82a1",
          3120 => x"f451ffb2",
          3121 => x"933f963d",
          3122 => x"70465a80",
          3123 => x"f8527951",
          3124 => x"fdf33fb4",
          3125 => x"3dff8405",
          3126 => x"51f3c23f",
          3127 => x"82b5c808",
          3128 => x"902b7090",
          3129 => x"2c515978",
          3130 => x"80c22e87",
          3131 => x"a3387880",
          3132 => x"c224b238",
          3133 => x"78bd2e81",
          3134 => x"d23878bd",
          3135 => x"24903878",
          3136 => x"802effba",
          3137 => x"3878bc2e",
          3138 => x"80da388a",
          3139 => x"d4397880",
          3140 => x"c02e8399",
          3141 => x"387880c0",
          3142 => x"2485cd38",
          3143 => x"78bf2e82",
          3144 => x"8c388abd",
          3145 => x"397880f9",
          3146 => x"2e89d938",
          3147 => x"7880f924",
          3148 => x"92387880",
          3149 => x"c32e8888",
          3150 => x"387880f8",
          3151 => x"2e89a138",
          3152 => x"8a9f3978",
          3153 => x"81832e8a",
          3154 => x"86387881",
          3155 => x"83248b38",
          3156 => x"7881822e",
          3157 => x"89eb388a",
          3158 => x"88397881",
          3159 => x"852e89fb",
          3160 => x"3889fe39",
          3161 => x"b43dff80",
          3162 => x"1153ff84",
          3163 => x"0551ecdc",
          3164 => x"3f82b5c8",
          3165 => x"08802efe",
          3166 => x"c538b43d",
          3167 => x"fefc1153",
          3168 => x"ff840551",
          3169 => x"ecc63f82",
          3170 => x"b5c80880",
          3171 => x"2efeaf38",
          3172 => x"b43dfef8",
          3173 => x"1153ff84",
          3174 => x"0551ecb0",
          3175 => x"3f82b5c8",
          3176 => x"08863882",
          3177 => x"b5c80842",
          3178 => x"82a1f851",
          3179 => x"ffb0a93f",
          3180 => x"63635c5a",
          3181 => x"797b2781",
          3182 => x"ec386159",
          3183 => x"787a7084",
          3184 => x"055c0c7a",
          3185 => x"7a26f538",
          3186 => x"81db39b4",
          3187 => x"3dff8011",
          3188 => x"53ff8405",
          3189 => x"51ebf53f",
          3190 => x"82b5c808",
          3191 => x"802efdde",
          3192 => x"38b43dfe",
          3193 => x"fc1153ff",
          3194 => x"840551eb",
          3195 => x"df3f82b5",
          3196 => x"c808802e",
          3197 => x"fdc838b4",
          3198 => x"3dfef811",
          3199 => x"53ff8405",
          3200 => x"51ebc93f",
          3201 => x"82b5c808",
          3202 => x"802efdb2",
          3203 => x"3882a288",
          3204 => x"51ffafc4",
          3205 => x"3f635a79",
          3206 => x"63278189",
          3207 => x"38615979",
          3208 => x"7081055b",
          3209 => x"33793461",
          3210 => x"810542eb",
          3211 => x"39b43dff",
          3212 => x"801153ff",
          3213 => x"840551eb",
          3214 => x"933f82b5",
          3215 => x"c808802e",
          3216 => x"fcfc38b4",
          3217 => x"3dfefc11",
          3218 => x"53ff8405",
          3219 => x"51eafd3f",
          3220 => x"82b5c808",
          3221 => x"802efce6",
          3222 => x"38b43dfe",
          3223 => x"f81153ff",
          3224 => x"840551ea",
          3225 => x"e73f82b5",
          3226 => x"c808802e",
          3227 => x"fcd03882",
          3228 => x"a29451ff",
          3229 => x"aee23f63",
          3230 => x"5a796327",
          3231 => x"a8386170",
          3232 => x"337b335e",
          3233 => x"5a5b787c",
          3234 => x"2e923878",
          3235 => x"557a5479",
          3236 => x"33537952",
          3237 => x"82a2a451",
          3238 => x"ffaebd3f",
          3239 => x"811a6281",
          3240 => x"05435ad5",
          3241 => x"398a51cd",
          3242 => x"dc3ffc92",
          3243 => x"39b43dff",
          3244 => x"801153ff",
          3245 => x"840551ea",
          3246 => x"933f82b5",
          3247 => x"c80880df",
          3248 => x"3882b4b4",
          3249 => x"33597880",
          3250 => x"2e893882",
          3251 => x"b3ec0844",
          3252 => x"80cd3982",
          3253 => x"b4b53359",
          3254 => x"78802e88",
          3255 => x"3882b3f4",
          3256 => x"0844bc39",
          3257 => x"82b4b633",
          3258 => x"5978802e",
          3259 => x"883882b3",
          3260 => x"fc0844ab",
          3261 => x"3982b4b7",
          3262 => x"33597880",
          3263 => x"2e883882",
          3264 => x"b4840844",
          3265 => x"9a3982b4",
          3266 => x"b2335978",
          3267 => x"802e8838",
          3268 => x"82b48c08",
          3269 => x"44893982",
          3270 => x"b49c08fc",
          3271 => x"800544b4",
          3272 => x"3dfefc11",
          3273 => x"53ff8405",
          3274 => x"51e9a13f",
          3275 => x"82b5c808",
          3276 => x"80de3882",
          3277 => x"b4b43359",
          3278 => x"78802e89",
          3279 => x"3882b3f0",
          3280 => x"084380cc",
          3281 => x"3982b4b5",
          3282 => x"33597880",
          3283 => x"2e883882",
          3284 => x"b3f80843",
          3285 => x"bb3982b4",
          3286 => x"b6335978",
          3287 => x"802e8838",
          3288 => x"82b48008",
          3289 => x"43aa3982",
          3290 => x"b4b73359",
          3291 => x"78802e88",
          3292 => x"3882b488",
          3293 => x"08439939",
          3294 => x"82b4b233",
          3295 => x"5978802e",
          3296 => x"883882b4",
          3297 => x"90084388",
          3298 => x"3982b49c",
          3299 => x"08880543",
          3300 => x"b43dfef8",
          3301 => x"1153ff84",
          3302 => x"0551e8b0",
          3303 => x"3f82b5c8",
          3304 => x"08802ea7",
          3305 => x"3880625c",
          3306 => x"5c7a882e",
          3307 => x"8338815c",
          3308 => x"7a903270",
          3309 => x"30707207",
          3310 => x"9f2a707f",
          3311 => x"0651515a",
          3312 => x"5a78802e",
          3313 => x"88387aa0",
          3314 => x"2e833888",
          3315 => x"4282a2c0",
          3316 => x"51c8903f",
          3317 => x"a0556354",
          3318 => x"61536252",
          3319 => x"6351f2a2",
          3320 => x"3f82a2cc",
          3321 => x"5186f539",
          3322 => x"b43dff80",
          3323 => x"1153ff84",
          3324 => x"0551e7d8",
          3325 => x"3f82b5c8",
          3326 => x"08802ef9",
          3327 => x"c138b43d",
          3328 => x"fefc1153",
          3329 => x"ff840551",
          3330 => x"e7c23f82",
          3331 => x"b5c80880",
          3332 => x"2ea43863",
          3333 => x"590280cb",
          3334 => x"05337934",
          3335 => x"63810544",
          3336 => x"b43dfefc",
          3337 => x"1153ff84",
          3338 => x"0551e7a0",
          3339 => x"3f82b5c8",
          3340 => x"08e138f9",
          3341 => x"89396370",
          3342 => x"33545282",
          3343 => x"a2d851ff",
          3344 => x"ab963f82",
          3345 => x"cd980853",
          3346 => x"80f85279",
          3347 => x"51ffabdd",
          3348 => x"3f794579",
          3349 => x"335978ae",
          3350 => x"2ef8e338",
          3351 => x"9f79279f",
          3352 => x"38b43dfe",
          3353 => x"fc1153ff",
          3354 => x"840551e6",
          3355 => x"df3f82b5",
          3356 => x"c808802e",
          3357 => x"91386359",
          3358 => x"0280cb05",
          3359 => x"33793463",
          3360 => x"810544ff",
          3361 => x"b13982a2",
          3362 => x"e451c6d7",
          3363 => x"3fffa739",
          3364 => x"b43dfef4",
          3365 => x"1153ff84",
          3366 => x"0551e0df",
          3367 => x"3f82b5c8",
          3368 => x"08802ef8",
          3369 => x"9938b43d",
          3370 => x"fef01153",
          3371 => x"ff840551",
          3372 => x"e0c93f82",
          3373 => x"b5c80880",
          3374 => x"2ea53860",
          3375 => x"5902be05",
          3376 => x"22797082",
          3377 => x"055b2378",
          3378 => x"41b43dfe",
          3379 => x"f01153ff",
          3380 => x"840551e0",
          3381 => x"a63f82b5",
          3382 => x"c808e038",
          3383 => x"f7e03960",
          3384 => x"70225452",
          3385 => x"82a2e851",
          3386 => x"ffa9ed3f",
          3387 => x"82cd9808",
          3388 => x"5380f852",
          3389 => x"7951ffaa",
          3390 => x"b43f7945",
          3391 => x"79335978",
          3392 => x"ae2ef7ba",
          3393 => x"38789f26",
          3394 => x"87386082",
          3395 => x"0541d039",
          3396 => x"b43dfef0",
          3397 => x"1153ff84",
          3398 => x"0551dfdf",
          3399 => x"3f82b5c8",
          3400 => x"08802e92",
          3401 => x"38605902",
          3402 => x"be052279",
          3403 => x"7082055b",
          3404 => x"237841ff",
          3405 => x"aa3982a2",
          3406 => x"e451c5a7",
          3407 => x"3fffa039",
          3408 => x"b43dfef4",
          3409 => x"1153ff84",
          3410 => x"0551dfaf",
          3411 => x"3f82b5c8",
          3412 => x"08802ef6",
          3413 => x"e938b43d",
          3414 => x"fef01153",
          3415 => x"ff840551",
          3416 => x"df993f82",
          3417 => x"b5c80880",
          3418 => x"2ea03860",
          3419 => x"60710c59",
          3420 => x"60840541",
          3421 => x"b43dfef0",
          3422 => x"1153ff84",
          3423 => x"0551defb",
          3424 => x"3f82b5c8",
          3425 => x"08e538f6",
          3426 => x"b5396070",
          3427 => x"08545282",
          3428 => x"a2f451ff",
          3429 => x"a8c23f82",
          3430 => x"cd980853",
          3431 => x"80f85279",
          3432 => x"51ffa989",
          3433 => x"3f794579",
          3434 => x"335978ae",
          3435 => x"2ef68f38",
          3436 => x"9f79279b",
          3437 => x"38b43dfe",
          3438 => x"f01153ff",
          3439 => x"840551de",
          3440 => x"ba3f82b5",
          3441 => x"c808802e",
          3442 => x"8d386060",
          3443 => x"710c5960",
          3444 => x"840541ff",
          3445 => x"b53982a2",
          3446 => x"e451c487",
          3447 => x"3fffab39",
          3448 => x"b43dff80",
          3449 => x"1153ff84",
          3450 => x"0551e3e0",
          3451 => x"3f82b5c8",
          3452 => x"08802ef5",
          3453 => x"c9386352",
          3454 => x"82a38451",
          3455 => x"ffa7d93f",
          3456 => x"63597804",
          3457 => x"b43dff80",
          3458 => x"1153ff84",
          3459 => x"0551e3bc",
          3460 => x"3f82b5c8",
          3461 => x"08802ef5",
          3462 => x"a5386352",
          3463 => x"82a3a051",
          3464 => x"ffa7b53f",
          3465 => x"6359782d",
          3466 => x"82b5c808",
          3467 => x"802ef58e",
          3468 => x"3882b5c8",
          3469 => x"085282a3",
          3470 => x"bc51ffa7",
          3471 => x"9b3ff4fe",
          3472 => x"3982a3d8",
          3473 => x"51c39c3f",
          3474 => x"ffa6ee3f",
          3475 => x"f4f03982",
          3476 => x"a3f451c3",
          3477 => x"8e3f8059",
          3478 => x"ffa83991",
          3479 => x"a73ff4de",
          3480 => x"39794579",
          3481 => x"33597880",
          3482 => x"2ef4d338",
          3483 => x"7d7d0659",
          3484 => x"78802e81",
          3485 => x"cf38b43d",
          3486 => x"ff840551",
          3487 => x"83ca3f82",
          3488 => x"b5c8085c",
          3489 => x"815b7a82",
          3490 => x"2eb2387a",
          3491 => x"82248938",
          3492 => x"7a812e8c",
          3493 => x"3880ca39",
          3494 => x"7a832ead",
          3495 => x"3880c239",
          3496 => x"82a48856",
          3497 => x"7b5582a4",
          3498 => x"8c548053",
          3499 => x"82a49052",
          3500 => x"b43dffb0",
          3501 => x"0551ffa9",
          3502 => x"873fb839",
          3503 => x"7b52b43d",
          3504 => x"ffb00551",
          3505 => x"cfad3fab",
          3506 => x"397b5582",
          3507 => x"a48c5480",
          3508 => x"5382a4a0",
          3509 => x"52b43dff",
          3510 => x"b00551ff",
          3511 => x"a8e23f93",
          3512 => x"397b5480",
          3513 => x"5382a4ac",
          3514 => x"52b43dff",
          3515 => x"b00551ff",
          3516 => x"a8ce3f82",
          3517 => x"b3ec5882",
          3518 => x"b5f85780",
          3519 => x"56645580",
          3520 => x"5482d080",
          3521 => x"5382d080",
          3522 => x"52b43dff",
          3523 => x"b00551eb",
          3524 => x"a43f82b5",
          3525 => x"c80882b5",
          3526 => x"c8080970",
          3527 => x"30707207",
          3528 => x"8025515b",
          3529 => x"5b5f805a",
          3530 => x"7a832683",
          3531 => x"38815a78",
          3532 => x"7a065978",
          3533 => x"802e8d38",
          3534 => x"811b7081",
          3535 => x"ff065c59",
          3536 => x"7afec338",
          3537 => x"7d81327d",
          3538 => x"81320759",
          3539 => x"788a387e",
          3540 => x"ff2e0981",
          3541 => x"06f2e738",
          3542 => x"82a4b451",
          3543 => x"c1853ff2",
          3544 => x"dd39f53d",
          3545 => x"0d800b82",
          3546 => x"b5f83487",
          3547 => x"c0948c70",
          3548 => x"08545587",
          3549 => x"84805272",
          3550 => x"51d8883f",
          3551 => x"82b5c808",
          3552 => x"902b7508",
          3553 => x"55538784",
          3554 => x"80527351",
          3555 => x"d7f53f72",
          3556 => x"82b5c808",
          3557 => x"07750c87",
          3558 => x"c0949c70",
          3559 => x"08545587",
          3560 => x"84805272",
          3561 => x"51d7dc3f",
          3562 => x"82b5c808",
          3563 => x"902b7508",
          3564 => x"55538784",
          3565 => x"80527351",
          3566 => x"d7c93f72",
          3567 => x"82b5c808",
          3568 => x"07750c8c",
          3569 => x"80830b87",
          3570 => x"c094840c",
          3571 => x"8c80830b",
          3572 => x"87c09494",
          3573 => x"0c80f5e7",
          3574 => x"5a80f8d3",
          3575 => x"5b830284",
          3576 => x"05990534",
          3577 => x"805c82cd",
          3578 => x"980b873d",
          3579 => x"7088130c",
          3580 => x"70720c82",
          3581 => x"cd9c0c54",
          3582 => x"89be3f93",
          3583 => x"813f82a4",
          3584 => x"c451ffbf",
          3585 => x"de3f82a4",
          3586 => x"d051ffbf",
          3587 => x"d63f80dd",
          3588 => x"b15192e5",
          3589 => x"3f8151ec",
          3590 => x"db3ff0d1",
          3591 => x"3f8004fe",
          3592 => x"3d0d8052",
          3593 => x"83537188",
          3594 => x"2b5287d8",
          3595 => x"3f82b5c8",
          3596 => x"0881ff06",
          3597 => x"7207ff14",
          3598 => x"54527280",
          3599 => x"25e83871",
          3600 => x"82b5c80c",
          3601 => x"843d0d04",
          3602 => x"fc3d0d76",
          3603 => x"70085455",
          3604 => x"80735254",
          3605 => x"72742e81",
          3606 => x"8a387233",
          3607 => x"5170a02e",
          3608 => x"09810686",
          3609 => x"38811353",
          3610 => x"f1397233",
          3611 => x"5170a22e",
          3612 => x"09810686",
          3613 => x"38811353",
          3614 => x"81547252",
          3615 => x"73812e09",
          3616 => x"81069f38",
          3617 => x"84398112",
          3618 => x"52807233",
          3619 => x"525470a2",
          3620 => x"2e833881",
          3621 => x"5470802e",
          3622 => x"9d3873ea",
          3623 => x"38983981",
          3624 => x"12528072",
          3625 => x"33525470",
          3626 => x"a02e8338",
          3627 => x"81547080",
          3628 => x"2e843873",
          3629 => x"ea388072",
          3630 => x"33525470",
          3631 => x"a02e0981",
          3632 => x"06833881",
          3633 => x"5470a232",
          3634 => x"70307080",
          3635 => x"25760751",
          3636 => x"51517080",
          3637 => x"2e883880",
          3638 => x"72708105",
          3639 => x"54347175",
          3640 => x"0c725170",
          3641 => x"82b5c80c",
          3642 => x"863d0d04",
          3643 => x"fc3d0d76",
          3644 => x"53720880",
          3645 => x"2e913886",
          3646 => x"3dfc0552",
          3647 => x"7251d7fb",
          3648 => x"3f82b5c8",
          3649 => x"08853880",
          3650 => x"53833974",
          3651 => x"537282b5",
          3652 => x"c80c863d",
          3653 => x"0d04fc3d",
          3654 => x"0d768211",
          3655 => x"33ff0552",
          3656 => x"53815270",
          3657 => x"8b268198",
          3658 => x"38831333",
          3659 => x"ff055182",
          3660 => x"52709e26",
          3661 => x"818a3884",
          3662 => x"13335183",
          3663 => x"52709726",
          3664 => x"80fe3885",
          3665 => x"13335184",
          3666 => x"5270bb26",
          3667 => x"80f23886",
          3668 => x"13335185",
          3669 => x"5270bb26",
          3670 => x"80e63888",
          3671 => x"13225586",
          3672 => x"527487e7",
          3673 => x"2680d938",
          3674 => x"8a132254",
          3675 => x"87527387",
          3676 => x"e72680cc",
          3677 => x"38810b87",
          3678 => x"c0989c0c",
          3679 => x"722287c0",
          3680 => x"98bc0c82",
          3681 => x"133387c0",
          3682 => x"98b80c83",
          3683 => x"133387c0",
          3684 => x"98b40c84",
          3685 => x"133387c0",
          3686 => x"98b00c85",
          3687 => x"133387c0",
          3688 => x"98ac0c86",
          3689 => x"133387c0",
          3690 => x"98a80c74",
          3691 => x"87c098a4",
          3692 => x"0c7387c0",
          3693 => x"98a00c80",
          3694 => x"0b87c098",
          3695 => x"9c0c8052",
          3696 => x"7182b5c8",
          3697 => x"0c863d0d",
          3698 => x"04f33d0d",
          3699 => x"7f5b87c0",
          3700 => x"989c5d81",
          3701 => x"7d0c87c0",
          3702 => x"98bc085e",
          3703 => x"7d7b2387",
          3704 => x"c098b808",
          3705 => x"5a79821c",
          3706 => x"3487c098",
          3707 => x"b4085a79",
          3708 => x"831c3487",
          3709 => x"c098b008",
          3710 => x"5a79841c",
          3711 => x"3487c098",
          3712 => x"ac085a79",
          3713 => x"851c3487",
          3714 => x"c098a808",
          3715 => x"5a79861c",
          3716 => x"3487c098",
          3717 => x"a4085c7b",
          3718 => x"881c2387",
          3719 => x"c098a008",
          3720 => x"5a798a1c",
          3721 => x"23807d0c",
          3722 => x"7983ffff",
          3723 => x"06597b83",
          3724 => x"ffff0658",
          3725 => x"861b3357",
          3726 => x"851b3356",
          3727 => x"841b3355",
          3728 => x"831b3354",
          3729 => x"821b3353",
          3730 => x"7d83ffff",
          3731 => x"065282a4",
          3732 => x"e851ff9f",
          3733 => x"833f8f3d",
          3734 => x"0d04fb3d",
          3735 => x"0d029f05",
          3736 => x"3382b3e8",
          3737 => x"337081ff",
          3738 => x"06585555",
          3739 => x"87c09484",
          3740 => x"5175802e",
          3741 => x"863887c0",
          3742 => x"94945170",
          3743 => x"0870962a",
          3744 => x"70810653",
          3745 => x"54527080",
          3746 => x"2e8c3871",
          3747 => x"912a7081",
          3748 => x"06515170",
          3749 => x"d7387281",
          3750 => x"32708106",
          3751 => x"51517080",
          3752 => x"2e8d3871",
          3753 => x"932a7081",
          3754 => x"06515170",
          3755 => x"ffbe3873",
          3756 => x"81ff0651",
          3757 => x"87c09480",
          3758 => x"5270802e",
          3759 => x"863887c0",
          3760 => x"94905274",
          3761 => x"720c7482",
          3762 => x"b5c80c87",
          3763 => x"3d0d04ff",
          3764 => x"3d0d028f",
          3765 => x"05337030",
          3766 => x"709f2a51",
          3767 => x"52527082",
          3768 => x"b3e83483",
          3769 => x"3d0d04f9",
          3770 => x"3d0d02a7",
          3771 => x"05335877",
          3772 => x"8a2e0981",
          3773 => x"0687387a",
          3774 => x"528d51eb",
          3775 => x"3f82b3e8",
          3776 => x"337081ff",
          3777 => x"06585687",
          3778 => x"c0948453",
          3779 => x"76802e86",
          3780 => x"3887c094",
          3781 => x"94537208",
          3782 => x"70962a70",
          3783 => x"81065556",
          3784 => x"5472802e",
          3785 => x"8c387391",
          3786 => x"2a708106",
          3787 => x"515372d7",
          3788 => x"38748132",
          3789 => x"70810651",
          3790 => x"5372802e",
          3791 => x"8d387393",
          3792 => x"2a708106",
          3793 => x"515372ff",
          3794 => x"be387581",
          3795 => x"ff065387",
          3796 => x"c0948054",
          3797 => x"72802e86",
          3798 => x"3887c094",
          3799 => x"90547774",
          3800 => x"0c800b82",
          3801 => x"b5c80c89",
          3802 => x"3d0d04f9",
          3803 => x"3d0d7954",
          3804 => x"80743370",
          3805 => x"81ff0653",
          3806 => x"53577077",
          3807 => x"2e80fc38",
          3808 => x"7181ff06",
          3809 => x"811582b3",
          3810 => x"e8337081",
          3811 => x"ff065957",
          3812 => x"555887c0",
          3813 => x"94845175",
          3814 => x"802e8638",
          3815 => x"87c09494",
          3816 => x"51700870",
          3817 => x"962a7081",
          3818 => x"06535452",
          3819 => x"70802e8c",
          3820 => x"3871912a",
          3821 => x"70810651",
          3822 => x"5170d738",
          3823 => x"72813270",
          3824 => x"81065151",
          3825 => x"70802e8d",
          3826 => x"3871932a",
          3827 => x"70810651",
          3828 => x"5170ffbe",
          3829 => x"387481ff",
          3830 => x"065187c0",
          3831 => x"94805270",
          3832 => x"802e8638",
          3833 => x"87c09490",
          3834 => x"5277720c",
          3835 => x"81177433",
          3836 => x"7081ff06",
          3837 => x"53535770",
          3838 => x"ff863876",
          3839 => x"82b5c80c",
          3840 => x"893d0d04",
          3841 => x"fe3d0d82",
          3842 => x"b3e83370",
          3843 => x"81ff0654",
          3844 => x"5287c094",
          3845 => x"84517280",
          3846 => x"2e863887",
          3847 => x"c0949451",
          3848 => x"70087082",
          3849 => x"2a708106",
          3850 => x"51515170",
          3851 => x"802ee238",
          3852 => x"7181ff06",
          3853 => x"5187c094",
          3854 => x"80527080",
          3855 => x"2e863887",
          3856 => x"c0949052",
          3857 => x"71087081",
          3858 => x"ff0682b5",
          3859 => x"c80c5184",
          3860 => x"3d0d04ff",
          3861 => x"af3f82b5",
          3862 => x"c80881ff",
          3863 => x"0682b5c8",
          3864 => x"0c04fe3d",
          3865 => x"0d82b3e8",
          3866 => x"337081ff",
          3867 => x"06525387",
          3868 => x"c0948452",
          3869 => x"70802e86",
          3870 => x"3887c094",
          3871 => x"94527108",
          3872 => x"70822a70",
          3873 => x"81065151",
          3874 => x"51ff5270",
          3875 => x"802ea038",
          3876 => x"7281ff06",
          3877 => x"5187c094",
          3878 => x"80527080",
          3879 => x"2e863887",
          3880 => x"c0949052",
          3881 => x"71087098",
          3882 => x"2b70982c",
          3883 => x"51535171",
          3884 => x"82b5c80c",
          3885 => x"843d0d04",
          3886 => x"ff3d0d87",
          3887 => x"c09e8008",
          3888 => x"709c2a8a",
          3889 => x"06515170",
          3890 => x"802e84b4",
          3891 => x"3887c09e",
          3892 => x"a40882b3",
          3893 => x"ec0c87c0",
          3894 => x"9ea80882",
          3895 => x"b3f00c87",
          3896 => x"c09e9408",
          3897 => x"82b3f40c",
          3898 => x"87c09e98",
          3899 => x"0882b3f8",
          3900 => x"0c87c09e",
          3901 => x"9c0882b3",
          3902 => x"fc0c87c0",
          3903 => x"9ea00882",
          3904 => x"b4800c87",
          3905 => x"c09eac08",
          3906 => x"82b4840c",
          3907 => x"87c09eb0",
          3908 => x"0882b488",
          3909 => x"0c87c09e",
          3910 => x"b40882b4",
          3911 => x"8c0c87c0",
          3912 => x"9eb80882",
          3913 => x"b4900c87",
          3914 => x"c09ebc08",
          3915 => x"82b4940c",
          3916 => x"87c09ec0",
          3917 => x"0882b498",
          3918 => x"0c87c09e",
          3919 => x"c40882b4",
          3920 => x"9c0c87c0",
          3921 => x"9e800851",
          3922 => x"7082b4a0",
          3923 => x"2387c09e",
          3924 => x"840882b4",
          3925 => x"a40c87c0",
          3926 => x"9e880882",
          3927 => x"b4a80c87",
          3928 => x"c09e8c08",
          3929 => x"82b4ac0c",
          3930 => x"810b82b4",
          3931 => x"b034800b",
          3932 => x"87c09e90",
          3933 => x"08708480",
          3934 => x"0a065152",
          3935 => x"5270802e",
          3936 => x"83388152",
          3937 => x"7182b4b1",
          3938 => x"34800b87",
          3939 => x"c09e9008",
          3940 => x"7088800a",
          3941 => x"06515252",
          3942 => x"70802e83",
          3943 => x"38815271",
          3944 => x"82b4b234",
          3945 => x"800b87c0",
          3946 => x"9e900870",
          3947 => x"90800a06",
          3948 => x"51525270",
          3949 => x"802e8338",
          3950 => x"81527182",
          3951 => x"b4b33480",
          3952 => x"0b87c09e",
          3953 => x"90087088",
          3954 => x"80800651",
          3955 => x"52527080",
          3956 => x"2e833881",
          3957 => x"527182b4",
          3958 => x"b434800b",
          3959 => x"87c09e90",
          3960 => x"0870a080",
          3961 => x"80065152",
          3962 => x"5270802e",
          3963 => x"83388152",
          3964 => x"7182b4b5",
          3965 => x"34800b87",
          3966 => x"c09e9008",
          3967 => x"70908080",
          3968 => x"06515252",
          3969 => x"70802e83",
          3970 => x"38815271",
          3971 => x"82b4b634",
          3972 => x"800b87c0",
          3973 => x"9e900870",
          3974 => x"84808006",
          3975 => x"51525270",
          3976 => x"802e8338",
          3977 => x"81527182",
          3978 => x"b4b73480",
          3979 => x"0b87c09e",
          3980 => x"90087082",
          3981 => x"80800651",
          3982 => x"52527080",
          3983 => x"2e833881",
          3984 => x"527182b4",
          3985 => x"b834800b",
          3986 => x"87c09e90",
          3987 => x"08708180",
          3988 => x"80065152",
          3989 => x"5270802e",
          3990 => x"83388152",
          3991 => x"7182b4b9",
          3992 => x"34800b87",
          3993 => x"c09e9008",
          3994 => x"7080c080",
          3995 => x"06515252",
          3996 => x"70802e83",
          3997 => x"38815271",
          3998 => x"82b4ba34",
          3999 => x"800b87c0",
          4000 => x"9e900870",
          4001 => x"a0800651",
          4002 => x"52527080",
          4003 => x"2e833881",
          4004 => x"527182b4",
          4005 => x"bb3487c0",
          4006 => x"9e900870",
          4007 => x"98800670",
          4008 => x"8a2a5151",
          4009 => x"517082b4",
          4010 => x"bc34800b",
          4011 => x"87c09e90",
          4012 => x"08708480",
          4013 => x"06515252",
          4014 => x"70802e83",
          4015 => x"38815271",
          4016 => x"82b4bd34",
          4017 => x"87c09e90",
          4018 => x"087083f0",
          4019 => x"0670842a",
          4020 => x"51515170",
          4021 => x"82b4be34",
          4022 => x"800b87c0",
          4023 => x"9e900870",
          4024 => x"88065152",
          4025 => x"5270802e",
          4026 => x"83388152",
          4027 => x"7182b4bf",
          4028 => x"3487c09e",
          4029 => x"90087087",
          4030 => x"06515170",
          4031 => x"82b4c034",
          4032 => x"833d0d04",
          4033 => x"fb3d0d82",
          4034 => x"a58051ff",
          4035 => x"b1d53f82",
          4036 => x"b4b03354",
          4037 => x"73802e89",
          4038 => x"3882a594",
          4039 => x"51ffb1c3",
          4040 => x"3f82a5a8",
          4041 => x"51ffb1bb",
          4042 => x"3f82b4b2",
          4043 => x"33547380",
          4044 => x"2e943882",
          4045 => x"b48c0882",
          4046 => x"b4900811",
          4047 => x"545282a5",
          4048 => x"c051ff95",
          4049 => x"933f82b4",
          4050 => x"b7335473",
          4051 => x"802e9438",
          4052 => x"82b48408",
          4053 => x"82b48808",
          4054 => x"11545282",
          4055 => x"a5dc51ff",
          4056 => x"94f63f82",
          4057 => x"b4b43354",
          4058 => x"73802e94",
          4059 => x"3882b3ec",
          4060 => x"0882b3f0",
          4061 => x"08115452",
          4062 => x"82a5f851",
          4063 => x"ff94d93f",
          4064 => x"82b4b533",
          4065 => x"5473802e",
          4066 => x"943882b3",
          4067 => x"f40882b3",
          4068 => x"f8081154",
          4069 => x"5282a694",
          4070 => x"51ff94bc",
          4071 => x"3f82b4b6",
          4072 => x"33547380",
          4073 => x"2e943882",
          4074 => x"b3fc0882",
          4075 => x"b4800811",
          4076 => x"545282a6",
          4077 => x"b051ff94",
          4078 => x"9f3f82b4",
          4079 => x"bb335473",
          4080 => x"802e8e38",
          4081 => x"82b4bc33",
          4082 => x"5282a6cc",
          4083 => x"51ff9488",
          4084 => x"3f82b4bf",
          4085 => x"33547380",
          4086 => x"2e8e3882",
          4087 => x"b4c03352",
          4088 => x"82a6ec51",
          4089 => x"ff93f13f",
          4090 => x"82b4bd33",
          4091 => x"5473802e",
          4092 => x"8e3882b4",
          4093 => x"be335282",
          4094 => x"a78c51ff",
          4095 => x"93da3f82",
          4096 => x"b4b13354",
          4097 => x"73802e89",
          4098 => x"3882a7ac",
          4099 => x"51ffafd3",
          4100 => x"3f82b4b3",
          4101 => x"33547380",
          4102 => x"2e893882",
          4103 => x"a7c051ff",
          4104 => x"afc13f82",
          4105 => x"b4b83354",
          4106 => x"73802e89",
          4107 => x"3882a7cc",
          4108 => x"51ffafaf",
          4109 => x"3f82b4b9",
          4110 => x"33547380",
          4111 => x"2e893882",
          4112 => x"a7d851ff",
          4113 => x"af9d3f82",
          4114 => x"b4ba3354",
          4115 => x"73802e89",
          4116 => x"3882a7e4",
          4117 => x"51ffaf8b",
          4118 => x"3f82a7f0",
          4119 => x"51ffaf83",
          4120 => x"3f82b494",
          4121 => x"085282a7",
          4122 => x"fc51ff92",
          4123 => x"eb3f82b4",
          4124 => x"98085282",
          4125 => x"a8a451ff",
          4126 => x"92de3f82",
          4127 => x"b49c0852",
          4128 => x"82a8cc51",
          4129 => x"ff92d13f",
          4130 => x"82a8f451",
          4131 => x"ffaed43f",
          4132 => x"82b4a022",
          4133 => x"5282a8fc",
          4134 => x"51ff92bc",
          4135 => x"3f82b4a4",
          4136 => x"0856bd84",
          4137 => x"c0527551",
          4138 => x"c5d93f82",
          4139 => x"b5c808bd",
          4140 => x"84c02976",
          4141 => x"71315454",
          4142 => x"82b5c808",
          4143 => x"5282a9a4",
          4144 => x"51ff9294",
          4145 => x"3f82b4b7",
          4146 => x"33547380",
          4147 => x"2ea93882",
          4148 => x"b4a80856",
          4149 => x"bd84c052",
          4150 => x"7551c5a7",
          4151 => x"3f82b5c8",
          4152 => x"08bd84c0",
          4153 => x"29767131",
          4154 => x"545482b5",
          4155 => x"c8085282",
          4156 => x"a9d051ff",
          4157 => x"91e23f82",
          4158 => x"b4b23354",
          4159 => x"73802ea9",
          4160 => x"3882b4ac",
          4161 => x"0856bd84",
          4162 => x"c0527551",
          4163 => x"c4f53f82",
          4164 => x"b5c808bd",
          4165 => x"84c02976",
          4166 => x"71315454",
          4167 => x"82b5c808",
          4168 => x"5282a9fc",
          4169 => x"51ff91b0",
          4170 => x"3f82a2bc",
          4171 => x"51ffadb3",
          4172 => x"3f873d0d",
          4173 => x"04fe3d0d",
          4174 => x"02920533",
          4175 => x"ff055271",
          4176 => x"8426aa38",
          4177 => x"71842982",
          4178 => x"95f80552",
          4179 => x"71080482",
          4180 => x"aaa8519d",
          4181 => x"3982aab0",
          4182 => x"51973982",
          4183 => x"aab85191",
          4184 => x"3982aac0",
          4185 => x"518b3982",
          4186 => x"aac45185",
          4187 => x"3982aacc",
          4188 => x"51ffacef",
          4189 => x"3f843d0d",
          4190 => x"04718880",
          4191 => x"0c04800b",
          4192 => x"87c09684",
          4193 => x"0c0482b4",
          4194 => x"c40887c0",
          4195 => x"96840c04",
          4196 => x"fd3d0d76",
          4197 => x"982b7098",
          4198 => x"2c79982b",
          4199 => x"70982c72",
          4200 => x"10137082",
          4201 => x"2b515351",
          4202 => x"54515180",
          4203 => x"0b82aad8",
          4204 => x"12335553",
          4205 => x"7174259c",
          4206 => x"3882aad4",
          4207 => x"11081202",
          4208 => x"84059705",
          4209 => x"33713352",
          4210 => x"52527072",
          4211 => x"2e098106",
          4212 => x"83388153",
          4213 => x"7282b5c8",
          4214 => x"0c853d0d",
          4215 => x"04fb3d0d",
          4216 => x"79028405",
          4217 => x"a3053371",
          4218 => x"33555654",
          4219 => x"72802eb1",
          4220 => x"3882cd9c",
          4221 => x"08528851",
          4222 => x"ffafb73f",
          4223 => x"82cd9c08",
          4224 => x"52a051ff",
          4225 => x"afac3f82",
          4226 => x"cd9c0852",
          4227 => x"8851ffaf",
          4228 => x"a13f7333",
          4229 => x"ff055372",
          4230 => x"74347281",
          4231 => x"ff0653cc",
          4232 => x"397751ff",
          4233 => x"8fb23f74",
          4234 => x"7434873d",
          4235 => x"0d04f63d",
          4236 => x"0d7c0284",
          4237 => x"05b70533",
          4238 => x"028805bb",
          4239 => x"053382b5",
          4240 => x"a0337084",
          4241 => x"2982b4c8",
          4242 => x"05700851",
          4243 => x"59595a58",
          4244 => x"5974802e",
          4245 => x"86387451",
          4246 => x"9afa3f82",
          4247 => x"b5a03370",
          4248 => x"842982b4",
          4249 => x"c8058119",
          4250 => x"70545856",
          4251 => x"5a9dfb3f",
          4252 => x"82b5c808",
          4253 => x"750c82b5",
          4254 => x"a0337084",
          4255 => x"2982b4c8",
          4256 => x"05700851",
          4257 => x"565a7480",
          4258 => x"2ea73875",
          4259 => x"53785274",
          4260 => x"51ffb8d1",
          4261 => x"3f82b5a0",
          4262 => x"33810555",
          4263 => x"7482b5a0",
          4264 => x"347481ff",
          4265 => x"06559375",
          4266 => x"27873880",
          4267 => x"0b82b5a0",
          4268 => x"3477802e",
          4269 => x"b63882b5",
          4270 => x"9c085675",
          4271 => x"802eac38",
          4272 => x"82b59833",
          4273 => x"5574a438",
          4274 => x"8c3dfc05",
          4275 => x"54765378",
          4276 => x"52755180",
          4277 => x"da883f82",
          4278 => x"b59c0852",
          4279 => x"8a51818f",
          4280 => x"953f82b5",
          4281 => x"9c085180",
          4282 => x"dde53f8c",
          4283 => x"3d0d04fd",
          4284 => x"3d0d82b4",
          4285 => x"c8539354",
          4286 => x"72085271",
          4287 => x"802e8938",
          4288 => x"715199d0",
          4289 => x"3f80730c",
          4290 => x"ff148414",
          4291 => x"54547380",
          4292 => x"25e63880",
          4293 => x"0b82b5a0",
          4294 => x"3482b59c",
          4295 => x"08527180",
          4296 => x"2e953871",
          4297 => x"5180dec5",
          4298 => x"3f82b59c",
          4299 => x"085199a4",
          4300 => x"3f800b82",
          4301 => x"b59c0c85",
          4302 => x"3d0d04dc",
          4303 => x"3d0d8157",
          4304 => x"805282b5",
          4305 => x"9c085180",
          4306 => x"e3b23f82",
          4307 => x"b5c80880",
          4308 => x"d33882b5",
          4309 => x"9c085380",
          4310 => x"f852883d",
          4311 => x"70525681",
          4312 => x"8c803f82",
          4313 => x"b5c80880",
          4314 => x"2eba3875",
          4315 => x"51ffb595",
          4316 => x"3f82b5c8",
          4317 => x"0855800b",
          4318 => x"82b5c808",
          4319 => x"259d3882",
          4320 => x"b5c808ff",
          4321 => x"05701755",
          4322 => x"55807434",
          4323 => x"75537652",
          4324 => x"811782ad",
          4325 => x"c85257ff",
          4326 => x"8cbe3f74",
          4327 => x"ff2e0981",
          4328 => x"06ffaf38",
          4329 => x"a63d0d04",
          4330 => x"d93d0daa",
          4331 => x"3d08ad3d",
          4332 => x"085a5a81",
          4333 => x"70585880",
          4334 => x"5282b59c",
          4335 => x"085180e2",
          4336 => x"bb3f82b5",
          4337 => x"c8088195",
          4338 => x"38ff0b82",
          4339 => x"b59c0854",
          4340 => x"5580f852",
          4341 => x"8b3d7052",
          4342 => x"56818b86",
          4343 => x"3f82b5c8",
          4344 => x"08802ea5",
          4345 => x"387551ff",
          4346 => x"b49b3f82",
          4347 => x"b5c80881",
          4348 => x"18585580",
          4349 => x"0b82b5c8",
          4350 => x"08258e38",
          4351 => x"82b5c808",
          4352 => x"ff057017",
          4353 => x"55558074",
          4354 => x"34740970",
          4355 => x"30707207",
          4356 => x"9f2a5155",
          4357 => x"5578772e",
          4358 => x"853873ff",
          4359 => x"ac3882b5",
          4360 => x"9c088c11",
          4361 => x"08535180",
          4362 => x"e1d23f82",
          4363 => x"b5c80880",
          4364 => x"2e893882",
          4365 => x"add451ff",
          4366 => x"8b9e3f78",
          4367 => x"772e0981",
          4368 => x"069b3875",
          4369 => x"527951ff",
          4370 => x"b4a93f79",
          4371 => x"51ffb3b5",
          4372 => x"3fab3d08",
          4373 => x"5482b5c8",
          4374 => x"08743480",
          4375 => x"587782b5",
          4376 => x"c80ca93d",
          4377 => x"0d04f63d",
          4378 => x"0d7c7e71",
          4379 => x"5c717233",
          4380 => x"57595a58",
          4381 => x"73a02e09",
          4382 => x"8106a238",
          4383 => x"78337805",
          4384 => x"56777627",
          4385 => x"98388117",
          4386 => x"705b7071",
          4387 => x"33565855",
          4388 => x"73a02e09",
          4389 => x"81068638",
          4390 => x"757526ea",
          4391 => x"38805473",
          4392 => x"882982b5",
          4393 => x"a4057008",
          4394 => x"5255ffb2",
          4395 => x"d83f82b5",
          4396 => x"c8085379",
          4397 => x"52740851",
          4398 => x"ffb5d73f",
          4399 => x"82b5c808",
          4400 => x"80c53884",
          4401 => x"15335574",
          4402 => x"812e8838",
          4403 => x"74822e88",
          4404 => x"38b539fc",
          4405 => x"e63fac39",
          4406 => x"811a5a8c",
          4407 => x"3dfc1153",
          4408 => x"f80551c5",
          4409 => x"e73f82b5",
          4410 => x"c808802e",
          4411 => x"9a38ff1b",
          4412 => x"53785277",
          4413 => x"51fdb13f",
          4414 => x"82b5c808",
          4415 => x"81ff0655",
          4416 => x"74853874",
          4417 => x"54913981",
          4418 => x"147081ff",
          4419 => x"06515482",
          4420 => x"7427ff8b",
          4421 => x"38805473",
          4422 => x"82b5c80c",
          4423 => x"8c3d0d04",
          4424 => x"d33d0db0",
          4425 => x"3d08b23d",
          4426 => x"08b43d08",
          4427 => x"595f5a80",
          4428 => x"0baf3d34",
          4429 => x"82b5a033",
          4430 => x"82b59c08",
          4431 => x"555b7381",
          4432 => x"cb387382",
          4433 => x"b5983355",
          4434 => x"55738338",
          4435 => x"81557680",
          4436 => x"2e81bc38",
          4437 => x"81707606",
          4438 => x"55567380",
          4439 => x"2e81ad38",
          4440 => x"a8519886",
          4441 => x"3f82b5c8",
          4442 => x"0882b59c",
          4443 => x"0c82b5c8",
          4444 => x"08802e81",
          4445 => x"92389353",
          4446 => x"765282b5",
          4447 => x"c8085180",
          4448 => x"ccfa3f82",
          4449 => x"b5c80880",
          4450 => x"2e8c3882",
          4451 => x"ae8051ff",
          4452 => x"a4d13f80",
          4453 => x"f73982b5",
          4454 => x"c8085b82",
          4455 => x"b59c0853",
          4456 => x"80f85290",
          4457 => x"3d705254",
          4458 => x"8187b73f",
          4459 => x"82b5c808",
          4460 => x"5682b5c8",
          4461 => x"08742e09",
          4462 => x"810680d0",
          4463 => x"3882b5c8",
          4464 => x"0851ffb0",
          4465 => x"c03f82b5",
          4466 => x"c8085580",
          4467 => x"0b82b5c8",
          4468 => x"0825a938",
          4469 => x"82b5c808",
          4470 => x"ff057017",
          4471 => x"55558074",
          4472 => x"34805374",
          4473 => x"81ff0652",
          4474 => x"7551f8c2",
          4475 => x"3f811b70",
          4476 => x"81ff065c",
          4477 => x"54937b27",
          4478 => x"8338805b",
          4479 => x"74ff2e09",
          4480 => x"8106ff97",
          4481 => x"38863975",
          4482 => x"82b59834",
          4483 => x"768c3882",
          4484 => x"b59c0880",
          4485 => x"2e8438f9",
          4486 => x"d63f8f3d",
          4487 => x"5decc33f",
          4488 => x"82b5c808",
          4489 => x"982b7098",
          4490 => x"2c515978",
          4491 => x"ff2eee38",
          4492 => x"7881ff06",
          4493 => x"82ccf433",
          4494 => x"70982b70",
          4495 => x"982c82cc",
          4496 => x"f0337098",
          4497 => x"2b70972c",
          4498 => x"71982c05",
          4499 => x"70842982",
          4500 => x"aad40570",
          4501 => x"08157033",
          4502 => x"51515151",
          4503 => x"59595159",
          4504 => x"5d588156",
          4505 => x"73782e80",
          4506 => x"e9387774",
          4507 => x"27b43874",
          4508 => x"81800a29",
          4509 => x"81ff0a05",
          4510 => x"70982c51",
          4511 => x"55807524",
          4512 => x"80ce3876",
          4513 => x"53745277",
          4514 => x"51f6853f",
          4515 => x"82b5c808",
          4516 => x"81ff0654",
          4517 => x"73802ed7",
          4518 => x"387482cc",
          4519 => x"f0348156",
          4520 => x"b1397481",
          4521 => x"800a2981",
          4522 => x"800a0570",
          4523 => x"982c7081",
          4524 => x"ff065651",
          4525 => x"55739526",
          4526 => x"97387653",
          4527 => x"74527751",
          4528 => x"f5ce3f82",
          4529 => x"b5c80881",
          4530 => x"ff065473",
          4531 => x"cc38d339",
          4532 => x"80567580",
          4533 => x"2e80ca38",
          4534 => x"811c5574",
          4535 => x"82ccf434",
          4536 => x"74982b70",
          4537 => x"982c82cc",
          4538 => x"f0337098",
          4539 => x"2b70982c",
          4540 => x"70101170",
          4541 => x"822b82aa",
          4542 => x"d811335e",
          4543 => x"51515157",
          4544 => x"58515574",
          4545 => x"772e0981",
          4546 => x"06fe9238",
          4547 => x"82aadc14",
          4548 => x"087d0c80",
          4549 => x"0b82ccf4",
          4550 => x"34800b82",
          4551 => x"ccf03492",
          4552 => x"397582cc",
          4553 => x"f4347582",
          4554 => x"ccf03478",
          4555 => x"af3d3475",
          4556 => x"7d0c7e54",
          4557 => x"739526fd",
          4558 => x"e1387384",
          4559 => x"2982968c",
          4560 => x"05547308",
          4561 => x"0482ccfc",
          4562 => x"3354737e",
          4563 => x"2efdcb38",
          4564 => x"82ccf833",
          4565 => x"55737527",
          4566 => x"ab387498",
          4567 => x"2b70982c",
          4568 => x"51557375",
          4569 => x"249e3874",
          4570 => x"1a547333",
          4571 => x"81153474",
          4572 => x"81800a29",
          4573 => x"81ff0a05",
          4574 => x"70982c82",
          4575 => x"ccfc3356",
          4576 => x"5155df39",
          4577 => x"82ccfc33",
          4578 => x"81115654",
          4579 => x"7482ccfc",
          4580 => x"34731a54",
          4581 => x"ae3d3374",
          4582 => x"3482ccf8",
          4583 => x"3354737e",
          4584 => x"25893881",
          4585 => x"14547382",
          4586 => x"ccf83482",
          4587 => x"ccfc3370",
          4588 => x"81800a29",
          4589 => x"81ff0a05",
          4590 => x"70982c82",
          4591 => x"ccf8335a",
          4592 => x"51565674",
          4593 => x"7725a838",
          4594 => x"82cd9c08",
          4595 => x"52741a70",
          4596 => x"335254ff",
          4597 => x"a3dc3f74",
          4598 => x"81800a29",
          4599 => x"81800a05",
          4600 => x"70982c82",
          4601 => x"ccf83356",
          4602 => x"51557375",
          4603 => x"24da3882",
          4604 => x"ccfc3370",
          4605 => x"982b7098",
          4606 => x"2c82ccf8",
          4607 => x"335a5156",
          4608 => x"56747725",
          4609 => x"fc943882",
          4610 => x"cd9c0852",
          4611 => x"8851ffa3",
          4612 => x"a13f7481",
          4613 => x"800a2981",
          4614 => x"800a0570",
          4615 => x"982c82cc",
          4616 => x"f8335651",
          4617 => x"55737524",
          4618 => x"de38fbee",
          4619 => x"39837a34",
          4620 => x"800b811b",
          4621 => x"3482ccfc",
          4622 => x"53805282",
          4623 => x"9ec851f3",
          4624 => x"9c3f81fd",
          4625 => x"3982ccfc",
          4626 => x"337081ff",
          4627 => x"06555573",
          4628 => x"802efbc6",
          4629 => x"3882ccf8",
          4630 => x"33ff0554",
          4631 => x"7382ccf8",
          4632 => x"34ff1554",
          4633 => x"7382ccfc",
          4634 => x"3482cd9c",
          4635 => x"08528851",
          4636 => x"ffa2bf3f",
          4637 => x"82ccfc33",
          4638 => x"70982b70",
          4639 => x"982c82cc",
          4640 => x"f8335751",
          4641 => x"56577474",
          4642 => x"25ad3874",
          4643 => x"1a548114",
          4644 => x"33743482",
          4645 => x"cd9c0852",
          4646 => x"733351ff",
          4647 => x"a2943f74",
          4648 => x"81800a29",
          4649 => x"81800a05",
          4650 => x"70982c82",
          4651 => x"ccf83358",
          4652 => x"51557575",
          4653 => x"24d53882",
          4654 => x"cd9c0852",
          4655 => x"a051ffa1",
          4656 => x"f13f82cc",
          4657 => x"fc337098",
          4658 => x"2b70982c",
          4659 => x"82ccf833",
          4660 => x"57515657",
          4661 => x"747424fa",
          4662 => x"c13882cd",
          4663 => x"9c085288",
          4664 => x"51ffa1ce",
          4665 => x"3f748180",
          4666 => x"0a298180",
          4667 => x"0a057098",
          4668 => x"2c82ccf8",
          4669 => x"33585155",
          4670 => x"757525de",
          4671 => x"38fa9b39",
          4672 => x"82ccf833",
          4673 => x"7a055480",
          4674 => x"743482cd",
          4675 => x"9c08528a",
          4676 => x"51ffa19e",
          4677 => x"3f82ccf8",
          4678 => x"527951f6",
          4679 => x"c93f82b5",
          4680 => x"c80881ff",
          4681 => x"06547396",
          4682 => x"3882ccf8",
          4683 => x"33547380",
          4684 => x"2e8f3881",
          4685 => x"53735279",
          4686 => x"51f1f33f",
          4687 => x"8439807a",
          4688 => x"34800b82",
          4689 => x"ccfc3480",
          4690 => x"0b82ccf8",
          4691 => x"347982b5",
          4692 => x"c80caf3d",
          4693 => x"0d0482cc",
          4694 => x"fc335473",
          4695 => x"802ef9ba",
          4696 => x"3882cd9c",
          4697 => x"08528851",
          4698 => x"ffa0c73f",
          4699 => x"82ccfc33",
          4700 => x"ff055473",
          4701 => x"82ccfc34",
          4702 => x"7381ff06",
          4703 => x"54dd3982",
          4704 => x"ccfc3382",
          4705 => x"ccf83355",
          4706 => x"5573752e",
          4707 => x"f98c38ff",
          4708 => x"14547382",
          4709 => x"ccf83474",
          4710 => x"982b7098",
          4711 => x"2c7581ff",
          4712 => x"06565155",
          4713 => x"747425ad",
          4714 => x"38741a54",
          4715 => x"81143374",
          4716 => x"3482cd9c",
          4717 => x"08527333",
          4718 => x"51ff9ff6",
          4719 => x"3f748180",
          4720 => x"0a298180",
          4721 => x"0a057098",
          4722 => x"2c82ccf8",
          4723 => x"33585155",
          4724 => x"757524d5",
          4725 => x"3882cd9c",
          4726 => x"0852a051",
          4727 => x"ff9fd33f",
          4728 => x"82ccfc33",
          4729 => x"70982b70",
          4730 => x"982c82cc",
          4731 => x"f8335751",
          4732 => x"56577474",
          4733 => x"24f8a338",
          4734 => x"82cd9c08",
          4735 => x"528851ff",
          4736 => x"9fb03f74",
          4737 => x"81800a29",
          4738 => x"81800a05",
          4739 => x"70982c82",
          4740 => x"ccf83358",
          4741 => x"51557575",
          4742 => x"25de38f7",
          4743 => x"fd3982cc",
          4744 => x"fc337081",
          4745 => x"ff0682cc",
          4746 => x"f8335956",
          4747 => x"54747727",
          4748 => x"f7e83882",
          4749 => x"cd9c0852",
          4750 => x"81145473",
          4751 => x"82ccfc34",
          4752 => x"741a7033",
          4753 => x"5254ff9e",
          4754 => x"e93f82cc",
          4755 => x"fc337081",
          4756 => x"ff0682cc",
          4757 => x"f8335856",
          4758 => x"54757526",
          4759 => x"d638f7ba",
          4760 => x"3982ccfc",
          4761 => x"53805282",
          4762 => x"9ec851ee",
          4763 => x"f03f800b",
          4764 => x"82ccfc34",
          4765 => x"800b82cc",
          4766 => x"f834f79e",
          4767 => x"397ab038",
          4768 => x"82b59408",
          4769 => x"5574802e",
          4770 => x"a6387451",
          4771 => x"ffa6f63f",
          4772 => x"82b5c808",
          4773 => x"82ccf834",
          4774 => x"82b5c808",
          4775 => x"81ff0681",
          4776 => x"05537452",
          4777 => x"7951ffa8",
          4778 => x"bc3f935b",
          4779 => x"81c0397a",
          4780 => x"842982b4",
          4781 => x"c805fc11",
          4782 => x"08565474",
          4783 => x"802ea738",
          4784 => x"7451ffa6",
          4785 => x"c03f82b5",
          4786 => x"c80882cc",
          4787 => x"f83482b5",
          4788 => x"c80881ff",
          4789 => x"06810553",
          4790 => x"74527951",
          4791 => x"ffa8863f",
          4792 => x"ff1b5480",
          4793 => x"fa397308",
          4794 => x"5574802e",
          4795 => x"f6ac3874",
          4796 => x"51ffa691",
          4797 => x"3f99397a",
          4798 => x"932e0981",
          4799 => x"06ae3882",
          4800 => x"b4c80855",
          4801 => x"74802ea4",
          4802 => x"387451ff",
          4803 => x"a5f73f82",
          4804 => x"b5c80882",
          4805 => x"ccf83482",
          4806 => x"b5c80881",
          4807 => x"ff068105",
          4808 => x"53745279",
          4809 => x"51ffa7bd",
          4810 => x"3f80c339",
          4811 => x"7a842982",
          4812 => x"b4cc0570",
          4813 => x"08565474",
          4814 => x"802eab38",
          4815 => x"7451ffa5",
          4816 => x"c43f82b5",
          4817 => x"c80882cc",
          4818 => x"f83482b5",
          4819 => x"c80881ff",
          4820 => x"06810553",
          4821 => x"74527951",
          4822 => x"ffa78a3f",
          4823 => x"811b5473",
          4824 => x"81ff065b",
          4825 => x"89397482",
          4826 => x"ccf83474",
          4827 => x"7a3482cc",
          4828 => x"fc5382cc",
          4829 => x"f8335279",
          4830 => x"51ece23f",
          4831 => x"f59c3982",
          4832 => x"ccfc3370",
          4833 => x"81ff0682",
          4834 => x"ccf83359",
          4835 => x"56547477",
          4836 => x"27f58738",
          4837 => x"82cd9c08",
          4838 => x"52811454",
          4839 => x"7382ccfc",
          4840 => x"34741a70",
          4841 => x"335254ff",
          4842 => x"9c883ff4",
          4843 => x"ed3982cc",
          4844 => x"fc335473",
          4845 => x"802ef4e2",
          4846 => x"3882cd9c",
          4847 => x"08528851",
          4848 => x"ff9bef3f",
          4849 => x"82ccfc33",
          4850 => x"ff055473",
          4851 => x"82ccfc34",
          4852 => x"f4c839f9",
          4853 => x"3d0d83bf",
          4854 => x"f40b82b5",
          4855 => x"c00c8480",
          4856 => x"0b82b5bc",
          4857 => x"23a08053",
          4858 => x"805283bf",
          4859 => x"f451ffaa",
          4860 => x"f53f82b5",
          4861 => x"c0085480",
          4862 => x"58777434",
          4863 => x"81577681",
          4864 => x"153482b5",
          4865 => x"c0085477",
          4866 => x"84153476",
          4867 => x"85153482",
          4868 => x"b5c00854",
          4869 => x"77861534",
          4870 => x"76871534",
          4871 => x"82b5c008",
          4872 => x"82b5bc22",
          4873 => x"ff05fe80",
          4874 => x"80077083",
          4875 => x"ffff0670",
          4876 => x"882a5851",
          4877 => x"55567488",
          4878 => x"17347389",
          4879 => x"173482b5",
          4880 => x"bc227088",
          4881 => x"2982b5c0",
          4882 => x"0805f811",
          4883 => x"51555577",
          4884 => x"82153476",
          4885 => x"83153489",
          4886 => x"3d0d04ff",
          4887 => x"3d0d7352",
          4888 => x"81518472",
          4889 => x"278f38fb",
          4890 => x"12832a82",
          4891 => x"117083ff",
          4892 => x"ff065151",
          4893 => x"517082b5",
          4894 => x"c80c833d",
          4895 => x"0d04f93d",
          4896 => x"0d02a605",
          4897 => x"22028405",
          4898 => x"aa052271",
          4899 => x"0582b5c0",
          4900 => x"0871832b",
          4901 => x"71117483",
          4902 => x"2b731170",
          4903 => x"33811233",
          4904 => x"71882b07",
          4905 => x"02a405ae",
          4906 => x"05227181",
          4907 => x"ffff0607",
          4908 => x"70882a53",
          4909 => x"51525954",
          4910 => x"5b5b5753",
          4911 => x"54557177",
          4912 => x"34708118",
          4913 => x"3482b5c0",
          4914 => x"08147588",
          4915 => x"2a525470",
          4916 => x"82153474",
          4917 => x"83153482",
          4918 => x"b5c00870",
          4919 => x"17703381",
          4920 => x"12337188",
          4921 => x"2b077083",
          4922 => x"2b8ffff8",
          4923 => x"06515256",
          4924 => x"52710573",
          4925 => x"83ffff06",
          4926 => x"70882a54",
          4927 => x"54517182",
          4928 => x"12347281",
          4929 => x"ff065372",
          4930 => x"83123482",
          4931 => x"b5c00816",
          4932 => x"56717634",
          4933 => x"72811734",
          4934 => x"893d0d04",
          4935 => x"fb3d0d82",
          4936 => x"b5c00802",
          4937 => x"84059e05",
          4938 => x"2270832b",
          4939 => x"72118611",
          4940 => x"33871233",
          4941 => x"718b2b71",
          4942 => x"832b0758",
          4943 => x"5b595255",
          4944 => x"52720584",
          4945 => x"12338513",
          4946 => x"3371882b",
          4947 => x"0770882a",
          4948 => x"54565652",
          4949 => x"70841334",
          4950 => x"73851334",
          4951 => x"82b5c008",
          4952 => x"70148411",
          4953 => x"33851233",
          4954 => x"718b2b71",
          4955 => x"832b0756",
          4956 => x"59575272",
          4957 => x"05861233",
          4958 => x"87133371",
          4959 => x"882b0770",
          4960 => x"882a5456",
          4961 => x"56527086",
          4962 => x"13347387",
          4963 => x"133482b5",
          4964 => x"c0081370",
          4965 => x"33811233",
          4966 => x"71882b07",
          4967 => x"7081ffff",
          4968 => x"0670882a",
          4969 => x"53515353",
          4970 => x"53717334",
          4971 => x"70811434",
          4972 => x"873d0d04",
          4973 => x"fa3d0d02",
          4974 => x"a2052282",
          4975 => x"b5c00871",
          4976 => x"832b7111",
          4977 => x"70338112",
          4978 => x"3371882b",
          4979 => x"07708829",
          4980 => x"15703381",
          4981 => x"12337198",
          4982 => x"2b71902b",
          4983 => x"07535f53",
          4984 => x"55525a56",
          4985 => x"57535471",
          4986 => x"802580f6",
          4987 => x"387251fe",
          4988 => x"ab3f82b5",
          4989 => x"c0087016",
          4990 => x"70338112",
          4991 => x"33718b2b",
          4992 => x"71832b07",
          4993 => x"74117033",
          4994 => x"81123371",
          4995 => x"882b0770",
          4996 => x"832b8fff",
          4997 => x"f8065152",
          4998 => x"5451535a",
          4999 => x"58537205",
          5000 => x"74882a54",
          5001 => x"52728213",
          5002 => x"34738313",
          5003 => x"3482b5c0",
          5004 => x"08701670",
          5005 => x"33811233",
          5006 => x"718b2b71",
          5007 => x"832b0756",
          5008 => x"59575572",
          5009 => x"05703381",
          5010 => x"12337188",
          5011 => x"2b077081",
          5012 => x"ffff0670",
          5013 => x"882a5751",
          5014 => x"52585272",
          5015 => x"74347181",
          5016 => x"1534883d",
          5017 => x"0d04fb3d",
          5018 => x"0d82b5c0",
          5019 => x"08028405",
          5020 => x"9e052270",
          5021 => x"832b7211",
          5022 => x"82113383",
          5023 => x"1233718b",
          5024 => x"2b71832b",
          5025 => x"07595b59",
          5026 => x"52565273",
          5027 => x"05713381",
          5028 => x"13337188",
          5029 => x"2b07028c",
          5030 => x"05a20522",
          5031 => x"71077088",
          5032 => x"2a535153",
          5033 => x"53537173",
          5034 => x"34708114",
          5035 => x"3482b5c0",
          5036 => x"08701570",
          5037 => x"33811233",
          5038 => x"718b2b71",
          5039 => x"832b0756",
          5040 => x"59575272",
          5041 => x"05821233",
          5042 => x"83133371",
          5043 => x"882b0770",
          5044 => x"882a5455",
          5045 => x"56527082",
          5046 => x"13347283",
          5047 => x"133482b5",
          5048 => x"c0081482",
          5049 => x"11338312",
          5050 => x"3371882b",
          5051 => x"0782b5c8",
          5052 => x"0c525487",
          5053 => x"3d0d04f7",
          5054 => x"3d0d7b82",
          5055 => x"b5c00831",
          5056 => x"832a7083",
          5057 => x"ffff0670",
          5058 => x"535753fd",
          5059 => x"a73f82b5",
          5060 => x"c0087683",
          5061 => x"2b711182",
          5062 => x"11338312",
          5063 => x"33718b2b",
          5064 => x"71832b07",
          5065 => x"75117033",
          5066 => x"81123371",
          5067 => x"982b7190",
          5068 => x"2b075342",
          5069 => x"4051535b",
          5070 => x"58555954",
          5071 => x"7280258d",
          5072 => x"38828080",
          5073 => x"527551fe",
          5074 => x"9d3f8184",
          5075 => x"39841433",
          5076 => x"85153371",
          5077 => x"8b2b7183",
          5078 => x"2b077611",
          5079 => x"79882a53",
          5080 => x"51555855",
          5081 => x"76861434",
          5082 => x"7581ff06",
          5083 => x"56758714",
          5084 => x"3482b5c0",
          5085 => x"08701984",
          5086 => x"12338513",
          5087 => x"3371882b",
          5088 => x"0770882a",
          5089 => x"54575b56",
          5090 => x"53728416",
          5091 => x"34738516",
          5092 => x"3482b5c0",
          5093 => x"08185380",
          5094 => x"0b861434",
          5095 => x"800b8714",
          5096 => x"3482b5c0",
          5097 => x"08537684",
          5098 => x"14347585",
          5099 => x"143482b5",
          5100 => x"c0081870",
          5101 => x"33811233",
          5102 => x"71882b07",
          5103 => x"70828080",
          5104 => x"0770882a",
          5105 => x"53515556",
          5106 => x"54747434",
          5107 => x"72811534",
          5108 => x"8b3d0d04",
          5109 => x"ff3d0d73",
          5110 => x"5282b5c0",
          5111 => x"088438f7",
          5112 => x"f23f7180",
          5113 => x"2e863871",
          5114 => x"51fe8c3f",
          5115 => x"833d0d04",
          5116 => x"f53d0d80",
          5117 => x"7e5258f8",
          5118 => x"e23f82b5",
          5119 => x"c80883ff",
          5120 => x"ff0682b5",
          5121 => x"c0088411",
          5122 => x"33851233",
          5123 => x"71882b07",
          5124 => x"705f5956",
          5125 => x"585a81ff",
          5126 => x"ff597578",
          5127 => x"2e80cb38",
          5128 => x"75882917",
          5129 => x"70338112",
          5130 => x"3371882b",
          5131 => x"077081ff",
          5132 => x"ff067931",
          5133 => x"7083ffff",
          5134 => x"06707f27",
          5135 => x"52535156",
          5136 => x"59557779",
          5137 => x"278a3873",
          5138 => x"802e8538",
          5139 => x"75785a5b",
          5140 => x"84153385",
          5141 => x"16337188",
          5142 => x"2b075754",
          5143 => x"75c23878",
          5144 => x"81ffff2e",
          5145 => x"85387a79",
          5146 => x"59568076",
          5147 => x"832b82b5",
          5148 => x"c0081170",
          5149 => x"33811233",
          5150 => x"71882b07",
          5151 => x"7081ffff",
          5152 => x"0651525a",
          5153 => x"565c5573",
          5154 => x"752e8338",
          5155 => x"81558054",
          5156 => x"79782681",
          5157 => x"cc387454",
          5158 => x"74802e81",
          5159 => x"c438777a",
          5160 => x"2e098106",
          5161 => x"89387551",
          5162 => x"f8f23f81",
          5163 => x"ac398280",
          5164 => x"80537952",
          5165 => x"7551f7c6",
          5166 => x"3f82b5c0",
          5167 => x"08701c86",
          5168 => x"11338712",
          5169 => x"33718b2b",
          5170 => x"71832b07",
          5171 => x"535a5e55",
          5172 => x"74057a17",
          5173 => x"7083ffff",
          5174 => x"0670882a",
          5175 => x"5c595654",
          5176 => x"78841534",
          5177 => x"7681ff06",
          5178 => x"57768515",
          5179 => x"3482b5c0",
          5180 => x"0875832b",
          5181 => x"7111721e",
          5182 => x"86113387",
          5183 => x"12337188",
          5184 => x"2b077088",
          5185 => x"2a535b5e",
          5186 => x"535a5654",
          5187 => x"73861934",
          5188 => x"75871934",
          5189 => x"82b5c008",
          5190 => x"701c8411",
          5191 => x"33851233",
          5192 => x"718b2b71",
          5193 => x"832b0753",
          5194 => x"5d5a5574",
          5195 => x"05547886",
          5196 => x"15347687",
          5197 => x"153482b5",
          5198 => x"c0087016",
          5199 => x"711d8411",
          5200 => x"33851233",
          5201 => x"71882b07",
          5202 => x"70882a53",
          5203 => x"5a5f5256",
          5204 => x"54738416",
          5205 => x"34758516",
          5206 => x"3482b5c0",
          5207 => x"081b8405",
          5208 => x"547382b5",
          5209 => x"c80c8d3d",
          5210 => x"0d04fe3d",
          5211 => x"0d745282",
          5212 => x"b5c00884",
          5213 => x"38f4dc3f",
          5214 => x"71537180",
          5215 => x"2e8b3871",
          5216 => x"51fced3f",
          5217 => x"82b5c808",
          5218 => x"537282b5",
          5219 => x"c80c843d",
          5220 => x"0d04ee3d",
          5221 => x"0d646640",
          5222 => x"5c807042",
          5223 => x"4082b5c0",
          5224 => x"08602e09",
          5225 => x"81068438",
          5226 => x"f4a93f7b",
          5227 => x"8e387e51",
          5228 => x"ffb83f82",
          5229 => x"b5c80854",
          5230 => x"83c7397e",
          5231 => x"8b387b51",
          5232 => x"fc923f7e",
          5233 => x"5483ba39",
          5234 => x"7e51f58f",
          5235 => x"3f82b5c8",
          5236 => x"0883ffff",
          5237 => x"0682b5c0",
          5238 => x"087d7131",
          5239 => x"832a7083",
          5240 => x"ffff0670",
          5241 => x"832b7311",
          5242 => x"70338112",
          5243 => x"3371882b",
          5244 => x"07707531",
          5245 => x"7083ffff",
          5246 => x"06708829",
          5247 => x"fc057388",
          5248 => x"291a7033",
          5249 => x"81123371",
          5250 => x"882b0770",
          5251 => x"902b5344",
          5252 => x"4e534841",
          5253 => x"525c545b",
          5254 => x"415c565b",
          5255 => x"5b738025",
          5256 => x"8f387681",
          5257 => x"ffff0675",
          5258 => x"317083ff",
          5259 => x"ff064254",
          5260 => x"82163383",
          5261 => x"17337188",
          5262 => x"2b077088",
          5263 => x"291c7033",
          5264 => x"81123371",
          5265 => x"982b7190",
          5266 => x"2b075347",
          5267 => x"45525654",
          5268 => x"7380258b",
          5269 => x"38787531",
          5270 => x"7083ffff",
          5271 => x"06415477",
          5272 => x"7b2781fe",
          5273 => x"38601854",
          5274 => x"737b2e09",
          5275 => x"81068f38",
          5276 => x"7851f6c0",
          5277 => x"3f7a83ff",
          5278 => x"ff065881",
          5279 => x"e5397f8e",
          5280 => x"387a7424",
          5281 => x"89387851",
          5282 => x"f6aa3f81",
          5283 => x"a5397f18",
          5284 => x"557a7524",
          5285 => x"80c83879",
          5286 => x"1d821133",
          5287 => x"83123371",
          5288 => x"882b0753",
          5289 => x"5754f4f4",
          5290 => x"3f805278",
          5291 => x"51f7b73f",
          5292 => x"82b5c808",
          5293 => x"83ffff06",
          5294 => x"7e547c53",
          5295 => x"70832b82",
          5296 => x"b5c00811",
          5297 => x"84055355",
          5298 => x"59ff93cf",
          5299 => x"3f82b5c0",
          5300 => x"08148405",
          5301 => x"7583ffff",
          5302 => x"06595c81",
          5303 => x"85396015",
          5304 => x"547a7424",
          5305 => x"80d43878",
          5306 => x"51f5c93f",
          5307 => x"82b5c008",
          5308 => x"1d821133",
          5309 => x"83123371",
          5310 => x"882b0753",
          5311 => x"4354f49c",
          5312 => x"3f805278",
          5313 => x"51f6df3f",
          5314 => x"82b5c808",
          5315 => x"83ffff06",
          5316 => x"7e547c53",
          5317 => x"70832b82",
          5318 => x"b5c00811",
          5319 => x"84055355",
          5320 => x"59ff92f7",
          5321 => x"3f82b5c0",
          5322 => x"08148405",
          5323 => x"60620519",
          5324 => x"555c7383",
          5325 => x"ffff0658",
          5326 => x"a9397b7f",
          5327 => x"5254f9b0",
          5328 => x"3f82b5c8",
          5329 => x"085c82b5",
          5330 => x"c808802e",
          5331 => x"93387d53",
          5332 => x"735282b5",
          5333 => x"c80851ff",
          5334 => x"978b3f73",
          5335 => x"51f7983f",
          5336 => x"7a587a78",
          5337 => x"27993880",
          5338 => x"537a5278",
          5339 => x"51f28f3f",
          5340 => x"7a19832b",
          5341 => x"82b5c008",
          5342 => x"05840551",
          5343 => x"f6f93f7b",
          5344 => x"547382b5",
          5345 => x"c80c943d",
          5346 => x"0d04fc3d",
          5347 => x"0d777729",
          5348 => x"705254fb",
          5349 => x"d53f82b5",
          5350 => x"c8085582",
          5351 => x"b5c80880",
          5352 => x"2e8e3873",
          5353 => x"53805282",
          5354 => x"b5c80851",
          5355 => x"ff9bb73f",
          5356 => x"7482b5c8",
          5357 => x"0c863d0d",
          5358 => x"04ff3d0d",
          5359 => x"028f0533",
          5360 => x"51815270",
          5361 => x"72268738",
          5362 => x"82b5c411",
          5363 => x"33527182",
          5364 => x"b5c80c83",
          5365 => x"3d0d04fc",
          5366 => x"3d0d029b",
          5367 => x"05330284",
          5368 => x"059f0533",
          5369 => x"56538351",
          5370 => x"72812680",
          5371 => x"e0387284",
          5372 => x"2b87c092",
          5373 => x"8c115351",
          5374 => x"88547480",
          5375 => x"2e843881",
          5376 => x"88547372",
          5377 => x"0c87c092",
          5378 => x"8c115181",
          5379 => x"710c850b",
          5380 => x"87c0988c",
          5381 => x"0c705271",
          5382 => x"08708206",
          5383 => x"51517080",
          5384 => x"2e8a3887",
          5385 => x"c0988c08",
          5386 => x"5170ec38",
          5387 => x"7108fc80",
          5388 => x"80065271",
          5389 => x"923887c0",
          5390 => x"988c0851",
          5391 => x"70802e87",
          5392 => x"387182b5",
          5393 => x"c4143482",
          5394 => x"b5c41333",
          5395 => x"517082b5",
          5396 => x"c80c863d",
          5397 => x"0d04f33d",
          5398 => x"0d606264",
          5399 => x"028c05bf",
          5400 => x"05335740",
          5401 => x"585b8374",
          5402 => x"525afecd",
          5403 => x"3f82b5c8",
          5404 => x"0881067a",
          5405 => x"54527181",
          5406 => x"be387172",
          5407 => x"75842b87",
          5408 => x"c0928011",
          5409 => x"87c0928c",
          5410 => x"1287c092",
          5411 => x"8413415a",
          5412 => x"40575a58",
          5413 => x"850b87c0",
          5414 => x"988c0c76",
          5415 => x"7d0c8476",
          5416 => x"0c750870",
          5417 => x"852a7081",
          5418 => x"06515354",
          5419 => x"71802e8e",
          5420 => x"387b0852",
          5421 => x"717b7081",
          5422 => x"055d3481",
          5423 => x"19598074",
          5424 => x"a2065353",
          5425 => x"71732e83",
          5426 => x"38815378",
          5427 => x"83ff268f",
          5428 => x"3872802e",
          5429 => x"8a3887c0",
          5430 => x"988c0852",
          5431 => x"71c33887",
          5432 => x"c0988c08",
          5433 => x"5271802e",
          5434 => x"87387884",
          5435 => x"802e9938",
          5436 => x"81760c87",
          5437 => x"c0928c15",
          5438 => x"53720870",
          5439 => x"82065152",
          5440 => x"71f738ff",
          5441 => x"1a5a8d39",
          5442 => x"84801781",
          5443 => x"197081ff",
          5444 => x"065a5357",
          5445 => x"79802e90",
          5446 => x"3873fc80",
          5447 => x"80065271",
          5448 => x"87387d78",
          5449 => x"26feed38",
          5450 => x"73fc8080",
          5451 => x"06527180",
          5452 => x"2e833881",
          5453 => x"52715372",
          5454 => x"82b5c80c",
          5455 => x"8f3d0d04",
          5456 => x"f33d0d60",
          5457 => x"6264028c",
          5458 => x"05bf0533",
          5459 => x"5740585b",
          5460 => x"83598074",
          5461 => x"5258fce1",
          5462 => x"3f82b5c8",
          5463 => x"08810679",
          5464 => x"54527178",
          5465 => x"2e098106",
          5466 => x"81b13877",
          5467 => x"74842b87",
          5468 => x"c0928011",
          5469 => x"87c0928c",
          5470 => x"1287c092",
          5471 => x"84134059",
          5472 => x"5f565a85",
          5473 => x"0b87c098",
          5474 => x"8c0c767d",
          5475 => x"0c82760c",
          5476 => x"80587508",
          5477 => x"70842a70",
          5478 => x"81065153",
          5479 => x"5471802e",
          5480 => x"8c387a70",
          5481 => x"81055c33",
          5482 => x"7c0c8118",
          5483 => x"5873812a",
          5484 => x"70810651",
          5485 => x"5271802e",
          5486 => x"8a3887c0",
          5487 => x"988c0852",
          5488 => x"71d03887",
          5489 => x"c0988c08",
          5490 => x"5271802e",
          5491 => x"87387784",
          5492 => x"802e9938",
          5493 => x"81760c87",
          5494 => x"c0928c15",
          5495 => x"53720870",
          5496 => x"82065152",
          5497 => x"71f738ff",
          5498 => x"19598d39",
          5499 => x"811a7081",
          5500 => x"ff068480",
          5501 => x"19595b52",
          5502 => x"78802e90",
          5503 => x"3873fc80",
          5504 => x"80065271",
          5505 => x"87387d7a",
          5506 => x"26fef838",
          5507 => x"73fc8080",
          5508 => x"06527180",
          5509 => x"2e833881",
          5510 => x"52715372",
          5511 => x"82b5c80c",
          5512 => x"8f3d0d04",
          5513 => x"fa3d0d7a",
          5514 => x"028405a3",
          5515 => x"05330288",
          5516 => x"05a70533",
          5517 => x"71545456",
          5518 => x"57fafe3f",
          5519 => x"82b5c808",
          5520 => x"81065383",
          5521 => x"547280fe",
          5522 => x"38850b87",
          5523 => x"c0988c0c",
          5524 => x"81567176",
          5525 => x"2e80dc38",
          5526 => x"71762493",
          5527 => x"3874842b",
          5528 => x"87c0928c",
          5529 => x"11545471",
          5530 => x"802e8d38",
          5531 => x"80d43971",
          5532 => x"832e80c6",
          5533 => x"3880cb39",
          5534 => x"72087081",
          5535 => x"2a708106",
          5536 => x"51515271",
          5537 => x"802e8a38",
          5538 => x"87c0988c",
          5539 => x"085271e8",
          5540 => x"3887c098",
          5541 => x"8c085271",
          5542 => x"96388173",
          5543 => x"0c87c092",
          5544 => x"8c145372",
          5545 => x"08708206",
          5546 => x"515271f7",
          5547 => x"38963980",
          5548 => x"56923988",
          5549 => x"800a770c",
          5550 => x"85398180",
          5551 => x"770c7256",
          5552 => x"83398456",
          5553 => x"75547382",
          5554 => x"b5c80c88",
          5555 => x"3d0d04fe",
          5556 => x"3d0d7481",
          5557 => x"11337133",
          5558 => x"71882b07",
          5559 => x"82b5c80c",
          5560 => x"5351843d",
          5561 => x"0d04fd3d",
          5562 => x"0d758311",
          5563 => x"33821233",
          5564 => x"71902b71",
          5565 => x"882b0781",
          5566 => x"14337072",
          5567 => x"07882b75",
          5568 => x"33710782",
          5569 => x"b5c80c52",
          5570 => x"53545654",
          5571 => x"52853d0d",
          5572 => x"04ff3d0d",
          5573 => x"73028405",
          5574 => x"92052252",
          5575 => x"52707270",
          5576 => x"81055434",
          5577 => x"70882a51",
          5578 => x"70723483",
          5579 => x"3d0d04ff",
          5580 => x"3d0d7375",
          5581 => x"52527072",
          5582 => x"70810554",
          5583 => x"3470882a",
          5584 => x"51707270",
          5585 => x"81055434",
          5586 => x"70882a51",
          5587 => x"70727081",
          5588 => x"05543470",
          5589 => x"882a5170",
          5590 => x"7234833d",
          5591 => x"0d04fe3d",
          5592 => x"0d767577",
          5593 => x"54545170",
          5594 => x"802e9238",
          5595 => x"71708105",
          5596 => x"53337370",
          5597 => x"81055534",
          5598 => x"ff1151eb",
          5599 => x"39843d0d",
          5600 => x"04fe3d0d",
          5601 => x"75777654",
          5602 => x"52537272",
          5603 => x"70810554",
          5604 => x"34ff1151",
          5605 => x"70f43884",
          5606 => x"3d0d04fc",
          5607 => x"3d0d7877",
          5608 => x"79565653",
          5609 => x"74708105",
          5610 => x"56337470",
          5611 => x"81055633",
          5612 => x"717131ff",
          5613 => x"16565252",
          5614 => x"5272802e",
          5615 => x"86387180",
          5616 => x"2ee23871",
          5617 => x"82b5c80c",
          5618 => x"863d0d04",
          5619 => x"fe3d0d74",
          5620 => x"76545189",
          5621 => x"3971732e",
          5622 => x"8a388111",
          5623 => x"51703352",
          5624 => x"71f33870",
          5625 => x"3382b5c8",
          5626 => x"0c843d0d",
          5627 => x"04800b82",
          5628 => x"b5c80c04",
          5629 => x"800b82b5",
          5630 => x"c80c04f7",
          5631 => x"3d0d7b56",
          5632 => x"800b8317",
          5633 => x"33565a74",
          5634 => x"7a2e80d6",
          5635 => x"388154b0",
          5636 => x"160853b4",
          5637 => x"16705381",
          5638 => x"17335259",
          5639 => x"faa23f82",
          5640 => x"b5c8087a",
          5641 => x"2e098106",
          5642 => x"b73882b5",
          5643 => x"c8088317",
          5644 => x"34b01608",
          5645 => x"70a41808",
          5646 => x"319c1808",
          5647 => x"59565874",
          5648 => x"77279f38",
          5649 => x"82163355",
          5650 => x"74822e09",
          5651 => x"81069338",
          5652 => x"81547618",
          5653 => x"53785281",
          5654 => x"163351f9",
          5655 => x"e33f8339",
          5656 => x"815a7982",
          5657 => x"b5c80c8b",
          5658 => x"3d0d04fa",
          5659 => x"3d0d787a",
          5660 => x"56568057",
          5661 => x"74b01708",
          5662 => x"2eaf3875",
          5663 => x"51fefc3f",
          5664 => x"82b5c808",
          5665 => x"5782b5c8",
          5666 => x"089f3881",
          5667 => x"547453b4",
          5668 => x"16528116",
          5669 => x"3351f7be",
          5670 => x"3f82b5c8",
          5671 => x"08802e85",
          5672 => x"38ff5581",
          5673 => x"5774b017",
          5674 => x"0c7682b5",
          5675 => x"c80c883d",
          5676 => x"0d04f83d",
          5677 => x"0d7a7052",
          5678 => x"57fec03f",
          5679 => x"82b5c808",
          5680 => x"5882b5c8",
          5681 => x"08819138",
          5682 => x"76335574",
          5683 => x"832e0981",
          5684 => x"0680f038",
          5685 => x"84173359",
          5686 => x"78812e09",
          5687 => x"810680e3",
          5688 => x"38848053",
          5689 => x"82b5c808",
          5690 => x"52b41770",
          5691 => x"5256fd91",
          5692 => x"3f82d4d5",
          5693 => x"5284b217",
          5694 => x"51fc963f",
          5695 => x"848b85a4",
          5696 => x"d2527551",
          5697 => x"fca93f86",
          5698 => x"8a85e4f2",
          5699 => x"52849817",
          5700 => x"51fc9c3f",
          5701 => x"90170852",
          5702 => x"849c1751",
          5703 => x"fc913f8c",
          5704 => x"17085284",
          5705 => x"a01751fc",
          5706 => x"863fa017",
          5707 => x"08810570",
          5708 => x"b0190c79",
          5709 => x"55537552",
          5710 => x"81173351",
          5711 => x"f8823f77",
          5712 => x"84183480",
          5713 => x"53805281",
          5714 => x"173351f9",
          5715 => x"d73f82b5",
          5716 => x"c808802e",
          5717 => x"83388158",
          5718 => x"7782b5c8",
          5719 => x"0c8a3d0d",
          5720 => x"04fb3d0d",
          5721 => x"77fe1a98",
          5722 => x"1208fe05",
          5723 => x"55565480",
          5724 => x"56747327",
          5725 => x"8d388a14",
          5726 => x"22757129",
          5727 => x"ac160805",
          5728 => x"57537582",
          5729 => x"b5c80c87",
          5730 => x"3d0d04f9",
          5731 => x"3d0d7a7a",
          5732 => x"70085654",
          5733 => x"57817727",
          5734 => x"81df3876",
          5735 => x"98150827",
          5736 => x"81d738ff",
          5737 => x"74335458",
          5738 => x"72822e80",
          5739 => x"f5387282",
          5740 => x"24893872",
          5741 => x"812e8d38",
          5742 => x"81bf3972",
          5743 => x"832e818e",
          5744 => x"3881b639",
          5745 => x"76812a17",
          5746 => x"70892aa4",
          5747 => x"16080553",
          5748 => x"745255fd",
          5749 => x"963f82b5",
          5750 => x"c808819f",
          5751 => x"387483ff",
          5752 => x"0614b411",
          5753 => x"33811770",
          5754 => x"892aa418",
          5755 => x"08055576",
          5756 => x"54575753",
          5757 => x"fcf53f82",
          5758 => x"b5c80880",
          5759 => x"fe387483",
          5760 => x"ff0614b4",
          5761 => x"11337088",
          5762 => x"2b780779",
          5763 => x"81067184",
          5764 => x"2a5c5258",
          5765 => x"51537280",
          5766 => x"e238759f",
          5767 => x"ff065880",
          5768 => x"da397688",
          5769 => x"2aa41508",
          5770 => x"05527351",
          5771 => x"fcbd3f82",
          5772 => x"b5c80880",
          5773 => x"c6387610",
          5774 => x"83fe0674",
          5775 => x"05b40551",
          5776 => x"f98d3f82",
          5777 => x"b5c80883",
          5778 => x"ffff0658",
          5779 => x"ae397687",
          5780 => x"2aa41508",
          5781 => x"05527351",
          5782 => x"fc913f82",
          5783 => x"b5c8089b",
          5784 => x"3876822b",
          5785 => x"83fc0674",
          5786 => x"05b40551",
          5787 => x"f8f83f82",
          5788 => x"b5c808f0",
          5789 => x"0a065883",
          5790 => x"39815877",
          5791 => x"82b5c80c",
          5792 => x"893d0d04",
          5793 => x"f83d0d7a",
          5794 => x"7c7e5a58",
          5795 => x"56825981",
          5796 => x"7727829e",
          5797 => x"38769817",
          5798 => x"08278296",
          5799 => x"38753353",
          5800 => x"72792e81",
          5801 => x"9d387279",
          5802 => x"24893872",
          5803 => x"812e8d38",
          5804 => x"82803972",
          5805 => x"832e81b8",
          5806 => x"3881f739",
          5807 => x"76812a17",
          5808 => x"70892aa4",
          5809 => x"18080553",
          5810 => x"765255fb",
          5811 => x"9e3f82b5",
          5812 => x"c8085982",
          5813 => x"b5c80881",
          5814 => x"d9387483",
          5815 => x"ff0616b4",
          5816 => x"05811678",
          5817 => x"81065956",
          5818 => x"54775376",
          5819 => x"802e8f38",
          5820 => x"77842b9f",
          5821 => x"f0067433",
          5822 => x"8f067107",
          5823 => x"51537274",
          5824 => x"34810b83",
          5825 => x"17347489",
          5826 => x"2aa41708",
          5827 => x"05527551",
          5828 => x"fad93f82",
          5829 => x"b5c80859",
          5830 => x"82b5c808",
          5831 => x"81943874",
          5832 => x"83ff0616",
          5833 => x"b4057884",
          5834 => x"2a545476",
          5835 => x"8f387788",
          5836 => x"2a743381",
          5837 => x"f006718f",
          5838 => x"06075153",
          5839 => x"72743480",
          5840 => x"ec397688",
          5841 => x"2aa41708",
          5842 => x"05527551",
          5843 => x"fa9d3f82",
          5844 => x"b5c80859",
          5845 => x"82b5c808",
          5846 => x"80d83877",
          5847 => x"83ffff06",
          5848 => x"52761083",
          5849 => x"fe067605",
          5850 => x"b40551f7",
          5851 => x"a43fbe39",
          5852 => x"76872aa4",
          5853 => x"17080552",
          5854 => x"7551f9ef",
          5855 => x"3f82b5c8",
          5856 => x"085982b5",
          5857 => x"c808ab38",
          5858 => x"77f00a06",
          5859 => x"77822b83",
          5860 => x"fc067018",
          5861 => x"b4057054",
          5862 => x"515454f6",
          5863 => x"c93f82b5",
          5864 => x"c8088f0a",
          5865 => x"06740752",
          5866 => x"7251f783",
          5867 => x"3f810b83",
          5868 => x"17347882",
          5869 => x"b5c80c8a",
          5870 => x"3d0d04f8",
          5871 => x"3d0d7a7c",
          5872 => x"7e720859",
          5873 => x"56565981",
          5874 => x"7527a438",
          5875 => x"74981708",
          5876 => x"279d3873",
          5877 => x"802eaa38",
          5878 => x"ff537352",
          5879 => x"7551fda4",
          5880 => x"3f82b5c8",
          5881 => x"085482b5",
          5882 => x"c80880f2",
          5883 => x"38933982",
          5884 => x"5480eb39",
          5885 => x"815480e6",
          5886 => x"3982b5c8",
          5887 => x"085480de",
          5888 => x"39745278",
          5889 => x"51fb843f",
          5890 => x"82b5c808",
          5891 => x"5882b5c8",
          5892 => x"08802e80",
          5893 => x"c73882b5",
          5894 => x"c808812e",
          5895 => x"d23882b5",
          5896 => x"c808ff2e",
          5897 => x"cf388053",
          5898 => x"74527551",
          5899 => x"fcd63f82",
          5900 => x"b5c808c5",
          5901 => x"38981608",
          5902 => x"fe119018",
          5903 => x"08575557",
          5904 => x"74742790",
          5905 => x"38811590",
          5906 => x"170c8416",
          5907 => x"33810754",
          5908 => x"73841734",
          5909 => x"77557678",
          5910 => x"26ffa638",
          5911 => x"80547382",
          5912 => x"b5c80c8a",
          5913 => x"3d0d04f6",
          5914 => x"3d0d7c7e",
          5915 => x"7108595b",
          5916 => x"5b799538",
          5917 => x"8c170858",
          5918 => x"77802e88",
          5919 => x"38981708",
          5920 => x"7826b238",
          5921 => x"8158ae39",
          5922 => x"79527a51",
          5923 => x"f9fd3f81",
          5924 => x"557482b5",
          5925 => x"c8082782",
          5926 => x"e03882b5",
          5927 => x"c8085582",
          5928 => x"b5c808ff",
          5929 => x"2e82d238",
          5930 => x"98170882",
          5931 => x"b5c80826",
          5932 => x"82c73879",
          5933 => x"58901708",
          5934 => x"70565473",
          5935 => x"802e82b9",
          5936 => x"38777a2e",
          5937 => x"09810680",
          5938 => x"e238811a",
          5939 => x"56981708",
          5940 => x"76268338",
          5941 => x"82567552",
          5942 => x"7a51f9af",
          5943 => x"3f805982",
          5944 => x"b5c80881",
          5945 => x"2e098106",
          5946 => x"863882b5",
          5947 => x"c8085982",
          5948 => x"b5c80809",
          5949 => x"70307072",
          5950 => x"07802570",
          5951 => x"7c0782b5",
          5952 => x"c8085451",
          5953 => x"51555573",
          5954 => x"81ef3882",
          5955 => x"b5c80880",
          5956 => x"2e95388c",
          5957 => x"17085481",
          5958 => x"74279038",
          5959 => x"73981808",
          5960 => x"27893873",
          5961 => x"58853975",
          5962 => x"80db3877",
          5963 => x"56811656",
          5964 => x"98170876",
          5965 => x"26893882",
          5966 => x"56757826",
          5967 => x"81ac3875",
          5968 => x"527a51f8",
          5969 => x"c63f82b5",
          5970 => x"c808802e",
          5971 => x"b8388059",
          5972 => x"82b5c808",
          5973 => x"812e0981",
          5974 => x"06863882",
          5975 => x"b5c80859",
          5976 => x"82b5c808",
          5977 => x"09703070",
          5978 => x"72078025",
          5979 => x"707c0751",
          5980 => x"51555573",
          5981 => x"80f83875",
          5982 => x"782e0981",
          5983 => x"06ffae38",
          5984 => x"735580f5",
          5985 => x"39ff5375",
          5986 => x"527651f9",
          5987 => x"f73f82b5",
          5988 => x"c80882b5",
          5989 => x"c8083070",
          5990 => x"82b5c808",
          5991 => x"07802551",
          5992 => x"55557980",
          5993 => x"2e943873",
          5994 => x"802e8f38",
          5995 => x"75537952",
          5996 => x"7651f9d0",
          5997 => x"3f82b5c8",
          5998 => x"085574a5",
          5999 => x"38758c18",
          6000 => x"0c981708",
          6001 => x"fe059018",
          6002 => x"08565474",
          6003 => x"74268638",
          6004 => x"ff159018",
          6005 => x"0c841733",
          6006 => x"81075473",
          6007 => x"84183497",
          6008 => x"39ff5674",
          6009 => x"812e9038",
          6010 => x"8c398055",
          6011 => x"8c3982b5",
          6012 => x"c8085585",
          6013 => x"39815675",
          6014 => x"557482b5",
          6015 => x"c80c8c3d",
          6016 => x"0d04f83d",
          6017 => x"0d7a7052",
          6018 => x"55f3f03f",
          6019 => x"82b5c808",
          6020 => x"58815682",
          6021 => x"b5c80880",
          6022 => x"d8387b52",
          6023 => x"7451f6c1",
          6024 => x"3f82b5c8",
          6025 => x"0882b5c8",
          6026 => x"08b0170c",
          6027 => x"59848053",
          6028 => x"7752b415",
          6029 => x"705257f2",
          6030 => x"c83f7756",
          6031 => x"84398116",
          6032 => x"568a1522",
          6033 => x"58757827",
          6034 => x"97388154",
          6035 => x"75195376",
          6036 => x"52811533",
          6037 => x"51ede93f",
          6038 => x"82b5c808",
          6039 => x"802edf38",
          6040 => x"8a152276",
          6041 => x"32703070",
          6042 => x"7207709f",
          6043 => x"2a535156",
          6044 => x"567582b5",
          6045 => x"c80c8a3d",
          6046 => x"0d04f83d",
          6047 => x"0d7a7c71",
          6048 => x"08585657",
          6049 => x"74f0800a",
          6050 => x"2680f138",
          6051 => x"749f0653",
          6052 => x"7280e938",
          6053 => x"7490180c",
          6054 => x"88170854",
          6055 => x"73aa3875",
          6056 => x"33538273",
          6057 => x"278838a8",
          6058 => x"16085473",
          6059 => x"9b387485",
          6060 => x"2a53820b",
          6061 => x"8817225a",
          6062 => x"58727927",
          6063 => x"80fe38a8",
          6064 => x"16089818",
          6065 => x"0c80cd39",
          6066 => x"8a162270",
          6067 => x"892b5458",
          6068 => x"727526b2",
          6069 => x"38735276",
          6070 => x"51f5b03f",
          6071 => x"82b5c808",
          6072 => x"5482b5c8",
          6073 => x"08ff2ebd",
          6074 => x"38810b82",
          6075 => x"b5c80827",
          6076 => x"8b389816",
          6077 => x"0882b5c8",
          6078 => x"08268538",
          6079 => x"8258bd39",
          6080 => x"74733155",
          6081 => x"cb397352",
          6082 => x"7551f4d5",
          6083 => x"3f82b5c8",
          6084 => x"0898180c",
          6085 => x"7394180c",
          6086 => x"98170853",
          6087 => x"82587280",
          6088 => x"2e9a3885",
          6089 => x"39815894",
          6090 => x"3974892a",
          6091 => x"1398180c",
          6092 => x"7483ff06",
          6093 => x"16b4059c",
          6094 => x"180c8058",
          6095 => x"7782b5c8",
          6096 => x"0c8a3d0d",
          6097 => x"04f83d0d",
          6098 => x"7a700890",
          6099 => x"1208a005",
          6100 => x"595754f0",
          6101 => x"800a7727",
          6102 => x"8638800b",
          6103 => x"98150c98",
          6104 => x"14085384",
          6105 => x"5572802e",
          6106 => x"81cb3876",
          6107 => x"83ff0658",
          6108 => x"7781b538",
          6109 => x"81139815",
          6110 => x"0c941408",
          6111 => x"55749238",
          6112 => x"76852a88",
          6113 => x"17225653",
          6114 => x"74732681",
          6115 => x"9b3880c0",
          6116 => x"398a1622",
          6117 => x"ff057789",
          6118 => x"2a065372",
          6119 => x"818a3874",
          6120 => x"527351f3",
          6121 => x"e63f82b5",
          6122 => x"c8085382",
          6123 => x"55810b82",
          6124 => x"b5c80827",
          6125 => x"80ff3881",
          6126 => x"5582b5c8",
          6127 => x"08ff2e80",
          6128 => x"f4389816",
          6129 => x"0882b5c8",
          6130 => x"082680ca",
          6131 => x"387b8a38",
          6132 => x"7798150c",
          6133 => x"845580dd",
          6134 => x"39941408",
          6135 => x"527351f9",
          6136 => x"863f82b5",
          6137 => x"c8085387",
          6138 => x"5582b5c8",
          6139 => x"08802e80",
          6140 => x"c4388255",
          6141 => x"82b5c808",
          6142 => x"812eba38",
          6143 => x"815582b5",
          6144 => x"c808ff2e",
          6145 => x"b03882b5",
          6146 => x"c8085275",
          6147 => x"51fbf33f",
          6148 => x"82b5c808",
          6149 => x"a0387294",
          6150 => x"150c7252",
          6151 => x"7551f2c1",
          6152 => x"3f82b5c8",
          6153 => x"0898150c",
          6154 => x"7690150c",
          6155 => x"7716b405",
          6156 => x"9c150c80",
          6157 => x"557482b5",
          6158 => x"c80c8a3d",
          6159 => x"0d04f73d",
          6160 => x"0d7b7d71",
          6161 => x"085b5b57",
          6162 => x"80527651",
          6163 => x"fcac3f82",
          6164 => x"b5c80854",
          6165 => x"82b5c808",
          6166 => x"80ec3882",
          6167 => x"b5c80856",
          6168 => x"98170852",
          6169 => x"7851f083",
          6170 => x"3f82b5c8",
          6171 => x"085482b5",
          6172 => x"c80880d2",
          6173 => x"3882b5c8",
          6174 => x"089c1808",
          6175 => x"70335154",
          6176 => x"587281e5",
          6177 => x"2e098106",
          6178 => x"83388158",
          6179 => x"82b5c808",
          6180 => x"55728338",
          6181 => x"81557775",
          6182 => x"07537280",
          6183 => x"2e8e3881",
          6184 => x"1656757a",
          6185 => x"2e098106",
          6186 => x"8838a539",
          6187 => x"82b5c808",
          6188 => x"56815276",
          6189 => x"51fd8e3f",
          6190 => x"82b5c808",
          6191 => x"5482b5c8",
          6192 => x"08802eff",
          6193 => x"9b387384",
          6194 => x"2e098106",
          6195 => x"83388754",
          6196 => x"7382b5c8",
          6197 => x"0c8b3d0d",
          6198 => x"04fd3d0d",
          6199 => x"769a1152",
          6200 => x"54ebec3f",
          6201 => x"82b5c808",
          6202 => x"83ffff06",
          6203 => x"76703351",
          6204 => x"53537183",
          6205 => x"2e098106",
          6206 => x"90389414",
          6207 => x"51ebd03f",
          6208 => x"82b5c808",
          6209 => x"902b7307",
          6210 => x"537282b5",
          6211 => x"c80c853d",
          6212 => x"0d04fc3d",
          6213 => x"0d777970",
          6214 => x"83ffff06",
          6215 => x"549a1253",
          6216 => x"5555ebed",
          6217 => x"3f767033",
          6218 => x"51537283",
          6219 => x"2e098106",
          6220 => x"8b387390",
          6221 => x"2a529415",
          6222 => x"51ebd63f",
          6223 => x"863d0d04",
          6224 => x"f73d0d7b",
          6225 => x"7d5b5584",
          6226 => x"75085a58",
          6227 => x"98150880",
          6228 => x"2e818a38",
          6229 => x"98150852",
          6230 => x"7851ee8f",
          6231 => x"3f82b5c8",
          6232 => x"085882b5",
          6233 => x"c80880f5",
          6234 => x"389c1508",
          6235 => x"70335553",
          6236 => x"73863884",
          6237 => x"5880e639",
          6238 => x"8b133370",
          6239 => x"bf067081",
          6240 => x"ff065851",
          6241 => x"53728616",
          6242 => x"3482b5c8",
          6243 => x"08537381",
          6244 => x"e52e8338",
          6245 => x"815373ae",
          6246 => x"2ea93881",
          6247 => x"70740654",
          6248 => x"5772802e",
          6249 => x"9e38758f",
          6250 => x"2e993882",
          6251 => x"b5c80876",
          6252 => x"df065454",
          6253 => x"72882e09",
          6254 => x"81068338",
          6255 => x"7654737a",
          6256 => x"2ea03880",
          6257 => x"527451fa",
          6258 => x"fc3f82b5",
          6259 => x"c8085882",
          6260 => x"b5c80889",
          6261 => x"38981508",
          6262 => x"fefa3886",
          6263 => x"39800b98",
          6264 => x"160c7782",
          6265 => x"b5c80c8b",
          6266 => x"3d0d04fb",
          6267 => x"3d0d7770",
          6268 => x"08575481",
          6269 => x"527351fc",
          6270 => x"c53f82b5",
          6271 => x"c8085582",
          6272 => x"b5c808b4",
          6273 => x"38981408",
          6274 => x"527551ec",
          6275 => x"de3f82b5",
          6276 => x"c8085582",
          6277 => x"b5c808a0",
          6278 => x"38a05382",
          6279 => x"b5c80852",
          6280 => x"9c140851",
          6281 => x"eadb3f8b",
          6282 => x"53a01452",
          6283 => x"9c140851",
          6284 => x"eaac3f81",
          6285 => x"0b831734",
          6286 => x"7482b5c8",
          6287 => x"0c873d0d",
          6288 => x"04fd3d0d",
          6289 => x"75700898",
          6290 => x"12085470",
          6291 => x"535553ec",
          6292 => x"9a3f82b5",
          6293 => x"c8088d38",
          6294 => x"9c130853",
          6295 => x"e5733481",
          6296 => x"0b831534",
          6297 => x"853d0d04",
          6298 => x"fa3d0d78",
          6299 => x"7a575780",
          6300 => x"0b891734",
          6301 => x"98170880",
          6302 => x"2e818238",
          6303 => x"80708918",
          6304 => x"5555559c",
          6305 => x"17081470",
          6306 => x"33811656",
          6307 => x"515271a0",
          6308 => x"2ea83871",
          6309 => x"852e0981",
          6310 => x"06843881",
          6311 => x"e5527389",
          6312 => x"2e098106",
          6313 => x"8b38ae73",
          6314 => x"70810555",
          6315 => x"34811555",
          6316 => x"71737081",
          6317 => x"05553481",
          6318 => x"15558a74",
          6319 => x"27c53875",
          6320 => x"15880552",
          6321 => x"800b8113",
          6322 => x"349c1708",
          6323 => x"528b1233",
          6324 => x"8817349c",
          6325 => x"17089c11",
          6326 => x"5252e88a",
          6327 => x"3f82b5c8",
          6328 => x"08760c96",
          6329 => x"1251e7e7",
          6330 => x"3f82b5c8",
          6331 => x"08861723",
          6332 => x"981251e7",
          6333 => x"da3f82b5",
          6334 => x"c8088417",
          6335 => x"23883d0d",
          6336 => x"04f33d0d",
          6337 => x"7f70085e",
          6338 => x"5b806170",
          6339 => x"33515555",
          6340 => x"73af2e83",
          6341 => x"38815573",
          6342 => x"80dc2e91",
          6343 => x"3874802e",
          6344 => x"8c38941d",
          6345 => x"08881c0c",
          6346 => x"aa398115",
          6347 => x"41806170",
          6348 => x"33565656",
          6349 => x"73af2e09",
          6350 => x"81068338",
          6351 => x"81567380",
          6352 => x"dc327030",
          6353 => x"70802578",
          6354 => x"07515154",
          6355 => x"73dc3873",
          6356 => x"881c0c60",
          6357 => x"70335154",
          6358 => x"739f2696",
          6359 => x"38ff800b",
          6360 => x"ab1c3480",
          6361 => x"527a51f6",
          6362 => x"913f82b5",
          6363 => x"c8085585",
          6364 => x"9839913d",
          6365 => x"61a01d5c",
          6366 => x"5a5e8b53",
          6367 => x"a0527951",
          6368 => x"e7ff3f80",
          6369 => x"70595788",
          6370 => x"7933555c",
          6371 => x"73ae2e09",
          6372 => x"810680d4",
          6373 => x"38781870",
          6374 => x"33811a71",
          6375 => x"ae327030",
          6376 => x"709f2a73",
          6377 => x"82260751",
          6378 => x"51535a57",
          6379 => x"54738c38",
          6380 => x"79175475",
          6381 => x"74348117",
          6382 => x"57db3975",
          6383 => x"af327030",
          6384 => x"709f2a51",
          6385 => x"51547580",
          6386 => x"dc2e8c38",
          6387 => x"73802e87",
          6388 => x"3875a026",
          6389 => x"82bd3877",
          6390 => x"197e0ca4",
          6391 => x"54a07627",
          6392 => x"82bd38a0",
          6393 => x"5482b839",
          6394 => x"78187033",
          6395 => x"811a5a57",
          6396 => x"54a07627",
          6397 => x"81fc3875",
          6398 => x"af327030",
          6399 => x"7780dc32",
          6400 => x"70307280",
          6401 => x"25718025",
          6402 => x"07515156",
          6403 => x"51557380",
          6404 => x"2eac3884",
          6405 => x"39811858",
          6406 => x"80781a70",
          6407 => x"33515555",
          6408 => x"73af2e09",
          6409 => x"81068338",
          6410 => x"81557380",
          6411 => x"dc327030",
          6412 => x"70802577",
          6413 => x"07515154",
          6414 => x"73db3881",
          6415 => x"b53975ae",
          6416 => x"2e098106",
          6417 => x"83388154",
          6418 => x"767c2774",
          6419 => x"07547380",
          6420 => x"2ea2387b",
          6421 => x"8b327030",
          6422 => x"77ae3270",
          6423 => x"30728025",
          6424 => x"719f2a07",
          6425 => x"53515651",
          6426 => x"557481a7",
          6427 => x"3888578b",
          6428 => x"5cfef539",
          6429 => x"75982b54",
          6430 => x"7380258c",
          6431 => x"387580ff",
          6432 => x"0682af90",
          6433 => x"11335754",
          6434 => x"7551e6e1",
          6435 => x"3f82b5c8",
          6436 => x"08802eb2",
          6437 => x"38781870",
          6438 => x"33811a71",
          6439 => x"545a5654",
          6440 => x"e6d23f82",
          6441 => x"b5c80880",
          6442 => x"2e80e838",
          6443 => x"ff1c5476",
          6444 => x"742780df",
          6445 => x"38791754",
          6446 => x"75743481",
          6447 => x"177a1155",
          6448 => x"57747434",
          6449 => x"a7397552",
          6450 => x"82aeb051",
          6451 => x"e5fe3f82",
          6452 => x"b5c808bf",
          6453 => x"38ff9f16",
          6454 => x"54739926",
          6455 => x"8938e016",
          6456 => x"7081ff06",
          6457 => x"57547917",
          6458 => x"54757434",
          6459 => x"811757fd",
          6460 => x"f7397719",
          6461 => x"7e0c7680",
          6462 => x"2e993879",
          6463 => x"33547381",
          6464 => x"e52e0981",
          6465 => x"06843885",
          6466 => x"7a348454",
          6467 => x"a076278f",
          6468 => x"388b3986",
          6469 => x"5581f239",
          6470 => x"845680f3",
          6471 => x"39805473",
          6472 => x"8b1b3480",
          6473 => x"7b085852",
          6474 => x"7a51f2ce",
          6475 => x"3f82b5c8",
          6476 => x"085682b5",
          6477 => x"c80880d7",
          6478 => x"38981b08",
          6479 => x"527651e6",
          6480 => x"aa3f82b5",
          6481 => x"c8085682",
          6482 => x"b5c80880",
          6483 => x"c2389c1b",
          6484 => x"08703355",
          6485 => x"5573802e",
          6486 => x"ffbe388b",
          6487 => x"1533bf06",
          6488 => x"5473861c",
          6489 => x"348b1533",
          6490 => x"70832a70",
          6491 => x"81065155",
          6492 => x"58739238",
          6493 => x"8b537952",
          6494 => x"7451e49f",
          6495 => x"3f82b5c8",
          6496 => x"08802e8b",
          6497 => x"3875527a",
          6498 => x"51f3ba3f",
          6499 => x"ff9f3975",
          6500 => x"ab1c3357",
          6501 => x"5574802e",
          6502 => x"bb387484",
          6503 => x"2e098106",
          6504 => x"80e73875",
          6505 => x"852a7081",
          6506 => x"0677822a",
          6507 => x"58515473",
          6508 => x"802e9638",
          6509 => x"75810654",
          6510 => x"73802efb",
          6511 => x"b538ff80",
          6512 => x"0bab1c34",
          6513 => x"805580c1",
          6514 => x"39758106",
          6515 => x"5473ba38",
          6516 => x"8555b639",
          6517 => x"75822a70",
          6518 => x"81065154",
          6519 => x"73ab3886",
          6520 => x"1b337084",
          6521 => x"2a708106",
          6522 => x"51555573",
          6523 => x"802ee138",
          6524 => x"901b0883",
          6525 => x"ff061db4",
          6526 => x"05527c51",
          6527 => x"f5db3f82",
          6528 => x"b5c80888",
          6529 => x"1c0cfaea",
          6530 => x"397482b5",
          6531 => x"c80c8f3d",
          6532 => x"0d04f63d",
          6533 => x"0d7c5bff",
          6534 => x"7b087071",
          6535 => x"7355595c",
          6536 => x"55597380",
          6537 => x"2e81c638",
          6538 => x"75708105",
          6539 => x"573370a0",
          6540 => x"26525271",
          6541 => x"ba2e8d38",
          6542 => x"70ee3871",
          6543 => x"ba2e0981",
          6544 => x"0681a538",
          6545 => x"7333d011",
          6546 => x"7081ff06",
          6547 => x"51525370",
          6548 => x"89269138",
          6549 => x"82147381",
          6550 => x"ff06d005",
          6551 => x"56527176",
          6552 => x"2e80f738",
          6553 => x"800b82af",
          6554 => x"80595577",
          6555 => x"087a5557",
          6556 => x"76708105",
          6557 => x"58337470",
          6558 => x"81055633",
          6559 => x"ff9f1253",
          6560 => x"53537099",
          6561 => x"268938e0",
          6562 => x"137081ff",
          6563 => x"065451ff",
          6564 => x"9f125170",
          6565 => x"99268938",
          6566 => x"e0127081",
          6567 => x"ff065351",
          6568 => x"7230709f",
          6569 => x"2a515172",
          6570 => x"722e0981",
          6571 => x"06853870",
          6572 => x"ffbe3872",
          6573 => x"30747732",
          6574 => x"70307072",
          6575 => x"079f2a73",
          6576 => x"9f2a0753",
          6577 => x"54545170",
          6578 => x"802e8f38",
          6579 => x"81158419",
          6580 => x"59558375",
          6581 => x"25ff9438",
          6582 => x"8b397483",
          6583 => x"24863874",
          6584 => x"767c0c59",
          6585 => x"78518639",
          6586 => x"82cd9433",
          6587 => x"517082b5",
          6588 => x"c80c8c3d",
          6589 => x"0d04fa3d",
          6590 => x"0d785680",
          6591 => x"0b831734",
          6592 => x"ff0bb017",
          6593 => x"0c795275",
          6594 => x"51e2e03f",
          6595 => x"845582b5",
          6596 => x"c8088180",
          6597 => x"3884b216",
          6598 => x"51dfb43f",
          6599 => x"82b5c808",
          6600 => x"83ffff06",
          6601 => x"54835573",
          6602 => x"82d4d52e",
          6603 => x"09810680",
          6604 => x"e338800b",
          6605 => x"b4173356",
          6606 => x"577481e9",
          6607 => x"2e098106",
          6608 => x"83388157",
          6609 => x"7481eb32",
          6610 => x"70307080",
          6611 => x"25790751",
          6612 => x"5154738a",
          6613 => x"387481e8",
          6614 => x"2e098106",
          6615 => x"b5388353",
          6616 => x"82aec052",
          6617 => x"80ea1651",
          6618 => x"e0b13f82",
          6619 => x"b5c80855",
          6620 => x"82b5c808",
          6621 => x"802e9d38",
          6622 => x"855382ae",
          6623 => x"c4528186",
          6624 => x"1651e097",
          6625 => x"3f82b5c8",
          6626 => x"085582b5",
          6627 => x"c808802e",
          6628 => x"83388255",
          6629 => x"7482b5c8",
          6630 => x"0c883d0d",
          6631 => x"04f23d0d",
          6632 => x"61028405",
          6633 => x"80cb0533",
          6634 => x"58558075",
          6635 => x"0c6051fc",
          6636 => x"e13f82b5",
          6637 => x"c808588b",
          6638 => x"56800b82",
          6639 => x"b5c80824",
          6640 => x"86fc3882",
          6641 => x"b5c80884",
          6642 => x"2982cd80",
          6643 => x"05700855",
          6644 => x"538c5673",
          6645 => x"802e86e6",
          6646 => x"3873750c",
          6647 => x"7681fe06",
          6648 => x"74335457",
          6649 => x"72802eae",
          6650 => x"38811433",
          6651 => x"51d7ca3f",
          6652 => x"82b5c808",
          6653 => x"81ff0670",
          6654 => x"81065455",
          6655 => x"72983876",
          6656 => x"802e86b8",
          6657 => x"3874822a",
          6658 => x"70810651",
          6659 => x"538a5672",
          6660 => x"86ac3886",
          6661 => x"a7398074",
          6662 => x"34778115",
          6663 => x"34815281",
          6664 => x"143351d7",
          6665 => x"b23f82b5",
          6666 => x"c80881ff",
          6667 => x"06708106",
          6668 => x"54558356",
          6669 => x"72868738",
          6670 => x"76802e8f",
          6671 => x"3874822a",
          6672 => x"70810651",
          6673 => x"538a5672",
          6674 => x"85f43880",
          6675 => x"70537452",
          6676 => x"5bfda33f",
          6677 => x"82b5c808",
          6678 => x"81ff0657",
          6679 => x"76822e09",
          6680 => x"810680e2",
          6681 => x"388c3d74",
          6682 => x"56588356",
          6683 => x"83f61533",
          6684 => x"70585372",
          6685 => x"802e8d38",
          6686 => x"83fa1551",
          6687 => x"dce83f82",
          6688 => x"b5c80857",
          6689 => x"76787084",
          6690 => x"055a0cff",
          6691 => x"16901656",
          6692 => x"56758025",
          6693 => x"d738800b",
          6694 => x"8d3d5456",
          6695 => x"72708405",
          6696 => x"54085b83",
          6697 => x"577a802e",
          6698 => x"95387a52",
          6699 => x"7351fcc6",
          6700 => x"3f82b5c8",
          6701 => x"0881ff06",
          6702 => x"57817727",
          6703 => x"89388116",
          6704 => x"56837627",
          6705 => x"d7388156",
          6706 => x"76842e84",
          6707 => x"f1388d56",
          6708 => x"76812684",
          6709 => x"e938bf14",
          6710 => x"51dbf43f",
          6711 => x"82b5c808",
          6712 => x"83ffff06",
          6713 => x"53728480",
          6714 => x"2e098106",
          6715 => x"84d03880",
          6716 => x"ca1451db",
          6717 => x"da3f82b5",
          6718 => x"c80883ff",
          6719 => x"ff065877",
          6720 => x"8d3880d8",
          6721 => x"1451dbde",
          6722 => x"3f82b5c8",
          6723 => x"0858779c",
          6724 => x"150c80c4",
          6725 => x"14338215",
          6726 => x"3480c414",
          6727 => x"33ff1170",
          6728 => x"81ff0651",
          6729 => x"54558d56",
          6730 => x"72812684",
          6731 => x"91387481",
          6732 => x"ff067871",
          6733 => x"2980c116",
          6734 => x"33525953",
          6735 => x"728a1523",
          6736 => x"72802e8b",
          6737 => x"38ff1373",
          6738 => x"06537280",
          6739 => x"2e86388d",
          6740 => x"5683eb39",
          6741 => x"80c51451",
          6742 => x"daf53f82",
          6743 => x"b5c80853",
          6744 => x"82b5c808",
          6745 => x"88152372",
          6746 => x"8f06578d",
          6747 => x"567683ce",
          6748 => x"3880c714",
          6749 => x"51dad83f",
          6750 => x"82b5c808",
          6751 => x"83ffff06",
          6752 => x"55748d38",
          6753 => x"80d41451",
          6754 => x"dadc3f82",
          6755 => x"b5c80855",
          6756 => x"80c21451",
          6757 => x"dab93f82",
          6758 => x"b5c80883",
          6759 => x"ffff0653",
          6760 => x"8d567280",
          6761 => x"2e839738",
          6762 => x"88142278",
          6763 => x"1471842a",
          6764 => x"055a5a78",
          6765 => x"75268386",
          6766 => x"388a1422",
          6767 => x"52747931",
          6768 => x"51fef3bf",
          6769 => x"3f82b5c8",
          6770 => x"085582b5",
          6771 => x"c808802e",
          6772 => x"82ec3882",
          6773 => x"b5c80880",
          6774 => x"fffffff5",
          6775 => x"26833883",
          6776 => x"577483ff",
          6777 => x"f5268338",
          6778 => x"8257749f",
          6779 => x"f5268538",
          6780 => x"81578939",
          6781 => x"8d567680",
          6782 => x"2e82c338",
          6783 => x"82157098",
          6784 => x"160c7ba0",
          6785 => x"160c731c",
          6786 => x"70a4170c",
          6787 => x"7a1dac17",
          6788 => x"0c545576",
          6789 => x"832e0981",
          6790 => x"06af3880",
          6791 => x"de1451d9",
          6792 => x"ae3f82b5",
          6793 => x"c80883ff",
          6794 => x"ff06538d",
          6795 => x"5672828e",
          6796 => x"3879828a",
          6797 => x"3880e014",
          6798 => x"51d9ab3f",
          6799 => x"82b5c808",
          6800 => x"a8150c74",
          6801 => x"822b53a2",
          6802 => x"398d5679",
          6803 => x"802e81ee",
          6804 => x"387713a8",
          6805 => x"150c7415",
          6806 => x"5376822e",
          6807 => x"8d387410",
          6808 => x"1570812a",
          6809 => x"76810605",
          6810 => x"515383ff",
          6811 => x"13892a53",
          6812 => x"8d56729c",
          6813 => x"15082681",
          6814 => x"c538ff0b",
          6815 => x"90150cff",
          6816 => x"0b8c150c",
          6817 => x"ff800b84",
          6818 => x"15347683",
          6819 => x"2e098106",
          6820 => x"81923880",
          6821 => x"e41451d8",
          6822 => x"b63f82b5",
          6823 => x"c80883ff",
          6824 => x"ff065372",
          6825 => x"812e0981",
          6826 => x"0680f938",
          6827 => x"811b5273",
          6828 => x"51dbb83f",
          6829 => x"82b5c808",
          6830 => x"80ea3882",
          6831 => x"b5c80884",
          6832 => x"153484b2",
          6833 => x"1451d887",
          6834 => x"3f82b5c8",
          6835 => x"0883ffff",
          6836 => x"06537282",
          6837 => x"d4d52e09",
          6838 => x"810680c8",
          6839 => x"38b41451",
          6840 => x"d8843f82",
          6841 => x"b5c80884",
          6842 => x"8b85a4d2",
          6843 => x"2e098106",
          6844 => x"b3388498",
          6845 => x"1451d7ee",
          6846 => x"3f82b5c8",
          6847 => x"08868a85",
          6848 => x"e4f22e09",
          6849 => x"81069d38",
          6850 => x"849c1451",
          6851 => x"d7d83f82",
          6852 => x"b5c80890",
          6853 => x"150c84a0",
          6854 => x"1451d7ca",
          6855 => x"3f82b5c8",
          6856 => x"088c150c",
          6857 => x"76743482",
          6858 => x"cd902281",
          6859 => x"05537282",
          6860 => x"cd902372",
          6861 => x"86152380",
          6862 => x"0b94150c",
          6863 => x"80567582",
          6864 => x"b5c80c90",
          6865 => x"3d0d04fb",
          6866 => x"3d0d7754",
          6867 => x"89557380",
          6868 => x"2eb93873",
          6869 => x"08537280",
          6870 => x"2eb13872",
          6871 => x"33527180",
          6872 => x"2ea93886",
          6873 => x"13228415",
          6874 => x"22575271",
          6875 => x"762e0981",
          6876 => x"06993881",
          6877 => x"133351d0",
          6878 => x"c03f82b5",
          6879 => x"c8088106",
          6880 => x"52718838",
          6881 => x"71740854",
          6882 => x"55833980",
          6883 => x"53787371",
          6884 => x"0c527482",
          6885 => x"b5c80c87",
          6886 => x"3d0d04fa",
          6887 => x"3d0d02ab",
          6888 => x"05337a58",
          6889 => x"893dfc05",
          6890 => x"5256f4e6",
          6891 => x"3f8b5480",
          6892 => x"0b82b5c8",
          6893 => x"0824bc38",
          6894 => x"82b5c808",
          6895 => x"842982cd",
          6896 => x"80057008",
          6897 => x"55557380",
          6898 => x"2e843880",
          6899 => x"74347854",
          6900 => x"73802e84",
          6901 => x"38807434",
          6902 => x"78750c75",
          6903 => x"5475802e",
          6904 => x"92388053",
          6905 => x"893d7053",
          6906 => x"840551f7",
          6907 => x"b03f82b5",
          6908 => x"c8085473",
          6909 => x"82b5c80c",
          6910 => x"883d0d04",
          6911 => x"eb3d0d67",
          6912 => x"02840580",
          6913 => x"e7053359",
          6914 => x"59895478",
          6915 => x"802e84c8",
          6916 => x"3877bf06",
          6917 => x"7054983d",
          6918 => x"d0055399",
          6919 => x"3d840552",
          6920 => x"58f6fa3f",
          6921 => x"82b5c808",
          6922 => x"5582b5c8",
          6923 => x"0884a438",
          6924 => x"7a5c6852",
          6925 => x"8c3d7052",
          6926 => x"56edc63f",
          6927 => x"82b5c808",
          6928 => x"5582b5c8",
          6929 => x"08923802",
          6930 => x"80d70533",
          6931 => x"70982b55",
          6932 => x"57738025",
          6933 => x"83388655",
          6934 => x"779c0654",
          6935 => x"73802e81",
          6936 => x"ab387480",
          6937 => x"2e953874",
          6938 => x"842e0981",
          6939 => x"06aa3875",
          6940 => x"51eaf83f",
          6941 => x"82b5c808",
          6942 => x"559e3902",
          6943 => x"b2053391",
          6944 => x"06547381",
          6945 => x"b8387782",
          6946 => x"2a708106",
          6947 => x"51547380",
          6948 => x"2e8e3888",
          6949 => x"5583bc39",
          6950 => x"77880758",
          6951 => x"7483b438",
          6952 => x"77832a70",
          6953 => x"81065154",
          6954 => x"73802e81",
          6955 => x"af386252",
          6956 => x"7a51e8a5",
          6957 => x"3f82b5c8",
          6958 => x"08568288",
          6959 => x"b20a5262",
          6960 => x"8e0551d4",
          6961 => x"ea3f6254",
          6962 => x"a00b8b15",
          6963 => x"34805362",
          6964 => x"527a51e8",
          6965 => x"bd3f8052",
          6966 => x"629c0551",
          6967 => x"d4d13f7a",
          6968 => x"54810b83",
          6969 => x"15347580",
          6970 => x"2e80f138",
          6971 => x"7ab01108",
          6972 => x"51548053",
          6973 => x"7552973d",
          6974 => x"d40551dd",
          6975 => x"be3f82b5",
          6976 => x"c8085582",
          6977 => x"b5c80882",
          6978 => x"ca38b739",
          6979 => x"7482c438",
          6980 => x"02b20533",
          6981 => x"70842a70",
          6982 => x"81065155",
          6983 => x"5673802e",
          6984 => x"86388455",
          6985 => x"82ad3977",
          6986 => x"812a7081",
          6987 => x"06515473",
          6988 => x"802ea938",
          6989 => x"75810654",
          6990 => x"73802ea0",
          6991 => x"38875582",
          6992 => x"92397352",
          6993 => x"7a51d6a3",
          6994 => x"3f82b5c8",
          6995 => x"087bff18",
          6996 => x"8c120c55",
          6997 => x"5582b5c8",
          6998 => x"0881f838",
          6999 => x"77832a70",
          7000 => x"81065154",
          7001 => x"73802e86",
          7002 => x"387780c0",
          7003 => x"07587ab0",
          7004 => x"1108a01b",
          7005 => x"0c63a41b",
          7006 => x"0c635370",
          7007 => x"5257e6d9",
          7008 => x"3f82b5c8",
          7009 => x"0882b5c8",
          7010 => x"08881b0c",
          7011 => x"639c0552",
          7012 => x"5ad2d33f",
          7013 => x"82b5c808",
          7014 => x"82b5c808",
          7015 => x"8c1b0c77",
          7016 => x"7a0c5686",
          7017 => x"1722841a",
          7018 => x"2377901a",
          7019 => x"34800b91",
          7020 => x"1a34800b",
          7021 => x"9c1a0c80",
          7022 => x"0b941a0c",
          7023 => x"77852a70",
          7024 => x"81065154",
          7025 => x"73802e81",
          7026 => x"8d3882b5",
          7027 => x"c808802e",
          7028 => x"81843882",
          7029 => x"b5c80894",
          7030 => x"1a0c8a17",
          7031 => x"2270892b",
          7032 => x"7b525957",
          7033 => x"a8397652",
          7034 => x"7851d79f",
          7035 => x"3f82b5c8",
          7036 => x"085782b5",
          7037 => x"c8088126",
          7038 => x"83388255",
          7039 => x"82b5c808",
          7040 => x"ff2e0981",
          7041 => x"06833879",
          7042 => x"55757831",
          7043 => x"56743070",
          7044 => x"76078025",
          7045 => x"51547776",
          7046 => x"278a3881",
          7047 => x"70750655",
          7048 => x"5a73c338",
          7049 => x"76981a0c",
          7050 => x"74a93875",
          7051 => x"83ff0654",
          7052 => x"73802ea2",
          7053 => x"3876527a",
          7054 => x"51d6a63f",
          7055 => x"82b5c808",
          7056 => x"85388255",
          7057 => x"8e397589",
          7058 => x"2a82b5c8",
          7059 => x"08059c1a",
          7060 => x"0c843980",
          7061 => x"790c7454",
          7062 => x"7382b5c8",
          7063 => x"0c973d0d",
          7064 => x"04f23d0d",
          7065 => x"60636564",
          7066 => x"40405d59",
          7067 => x"807e0c90",
          7068 => x"3dfc0552",
          7069 => x"7851f9cf",
          7070 => x"3f82b5c8",
          7071 => x"085582b5",
          7072 => x"c8088a38",
          7073 => x"91193355",
          7074 => x"74802e86",
          7075 => x"38745682",
          7076 => x"c4399019",
          7077 => x"33810655",
          7078 => x"87567480",
          7079 => x"2e82b638",
          7080 => x"9539820b",
          7081 => x"911a3482",
          7082 => x"5682aa39",
          7083 => x"810b911a",
          7084 => x"34815682",
          7085 => x"a0398c19",
          7086 => x"08941a08",
          7087 => x"3155747c",
          7088 => x"27833874",
          7089 => x"5c7b802e",
          7090 => x"82893894",
          7091 => x"19087083",
          7092 => x"ff065656",
          7093 => x"7481b238",
          7094 => x"7e8a1122",
          7095 => x"ff057789",
          7096 => x"2a065b55",
          7097 => x"79a83875",
          7098 => x"87388819",
          7099 => x"08558f39",
          7100 => x"98190852",
          7101 => x"7851d593",
          7102 => x"3f82b5c8",
          7103 => x"08558175",
          7104 => x"27ff9f38",
          7105 => x"74ff2eff",
          7106 => x"a3387498",
          7107 => x"1a0c9819",
          7108 => x"08527e51",
          7109 => x"d4cb3f82",
          7110 => x"b5c80880",
          7111 => x"2eff8338",
          7112 => x"82b5c808",
          7113 => x"1a7c892a",
          7114 => x"59577780",
          7115 => x"2e80d638",
          7116 => x"771a7f8a",
          7117 => x"1122585c",
          7118 => x"55757527",
          7119 => x"8538757a",
          7120 => x"31587754",
          7121 => x"76537c52",
          7122 => x"811b3351",
          7123 => x"ca883f82",
          7124 => x"b5c808fe",
          7125 => x"d7387e83",
          7126 => x"11335656",
          7127 => x"74802e9f",
          7128 => x"38b01608",
          7129 => x"77315574",
          7130 => x"78279438",
          7131 => x"848053b4",
          7132 => x"1652b016",
          7133 => x"08773189",
          7134 => x"2b7d0551",
          7135 => x"cfe03f77",
          7136 => x"892b56b9",
          7137 => x"39769c1a",
          7138 => x"0c941908",
          7139 => x"83ff0684",
          7140 => x"80713157",
          7141 => x"557b7627",
          7142 => x"83387b56",
          7143 => x"9c190852",
          7144 => x"7e51d1c7",
          7145 => x"3f82b5c8",
          7146 => x"08fe8138",
          7147 => x"75539419",
          7148 => x"0883ff06",
          7149 => x"1fb40552",
          7150 => x"7c51cfa2",
          7151 => x"3f7b7631",
          7152 => x"7e08177f",
          7153 => x"0c761e94",
          7154 => x"1b081894",
          7155 => x"1c0c5e5c",
          7156 => x"fdf33980",
          7157 => x"567582b5",
          7158 => x"c80c903d",
          7159 => x"0d04f23d",
          7160 => x"0d606365",
          7161 => x"6440405d",
          7162 => x"58807e0c",
          7163 => x"903dfc05",
          7164 => x"527751f6",
          7165 => x"d23f82b5",
          7166 => x"c8085582",
          7167 => x"b5c8088a",
          7168 => x"38911833",
          7169 => x"5574802e",
          7170 => x"86387456",
          7171 => x"83b83990",
          7172 => x"18337081",
          7173 => x"2a708106",
          7174 => x"51565687",
          7175 => x"5674802e",
          7176 => x"83a43895",
          7177 => x"39820b91",
          7178 => x"19348256",
          7179 => x"83983981",
          7180 => x"0b911934",
          7181 => x"8156838e",
          7182 => x"39941808",
          7183 => x"7c115656",
          7184 => x"74762784",
          7185 => x"3875095c",
          7186 => x"7b802e82",
          7187 => x"ec389418",
          7188 => x"087083ff",
          7189 => x"06565674",
          7190 => x"81fd387e",
          7191 => x"8a1122ff",
          7192 => x"0577892a",
          7193 => x"065c557a",
          7194 => x"bf38758c",
          7195 => x"38881808",
          7196 => x"55749c38",
          7197 => x"7a528539",
          7198 => x"98180852",
          7199 => x"7751d7e7",
          7200 => x"3f82b5c8",
          7201 => x"085582b5",
          7202 => x"c808802e",
          7203 => x"82ab3874",
          7204 => x"812eff91",
          7205 => x"3874ff2e",
          7206 => x"ff953874",
          7207 => x"98190c88",
          7208 => x"18088538",
          7209 => x"7488190c",
          7210 => x"7e55b015",
          7211 => x"089c1908",
          7212 => x"2e098106",
          7213 => x"8d387451",
          7214 => x"cec13f82",
          7215 => x"b5c808fe",
          7216 => x"ee389818",
          7217 => x"08527e51",
          7218 => x"d1973f82",
          7219 => x"b5c80880",
          7220 => x"2efed238",
          7221 => x"82b5c808",
          7222 => x"1b7c892a",
          7223 => x"5a577880",
          7224 => x"2e80d538",
          7225 => x"781b7f8a",
          7226 => x"1122585b",
          7227 => x"55757527",
          7228 => x"8538757b",
          7229 => x"31597854",
          7230 => x"76537c52",
          7231 => x"811a3351",
          7232 => x"c8be3f82",
          7233 => x"b5c808fe",
          7234 => x"a6387eb0",
          7235 => x"11087831",
          7236 => x"56567479",
          7237 => x"279b3884",
          7238 => x"8053b016",
          7239 => x"08773189",
          7240 => x"2b7d0552",
          7241 => x"b41651cc",
          7242 => x"b53f7e55",
          7243 => x"800b8316",
          7244 => x"3478892b",
          7245 => x"5680db39",
          7246 => x"8c180894",
          7247 => x"19082693",
          7248 => x"387e51cd",
          7249 => x"b63f82b5",
          7250 => x"c808fde3",
          7251 => x"387e77b0",
          7252 => x"120c5576",
          7253 => x"9c190c94",
          7254 => x"180883ff",
          7255 => x"06848071",
          7256 => x"3157557b",
          7257 => x"76278338",
          7258 => x"7b569c18",
          7259 => x"08527e51",
          7260 => x"cdf93f82",
          7261 => x"b5c808fd",
          7262 => x"b6387553",
          7263 => x"7c529418",
          7264 => x"0883ff06",
          7265 => x"1fb40551",
          7266 => x"cbd43f7e",
          7267 => x"55810b83",
          7268 => x"16347b76",
          7269 => x"317e0817",
          7270 => x"7f0c761e",
          7271 => x"941a0818",
          7272 => x"70941c0c",
          7273 => x"8c1b0858",
          7274 => x"585e5c74",
          7275 => x"76278338",
          7276 => x"7555748c",
          7277 => x"190cfd90",
          7278 => x"39901833",
          7279 => x"80c00755",
          7280 => x"74901934",
          7281 => x"80567582",
          7282 => x"b5c80c90",
          7283 => x"3d0d04f8",
          7284 => x"3d0d7a8b",
          7285 => x"3dfc0553",
          7286 => x"705256f2",
          7287 => x"ea3f82b5",
          7288 => x"c8085782",
          7289 => x"b5c80880",
          7290 => x"fb389016",
          7291 => x"3370862a",
          7292 => x"70810651",
          7293 => x"55557380",
          7294 => x"2e80e938",
          7295 => x"a0160852",
          7296 => x"7851cce7",
          7297 => x"3f82b5c8",
          7298 => x"085782b5",
          7299 => x"c80880d4",
          7300 => x"38a41608",
          7301 => x"8b1133a0",
          7302 => x"07555573",
          7303 => x"8b163488",
          7304 => x"16085374",
          7305 => x"52750851",
          7306 => x"dde83f8c",
          7307 => x"1608529c",
          7308 => x"1551c9fb",
          7309 => x"3f8288b2",
          7310 => x"0a529615",
          7311 => x"51c9f03f",
          7312 => x"76529215",
          7313 => x"51c9ca3f",
          7314 => x"7854810b",
          7315 => x"83153478",
          7316 => x"51ccdf3f",
          7317 => x"82b5c808",
          7318 => x"90173381",
          7319 => x"bf065557",
          7320 => x"73901734",
          7321 => x"7682b5c8",
          7322 => x"0c8a3d0d",
          7323 => x"04fc3d0d",
          7324 => x"76705254",
          7325 => x"fed93f82",
          7326 => x"b5c80853",
          7327 => x"82b5c808",
          7328 => x"9c38863d",
          7329 => x"fc055273",
          7330 => x"51f1bc3f",
          7331 => x"82b5c808",
          7332 => x"5382b5c8",
          7333 => x"08873882",
          7334 => x"b5c80874",
          7335 => x"0c7282b5",
          7336 => x"c80c863d",
          7337 => x"0d04ff3d",
          7338 => x"0d843d51",
          7339 => x"e6e43f8b",
          7340 => x"52800b82",
          7341 => x"b5c80824",
          7342 => x"8b3882b5",
          7343 => x"c80882cd",
          7344 => x"94348052",
          7345 => x"7182b5c8",
          7346 => x"0c833d0d",
          7347 => x"04ef3d0d",
          7348 => x"8053933d",
          7349 => x"d0055294",
          7350 => x"3d51e9c1",
          7351 => x"3f82b5c8",
          7352 => x"085582b5",
          7353 => x"c80880e0",
          7354 => x"38765863",
          7355 => x"52933dd4",
          7356 => x"0551e08d",
          7357 => x"3f82b5c8",
          7358 => x"085582b5",
          7359 => x"c808bc38",
          7360 => x"0280c705",
          7361 => x"3370982b",
          7362 => x"55567380",
          7363 => x"25893876",
          7364 => x"7a94120c",
          7365 => x"54b23902",
          7366 => x"a2053370",
          7367 => x"842a7081",
          7368 => x"06515556",
          7369 => x"73802e9e",
          7370 => x"38767f53",
          7371 => x"705254db",
          7372 => x"a83f82b5",
          7373 => x"c8089415",
          7374 => x"0c8e3982",
          7375 => x"b5c80884",
          7376 => x"2e098106",
          7377 => x"83388555",
          7378 => x"7482b5c8",
          7379 => x"0c933d0d",
          7380 => x"04e43d0d",
          7381 => x"6f6f5b5b",
          7382 => x"807a3480",
          7383 => x"539e3dff",
          7384 => x"b805529f",
          7385 => x"3d51e8b5",
          7386 => x"3f82b5c8",
          7387 => x"085782b5",
          7388 => x"c80882fc",
          7389 => x"387b437a",
          7390 => x"7c941108",
          7391 => x"47555864",
          7392 => x"5473802e",
          7393 => x"81ed38a0",
          7394 => x"52933d70",
          7395 => x"5255d5ea",
          7396 => x"3f82b5c8",
          7397 => x"085782b5",
          7398 => x"c80882d4",
          7399 => x"3868527b",
          7400 => x"51c9c83f",
          7401 => x"82b5c808",
          7402 => x"5782b5c8",
          7403 => x"0882c138",
          7404 => x"69527b51",
          7405 => x"daa33f82",
          7406 => x"b5c80845",
          7407 => x"76527451",
          7408 => x"d5b83f82",
          7409 => x"b5c80857",
          7410 => x"82b5c808",
          7411 => x"82a23880",
          7412 => x"527451da",
          7413 => x"eb3f82b5",
          7414 => x"c8085782",
          7415 => x"b5c808a4",
          7416 => x"3869527b",
          7417 => x"51d9f23f",
          7418 => x"7382b5c8",
          7419 => x"082ea638",
          7420 => x"76527451",
          7421 => x"d6cf3f82",
          7422 => x"b5c80857",
          7423 => x"82b5c808",
          7424 => x"802ecc38",
          7425 => x"76842e09",
          7426 => x"81068638",
          7427 => x"825781e0",
          7428 => x"397681dc",
          7429 => x"389e3dff",
          7430 => x"bc055274",
          7431 => x"51dcc93f",
          7432 => x"76903d78",
          7433 => x"11811133",
          7434 => x"51565a56",
          7435 => x"73802e91",
          7436 => x"3802b905",
          7437 => x"55811681",
          7438 => x"16703356",
          7439 => x"565673f5",
          7440 => x"38811654",
          7441 => x"73782681",
          7442 => x"90387580",
          7443 => x"2e993878",
          7444 => x"16810555",
          7445 => x"ff186f11",
          7446 => x"ff18ff18",
          7447 => x"58585558",
          7448 => x"74337434",
          7449 => x"75ee38ff",
          7450 => x"186f1155",
          7451 => x"58af7434",
          7452 => x"fe8d3977",
          7453 => x"7b2e0981",
          7454 => x"068a38ff",
          7455 => x"186f1155",
          7456 => x"58af7434",
          7457 => x"800b82cd",
          7458 => x"94337084",
          7459 => x"2982af80",
          7460 => x"05700870",
          7461 => x"33525c56",
          7462 => x"56567376",
          7463 => x"2e8d3881",
          7464 => x"16701a70",
          7465 => x"33515556",
          7466 => x"73f53882",
          7467 => x"16547378",
          7468 => x"26a73880",
          7469 => x"55747627",
          7470 => x"91387419",
          7471 => x"5473337a",
          7472 => x"7081055c",
          7473 => x"34811555",
          7474 => x"ec39ba7a",
          7475 => x"7081055c",
          7476 => x"3474ff2e",
          7477 => x"09810685",
          7478 => x"38915794",
          7479 => x"396e1881",
          7480 => x"19595473",
          7481 => x"337a7081",
          7482 => x"055c347a",
          7483 => x"7826ee38",
          7484 => x"807a3476",
          7485 => x"82b5c80c",
          7486 => x"9e3d0d04",
          7487 => x"f73d0d7b",
          7488 => x"7d8d3dfc",
          7489 => x"05547153",
          7490 => x"5755ecbb",
          7491 => x"3f82b5c8",
          7492 => x"085382b5",
          7493 => x"c80882fa",
          7494 => x"38911533",
          7495 => x"537282f2",
          7496 => x"388c1508",
          7497 => x"54737627",
          7498 => x"92389015",
          7499 => x"3370812a",
          7500 => x"70810651",
          7501 => x"54577283",
          7502 => x"38735694",
          7503 => x"15085480",
          7504 => x"7094170c",
          7505 => x"5875782e",
          7506 => x"82973879",
          7507 => x"8a112270",
          7508 => x"892b5951",
          7509 => x"5373782e",
          7510 => x"b7387652",
          7511 => x"ff1651fe",
          7512 => x"dca13f82",
          7513 => x"b5c808ff",
          7514 => x"15785470",
          7515 => x"535553fe",
          7516 => x"dc913f82",
          7517 => x"b5c80873",
          7518 => x"26963876",
          7519 => x"30707506",
          7520 => x"7094180c",
          7521 => x"77713198",
          7522 => x"18085758",
          7523 => x"5153b139",
          7524 => x"88150854",
          7525 => x"73a63873",
          7526 => x"527451cd",
          7527 => x"ca3f82b5",
          7528 => x"c8085482",
          7529 => x"b5c80881",
          7530 => x"2e819a38",
          7531 => x"82b5c808",
          7532 => x"ff2e819b",
          7533 => x"3882b5c8",
          7534 => x"0888160c",
          7535 => x"7398160c",
          7536 => x"73802e81",
          7537 => x"9c387676",
          7538 => x"2780dc38",
          7539 => x"75773194",
          7540 => x"16081894",
          7541 => x"170c9016",
          7542 => x"3370812a",
          7543 => x"70810651",
          7544 => x"555a5672",
          7545 => x"802e9a38",
          7546 => x"73527451",
          7547 => x"ccf93f82",
          7548 => x"b5c80854",
          7549 => x"82b5c808",
          7550 => x"943882b5",
          7551 => x"c80856a7",
          7552 => x"39735274",
          7553 => x"51c7843f",
          7554 => x"82b5c808",
          7555 => x"5473ff2e",
          7556 => x"be388174",
          7557 => x"27af3879",
          7558 => x"53739814",
          7559 => x"0827a638",
          7560 => x"7398160c",
          7561 => x"ffa03994",
          7562 => x"15081694",
          7563 => x"160c7583",
          7564 => x"ff065372",
          7565 => x"802eaa38",
          7566 => x"73527951",
          7567 => x"c6a33f82",
          7568 => x"b5c80894",
          7569 => x"38820b91",
          7570 => x"16348253",
          7571 => x"80c43981",
          7572 => x"0b911634",
          7573 => x"8153bb39",
          7574 => x"75892a82",
          7575 => x"b5c80805",
          7576 => x"58941508",
          7577 => x"548c1508",
          7578 => x"74279038",
          7579 => x"738c160c",
          7580 => x"90153380",
          7581 => x"c0075372",
          7582 => x"90163473",
          7583 => x"83ff0653",
          7584 => x"72802e8c",
          7585 => x"38779c16",
          7586 => x"082e8538",
          7587 => x"779c160c",
          7588 => x"80537282",
          7589 => x"b5c80c8b",
          7590 => x"3d0d04f9",
          7591 => x"3d0d7956",
          7592 => x"89547580",
          7593 => x"2e818a38",
          7594 => x"8053893d",
          7595 => x"fc05528a",
          7596 => x"3d840551",
          7597 => x"e1e73f82",
          7598 => x"b5c80855",
          7599 => x"82b5c808",
          7600 => x"80ea3877",
          7601 => x"760c7a52",
          7602 => x"7551d8b5",
          7603 => x"3f82b5c8",
          7604 => x"085582b5",
          7605 => x"c80880c3",
          7606 => x"38ab1633",
          7607 => x"70982b55",
          7608 => x"57807424",
          7609 => x"a2388616",
          7610 => x"3370842a",
          7611 => x"70810651",
          7612 => x"55577380",
          7613 => x"2ead389c",
          7614 => x"16085277",
          7615 => x"51d3da3f",
          7616 => x"82b5c808",
          7617 => x"88170c77",
          7618 => x"54861422",
          7619 => x"84172374",
          7620 => x"527551ce",
          7621 => x"e53f82b5",
          7622 => x"c8085574",
          7623 => x"842e0981",
          7624 => x"06853885",
          7625 => x"55863974",
          7626 => x"802e8438",
          7627 => x"80760c74",
          7628 => x"547382b5",
          7629 => x"c80c893d",
          7630 => x"0d04fc3d",
          7631 => x"0d76873d",
          7632 => x"fc055370",
          7633 => x"5253e7ff",
          7634 => x"3f82b5c8",
          7635 => x"08873882",
          7636 => x"b5c80873",
          7637 => x"0c863d0d",
          7638 => x"04fb3d0d",
          7639 => x"7779893d",
          7640 => x"fc055471",
          7641 => x"535654e7",
          7642 => x"de3f82b5",
          7643 => x"c8085382",
          7644 => x"b5c80880",
          7645 => x"df387493",
          7646 => x"3882b5c8",
          7647 => x"08527351",
          7648 => x"cdf83f82",
          7649 => x"b5c80853",
          7650 => x"80ca3982",
          7651 => x"b5c80852",
          7652 => x"7351d3ac",
          7653 => x"3f82b5c8",
          7654 => x"085382b5",
          7655 => x"c808842e",
          7656 => x"09810685",
          7657 => x"38805387",
          7658 => x"3982b5c8",
          7659 => x"08a63874",
          7660 => x"527351d5",
          7661 => x"b33f7252",
          7662 => x"7351cf89",
          7663 => x"3f82b5c8",
          7664 => x"08843270",
          7665 => x"30707207",
          7666 => x"9f2c7082",
          7667 => x"b5c80806",
          7668 => x"51515454",
          7669 => x"7282b5c8",
          7670 => x"0c873d0d",
          7671 => x"04ee3d0d",
          7672 => x"65578053",
          7673 => x"893d7053",
          7674 => x"963d5256",
          7675 => x"dfaf3f82",
          7676 => x"b5c80855",
          7677 => x"82b5c808",
          7678 => x"b2386452",
          7679 => x"7551d681",
          7680 => x"3f82b5c8",
          7681 => x"085582b5",
          7682 => x"c808a038",
          7683 => x"0280cb05",
          7684 => x"3370982b",
          7685 => x"55587380",
          7686 => x"25853886",
          7687 => x"558d3976",
          7688 => x"802e8838",
          7689 => x"76527551",
          7690 => x"d4be3f74",
          7691 => x"82b5c80c",
          7692 => x"943d0d04",
          7693 => x"f03d0d63",
          7694 => x"65555c80",
          7695 => x"53923dec",
          7696 => x"0552933d",
          7697 => x"51ded63f",
          7698 => x"82b5c808",
          7699 => x"5b82b5c8",
          7700 => x"08828038",
          7701 => x"7c740c73",
          7702 => x"08981108",
          7703 => x"fe119013",
          7704 => x"08595658",
          7705 => x"55757426",
          7706 => x"9138757c",
          7707 => x"0c81e439",
          7708 => x"815b81cc",
          7709 => x"39825b81",
          7710 => x"c73982b5",
          7711 => x"c8087533",
          7712 => x"55597381",
          7713 => x"2e098106",
          7714 => x"bf388275",
          7715 => x"5f577652",
          7716 => x"923df005",
          7717 => x"51c1f43f",
          7718 => x"82b5c808",
          7719 => x"ff2ed138",
          7720 => x"82b5c808",
          7721 => x"812ece38",
          7722 => x"82b5c808",
          7723 => x"307082b5",
          7724 => x"c8080780",
          7725 => x"257a0581",
          7726 => x"197f5359",
          7727 => x"5a549814",
          7728 => x"087726ca",
          7729 => x"3880f939",
          7730 => x"a4150882",
          7731 => x"b5c80857",
          7732 => x"58759838",
          7733 => x"77528118",
          7734 => x"7d5258ff",
          7735 => x"bf8d3f82",
          7736 => x"b5c8085b",
          7737 => x"82b5c808",
          7738 => x"80d6387c",
          7739 => x"70337712",
          7740 => x"ff1a5d52",
          7741 => x"56547482",
          7742 => x"2e098106",
          7743 => x"9e38b414",
          7744 => x"51ffbbcb",
          7745 => x"3f82b5c8",
          7746 => x"0883ffff",
          7747 => x"06703070",
          7748 => x"80251b82",
          7749 => x"19595b51",
          7750 => x"549b39b4",
          7751 => x"1451ffbb",
          7752 => x"c53f82b5",
          7753 => x"c808f00a",
          7754 => x"06703070",
          7755 => x"80251b84",
          7756 => x"19595b51",
          7757 => x"547583ff",
          7758 => x"067a5856",
          7759 => x"79ff9238",
          7760 => x"787c0c7c",
          7761 => x"7990120c",
          7762 => x"84113381",
          7763 => x"07565474",
          7764 => x"8415347a",
          7765 => x"82b5c80c",
          7766 => x"923d0d04",
          7767 => x"f93d0d79",
          7768 => x"8a3dfc05",
          7769 => x"53705257",
          7770 => x"e3dd3f82",
          7771 => x"b5c80856",
          7772 => x"82b5c808",
          7773 => x"81a83891",
          7774 => x"17335675",
          7775 => x"81a03890",
          7776 => x"17337081",
          7777 => x"2a708106",
          7778 => x"51555587",
          7779 => x"5573802e",
          7780 => x"818e3894",
          7781 => x"17085473",
          7782 => x"8c180827",
          7783 => x"81803873",
          7784 => x"9b3882b5",
          7785 => x"c8085388",
          7786 => x"17085276",
          7787 => x"51c48c3f",
          7788 => x"82b5c808",
          7789 => x"7488190c",
          7790 => x"5680c939",
          7791 => x"98170852",
          7792 => x"7651ffbf",
          7793 => x"c63f82b5",
          7794 => x"c808ff2e",
          7795 => x"09810683",
          7796 => x"38815682",
          7797 => x"b5c80881",
          7798 => x"2e098106",
          7799 => x"85388256",
          7800 => x"a33975a0",
          7801 => x"38775482",
          7802 => x"b5c80898",
          7803 => x"15082794",
          7804 => x"38981708",
          7805 => x"5382b5c8",
          7806 => x"08527651",
          7807 => x"c3bd3f82",
          7808 => x"b5c80856",
          7809 => x"9417088c",
          7810 => x"180c9017",
          7811 => x"3380c007",
          7812 => x"54739018",
          7813 => x"3475802e",
          7814 => x"85387591",
          7815 => x"18347555",
          7816 => x"7482b5c8",
          7817 => x"0c893d0d",
          7818 => x"04e23d0d",
          7819 => x"8253a03d",
          7820 => x"ffa40552",
          7821 => x"a13d51da",
          7822 => x"e43f82b5",
          7823 => x"c8085582",
          7824 => x"b5c80881",
          7825 => x"f5387845",
          7826 => x"a13d0852",
          7827 => x"953d7052",
          7828 => x"58d1ae3f",
          7829 => x"82b5c808",
          7830 => x"5582b5c8",
          7831 => x"0881db38",
          7832 => x"0280fb05",
          7833 => x"3370852a",
          7834 => x"70810651",
          7835 => x"55568655",
          7836 => x"7381c738",
          7837 => x"75982b54",
          7838 => x"80742481",
          7839 => x"bd380280",
          7840 => x"d6053370",
          7841 => x"81065854",
          7842 => x"87557681",
          7843 => x"ad386b52",
          7844 => x"7851ccc5",
          7845 => x"3f82b5c8",
          7846 => x"0874842a",
          7847 => x"70810651",
          7848 => x"55567380",
          7849 => x"2e80d438",
          7850 => x"785482b5",
          7851 => x"c8089415",
          7852 => x"082e8186",
          7853 => x"38735a82",
          7854 => x"b5c8085c",
          7855 => x"76528a3d",
          7856 => x"705254c7",
          7857 => x"b53f82b5",
          7858 => x"c8085582",
          7859 => x"b5c80880",
          7860 => x"e93882b5",
          7861 => x"c8085273",
          7862 => x"51cce53f",
          7863 => x"82b5c808",
          7864 => x"5582b5c8",
          7865 => x"08863887",
          7866 => x"5580cf39",
          7867 => x"82b5c808",
          7868 => x"842e8838",
          7869 => x"82b5c808",
          7870 => x"80c03877",
          7871 => x"51cec23f",
          7872 => x"82b5c808",
          7873 => x"82b5c808",
          7874 => x"307082b5",
          7875 => x"c8080780",
          7876 => x"25515555",
          7877 => x"75802e94",
          7878 => x"3873802e",
          7879 => x"8f388053",
          7880 => x"75527751",
          7881 => x"c1953f82",
          7882 => x"b5c80855",
          7883 => x"748c3878",
          7884 => x"51ffbafe",
          7885 => x"3f82b5c8",
          7886 => x"08557482",
          7887 => x"b5c80ca0",
          7888 => x"3d0d04e9",
          7889 => x"3d0d8253",
          7890 => x"993dc005",
          7891 => x"529a3d51",
          7892 => x"d8cb3f82",
          7893 => x"b5c80854",
          7894 => x"82b5c808",
          7895 => x"82b03878",
          7896 => x"5e69528e",
          7897 => x"3d705258",
          7898 => x"cf973f82",
          7899 => x"b5c80854",
          7900 => x"82b5c808",
          7901 => x"86388854",
          7902 => x"82943982",
          7903 => x"b5c80884",
          7904 => x"2e098106",
          7905 => x"82883802",
          7906 => x"80df0533",
          7907 => x"70852a81",
          7908 => x"06515586",
          7909 => x"547481f6",
          7910 => x"38785a74",
          7911 => x"528a3d70",
          7912 => x"5257c1c3",
          7913 => x"3f82b5c8",
          7914 => x"08755556",
          7915 => x"82b5c808",
          7916 => x"83388754",
          7917 => x"82b5c808",
          7918 => x"812e0981",
          7919 => x"06833882",
          7920 => x"5482b5c8",
          7921 => x"08ff2e09",
          7922 => x"81068638",
          7923 => x"815481b4",
          7924 => x"397381b0",
          7925 => x"3882b5c8",
          7926 => x"08527851",
          7927 => x"c4a43f82",
          7928 => x"b5c80854",
          7929 => x"82b5c808",
          7930 => x"819a388b",
          7931 => x"53a052b4",
          7932 => x"1951ffb7",
          7933 => x"8c3f7854",
          7934 => x"ae0bb415",
          7935 => x"34785490",
          7936 => x"0bbf1534",
          7937 => x"8288b20a",
          7938 => x"5280ca19",
          7939 => x"51ffb69f",
          7940 => x"3f755378",
          7941 => x"b4115351",
          7942 => x"c9f83fa0",
          7943 => x"5378b411",
          7944 => x"5380d405",
          7945 => x"51ffb6b6",
          7946 => x"3f7854ae",
          7947 => x"0b80d515",
          7948 => x"347f5378",
          7949 => x"80d41153",
          7950 => x"51c9d73f",
          7951 => x"7854810b",
          7952 => x"83153477",
          7953 => x"51cba43f",
          7954 => x"82b5c808",
          7955 => x"5482b5c8",
          7956 => x"08b23882",
          7957 => x"88b20a52",
          7958 => x"64960551",
          7959 => x"ffb5d03f",
          7960 => x"75536452",
          7961 => x"7851c9aa",
          7962 => x"3f645490",
          7963 => x"0b8b1534",
          7964 => x"7854810b",
          7965 => x"83153478",
          7966 => x"51ffb8b6",
          7967 => x"3f82b5c8",
          7968 => x"08548b39",
          7969 => x"80537552",
          7970 => x"7651ffbe",
          7971 => x"ae3f7382",
          7972 => x"b5c80c99",
          7973 => x"3d0d04da",
          7974 => x"3d0da93d",
          7975 => x"840551d2",
          7976 => x"f13f8253",
          7977 => x"a83dff84",
          7978 => x"0552a93d",
          7979 => x"51d5ee3f",
          7980 => x"82b5c808",
          7981 => x"5582b5c8",
          7982 => x"0882d338",
          7983 => x"784da93d",
          7984 => x"08529d3d",
          7985 => x"705258cc",
          7986 => x"b83f82b5",
          7987 => x"c8085582",
          7988 => x"b5c80882",
          7989 => x"b9380281",
          7990 => x"9b053381",
          7991 => x"a0065486",
          7992 => x"557382aa",
          7993 => x"38a053a4",
          7994 => x"3d0852a8",
          7995 => x"3dff8805",
          7996 => x"51ffb4ea",
          7997 => x"3fac5377",
          7998 => x"52923d70",
          7999 => x"5254ffb4",
          8000 => x"dd3faa3d",
          8001 => x"08527351",
          8002 => x"cbf73f82",
          8003 => x"b5c80855",
          8004 => x"82b5c808",
          8005 => x"9538636f",
          8006 => x"2e098106",
          8007 => x"883865a2",
          8008 => x"3d082e92",
          8009 => x"38885581",
          8010 => x"e53982b5",
          8011 => x"c808842e",
          8012 => x"09810681",
          8013 => x"b8387351",
          8014 => x"c9b13f82",
          8015 => x"b5c80855",
          8016 => x"82b5c808",
          8017 => x"81c83868",
          8018 => x"569353a8",
          8019 => x"3dff9505",
          8020 => x"528d1651",
          8021 => x"ffb4873f",
          8022 => x"02af0533",
          8023 => x"8b17348b",
          8024 => x"16337084",
          8025 => x"2a708106",
          8026 => x"51555573",
          8027 => x"893874a0",
          8028 => x"0754738b",
          8029 => x"17347854",
          8030 => x"810b8315",
          8031 => x"348b1633",
          8032 => x"70842a70",
          8033 => x"81065155",
          8034 => x"5573802e",
          8035 => x"80e5386e",
          8036 => x"642e80df",
          8037 => x"38755278",
          8038 => x"51c6be3f",
          8039 => x"82b5c808",
          8040 => x"527851ff",
          8041 => x"b7bb3f82",
          8042 => x"5582b5c8",
          8043 => x"08802e80",
          8044 => x"dd3882b5",
          8045 => x"c8085278",
          8046 => x"51ffb5af",
          8047 => x"3f82b5c8",
          8048 => x"087980d4",
          8049 => x"11585855",
          8050 => x"82b5c808",
          8051 => x"80c03881",
          8052 => x"16335473",
          8053 => x"ae2e0981",
          8054 => x"06993863",
          8055 => x"53755276",
          8056 => x"51c6af3f",
          8057 => x"7854810b",
          8058 => x"83153487",
          8059 => x"3982b5c8",
          8060 => x"089c3877",
          8061 => x"51c8ca3f",
          8062 => x"82b5c808",
          8063 => x"5582b5c8",
          8064 => x"088c3878",
          8065 => x"51ffb5aa",
          8066 => x"3f82b5c8",
          8067 => x"08557482",
          8068 => x"b5c80ca8",
          8069 => x"3d0d04ed",
          8070 => x"3d0d0280",
          8071 => x"db053302",
          8072 => x"840580df",
          8073 => x"05335757",
          8074 => x"8253953d",
          8075 => x"d0055296",
          8076 => x"3d51d2e9",
          8077 => x"3f82b5c8",
          8078 => x"085582b5",
          8079 => x"c80880cf",
          8080 => x"38785a65",
          8081 => x"52953dd4",
          8082 => x"0551c9b5",
          8083 => x"3f82b5c8",
          8084 => x"085582b5",
          8085 => x"c808b838",
          8086 => x"0280cf05",
          8087 => x"3381a006",
          8088 => x"54865573",
          8089 => x"aa3875a7",
          8090 => x"06617109",
          8091 => x"8b123371",
          8092 => x"067a7406",
          8093 => x"07515755",
          8094 => x"56748b15",
          8095 => x"34785481",
          8096 => x"0b831534",
          8097 => x"7851ffb4",
          8098 => x"a93f82b5",
          8099 => x"c8085574",
          8100 => x"82b5c80c",
          8101 => x"953d0d04",
          8102 => x"ef3d0d64",
          8103 => x"56825393",
          8104 => x"3dd00552",
          8105 => x"943d51d1",
          8106 => x"f43f82b5",
          8107 => x"c8085582",
          8108 => x"b5c80880",
          8109 => x"cb387658",
          8110 => x"6352933d",
          8111 => x"d40551c8",
          8112 => x"c03f82b5",
          8113 => x"c8085582",
          8114 => x"b5c808b4",
          8115 => x"380280c7",
          8116 => x"053381a0",
          8117 => x"06548655",
          8118 => x"73a63884",
          8119 => x"16228617",
          8120 => x"2271902b",
          8121 => x"07535496",
          8122 => x"1f51ffb0",
          8123 => x"c23f7654",
          8124 => x"810b8315",
          8125 => x"347651ff",
          8126 => x"b3b83f82",
          8127 => x"b5c80855",
          8128 => x"7482b5c8",
          8129 => x"0c933d0d",
          8130 => x"04ea3d0d",
          8131 => x"696b5c5a",
          8132 => x"8053983d",
          8133 => x"d0055299",
          8134 => x"3d51d181",
          8135 => x"3f82b5c8",
          8136 => x"0882b5c8",
          8137 => x"08307082",
          8138 => x"b5c80807",
          8139 => x"80255155",
          8140 => x"5779802e",
          8141 => x"81853881",
          8142 => x"70750655",
          8143 => x"5573802e",
          8144 => x"80f9387b",
          8145 => x"5d805f80",
          8146 => x"528d3d70",
          8147 => x"5254ffbe",
          8148 => x"a93f82b5",
          8149 => x"c8085782",
          8150 => x"b5c80880",
          8151 => x"d1387452",
          8152 => x"7351c3dc",
          8153 => x"3f82b5c8",
          8154 => x"085782b5",
          8155 => x"c808bf38",
          8156 => x"82b5c808",
          8157 => x"82b5c808",
          8158 => x"655b5956",
          8159 => x"78188119",
          8160 => x"7b185659",
          8161 => x"55743374",
          8162 => x"34811656",
          8163 => x"8a7827ec",
          8164 => x"388b5675",
          8165 => x"1a548074",
          8166 => x"3475802e",
          8167 => x"9e38ff16",
          8168 => x"701b7033",
          8169 => x"51555673",
          8170 => x"a02ee838",
          8171 => x"8e397684",
          8172 => x"2e098106",
          8173 => x"8638807a",
          8174 => x"34805776",
          8175 => x"30707807",
          8176 => x"80255154",
          8177 => x"7a802e80",
          8178 => x"c1387380",
          8179 => x"2ebc387b",
          8180 => x"a0110853",
          8181 => x"51ffb193",
          8182 => x"3f82b5c8",
          8183 => x"085782b5",
          8184 => x"c808a738",
          8185 => x"7b703355",
          8186 => x"5580c356",
          8187 => x"73832e8b",
          8188 => x"3880e456",
          8189 => x"73842e83",
          8190 => x"38a75675",
          8191 => x"15b40551",
          8192 => x"ffade33f",
          8193 => x"82b5c808",
          8194 => x"7b0c7682",
          8195 => x"b5c80c98",
          8196 => x"3d0d04e6",
          8197 => x"3d0d8253",
          8198 => x"9c3dffb8",
          8199 => x"05529d3d",
          8200 => x"51cefa3f",
          8201 => x"82b5c808",
          8202 => x"82b5c808",
          8203 => x"565482b5",
          8204 => x"c8088398",
          8205 => x"388b53a0",
          8206 => x"528b3d70",
          8207 => x"5259ffae",
          8208 => x"c03f736d",
          8209 => x"70337081",
          8210 => x"ff065257",
          8211 => x"55579f74",
          8212 => x"2781bc38",
          8213 => x"78587481",
          8214 => x"ff066d81",
          8215 => x"054e7052",
          8216 => x"55ffaf89",
          8217 => x"3f82b5c8",
          8218 => x"08802ea5",
          8219 => x"386c7033",
          8220 => x"70535754",
          8221 => x"ffaefd3f",
          8222 => x"82b5c808",
          8223 => x"802e8d38",
          8224 => x"74882b76",
          8225 => x"076d8105",
          8226 => x"4e558639",
          8227 => x"82b5c808",
          8228 => x"55ff9f15",
          8229 => x"7083ffff",
          8230 => x"06515473",
          8231 => x"99268a38",
          8232 => x"e0157083",
          8233 => x"ffff0656",
          8234 => x"5480ff75",
          8235 => x"27873882",
          8236 => x"ae901533",
          8237 => x"5574802e",
          8238 => x"a3387452",
          8239 => x"82b09051",
          8240 => x"ffae893f",
          8241 => x"82b5c808",
          8242 => x"933881ff",
          8243 => x"75278838",
          8244 => x"76892688",
          8245 => x"388b398a",
          8246 => x"77278638",
          8247 => x"865581ec",
          8248 => x"3981ff75",
          8249 => x"278f3874",
          8250 => x"882a5473",
          8251 => x"78708105",
          8252 => x"5a348117",
          8253 => x"57747870",
          8254 => x"81055a34",
          8255 => x"81176d70",
          8256 => x"337081ff",
          8257 => x"06525755",
          8258 => x"57739f26",
          8259 => x"fec8388b",
          8260 => x"3d335486",
          8261 => x"557381e5",
          8262 => x"2e81b138",
          8263 => x"76802e99",
          8264 => x"3802a705",
          8265 => x"55761570",
          8266 => x"33515473",
          8267 => x"a02e0981",
          8268 => x"068738ff",
          8269 => x"175776ed",
          8270 => x"38794180",
          8271 => x"43805291",
          8272 => x"3d705255",
          8273 => x"ffbab33f",
          8274 => x"82b5c808",
          8275 => x"5482b5c8",
          8276 => x"0880f738",
          8277 => x"81527451",
          8278 => x"ffbfe53f",
          8279 => x"82b5c808",
          8280 => x"5482b5c8",
          8281 => x"088d3876",
          8282 => x"80c43867",
          8283 => x"54e57434",
          8284 => x"80c63982",
          8285 => x"b5c80884",
          8286 => x"2e098106",
          8287 => x"80cc3880",
          8288 => x"5476742e",
          8289 => x"80c43881",
          8290 => x"527451ff",
          8291 => x"bdb03f82",
          8292 => x"b5c80854",
          8293 => x"82b5c808",
          8294 => x"b138a053",
          8295 => x"82b5c808",
          8296 => x"526751ff",
          8297 => x"abdb3f67",
          8298 => x"54880b8b",
          8299 => x"15348b53",
          8300 => x"78526751",
          8301 => x"ffaba73f",
          8302 => x"7954810b",
          8303 => x"83153479",
          8304 => x"51ffadee",
          8305 => x"3f82b5c8",
          8306 => x"08547355",
          8307 => x"7482b5c8",
          8308 => x"0c9c3d0d",
          8309 => x"04f23d0d",
          8310 => x"60620288",
          8311 => x"0580cb05",
          8312 => x"33933dfc",
          8313 => x"05557254",
          8314 => x"405e5ad2",
          8315 => x"da3f82b5",
          8316 => x"c8085882",
          8317 => x"b5c80882",
          8318 => x"bd38911a",
          8319 => x"33587782",
          8320 => x"b5387c80",
          8321 => x"2e97388c",
          8322 => x"1a085978",
          8323 => x"9038901a",
          8324 => x"3370812a",
          8325 => x"70810651",
          8326 => x"55557390",
          8327 => x"38875482",
          8328 => x"97398258",
          8329 => x"82903981",
          8330 => x"58828b39",
          8331 => x"7e8a1122",
          8332 => x"70892b70",
          8333 => x"557f5456",
          8334 => x"5656fec2",
          8335 => x"c63fff14",
          8336 => x"7d067030",
          8337 => x"7072079f",
          8338 => x"2a82b5c8",
          8339 => x"08058c19",
          8340 => x"087c405a",
          8341 => x"5d555581",
          8342 => x"77278838",
          8343 => x"98160877",
          8344 => x"26833882",
          8345 => x"57767756",
          8346 => x"59805674",
          8347 => x"527951ff",
          8348 => x"ae993f81",
          8349 => x"157f5555",
          8350 => x"98140875",
          8351 => x"26833882",
          8352 => x"5582b5c8",
          8353 => x"08812eff",
          8354 => x"993882b5",
          8355 => x"c808ff2e",
          8356 => x"ff953882",
          8357 => x"b5c8088e",
          8358 => x"38811656",
          8359 => x"757b2e09",
          8360 => x"81068738",
          8361 => x"93397459",
          8362 => x"80567477",
          8363 => x"2e098106",
          8364 => x"ffb93887",
          8365 => x"5880ff39",
          8366 => x"7d802eba",
          8367 => x"38787b55",
          8368 => x"557a802e",
          8369 => x"b4388115",
          8370 => x"5673812e",
          8371 => x"09810683",
          8372 => x"38ff5675",
          8373 => x"5374527e",
          8374 => x"51ffafa8",
          8375 => x"3f82b5c8",
          8376 => x"085882b5",
          8377 => x"c80880ce",
          8378 => x"38748116",
          8379 => x"ff165656",
          8380 => x"5c73d338",
          8381 => x"8439ff19",
          8382 => x"5c7e7c8c",
          8383 => x"120c557d",
          8384 => x"802eb338",
          8385 => x"78881b0c",
          8386 => x"7c8c1b0c",
          8387 => x"901a3380",
          8388 => x"c0075473",
          8389 => x"901b3498",
          8390 => x"1508fe05",
          8391 => x"90160857",
          8392 => x"54757426",
          8393 => x"9138757b",
          8394 => x"3190160c",
          8395 => x"84153381",
          8396 => x"07547384",
          8397 => x"16347754",
          8398 => x"7382b5c8",
          8399 => x"0c903d0d",
          8400 => x"04e93d0d",
          8401 => x"6b6d0288",
          8402 => x"0580eb05",
          8403 => x"339d3d54",
          8404 => x"5a5c59c5",
          8405 => x"bd3f8b56",
          8406 => x"800b82b5",
          8407 => x"c808248b",
          8408 => x"f83882b5",
          8409 => x"c8088429",
          8410 => x"82cd8005",
          8411 => x"70085155",
          8412 => x"74802e84",
          8413 => x"38807534",
          8414 => x"82b5c808",
          8415 => x"81ff065f",
          8416 => x"81527e51",
          8417 => x"ffa0d03f",
          8418 => x"82b5c808",
          8419 => x"81ff0670",
          8420 => x"81065657",
          8421 => x"8356748b",
          8422 => x"c0387682",
          8423 => x"2a708106",
          8424 => x"51558a56",
          8425 => x"748bb238",
          8426 => x"993dfc05",
          8427 => x"5383527e",
          8428 => x"51ffa4f0",
          8429 => x"3f82b5c8",
          8430 => x"08993867",
          8431 => x"5574802e",
          8432 => x"92387482",
          8433 => x"8080268b",
          8434 => x"38ff1575",
          8435 => x"06557480",
          8436 => x"2e833881",
          8437 => x"4878802e",
          8438 => x"87388480",
          8439 => x"79269238",
          8440 => x"7881800a",
          8441 => x"268b38ff",
          8442 => x"19790655",
          8443 => x"74802e86",
          8444 => x"3893568a",
          8445 => x"e4397889",
          8446 => x"2a6e892a",
          8447 => x"70892b77",
          8448 => x"59484359",
          8449 => x"7a833881",
          8450 => x"56613070",
          8451 => x"80257707",
          8452 => x"51559156",
          8453 => x"748ac238",
          8454 => x"993df805",
          8455 => x"5381527e",
          8456 => x"51ffa480",
          8457 => x"3f815682",
          8458 => x"b5c8088a",
          8459 => x"ac387783",
          8460 => x"2a707706",
          8461 => x"82b5c808",
          8462 => x"43564574",
          8463 => x"8338bf41",
          8464 => x"66558e56",
          8465 => x"6075268a",
          8466 => x"90387461",
          8467 => x"31704855",
          8468 => x"80ff7527",
          8469 => x"8a833893",
          8470 => x"56788180",
          8471 => x"2689fa38",
          8472 => x"77812a70",
          8473 => x"81065643",
          8474 => x"74802e95",
          8475 => x"38778706",
          8476 => x"5574822e",
          8477 => x"838d3877",
          8478 => x"81065574",
          8479 => x"802e8383",
          8480 => x"38778106",
          8481 => x"55935682",
          8482 => x"5e74802e",
          8483 => x"89cb3878",
          8484 => x"5a7d832e",
          8485 => x"09810680",
          8486 => x"e13878ae",
          8487 => x"3866912a",
          8488 => x"57810b82",
          8489 => x"b0b42256",
          8490 => x"5a74802e",
          8491 => x"9d387477",
          8492 => x"26983882",
          8493 => x"b0b45679",
          8494 => x"10821770",
          8495 => x"2257575a",
          8496 => x"74802e86",
          8497 => x"38767527",
          8498 => x"ee387952",
          8499 => x"6651febd",
          8500 => x"b23f82b5",
          8501 => x"c8088429",
          8502 => x"84870570",
          8503 => x"892a5e55",
          8504 => x"a05c800b",
          8505 => x"82b5c808",
          8506 => x"fc808a05",
          8507 => x"5644fdff",
          8508 => x"f00a7527",
          8509 => x"80ec3888",
          8510 => x"d33978ae",
          8511 => x"38668c2a",
          8512 => x"57810b82",
          8513 => x"b0a42256",
          8514 => x"5a74802e",
          8515 => x"9d387477",
          8516 => x"26983882",
          8517 => x"b0a45679",
          8518 => x"10821770",
          8519 => x"2257575a",
          8520 => x"74802e86",
          8521 => x"38767527",
          8522 => x"ee387952",
          8523 => x"6651febc",
          8524 => x"d23f82b5",
          8525 => x"c8081084",
          8526 => x"055782b5",
          8527 => x"c8089ff5",
          8528 => x"26963881",
          8529 => x"0b82b5c8",
          8530 => x"081082b5",
          8531 => x"c8080571",
          8532 => x"11722a83",
          8533 => x"0559565e",
          8534 => x"83ff1789",
          8535 => x"2a5d815c",
          8536 => x"a044601c",
          8537 => x"7d116505",
          8538 => x"697012ff",
          8539 => x"05713070",
          8540 => x"72067431",
          8541 => x"5c525957",
          8542 => x"59407d83",
          8543 => x"2e098106",
          8544 => x"8938761c",
          8545 => x"6018415c",
          8546 => x"8439761d",
          8547 => x"5d799029",
          8548 => x"18706231",
          8549 => x"68585155",
          8550 => x"74762687",
          8551 => x"af38757c",
          8552 => x"317d317a",
          8553 => x"53706531",
          8554 => x"5255febb",
          8555 => x"d63f82b5",
          8556 => x"c808587d",
          8557 => x"832e0981",
          8558 => x"069b3882",
          8559 => x"b5c80883",
          8560 => x"fff52680",
          8561 => x"dd387887",
          8562 => x"83387981",
          8563 => x"2a5978fd",
          8564 => x"be3886f8",
          8565 => x"397d822e",
          8566 => x"09810680",
          8567 => x"c53883ff",
          8568 => x"f50b82b5",
          8569 => x"c80827a0",
          8570 => x"38788f38",
          8571 => x"791a5574",
          8572 => x"80c02686",
          8573 => x"387459fd",
          8574 => x"96396281",
          8575 => x"06557480",
          8576 => x"2e8f3883",
          8577 => x"5efd8839",
          8578 => x"82b5c808",
          8579 => x"9ff52692",
          8580 => x"387886b8",
          8581 => x"38791a59",
          8582 => x"81807927",
          8583 => x"fcf13886",
          8584 => x"ab398055",
          8585 => x"7d812e09",
          8586 => x"81068338",
          8587 => x"7d559ff5",
          8588 => x"78278b38",
          8589 => x"74810655",
          8590 => x"8e567486",
          8591 => x"9c388480",
          8592 => x"5380527a",
          8593 => x"51ffa2b9",
          8594 => x"3f8b5382",
          8595 => x"aecc527a",
          8596 => x"51ffa28a",
          8597 => x"3f848052",
          8598 => x"8b1b51ff",
          8599 => x"a1b33f79",
          8600 => x"8d1c347b",
          8601 => x"83ffff06",
          8602 => x"528e1b51",
          8603 => x"ffa1a23f",
          8604 => x"810b901c",
          8605 => x"347d8332",
          8606 => x"70307096",
          8607 => x"2a848006",
          8608 => x"54515591",
          8609 => x"1b51ffa1",
          8610 => x"883f6655",
          8611 => x"7483ffff",
          8612 => x"26903874",
          8613 => x"83ffff06",
          8614 => x"52931b51",
          8615 => x"ffa0f23f",
          8616 => x"8a397452",
          8617 => x"a01b51ff",
          8618 => x"a1853ff8",
          8619 => x"0b951c34",
          8620 => x"bf52981b",
          8621 => x"51ffa0d9",
          8622 => x"3f81ff52",
          8623 => x"9a1b51ff",
          8624 => x"a0cf3f60",
          8625 => x"529c1b51",
          8626 => x"ffa0e43f",
          8627 => x"7d832e09",
          8628 => x"810680cb",
          8629 => x"388288b2",
          8630 => x"0a5280c3",
          8631 => x"1b51ffa0",
          8632 => x"ce3f7c52",
          8633 => x"a41b51ff",
          8634 => x"a0c53f82",
          8635 => x"52ac1b51",
          8636 => x"ffa0bc3f",
          8637 => x"8152b01b",
          8638 => x"51ffa095",
          8639 => x"3f8652b2",
          8640 => x"1b51ffa0",
          8641 => x"8c3fff80",
          8642 => x"0b80c01c",
          8643 => x"34a90b80",
          8644 => x"c21c3493",
          8645 => x"5382aed8",
          8646 => x"5280c71b",
          8647 => x"51ae3982",
          8648 => x"88b20a52",
          8649 => x"a71b51ff",
          8650 => x"a0853f7c",
          8651 => x"83ffff06",
          8652 => x"52961b51",
          8653 => x"ff9fda3f",
          8654 => x"ff800ba4",
          8655 => x"1c34a90b",
          8656 => x"a61c3493",
          8657 => x"5382aeec",
          8658 => x"52ab1b51",
          8659 => x"ffa08f3f",
          8660 => x"82d4d552",
          8661 => x"83fe1b70",
          8662 => x"5259ff9f",
          8663 => x"b43f8154",
          8664 => x"60537a52",
          8665 => x"7e51ff9b",
          8666 => x"d73f8156",
          8667 => x"82b5c808",
          8668 => x"83e7387d",
          8669 => x"832e0981",
          8670 => x"0680ee38",
          8671 => x"75546086",
          8672 => x"05537a52",
          8673 => x"7e51ff9b",
          8674 => x"b73f8480",
          8675 => x"5380527a",
          8676 => x"51ff9fed",
          8677 => x"3f848b85",
          8678 => x"a4d2527a",
          8679 => x"51ff9f8f",
          8680 => x"3f868a85",
          8681 => x"e4f25283",
          8682 => x"e41b51ff",
          8683 => x"9f813fff",
          8684 => x"185283e8",
          8685 => x"1b51ff9e",
          8686 => x"f63f8252",
          8687 => x"83ec1b51",
          8688 => x"ff9eec3f",
          8689 => x"82d4d552",
          8690 => x"7851ff9e",
          8691 => x"c43f7554",
          8692 => x"60870553",
          8693 => x"7a527e51",
          8694 => x"ff9ae53f",
          8695 => x"75546016",
          8696 => x"537a527e",
          8697 => x"51ff9ad8",
          8698 => x"3f655380",
          8699 => x"527a51ff",
          8700 => x"9f8f3f7f",
          8701 => x"5680587d",
          8702 => x"832e0981",
          8703 => x"069a38f8",
          8704 => x"527a51ff",
          8705 => x"9ea93fff",
          8706 => x"52841b51",
          8707 => x"ff9ea03f",
          8708 => x"f00a5288",
          8709 => x"1b519139",
          8710 => x"87fffff8",
          8711 => x"557d812e",
          8712 => x"8338f855",
          8713 => x"74527a51",
          8714 => x"ff9e843f",
          8715 => x"7c556157",
          8716 => x"74622683",
          8717 => x"38745776",
          8718 => x"5475537a",
          8719 => x"527e51ff",
          8720 => x"99fe3f82",
          8721 => x"b5c80882",
          8722 => x"87388480",
          8723 => x"5382b5c8",
          8724 => x"08527a51",
          8725 => x"ff9eaa3f",
          8726 => x"76167578",
          8727 => x"31565674",
          8728 => x"cd388118",
          8729 => x"5877802e",
          8730 => x"ff8d3879",
          8731 => x"557d832e",
          8732 => x"83386355",
          8733 => x"61577462",
          8734 => x"26833874",
          8735 => x"57765475",
          8736 => x"537a527e",
          8737 => x"51ff99b8",
          8738 => x"3f82b5c8",
          8739 => x"0881c138",
          8740 => x"76167578",
          8741 => x"31565674",
          8742 => x"db388c56",
          8743 => x"7d832e93",
          8744 => x"38865666",
          8745 => x"83ffff26",
          8746 => x"8a388456",
          8747 => x"7d822e83",
          8748 => x"38815664",
          8749 => x"81065877",
          8750 => x"80fe3884",
          8751 => x"80537752",
          8752 => x"7a51ff9d",
          8753 => x"bc3f82d4",
          8754 => x"d5527851",
          8755 => x"ff9cc23f",
          8756 => x"83be1b55",
          8757 => x"77753481",
          8758 => x"0b811634",
          8759 => x"810b8216",
          8760 => x"34778316",
          8761 => x"34758416",
          8762 => x"34606705",
          8763 => x"5680fdc1",
          8764 => x"527551fe",
          8765 => x"b58d3ffe",
          8766 => x"0b851634",
          8767 => x"82b5c808",
          8768 => x"822abf07",
          8769 => x"56758616",
          8770 => x"3482b5c8",
          8771 => x"08871634",
          8772 => x"605283c6",
          8773 => x"1b51ff9c",
          8774 => x"963f6652",
          8775 => x"83ca1b51",
          8776 => x"ff9c8c3f",
          8777 => x"81547753",
          8778 => x"7a527e51",
          8779 => x"ff98913f",
          8780 => x"815682b5",
          8781 => x"c808a238",
          8782 => x"80538052",
          8783 => x"7e51ff99",
          8784 => x"e33f8156",
          8785 => x"82b5c808",
          8786 => x"90388939",
          8787 => x"8e568a39",
          8788 => x"81568639",
          8789 => x"82b5c808",
          8790 => x"567582b5",
          8791 => x"c80c993d",
          8792 => x"0d04f53d",
          8793 => x"0d7d605b",
          8794 => x"59807960",
          8795 => x"ff055a57",
          8796 => x"57767825",
          8797 => x"b4388d3d",
          8798 => x"f8115555",
          8799 => x"8153fc15",
          8800 => x"527951c9",
          8801 => x"dc3f7a81",
          8802 => x"2e098106",
          8803 => x"9c388c3d",
          8804 => x"3355748d",
          8805 => x"2edb3874",
          8806 => x"76708105",
          8807 => x"58348117",
          8808 => x"57748a2e",
          8809 => x"098106c9",
          8810 => x"38807634",
          8811 => x"78557683",
          8812 => x"38765574",
          8813 => x"82b5c80c",
          8814 => x"8d3d0d04",
          8815 => x"f73d0d7b",
          8816 => x"028405b3",
          8817 => x"05335957",
          8818 => x"778a2e09",
          8819 => x"81068738",
          8820 => x"8d527651",
          8821 => x"e73f8417",
          8822 => x"08568076",
          8823 => x"24be3888",
          8824 => x"17087717",
          8825 => x"8c055659",
          8826 => x"77753481",
          8827 => x"1656bb76",
          8828 => x"25a1388b",
          8829 => x"3dfc0554",
          8830 => x"75538c17",
          8831 => x"52760851",
          8832 => x"cbdc3f79",
          8833 => x"76327030",
          8834 => x"7072079f",
          8835 => x"2a703053",
          8836 => x"51565675",
          8837 => x"84180c81",
          8838 => x"1988180c",
          8839 => x"8b3d0d04",
          8840 => x"f93d0d79",
          8841 => x"84110856",
          8842 => x"56807524",
          8843 => x"a738893d",
          8844 => x"fc055474",
          8845 => x"538c1652",
          8846 => x"750851cb",
          8847 => x"a13f82b5",
          8848 => x"c8089138",
          8849 => x"84160878",
          8850 => x"2e098106",
          8851 => x"87388816",
          8852 => x"08558339",
          8853 => x"ff557482",
          8854 => x"b5c80c89",
          8855 => x"3d0d04fd",
          8856 => x"3d0d7554",
          8857 => x"80cc5380",
          8858 => x"527351ff",
          8859 => x"9a933f76",
          8860 => x"740c853d",
          8861 => x"0d04ea3d",
          8862 => x"0d0280e3",
          8863 => x"05336a53",
          8864 => x"863d7053",
          8865 => x"5454d83f",
          8866 => x"73527251",
          8867 => x"feae3f72",
          8868 => x"51ff8d3f",
          8869 => x"983d0d04",
          8870 => x"00ffffff",
          8871 => x"ff00ffff",
          8872 => x"ffff00ff",
          8873 => x"ffffff00",
          8874 => x"00002baa",
          8875 => x"00002b2e",
          8876 => x"00002b35",
          8877 => x"00002b3c",
          8878 => x"00002b43",
          8879 => x"00002b4a",
          8880 => x"00002b51",
          8881 => x"00002b58",
          8882 => x"00002b5f",
          8883 => x"00002b66",
          8884 => x"00002b6d",
          8885 => x"00002b74",
          8886 => x"00002b7a",
          8887 => x"00002b80",
          8888 => x"00002b86",
          8889 => x"00002b8c",
          8890 => x"00002b92",
          8891 => x"00002b98",
          8892 => x"00002b9e",
          8893 => x"00002ba4",
          8894 => x"0000414f",
          8895 => x"00004155",
          8896 => x"0000415b",
          8897 => x"00004161",
          8898 => x"00004167",
          8899 => x"00004745",
          8900 => x"00004845",
          8901 => x"00004956",
          8902 => x"00004bae",
          8903 => x"0000482d",
          8904 => x"0000461a",
          8905 => x"00004a1e",
          8906 => x"00004b7f",
          8907 => x"00004a61",
          8908 => x"00004af7",
          8909 => x"00004a7d",
          8910 => x"00004900",
          8911 => x"0000461a",
          8912 => x"00004956",
          8913 => x"0000497f",
          8914 => x"00004a1e",
          8915 => x"0000461a",
          8916 => x"0000461a",
          8917 => x"00004a7d",
          8918 => x"00004af7",
          8919 => x"00004b7f",
          8920 => x"00004bae",
          8921 => x"00000e31",
          8922 => x"0000171a",
          8923 => x"0000171a",
          8924 => x"00000e60",
          8925 => x"0000171a",
          8926 => x"0000171a",
          8927 => x"0000171a",
          8928 => x"0000171a",
          8929 => x"0000171a",
          8930 => x"0000171a",
          8931 => x"0000171a",
          8932 => x"00000e1d",
          8933 => x"0000171a",
          8934 => x"00000e48",
          8935 => x"00000e78",
          8936 => x"0000171a",
          8937 => x"0000171a",
          8938 => x"0000171a",
          8939 => x"0000171a",
          8940 => x"0000171a",
          8941 => x"0000171a",
          8942 => x"0000171a",
          8943 => x"0000171a",
          8944 => x"0000171a",
          8945 => x"0000171a",
          8946 => x"0000171a",
          8947 => x"0000171a",
          8948 => x"0000171a",
          8949 => x"0000171a",
          8950 => x"0000171a",
          8951 => x"0000171a",
          8952 => x"0000171a",
          8953 => x"0000171a",
          8954 => x"0000171a",
          8955 => x"0000171a",
          8956 => x"0000171a",
          8957 => x"0000171a",
          8958 => x"0000171a",
          8959 => x"0000171a",
          8960 => x"0000171a",
          8961 => x"0000171a",
          8962 => x"0000171a",
          8963 => x"0000171a",
          8964 => x"0000171a",
          8965 => x"0000171a",
          8966 => x"0000171a",
          8967 => x"0000171a",
          8968 => x"0000171a",
          8969 => x"0000171a",
          8970 => x"0000171a",
          8971 => x"0000171a",
          8972 => x"00000fa8",
          8973 => x"0000171a",
          8974 => x"0000171a",
          8975 => x"0000171a",
          8976 => x"0000171a",
          8977 => x"00001116",
          8978 => x"0000171a",
          8979 => x"0000171a",
          8980 => x"0000171a",
          8981 => x"0000171a",
          8982 => x"0000171a",
          8983 => x"0000171a",
          8984 => x"0000171a",
          8985 => x"0000171a",
          8986 => x"0000171a",
          8987 => x"0000171a",
          8988 => x"00000ed8",
          8989 => x"0000103f",
          8990 => x"00000eaf",
          8991 => x"00000eaf",
          8992 => x"00000eaf",
          8993 => x"0000171a",
          8994 => x"0000103f",
          8995 => x"0000171a",
          8996 => x"0000171a",
          8997 => x"00000e98",
          8998 => x"0000171a",
          8999 => x"0000171a",
          9000 => x"000010ec",
          9001 => x"000010f7",
          9002 => x"0000171a",
          9003 => x"0000171a",
          9004 => x"00000f11",
          9005 => x"0000171a",
          9006 => x"0000111f",
          9007 => x"0000171a",
          9008 => x"0000171a",
          9009 => x"00001116",
          9010 => x"64696e69",
          9011 => x"74000000",
          9012 => x"64696f63",
          9013 => x"746c0000",
          9014 => x"66696e69",
          9015 => x"74000000",
          9016 => x"666c6f61",
          9017 => x"64000000",
          9018 => x"66657865",
          9019 => x"63000000",
          9020 => x"6d636c65",
          9021 => x"61720000",
          9022 => x"6d636f70",
          9023 => x"79000000",
          9024 => x"6d646966",
          9025 => x"66000000",
          9026 => x"6d64756d",
          9027 => x"70000000",
          9028 => x"6d656200",
          9029 => x"6d656800",
          9030 => x"6d657700",
          9031 => x"68696400",
          9032 => x"68696500",
          9033 => x"68666400",
          9034 => x"68666500",
          9035 => x"63616c6c",
          9036 => x"00000000",
          9037 => x"6a6d7000",
          9038 => x"72657374",
          9039 => x"61727400",
          9040 => x"72657365",
          9041 => x"74000000",
          9042 => x"696e666f",
          9043 => x"00000000",
          9044 => x"74657374",
          9045 => x"00000000",
          9046 => x"74626173",
          9047 => x"69630000",
          9048 => x"6d626173",
          9049 => x"69630000",
          9050 => x"6b696c6f",
          9051 => x"00000000",
          9052 => x"65640000",
          9053 => x"4469736b",
          9054 => x"20457272",
          9055 => x"6f720000",
          9056 => x"496e7465",
          9057 => x"726e616c",
          9058 => x"20657272",
          9059 => x"6f722e00",
          9060 => x"4469736b",
          9061 => x"206e6f74",
          9062 => x"20726561",
          9063 => x"64792e00",
          9064 => x"4e6f2066",
          9065 => x"696c6520",
          9066 => x"666f756e",
          9067 => x"642e0000",
          9068 => x"4e6f2070",
          9069 => x"61746820",
          9070 => x"666f756e",
          9071 => x"642e0000",
          9072 => x"496e7661",
          9073 => x"6c696420",
          9074 => x"66696c65",
          9075 => x"6e616d65",
          9076 => x"2e000000",
          9077 => x"41636365",
          9078 => x"73732064",
          9079 => x"656e6965",
          9080 => x"642e0000",
          9081 => x"46696c65",
          9082 => x"20616c72",
          9083 => x"65616479",
          9084 => x"20657869",
          9085 => x"7374732e",
          9086 => x"00000000",
          9087 => x"46696c65",
          9088 => x"2068616e",
          9089 => x"646c6520",
          9090 => x"696e7661",
          9091 => x"6c69642e",
          9092 => x"00000000",
          9093 => x"53442069",
          9094 => x"73207772",
          9095 => x"69746520",
          9096 => x"70726f74",
          9097 => x"65637465",
          9098 => x"642e0000",
          9099 => x"44726976",
          9100 => x"65206e75",
          9101 => x"6d626572",
          9102 => x"20697320",
          9103 => x"696e7661",
          9104 => x"6c69642e",
          9105 => x"00000000",
          9106 => x"4469736b",
          9107 => x"206e6f74",
          9108 => x"20656e61",
          9109 => x"626c6564",
          9110 => x"2e000000",
          9111 => x"4e6f2063",
          9112 => x"6f6d7061",
          9113 => x"7469626c",
          9114 => x"65206669",
          9115 => x"6c657379",
          9116 => x"7374656d",
          9117 => x"20666f75",
          9118 => x"6e64206f",
          9119 => x"6e206469",
          9120 => x"736b2e00",
          9121 => x"466f726d",
          9122 => x"61742061",
          9123 => x"626f7274",
          9124 => x"65642e00",
          9125 => x"54696d65",
          9126 => x"6f75742c",
          9127 => x"206f7065",
          9128 => x"72617469",
          9129 => x"6f6e2063",
          9130 => x"616e6365",
          9131 => x"6c6c6564",
          9132 => x"2e000000",
          9133 => x"46696c65",
          9134 => x"20697320",
          9135 => x"6c6f636b",
          9136 => x"65642e00",
          9137 => x"496e7375",
          9138 => x"66666963",
          9139 => x"69656e74",
          9140 => x"206d656d",
          9141 => x"6f72792e",
          9142 => x"00000000",
          9143 => x"546f6f20",
          9144 => x"6d616e79",
          9145 => x"206f7065",
          9146 => x"6e206669",
          9147 => x"6c65732e",
          9148 => x"00000000",
          9149 => x"50617261",
          9150 => x"6d657465",
          9151 => x"72732069",
          9152 => x"6e636f72",
          9153 => x"72656374",
          9154 => x"2e000000",
          9155 => x"53756363",
          9156 => x"6573732e",
          9157 => x"00000000",
          9158 => x"556e6b6e",
          9159 => x"6f776e20",
          9160 => x"6572726f",
          9161 => x"722e0000",
          9162 => x"0a256c75",
          9163 => x"20627974",
          9164 => x"65732025",
          9165 => x"73206174",
          9166 => x"20256c75",
          9167 => x"20627974",
          9168 => x"65732f73",
          9169 => x"65632e0a",
          9170 => x"00000000",
          9171 => x"72656164",
          9172 => x"00000000",
          9173 => x"2530386c",
          9174 => x"58000000",
          9175 => x"3a202000",
          9176 => x"25303458",
          9177 => x"00000000",
          9178 => x"20202020",
          9179 => x"20202020",
          9180 => x"00000000",
          9181 => x"25303258",
          9182 => x"00000000",
          9183 => x"20200000",
          9184 => x"207c0000",
          9185 => x"7c000000",
          9186 => x"7a4f5300",
          9187 => x"0a2a2a20",
          9188 => x"25732028",
          9189 => x"00000000",
          9190 => x"30322f30",
          9191 => x"352f3230",
          9192 => x"32300000",
          9193 => x"76312e30",
          9194 => x"32000000",
          9195 => x"205a5055",
          9196 => x"2c207265",
          9197 => x"76202530",
          9198 => x"32782920",
          9199 => x"25732025",
          9200 => x"73202a2a",
          9201 => x"0a0a0000",
          9202 => x"5a505520",
          9203 => x"496e7465",
          9204 => x"72727570",
          9205 => x"74204861",
          9206 => x"6e646c65",
          9207 => x"72000000",
          9208 => x"54696d65",
          9209 => x"7220696e",
          9210 => x"74657272",
          9211 => x"75707400",
          9212 => x"50533220",
          9213 => x"696e7465",
          9214 => x"72727570",
          9215 => x"74000000",
          9216 => x"494f4354",
          9217 => x"4c205244",
          9218 => x"20696e74",
          9219 => x"65727275",
          9220 => x"70740000",
          9221 => x"494f4354",
          9222 => x"4c205752",
          9223 => x"20696e74",
          9224 => x"65727275",
          9225 => x"70740000",
          9226 => x"55415254",
          9227 => x"30205258",
          9228 => x"20696e74",
          9229 => x"65727275",
          9230 => x"70740000",
          9231 => x"55415254",
          9232 => x"30205458",
          9233 => x"20696e74",
          9234 => x"65727275",
          9235 => x"70740000",
          9236 => x"55415254",
          9237 => x"31205258",
          9238 => x"20696e74",
          9239 => x"65727275",
          9240 => x"70740000",
          9241 => x"55415254",
          9242 => x"31205458",
          9243 => x"20696e74",
          9244 => x"65727275",
          9245 => x"70740000",
          9246 => x"53657474",
          9247 => x"696e6720",
          9248 => x"75702074",
          9249 => x"696d6572",
          9250 => x"2e2e2e00",
          9251 => x"456e6162",
          9252 => x"6c696e67",
          9253 => x"2074696d",
          9254 => x"65722e2e",
          9255 => x"2e000000",
          9256 => x"6175746f",
          9257 => x"65786563",
          9258 => x"2e626174",
          9259 => x"00000000",
          9260 => x"7a4f532e",
          9261 => x"68737400",
          9262 => x"303a0000",
          9263 => x"4661696c",
          9264 => x"65642074",
          9265 => x"6f20696e",
          9266 => x"69746961",
          9267 => x"6c697365",
          9268 => x"20736420",
          9269 => x"63617264",
          9270 => x"20302c20",
          9271 => x"706c6561",
          9272 => x"73652069",
          9273 => x"6e697420",
          9274 => x"6d616e75",
          9275 => x"616c6c79",
          9276 => x"2e000000",
          9277 => x"2a200000",
          9278 => x"436c6561",
          9279 => x"72696e67",
          9280 => x"2e2e2e2e",
          9281 => x"00000000",
          9282 => x"436f7079",
          9283 => x"696e672e",
          9284 => x"2e2e0000",
          9285 => x"436f6d70",
          9286 => x"6172696e",
          9287 => x"672e2e2e",
          9288 => x"00000000",
          9289 => x"2530386c",
          9290 => x"78282530",
          9291 => x"3878292d",
          9292 => x"3e253038",
          9293 => x"6c782825",
          9294 => x"30387829",
          9295 => x"0a000000",
          9296 => x"44756d70",
          9297 => x"204d656d",
          9298 => x"6f727900",
          9299 => x"0a436f6d",
          9300 => x"706c6574",
          9301 => x"652e0000",
          9302 => x"2530386c",
          9303 => x"58202530",
          9304 => x"32582d00",
          9305 => x"3f3f3f00",
          9306 => x"2530386c",
          9307 => x"58202530",
          9308 => x"34582d00",
          9309 => x"2530386c",
          9310 => x"58202530",
          9311 => x"386c582d",
          9312 => x"00000000",
          9313 => x"45786563",
          9314 => x"7574696e",
          9315 => x"6720636f",
          9316 => x"64652040",
          9317 => x"20253038",
          9318 => x"6c78202e",
          9319 => x"2e2e0a00",
          9320 => x"43616c6c",
          9321 => x"696e6720",
          9322 => x"636f6465",
          9323 => x"20402025",
          9324 => x"30386c78",
          9325 => x"202e2e2e",
          9326 => x"0a000000",
          9327 => x"43616c6c",
          9328 => x"20726574",
          9329 => x"75726e65",
          9330 => x"6420636f",
          9331 => x"64652028",
          9332 => x"2564292e",
          9333 => x"0a000000",
          9334 => x"52657374",
          9335 => x"61727469",
          9336 => x"6e672061",
          9337 => x"70706c69",
          9338 => x"63617469",
          9339 => x"6f6e2e2e",
          9340 => x"2e000000",
          9341 => x"436f6c64",
          9342 => x"20726562",
          9343 => x"6f6f7469",
          9344 => x"6e672e2e",
          9345 => x"2e000000",
          9346 => x"5a505500",
          9347 => x"62696e00",
          9348 => x"25643a5c",
          9349 => x"25735c25",
          9350 => x"732e2573",
          9351 => x"00000000",
          9352 => x"25643a5c",
          9353 => x"25735c25",
          9354 => x"73000000",
          9355 => x"25643a5c",
          9356 => x"25730000",
          9357 => x"42616420",
          9358 => x"636f6d6d",
          9359 => x"616e642e",
          9360 => x"00000000",
          9361 => x"52756e6e",
          9362 => x"696e672e",
          9363 => x"2e2e0000",
          9364 => x"456e6162",
          9365 => x"6c696e67",
          9366 => x"20696e74",
          9367 => x"65727275",
          9368 => x"7074732e",
          9369 => x"2e2e0000",
          9370 => x"25642f25",
          9371 => x"642f2564",
          9372 => x"2025643a",
          9373 => x"25643a25",
          9374 => x"642e2564",
          9375 => x"25640a00",
          9376 => x"536f4320",
          9377 => x"436f6e66",
          9378 => x"69677572",
          9379 => x"6174696f",
          9380 => x"6e000000",
          9381 => x"20286672",
          9382 => x"6f6d2053",
          9383 => x"6f432063",
          9384 => x"6f6e6669",
          9385 => x"67290000",
          9386 => x"3a0a4465",
          9387 => x"76696365",
          9388 => x"7320696d",
          9389 => x"706c656d",
          9390 => x"656e7465",
          9391 => x"643a0a00",
          9392 => x"20202020",
          9393 => x"57422053",
          9394 => x"4452414d",
          9395 => x"20202825",
          9396 => x"3038583a",
          9397 => x"25303858",
          9398 => x"292e0a00",
          9399 => x"20202020",
          9400 => x"53445241",
          9401 => x"4d202020",
          9402 => x"20202825",
          9403 => x"3038583a",
          9404 => x"25303858",
          9405 => x"292e0a00",
          9406 => x"20202020",
          9407 => x"494e534e",
          9408 => x"20425241",
          9409 => x"4d202825",
          9410 => x"3038583a",
          9411 => x"25303858",
          9412 => x"292e0a00",
          9413 => x"20202020",
          9414 => x"4252414d",
          9415 => x"20202020",
          9416 => x"20202825",
          9417 => x"3038583a",
          9418 => x"25303858",
          9419 => x"292e0a00",
          9420 => x"20202020",
          9421 => x"52414d20",
          9422 => x"20202020",
          9423 => x"20202825",
          9424 => x"3038583a",
          9425 => x"25303858",
          9426 => x"292e0a00",
          9427 => x"20202020",
          9428 => x"53442043",
          9429 => x"41524420",
          9430 => x"20202844",
          9431 => x"65766963",
          9432 => x"6573203d",
          9433 => x"25303264",
          9434 => x"292e0a00",
          9435 => x"20202020",
          9436 => x"54494d45",
          9437 => x"52312020",
          9438 => x"20202854",
          9439 => x"696d6572",
          9440 => x"7320203d",
          9441 => x"25303264",
          9442 => x"292e0a00",
          9443 => x"20202020",
          9444 => x"494e5452",
          9445 => x"20435452",
          9446 => x"4c202843",
          9447 => x"68616e6e",
          9448 => x"656c733d",
          9449 => x"25303264",
          9450 => x"292e0a00",
          9451 => x"20202020",
          9452 => x"57495348",
          9453 => x"424f4e45",
          9454 => x"20425553",
          9455 => x"0a000000",
          9456 => x"20202020",
          9457 => x"57422049",
          9458 => x"32430a00",
          9459 => x"20202020",
          9460 => x"494f4354",
          9461 => x"4c0a0000",
          9462 => x"20202020",
          9463 => x"5053320a",
          9464 => x"00000000",
          9465 => x"20202020",
          9466 => x"5350490a",
          9467 => x"00000000",
          9468 => x"41646472",
          9469 => x"65737365",
          9470 => x"733a0a00",
          9471 => x"20202020",
          9472 => x"43505520",
          9473 => x"52657365",
          9474 => x"74205665",
          9475 => x"63746f72",
          9476 => x"20416464",
          9477 => x"72657373",
          9478 => x"203d2025",
          9479 => x"3038580a",
          9480 => x"00000000",
          9481 => x"20202020",
          9482 => x"43505520",
          9483 => x"4d656d6f",
          9484 => x"72792053",
          9485 => x"74617274",
          9486 => x"20416464",
          9487 => x"72657373",
          9488 => x"203d2025",
          9489 => x"3038580a",
          9490 => x"00000000",
          9491 => x"20202020",
          9492 => x"53746163",
          9493 => x"6b205374",
          9494 => x"61727420",
          9495 => x"41646472",
          9496 => x"65737320",
          9497 => x"20202020",
          9498 => x"203d2025",
          9499 => x"3038580a",
          9500 => x"00000000",
          9501 => x"4d697363",
          9502 => x"3a0a0000",
          9503 => x"20202020",
          9504 => x"5a505520",
          9505 => x"49642020",
          9506 => x"20202020",
          9507 => x"20202020",
          9508 => x"20202020",
          9509 => x"20202020",
          9510 => x"203d2025",
          9511 => x"3034580a",
          9512 => x"00000000",
          9513 => x"20202020",
          9514 => x"53797374",
          9515 => x"656d2043",
          9516 => x"6c6f636b",
          9517 => x"20467265",
          9518 => x"71202020",
          9519 => x"20202020",
          9520 => x"203d2025",
          9521 => x"642e2530",
          9522 => x"34644d48",
          9523 => x"7a0a0000",
          9524 => x"20202020",
          9525 => x"53445241",
          9526 => x"4d20436c",
          9527 => x"6f636b20",
          9528 => x"46726571",
          9529 => x"20202020",
          9530 => x"20202020",
          9531 => x"203d2025",
          9532 => x"642e2530",
          9533 => x"34644d48",
          9534 => x"7a0a0000",
          9535 => x"20202020",
          9536 => x"57697368",
          9537 => x"626f6e65",
          9538 => x"20534452",
          9539 => x"414d2043",
          9540 => x"6c6f636b",
          9541 => x"20467265",
          9542 => x"713d2025",
          9543 => x"642e2530",
          9544 => x"34644d48",
          9545 => x"7a0a0000",
          9546 => x"536d616c",
          9547 => x"6c000000",
          9548 => x"4d656469",
          9549 => x"756d0000",
          9550 => x"466c6578",
          9551 => x"00000000",
          9552 => x"45564f00",
          9553 => x"45564f6d",
          9554 => x"696e0000",
          9555 => x"556e6b6e",
          9556 => x"6f776e00",
          9557 => x"000096b0",
          9558 => x"01000000",
          9559 => x"00000002",
          9560 => x"000096ac",
          9561 => x"01000000",
          9562 => x"00000003",
          9563 => x"000096a8",
          9564 => x"01000000",
          9565 => x"00000004",
          9566 => x"000096a4",
          9567 => x"01000000",
          9568 => x"00000005",
          9569 => x"000096a0",
          9570 => x"01000000",
          9571 => x"00000006",
          9572 => x"0000969c",
          9573 => x"01000000",
          9574 => x"00000007",
          9575 => x"00009698",
          9576 => x"01000000",
          9577 => x"00000001",
          9578 => x"00009694",
          9579 => x"01000000",
          9580 => x"00000008",
          9581 => x"00009690",
          9582 => x"01000000",
          9583 => x"0000000b",
          9584 => x"0000968c",
          9585 => x"01000000",
          9586 => x"00000009",
          9587 => x"00009688",
          9588 => x"01000000",
          9589 => x"0000000a",
          9590 => x"00009684",
          9591 => x"04000000",
          9592 => x"0000000d",
          9593 => x"00009680",
          9594 => x"04000000",
          9595 => x"0000000c",
          9596 => x"0000967c",
          9597 => x"04000000",
          9598 => x"0000000e",
          9599 => x"00009678",
          9600 => x"03000000",
          9601 => x"0000000f",
          9602 => x"00009674",
          9603 => x"04000000",
          9604 => x"0000000f",
          9605 => x"00009670",
          9606 => x"04000000",
          9607 => x"00000010",
          9608 => x"0000966c",
          9609 => x"04000000",
          9610 => x"00000011",
          9611 => x"00009668",
          9612 => x"03000000",
          9613 => x"00000012",
          9614 => x"00009664",
          9615 => x"03000000",
          9616 => x"00000013",
          9617 => x"00009660",
          9618 => x"03000000",
          9619 => x"00000014",
          9620 => x"0000965c",
          9621 => x"03000000",
          9622 => x"00000015",
          9623 => x"1b5b4400",
          9624 => x"1b5b4300",
          9625 => x"1b5b4200",
          9626 => x"1b5b4100",
          9627 => x"1b5b367e",
          9628 => x"1b5b357e",
          9629 => x"1b5b347e",
          9630 => x"1b304600",
          9631 => x"1b5b337e",
          9632 => x"1b5b327e",
          9633 => x"1b5b317e",
          9634 => x"10000000",
          9635 => x"0e000000",
          9636 => x"0d000000",
          9637 => x"0b000000",
          9638 => x"08000000",
          9639 => x"06000000",
          9640 => x"05000000",
          9641 => x"04000000",
          9642 => x"03000000",
          9643 => x"02000000",
          9644 => x"01000000",
          9645 => x"68697374",
          9646 => x"6f727900",
          9647 => x"68697374",
          9648 => x"00000000",
          9649 => x"21000000",
          9650 => x"2530346c",
          9651 => x"75202025",
          9652 => x"730a0000",
          9653 => x"4661696c",
          9654 => x"65642074",
          9655 => x"6f207265",
          9656 => x"73657420",
          9657 => x"74686520",
          9658 => x"68697374",
          9659 => x"6f727920",
          9660 => x"66696c65",
          9661 => x"20746f20",
          9662 => x"454f462e",
          9663 => x"00000000",
          9664 => x"43616e6e",
          9665 => x"6f74206f",
          9666 => x"70656e2f",
          9667 => x"63726561",
          9668 => x"74652068",
          9669 => x"6973746f",
          9670 => x"72792066",
          9671 => x"696c652c",
          9672 => x"20646973",
          9673 => x"61626c69",
          9674 => x"6e672e00",
          9675 => x"53440000",
          9676 => x"222a2b2c",
          9677 => x"3a3b3c3d",
          9678 => x"3e3f5b5d",
          9679 => x"7c7f0000",
          9680 => x"46415400",
          9681 => x"46415433",
          9682 => x"32000000",
          9683 => x"ebfe904d",
          9684 => x"53444f53",
          9685 => x"352e3000",
          9686 => x"4e4f204e",
          9687 => x"414d4520",
          9688 => x"20202046",
          9689 => x"41543332",
          9690 => x"20202000",
          9691 => x"4e4f204e",
          9692 => x"414d4520",
          9693 => x"20202046",
          9694 => x"41542020",
          9695 => x"20202000",
          9696 => x"0000972c",
          9697 => x"00000000",
          9698 => x"00000000",
          9699 => x"00000000",
          9700 => x"809a4541",
          9701 => x"8e418f80",
          9702 => x"45454549",
          9703 => x"49498e8f",
          9704 => x"9092924f",
          9705 => x"994f5555",
          9706 => x"59999a9b",
          9707 => x"9c9d9e9f",
          9708 => x"41494f55",
          9709 => x"a5a5a6a7",
          9710 => x"a8a9aaab",
          9711 => x"acadaeaf",
          9712 => x"b0b1b2b3",
          9713 => x"b4b5b6b7",
          9714 => x"b8b9babb",
          9715 => x"bcbdbebf",
          9716 => x"c0c1c2c3",
          9717 => x"c4c5c6c7",
          9718 => x"c8c9cacb",
          9719 => x"cccdcecf",
          9720 => x"d0d1d2d3",
          9721 => x"d4d5d6d7",
          9722 => x"d8d9dadb",
          9723 => x"dcdddedf",
          9724 => x"e0e1e2e3",
          9725 => x"e4e5e6e7",
          9726 => x"e8e9eaeb",
          9727 => x"ecedeeef",
          9728 => x"f0f1f2f3",
          9729 => x"f4f5f6f7",
          9730 => x"f8f9fafb",
          9731 => x"fcfdfeff",
          9732 => x"2b2e2c3b",
          9733 => x"3d5b5d2f",
          9734 => x"5c222a3a",
          9735 => x"3c3e3f7c",
          9736 => x"7f000000",
          9737 => x"00010004",
          9738 => x"00100040",
          9739 => x"01000200",
          9740 => x"00000000",
          9741 => x"00010002",
          9742 => x"00040008",
          9743 => x"00100020",
          9744 => x"00000000",
          9745 => x"00000000",
          9746 => x"00008cc8",
          9747 => x"01020100",
          9748 => x"00000000",
          9749 => x"00000000",
          9750 => x"00008cd0",
          9751 => x"01040100",
          9752 => x"00000000",
          9753 => x"00000000",
          9754 => x"00008cd8",
          9755 => x"01140300",
          9756 => x"00000000",
          9757 => x"00000000",
          9758 => x"00008ce0",
          9759 => x"012b0300",
          9760 => x"00000000",
          9761 => x"00000000",
          9762 => x"00008ce8",
          9763 => x"01300300",
          9764 => x"00000000",
          9765 => x"00000000",
          9766 => x"00008cf0",
          9767 => x"013c0400",
          9768 => x"00000000",
          9769 => x"00000000",
          9770 => x"00008cf8",
          9771 => x"013d0400",
          9772 => x"00000000",
          9773 => x"00000000",
          9774 => x"00008d00",
          9775 => x"013f0400",
          9776 => x"00000000",
          9777 => x"00000000",
          9778 => x"00008d08",
          9779 => x"01400400",
          9780 => x"00000000",
          9781 => x"00000000",
          9782 => x"00008d10",
          9783 => x"01410400",
          9784 => x"00000000",
          9785 => x"00000000",
          9786 => x"00008d14",
          9787 => x"01420400",
          9788 => x"00000000",
          9789 => x"00000000",
          9790 => x"00008d18",
          9791 => x"01430400",
          9792 => x"00000000",
          9793 => x"00000000",
          9794 => x"00008d1c",
          9795 => x"01500500",
          9796 => x"00000000",
          9797 => x"00000000",
          9798 => x"00008d20",
          9799 => x"01510500",
          9800 => x"00000000",
          9801 => x"00000000",
          9802 => x"00008d24",
          9803 => x"01540500",
          9804 => x"00000000",
          9805 => x"00000000",
          9806 => x"00008d28",
          9807 => x"01550500",
          9808 => x"00000000",
          9809 => x"00000000",
          9810 => x"00008d2c",
          9811 => x"01790700",
          9812 => x"00000000",
          9813 => x"00000000",
          9814 => x"00008d34",
          9815 => x"01780700",
          9816 => x"00000000",
          9817 => x"00000000",
          9818 => x"00008d38",
          9819 => x"01820800",
          9820 => x"00000000",
          9821 => x"00000000",
          9822 => x"00008d40",
          9823 => x"01830800",
          9824 => x"00000000",
          9825 => x"00000000",
          9826 => x"00008d48",
          9827 => x"01850800",
          9828 => x"00000000",
          9829 => x"00000000",
          9830 => x"00008d50",
          9831 => x"01870800",
          9832 => x"00000000",
          9833 => x"00000000",
          9834 => x"00008d58",
          9835 => x"018c0900",
          9836 => x"00000000",
          9837 => x"00000000",
          9838 => x"00008d60",
          9839 => x"018d0900",
          9840 => x"00000000",
          9841 => x"00000000",
          9842 => x"00008d68",
          9843 => x"018e0900",
          9844 => x"00000000",
          9845 => x"00000000",
          9846 => x"00008d70",
          9847 => x"018f0900",
          9848 => x"00000000",
          9849 => x"00000000",
          9850 => x"00000000",
          9851 => x"00000000",
          9852 => x"00007fff",
          9853 => x"00000000",
          9854 => x"00007fff",
          9855 => x"00010000",
          9856 => x"00007fff",
          9857 => x"00010000",
          9858 => x"00810000",
          9859 => x"01000000",
          9860 => x"017fffff",
          9861 => x"00000000",
          9862 => x"00000000",
          9863 => x"00007800",
          9864 => x"00000000",
          9865 => x"05f5e100",
          9866 => x"05f5e100",
          9867 => x"05f5e100",
          9868 => x"00000000",
          9869 => x"01010101",
          9870 => x"01010101",
          9871 => x"01011001",
          9872 => x"01000000",
          9873 => x"00000000",
          9874 => x"00000000",
          9875 => x"00000000",
          9876 => x"00000000",
          9877 => x"00000000",
          9878 => x"00000000",
          9879 => x"00000000",
          9880 => x"00000000",
          9881 => x"00000000",
          9882 => x"00000000",
          9883 => x"00000000",
          9884 => x"00000000",
          9885 => x"00000000",
          9886 => x"00000000",
          9887 => x"00000000",
          9888 => x"00000000",
          9889 => x"00000000",
          9890 => x"00000000",
          9891 => x"00000000",
          9892 => x"00000000",
          9893 => x"00000000",
          9894 => x"00000000",
          9895 => x"00000000",
          9896 => x"00000000",
          9897 => x"000096b4",
          9898 => x"01000000",
          9899 => x"000096bc",
          9900 => x"01000000",
          9901 => x"000096c4",
          9902 => x"02000000",
          9903 => x"00000000",
          9904 => x"00000000",
          9905 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

