-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b87fa",
             1 => x"f80d0b0b",
             2 => x"0b93e904",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"cd040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b93b0",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b83bf",
           162 => x"84738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93b50400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0bac",
           171 => x"cc2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0bab",
           179 => x"ab2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"96040b0b",
           269 => x"0b8ca604",
           270 => x"0b0b0b8c",
           271 => x"b6040b0b",
           272 => x"0b8cc604",
           273 => x"0b0b0b8c",
           274 => x"d6040b0b",
           275 => x"0b8ce604",
           276 => x"0b0b0b8c",
           277 => x"f6040b0b",
           278 => x"0b8d8604",
           279 => x"0b0b0b8d",
           280 => x"96040b0b",
           281 => x"0b8da604",
           282 => x"0b0b0b8d",
           283 => x"b6040b0b",
           284 => x"0b8dc604",
           285 => x"0b0b0b8d",
           286 => x"d7040b0b",
           287 => x"0b8de804",
           288 => x"0b0b0b8d",
           289 => x"f9040b0b",
           290 => x"0b8e8a04",
           291 => x"0b0b0b8e",
           292 => x"9b040b0b",
           293 => x"0b8eac04",
           294 => x"0b0b0b8e",
           295 => x"bd040b0b",
           296 => x"0b8ece04",
           297 => x"0b0b0b8e",
           298 => x"df040b0b",
           299 => x"0b8ef004",
           300 => x"0b0b0b8f",
           301 => x"81040b0b",
           302 => x"0b8f9204",
           303 => x"0b0b0b8f",
           304 => x"a3040b0b",
           305 => x"0b8fb404",
           306 => x"0b0b0b8f",
           307 => x"c5040b0b",
           308 => x"0b8fd604",
           309 => x"0b0b0b8f",
           310 => x"e7040b0b",
           311 => x"0b8ff804",
           312 => x"0b0b0b90",
           313 => x"89040b0b",
           314 => x"0b909a04",
           315 => x"0b0b0b90",
           316 => x"ab040b0b",
           317 => x"0b90bc04",
           318 => x"0b0b0b90",
           319 => x"cd040b0b",
           320 => x"0b90de04",
           321 => x"0b0b0b90",
           322 => x"ef040b0b",
           323 => x"0b918004",
           324 => x"0b0b0b91",
           325 => x"91040b0b",
           326 => x"0b91a204",
           327 => x"0b0b0b91",
           328 => x"b3040b0b",
           329 => x"0b91c404",
           330 => x"0b0b0b91",
           331 => x"d5040b0b",
           332 => x"0b91e604",
           333 => x"0b0b0b91",
           334 => x"f7040b0b",
           335 => x"0b928804",
           336 => x"0b0b0b92",
           337 => x"99040b0b",
           338 => x"0b92aa04",
           339 => x"0b0b0b92",
           340 => x"bb040b0b",
           341 => x"0b92cb04",
           342 => x"0b0b0b92",
           343 => x"dc040b0b",
           344 => x"0b92ed04",
           345 => x"0b0b0b92",
           346 => x"fe04ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0484bb90",
           386 => x"0c80d697",
           387 => x"2d84bb90",
           388 => x"0880c080",
           389 => x"900484bb",
           390 => x"900ca2ee",
           391 => x"2d84bb90",
           392 => x"0880c080",
           393 => x"900484bb",
           394 => x"900ca0f3",
           395 => x"2d84bb90",
           396 => x"0880c080",
           397 => x"900484bb",
           398 => x"900ca0e0",
           399 => x"2d84bb90",
           400 => x"0880c080",
           401 => x"900484bb",
           402 => x"900c94a3",
           403 => x"2d84bb90",
           404 => x"0880c080",
           405 => x"900484bb",
           406 => x"900ca1f6",
           407 => x"2d84bb90",
           408 => x"0880c080",
           409 => x"900484bb",
           410 => x"900caf86",
           411 => x"2d84bb90",
           412 => x"0880c080",
           413 => x"900484bb",
           414 => x"900cad82",
           415 => x"2d84bb90",
           416 => x"0880c080",
           417 => x"900484bb",
           418 => x"900c9488",
           419 => x"2d84bb90",
           420 => x"0880c080",
           421 => x"900484bb",
           422 => x"900c95a8",
           423 => x"2d84bb90",
           424 => x"0880c080",
           425 => x"900484bb",
           426 => x"900c95d1",
           427 => x"2d84bb90",
           428 => x"0880c080",
           429 => x"900484bb",
           430 => x"900cb18a",
           431 => x"2d84bb90",
           432 => x"0880c080",
           433 => x"900484bb",
           434 => x"900c80d4",
           435 => x"fc2d84bb",
           436 => x"900880c0",
           437 => x"80900484",
           438 => x"bb900c80",
           439 => x"d5e12d84",
           440 => x"bb900880",
           441 => x"c0809004",
           442 => x"84bb900c",
           443 => x"80d2b82d",
           444 => x"84bb9008",
           445 => x"80c08090",
           446 => x"0484bb90",
           447 => x"0c80d3eb",
           448 => x"2d84bb90",
           449 => x"0880c080",
           450 => x"900484bb",
           451 => x"900c82ca",
           452 => x"f62d84bb",
           453 => x"900880c0",
           454 => x"80900484",
           455 => x"bb900c82",
           456 => x"e3892d84",
           457 => x"bb900880",
           458 => x"c0809004",
           459 => x"84bb900c",
           460 => x"82d4c52d",
           461 => x"84bb9008",
           462 => x"80c08090",
           463 => x"0484bb90",
           464 => x"0c82d9a5",
           465 => x"2d84bb90",
           466 => x"0880c080",
           467 => x"900484bb",
           468 => x"900c82ed",
           469 => x"a62d84bb",
           470 => x"900880c0",
           471 => x"80900484",
           472 => x"bb900c82",
           473 => x"fafc2d84",
           474 => x"bb900880",
           475 => x"c0809004",
           476 => x"84bb900c",
           477 => x"82deb82d",
           478 => x"84bb9008",
           479 => x"80c08090",
           480 => x"0484bb90",
           481 => x"0c82f295",
           482 => x"2d84bb90",
           483 => x"0880c080",
           484 => x"900484bb",
           485 => x"900c82f3",
           486 => x"e22d84bb",
           487 => x"900880c0",
           488 => x"80900484",
           489 => x"bb900c82",
           490 => x"f4b72d84",
           491 => x"bb900880",
           492 => x"c0809004",
           493 => x"84bb900c",
           494 => x"8385b12d",
           495 => x"84bb9008",
           496 => x"80c08090",
           497 => x"0484bb90",
           498 => x"0c82fff6",
           499 => x"2d84bb90",
           500 => x"0880c080",
           501 => x"900484bb",
           502 => x"900c838c",
           503 => x"952d84bb",
           504 => x"900880c0",
           505 => x"80900484",
           506 => x"bb900c82",
           507 => x"f6942d84",
           508 => x"bb900880",
           509 => x"c0809004",
           510 => x"84bb900c",
           511 => x"83958c2d",
           512 => x"84bb9008",
           513 => x"80c08090",
           514 => x"0484bb90",
           515 => x"0c839697",
           516 => x"2d84bb90",
           517 => x"0880c080",
           518 => x"900484bb",
           519 => x"900c82e5",
           520 => x"d92d84bb",
           521 => x"900880c0",
           522 => x"80900484",
           523 => x"bb900c82",
           524 => x"e3f02d84",
           525 => x"bb900880",
           526 => x"c0809004",
           527 => x"84bb900c",
           528 => x"82e7972d",
           529 => x"84bb9008",
           530 => x"80c08090",
           531 => x"0484bb90",
           532 => x"0c82f6fe",
           533 => x"2d84bb90",
           534 => x"0880c080",
           535 => x"900484bb",
           536 => x"900c8397",
           537 => x"a92d84bb",
           538 => x"900880c0",
           539 => x"80900484",
           540 => x"bb900c83",
           541 => x"9b862d84",
           542 => x"bb900880",
           543 => x"c0809004",
           544 => x"84bb900c",
           545 => x"83a1f82d",
           546 => x"84bb9008",
           547 => x"80c08090",
           548 => x"0484bb90",
           549 => x"0c82c8c7",
           550 => x"2d84bb90",
           551 => x"0880c080",
           552 => x"900484bb",
           553 => x"900c83a5",
           554 => x"a12d84bb",
           555 => x"900880c0",
           556 => x"80900484",
           557 => x"bb900c83",
           558 => x"baa22d84",
           559 => x"bb900880",
           560 => x"c0809004",
           561 => x"84bb900c",
           562 => x"83b8d42d",
           563 => x"84bb9008",
           564 => x"80c08090",
           565 => x"0484bb90",
           566 => x"0c81f5ab",
           567 => x"2d84bb90",
           568 => x"0880c080",
           569 => x"900484bb",
           570 => x"900c81f6",
           571 => x"aa2d84bb",
           572 => x"900880c0",
           573 => x"80900484",
           574 => x"bb900c81",
           575 => x"f7a92d84",
           576 => x"bb900880",
           577 => x"c0809004",
           578 => x"84bb900c",
           579 => x"80d0ba2d",
           580 => x"84bb9008",
           581 => x"80c08090",
           582 => x"0484bb90",
           583 => x"0c80d28a",
           584 => x"2d84bb90",
           585 => x"0880c080",
           586 => x"900484bb",
           587 => x"900c80d7",
           588 => x"b52d84bb",
           589 => x"900880c0",
           590 => x"80900484",
           591 => x"bb900cb1",
           592 => x"9a2d84bb",
           593 => x"900880c0",
           594 => x"80900484",
           595 => x"bb900c81",
           596 => x"dcc92d84",
           597 => x"bb900880",
           598 => x"c0809004",
           599 => x"84bb900c",
           600 => x"81de842d",
           601 => x"84bb9008",
           602 => x"80c08090",
           603 => x"0484bb90",
           604 => x"0c81f385",
           605 => x"2d84bb90",
           606 => x"0880c080",
           607 => x"900484bb",
           608 => x"900c81d6",
           609 => x"d92d84bb",
           610 => x"900880c0",
           611 => x"8090043c",
           612 => x"04101010",
           613 => x"10101010",
           614 => x"10101010",
           615 => x"10101010",
           616 => x"10101010",
           617 => x"10101010",
           618 => x"10101010",
           619 => x"10101010",
           620 => x"53510400",
           621 => x"007381ff",
           622 => x"06738306",
           623 => x"09810583",
           624 => x"05101010",
           625 => x"2b0772fc",
           626 => x"060c5151",
           627 => x"04727280",
           628 => x"728106ff",
           629 => x"05097206",
           630 => x"05711052",
           631 => x"720a100a",
           632 => x"5372ed38",
           633 => x"51515351",
           634 => x"0484bb84",
           635 => x"7084e6f0",
           636 => x"278e3880",
           637 => x"71708405",
           638 => x"530c0b0b",
           639 => x"0b93ec04",
           640 => x"8c815180",
           641 => x"ceca0400",
           642 => x"fc3d0d87",
           643 => x"3d707084",
           644 => x"05520856",
           645 => x"53745284",
           646 => x"e6e80851",
           647 => x"81c53f86",
           648 => x"3d0d04fa",
           649 => x"3d0d787a",
           650 => x"7c851133",
           651 => x"81328106",
           652 => x"80732507",
           653 => x"56585557",
           654 => x"80527272",
           655 => x"2e098106",
           656 => x"80d338ff",
           657 => x"1477748a",
           658 => x"32703070",
           659 => x"72079f2a",
           660 => x"51555556",
           661 => x"54807425",
           662 => x"b7387180",
           663 => x"2eb23875",
           664 => x"518efa3f",
           665 => x"84bb8408",
           666 => x"5384bb84",
           667 => x"08ff2eae",
           668 => x"3884bb84",
           669 => x"08757081",
           670 => x"055734ff",
           671 => x"14738a32",
           672 => x"70307072",
           673 => x"079f2a51",
           674 => x"54545473",
           675 => x"8024cb38",
           676 => x"80753476",
           677 => x"527184bb",
           678 => x"840c883d",
           679 => x"0d04800b",
           680 => x"84bb840c",
           681 => x"883d0d04",
           682 => x"f53d0d7d",
           683 => x"54860284",
           684 => x"05990534",
           685 => x"7356fe0a",
           686 => x"588e3d88",
           687 => x"05537e52",
           688 => x"8d3de405",
           689 => x"519d3f73",
           690 => x"19548074",
           691 => x"348d3d0d",
           692 => x"04fd3d0d",
           693 => x"863d8805",
           694 => x"53765275",
           695 => x"51853f85",
           696 => x"3d0d04f1",
           697 => x"3d0d6163",
           698 => x"65425d5d",
           699 => x"80708c1f",
           700 => x"0c851e33",
           701 => x"70812a81",
           702 => x"32810655",
           703 => x"555bff54",
           704 => x"727b2e09",
           705 => x"810680d2",
           706 => x"387b3357",
           707 => x"767b2e80",
           708 => x"c538811c",
           709 => x"7b810654",
           710 => x"5c72802e",
           711 => x"818138d0",
           712 => x"175f7e89",
           713 => x"2681a338",
           714 => x"76b03270",
           715 => x"30708025",
           716 => x"51545578",
           717 => x"ae387280",
           718 => x"2ea9387a",
           719 => x"832a7081",
           720 => x"32810640",
           721 => x"547e802e",
           722 => x"9e387a82",
           723 => x"80075b7b",
           724 => x"335776ff",
           725 => x"bd388c1d",
           726 => x"08547384",
           727 => x"bb840c91",
           728 => x"3d0d047a",
           729 => x"832a5478",
           730 => x"10101079",
           731 => x"10057098",
           732 => x"2b70982c",
           733 => x"19708180",
           734 => x"0a298b0a",
           735 => x"0570982c",
           736 => x"525a5b56",
           737 => x"5f807924",
           738 => x"81863873",
           739 => x"81065372",
           740 => x"ffbd3878",
           741 => x"7c335858",
           742 => x"76fef738",
           743 => x"ffb83976",
           744 => x"a52e0981",
           745 => x"06933881",
           746 => x"73745a5a",
           747 => x"5b8a7c33",
           748 => x"585a76fe",
           749 => x"dd38ff9e",
           750 => x"397c5276",
           751 => x"518baf3f",
           752 => x"7b335776",
           753 => x"fecc38ff",
           754 => x"8d397a83",
           755 => x"2a708106",
           756 => x"5455788a",
           757 => x"38817074",
           758 => x"0640547e",
           759 => x"9538e017",
           760 => x"537280d8",
           761 => x"26973872",
           762 => x"101083cb",
           763 => x"94055473",
           764 => x"080473e0",
           765 => x"18545980",
           766 => x"d87327eb",
           767 => x"387c5276",
           768 => x"518aeb3f",
           769 => x"807c3358",
           770 => x"5b76fe86",
           771 => x"38fec739",
           772 => x"80ff59fe",
           773 => x"f639885a",
           774 => x"7f608405",
           775 => x"71087d83",
           776 => x"ffcf065e",
           777 => x"58415484",
           778 => x"bb945e79",
           779 => x"52755193",
           780 => x"9a3f84bb",
           781 => x"840881ff",
           782 => x"0684bb84",
           783 => x"0818df05",
           784 => x"56537289",
           785 => x"26883884",
           786 => x"bb8408b0",
           787 => x"0555747e",
           788 => x"70810540",
           789 => x"34795275",
           790 => x"5190ca3f",
           791 => x"84bb8408",
           792 => x"5684bb84",
           793 => x"08c5387d",
           794 => x"84bb9431",
           795 => x"982b7bb2",
           796 => x"0640567e",
           797 => x"802e8f38",
           798 => x"77848080",
           799 => x"29fc8080",
           800 => x"0570902c",
           801 => x"59557a86",
           802 => x"2a708106",
           803 => x"555f7380",
           804 => x"2e9e3877",
           805 => x"84808029",
           806 => x"f8808005",
           807 => x"5379902e",
           808 => x"8b387784",
           809 => x"808029fc",
           810 => x"80800553",
           811 => x"72902c58",
           812 => x"7a832a70",
           813 => x"81065455",
           814 => x"72802e9e",
           815 => x"3875982c",
           816 => x"7081ff06",
           817 => x"54547873",
           818 => x"2486cc38",
           819 => x"7a83fff7",
           820 => x"0670832a",
           821 => x"71862a41",
           822 => x"565b7481",
           823 => x"06547380",
           824 => x"2e85f038",
           825 => x"77793190",
           826 => x"2b70902c",
           827 => x"7c838006",
           828 => x"56595373",
           829 => x"802e8596",
           830 => x"387a812a",
           831 => x"81065473",
           832 => x"85eb387a",
           833 => x"842a8106",
           834 => x"54738698",
           835 => x"387a852a",
           836 => x"81065473",
           837 => x"8697387e",
           838 => x"81065473",
           839 => x"858f387a",
           840 => x"882a8106",
           841 => x"5f7e802e",
           842 => x"b2387778",
           843 => x"84808029",
           844 => x"fc808005",
           845 => x"70902c5a",
           846 => x"40548074",
           847 => x"259d387c",
           848 => x"52b05188",
           849 => x"a93f7778",
           850 => x"84808029",
           851 => x"fc808005",
           852 => x"70902c5a",
           853 => x"40547380",
           854 => x"24e53874",
           855 => x"81065372",
           856 => x"802eb238",
           857 => x"78798180",
           858 => x"0a2981ff",
           859 => x"0a057098",
           860 => x"2c5b5555",
           861 => x"8075259d",
           862 => x"387c52b0",
           863 => x"5187ef3f",
           864 => x"78798180",
           865 => x"0a2981ff",
           866 => x"0a057098",
           867 => x"2c5b5555",
           868 => x"748024e5",
           869 => x"387a872a",
           870 => x"7081065c",
           871 => x"557a802e",
           872 => x"81b93876",
           873 => x"80e32e84",
           874 => x"d8387680",
           875 => x"f32e81ca",
           876 => x"387680d3",
           877 => x"2e81e238",
           878 => x"7d84bb94",
           879 => x"2e96387c",
           880 => x"52ff1e70",
           881 => x"33525e87",
           882 => x"a53f7d84",
           883 => x"bb942e09",
           884 => x"8106ec38",
           885 => x"7481065b",
           886 => x"7a802efc",
           887 => x"a7387778",
           888 => x"84808029",
           889 => x"fc808005",
           890 => x"70902c5a",
           891 => x"40558075",
           892 => x"25fc9138",
           893 => x"7c52a051",
           894 => x"86f43fe2",
           895 => x"397a9007",
           896 => x"5b7aa007",
           897 => x"7c33585b",
           898 => x"76fa8738",
           899 => x"fac8397a",
           900 => x"80c0075b",
           901 => x"80f85790",
           902 => x"60618405",
           903 => x"71087e83",
           904 => x"ffcf065f",
           905 => x"5942555a",
           906 => x"fbfd397f",
           907 => x"60840577",
           908 => x"fe800a06",
           909 => x"83133370",
           910 => x"982b7207",
           911 => x"7c848080",
           912 => x"29fc8080",
           913 => x"0570902c",
           914 => x"5e525a56",
           915 => x"57415f7a",
           916 => x"872a7081",
           917 => x"065c557a",
           918 => x"fec93877",
           919 => x"78848080",
           920 => x"29fc8080",
           921 => x"0570902c",
           922 => x"5a545f80",
           923 => x"7f25feb3",
           924 => x"387c52a0",
           925 => x"5185f73f",
           926 => x"e239ff1a",
           927 => x"7083ffff",
           928 => x"065b5779",
           929 => x"83ffff2e",
           930 => x"feca387c",
           931 => x"52757081",
           932 => x"05573351",
           933 => x"85d83fe2",
           934 => x"39ff1a70",
           935 => x"83ffff06",
           936 => x"5b547983",
           937 => x"ffff2efe",
           938 => x"ab387c52",
           939 => x"75708105",
           940 => x"57335185",
           941 => x"b93fe239",
           942 => x"75fc0a06",
           943 => x"81fc0a07",
           944 => x"78848080",
           945 => x"29fc8080",
           946 => x"0570902c",
           947 => x"5a585680",
           948 => x"e37b872a",
           949 => x"7081065d",
           950 => x"56577afd",
           951 => x"c638fefb",
           952 => x"397f6084",
           953 => x"05710870",
           954 => x"53404156",
           955 => x"807e2482",
           956 => x"df387a83",
           957 => x"ffbf065b",
           958 => x"84bb945e",
           959 => x"faad397a",
           960 => x"84077c33",
           961 => x"585b76f8",
           962 => x"8938f8ca",
           963 => x"397a8807",
           964 => x"5b807c33",
           965 => x"585976f7",
           966 => x"f938f8ba",
           967 => x"397f6084",
           968 => x"05710877",
           969 => x"81065658",
           970 => x"415f7282",
           971 => x"8a387551",
           972 => x"87f63f84",
           973 => x"bb840883",
           974 => x"ffff0678",
           975 => x"7131902b",
           976 => x"545a7290",
           977 => x"2c58fe87",
           978 => x"397a80c0",
           979 => x"077c3358",
           980 => x"5b76f7be",
           981 => x"38f7ff39",
           982 => x"7f608405",
           983 => x"71087781",
           984 => x"065d5841",
           985 => x"547981cf",
           986 => x"38755187",
           987 => x"bb3f84bb",
           988 => x"840883ff",
           989 => x"ff067871",
           990 => x"31902b54",
           991 => x"5ac4397a",
           992 => x"8180077c",
           993 => x"33585b76",
           994 => x"f78838f7",
           995 => x"c9397778",
           996 => x"84808029",
           997 => x"fc808005",
           998 => x"70902c5a",
           999 => x"54548074",
          1000 => x"25fad638",
          1001 => x"7c52a051",
          1002 => x"83c43fe2",
          1003 => x"397c52b0",
          1004 => x"5183bb3f",
          1005 => x"79902e09",
          1006 => x"8106fae3",
          1007 => x"387c5276",
          1008 => x"5183ab3f",
          1009 => x"7a882a81",
          1010 => x"065f7e80",
          1011 => x"2efb8c38",
          1012 => x"fad83975",
          1013 => x"982c7871",
          1014 => x"31902b70",
          1015 => x"902c7d83",
          1016 => x"8006575a",
          1017 => x"515373fa",
          1018 => x"9038ffa2",
          1019 => x"397c52ad",
          1020 => x"5182fb3f",
          1021 => x"7e810654",
          1022 => x"73802efa",
          1023 => x"a238ffad",
          1024 => x"397c5275",
          1025 => x"982a5182",
          1026 => x"e53f7481",
          1027 => x"065b7a80",
          1028 => x"2ef7f138",
          1029 => x"fbc83978",
          1030 => x"7431982b",
          1031 => x"70982c5a",
          1032 => x"53f9b739",
          1033 => x"7c52ab51",
          1034 => x"82c43fc8",
          1035 => x"397c52a0",
          1036 => x"5182bb3f",
          1037 => x"ffbe3978",
          1038 => x"52755188",
          1039 => x"8b3f84bb",
          1040 => x"840883ff",
          1041 => x"ff067871",
          1042 => x"31902b54",
          1043 => x"5afdf339",
          1044 => x"7a82077e",
          1045 => x"307183ff",
          1046 => x"bf065257",
          1047 => x"5bfd9939",
          1048 => x"fe3d0d84",
          1049 => x"e6e40853",
          1050 => x"75527451",
          1051 => x"f3b53f84",
          1052 => x"3d0d04fa",
          1053 => x"3d0d7855",
          1054 => x"800b84e6",
          1055 => x"e8088511",
          1056 => x"3370812a",
          1057 => x"81327081",
          1058 => x"06515658",
          1059 => x"5557ff56",
          1060 => x"72772e09",
          1061 => x"810680d5",
          1062 => x"38747081",
          1063 => x"05563353",
          1064 => x"72772eb0",
          1065 => x"3884e6e8",
          1066 => x"08527251",
          1067 => x"90140853",
          1068 => x"722d84bb",
          1069 => x"8408802e",
          1070 => x"8338ff57",
          1071 => x"74708105",
          1072 => x"56335372",
          1073 => x"802e8838",
          1074 => x"84e6e808",
          1075 => x"54d73984",
          1076 => x"e6e80854",
          1077 => x"84e6e808",
          1078 => x"528a5190",
          1079 => x"14085574",
          1080 => x"2d84bb84",
          1081 => x"08802e83",
          1082 => x"38ff5776",
          1083 => x"567584bb",
          1084 => x"840c883d",
          1085 => x"0d04fa3d",
          1086 => x"0d787a56",
          1087 => x"54800b85",
          1088 => x"16337081",
          1089 => x"2a813270",
          1090 => x"81065155",
          1091 => x"5757ff56",
          1092 => x"72772e09",
          1093 => x"81069238",
          1094 => x"73708105",
          1095 => x"55335372",
          1096 => x"772e0981",
          1097 => x"06983876",
          1098 => x"567584bb",
          1099 => x"840c883d",
          1100 => x"0d047370",
          1101 => x"81055533",
          1102 => x"5372802e",
          1103 => x"ea387452",
          1104 => x"72519015",
          1105 => x"0853722d",
          1106 => x"84bb8408",
          1107 => x"802ee338",
          1108 => x"ff747081",
          1109 => x"05563354",
          1110 => x"5772e338",
          1111 => x"ca39ff3d",
          1112 => x"0d84e6e8",
          1113 => x"08527351",
          1114 => x"853f833d",
          1115 => x"0d04fa3d",
          1116 => x"0d787a85",
          1117 => x"11337081",
          1118 => x"2a813281",
          1119 => x"06565656",
          1120 => x"57ff5672",
          1121 => x"ae387382",
          1122 => x"2a810654",
          1123 => x"73802eac",
          1124 => x"388c1508",
          1125 => x"53728816",
          1126 => x"08259138",
          1127 => x"74085676",
          1128 => x"76347408",
          1129 => x"8105750c",
          1130 => x"8c150853",
          1131 => x"81138c16",
          1132 => x"0c765675",
          1133 => x"84bb840c",
          1134 => x"883d0d04",
          1135 => x"74527681",
          1136 => x"ff065190",
          1137 => x"15085473",
          1138 => x"2dff5684",
          1139 => x"bb8408e3",
          1140 => x"388c1508",
          1141 => x"81058c16",
          1142 => x"0c7656d7",
          1143 => x"39fb3d0d",
          1144 => x"77851133",
          1145 => x"7081ff06",
          1146 => x"70813281",
          1147 => x"06555556",
          1148 => x"56ff5471",
          1149 => x"b3387286",
          1150 => x"2a810652",
          1151 => x"71b33872",
          1152 => x"822a8106",
          1153 => x"5271802e",
          1154 => x"80c33875",
          1155 => x"08703353",
          1156 => x"5371802e",
          1157 => x"80f03881",
          1158 => x"13760c8c",
          1159 => x"16088105",
          1160 => x"8c170c71",
          1161 => x"81ff0654",
          1162 => x"7384bb84",
          1163 => x"0c873d0d",
          1164 => x"0474ffbf",
          1165 => x"06537285",
          1166 => x"17348c16",
          1167 => x"0881058c",
          1168 => x"170c8416",
          1169 => x"3384bb84",
          1170 => x"0c873d0d",
          1171 => x"04755194",
          1172 => x"16085574",
          1173 => x"2d84bb84",
          1174 => x"085284bb",
          1175 => x"84088025",
          1176 => x"ffb93885",
          1177 => x"16337090",
          1178 => x"07545284",
          1179 => x"bb8408ff",
          1180 => x"2e853871",
          1181 => x"a0075372",
          1182 => x"851734ff",
          1183 => x"547384bb",
          1184 => x"840c873d",
          1185 => x"0d0474a0",
          1186 => x"07537285",
          1187 => x"1734ff54",
          1188 => x"ec39fd3d",
          1189 => x"0d757771",
          1190 => x"54545471",
          1191 => x"70810553",
          1192 => x"335170f7",
          1193 => x"38ff1252",
          1194 => x"72708105",
          1195 => x"54335170",
          1196 => x"72708105",
          1197 => x"543470f0",
          1198 => x"387384bb",
          1199 => x"840c853d",
          1200 => x"0d04fc3d",
          1201 => x"0d767971",
          1202 => x"7a555552",
          1203 => x"5470802e",
          1204 => x"9d387372",
          1205 => x"27a13870",
          1206 => x"802e9338",
          1207 => x"71708105",
          1208 => x"53337370",
          1209 => x"81055534",
          1210 => x"ff115170",
          1211 => x"ef387384",
          1212 => x"bb840c86",
          1213 => x"3d0d0470",
          1214 => x"12557375",
          1215 => x"27d93870",
          1216 => x"14755353",
          1217 => x"ff13ff13",
          1218 => x"53537133",
          1219 => x"7334ff11",
          1220 => x"5170802e",
          1221 => x"d938ff13",
          1222 => x"ff135353",
          1223 => x"71337334",
          1224 => x"ff115170",
          1225 => x"df38c739",
          1226 => x"fe3d0d74",
          1227 => x"70535371",
          1228 => x"70810553",
          1229 => x"335170f7",
          1230 => x"38ff1270",
          1231 => x"743184bb",
          1232 => x"840c5184",
          1233 => x"3d0d04fd",
          1234 => x"3d0d7577",
          1235 => x"71545454",
          1236 => x"72708105",
          1237 => x"54335170",
          1238 => x"72708105",
          1239 => x"543470f0",
          1240 => x"387384bb",
          1241 => x"840c853d",
          1242 => x"0d04fd3d",
          1243 => x"0d757871",
          1244 => x"79555552",
          1245 => x"5470802e",
          1246 => x"93387170",
          1247 => x"81055333",
          1248 => x"73708105",
          1249 => x"5534ff11",
          1250 => x"5170ef38",
          1251 => x"7384bb84",
          1252 => x"0c853d0d",
          1253 => x"04fc3d0d",
          1254 => x"76787a55",
          1255 => x"56547280",
          1256 => x"2ea13873",
          1257 => x"33757081",
          1258 => x"05573352",
          1259 => x"5271712e",
          1260 => x"0981069a",
          1261 => x"38811454",
          1262 => x"71802eb7",
          1263 => x"38ff1353",
          1264 => x"72e13880",
          1265 => x"517084bb",
          1266 => x"840c863d",
          1267 => x"0d047280",
          1268 => x"2ef13873",
          1269 => x"3353ff51",
          1270 => x"72802ee9",
          1271 => x"38ff1533",
          1272 => x"52815171",
          1273 => x"802ede38",
          1274 => x"72723184",
          1275 => x"bb840c86",
          1276 => x"3d0d0471",
          1277 => x"84bb840c",
          1278 => x"863d0d04",
          1279 => x"fb3d0d77",
          1280 => x"79537052",
          1281 => x"5680c13f",
          1282 => x"84bb8408",
          1283 => x"84bb8408",
          1284 => x"81055255",
          1285 => x"81b4b23f",
          1286 => x"84bb8408",
          1287 => x"5484bb84",
          1288 => x"08802e9b",
          1289 => x"3884bb84",
          1290 => x"08155480",
          1291 => x"74347453",
          1292 => x"755284bb",
          1293 => x"840851fe",
          1294 => x"b13f84bb",
          1295 => x"84085473",
          1296 => x"84bb840c",
          1297 => x"873d0d04",
          1298 => x"fd3d0d75",
          1299 => x"77717154",
          1300 => x"55535471",
          1301 => x"802e9f38",
          1302 => x"72708105",
          1303 => x"54335170",
          1304 => x"802e8c38",
          1305 => x"ff125271",
          1306 => x"ff2e0981",
          1307 => x"06ea38ff",
          1308 => x"13707531",
          1309 => x"52527084",
          1310 => x"bb840c85",
          1311 => x"3d0d04fd",
          1312 => x"3d0d7577",
          1313 => x"79725553",
          1314 => x"54547080",
          1315 => x"2e8e3872",
          1316 => x"72708105",
          1317 => x"5434ff11",
          1318 => x"5170f438",
          1319 => x"7384bb84",
          1320 => x"0c853d0d",
          1321 => x"04fa3d0d",
          1322 => x"787a5854",
          1323 => x"a0527680",
          1324 => x"2e8b3876",
          1325 => x"5180f53f",
          1326 => x"84bb8408",
          1327 => x"52e01253",
          1328 => x"73802e8d",
          1329 => x"38735180",
          1330 => x"e33f7184",
          1331 => x"bb840831",
          1332 => x"53805272",
          1333 => x"9f2680cb",
          1334 => x"38735272",
          1335 => x"9f2e80c3",
          1336 => x"38811374",
          1337 => x"712aa072",
          1338 => x"3176712b",
          1339 => x"57545455",
          1340 => x"80567476",
          1341 => x"2ea83872",
          1342 => x"10749f2a",
          1343 => x"07741077",
          1344 => x"07787231",
          1345 => x"ff119f2c",
          1346 => x"7081067b",
          1347 => x"72067571",
          1348 => x"31ff1c5c",
          1349 => x"56525255",
          1350 => x"58555374",
          1351 => x"da387310",
          1352 => x"76075271",
          1353 => x"84bb840c",
          1354 => x"883d0d04",
          1355 => x"fc3d0d76",
          1356 => x"70fc8080",
          1357 => x"06703070",
          1358 => x"72078025",
          1359 => x"70842b90",
          1360 => x"71317571",
          1361 => x"2a7083fe",
          1362 => x"80067030",
          1363 => x"70802583",
          1364 => x"2b887131",
          1365 => x"74712a70",
          1366 => x"81f00670",
          1367 => x"30708025",
          1368 => x"822b8471",
          1369 => x"3174712a",
          1370 => x"5553751b",
          1371 => x"05738c06",
          1372 => x"70307080",
          1373 => x"25108271",
          1374 => x"3177712a",
          1375 => x"70812a81",
          1376 => x"32708106",
          1377 => x"70308274",
          1378 => x"31067519",
          1379 => x"0584bb84",
          1380 => x"0c515254",
          1381 => x"55515456",
          1382 => x"5a535555",
          1383 => x"55515656",
          1384 => x"56565158",
          1385 => x"56545286",
          1386 => x"3d0d04fd",
          1387 => x"3d0d7577",
          1388 => x"70547153",
          1389 => x"54548194",
          1390 => x"3f84bb84",
          1391 => x"08732974",
          1392 => x"713184bb",
          1393 => x"840c5385",
          1394 => x"3d0d04fa",
          1395 => x"3d0d787a",
          1396 => x"5854a053",
          1397 => x"76802e8b",
          1398 => x"387651fe",
          1399 => x"cf3f84bb",
          1400 => x"840853e0",
          1401 => x"13527380",
          1402 => x"2e8d3873",
          1403 => x"51febd3f",
          1404 => x"7284bb84",
          1405 => x"08315273",
          1406 => x"53719f26",
          1407 => x"80c53880",
          1408 => x"53719f2e",
          1409 => x"be388112",
          1410 => x"74712aa0",
          1411 => x"72317671",
          1412 => x"2b575454",
          1413 => x"55805674",
          1414 => x"762ea838",
          1415 => x"7210749f",
          1416 => x"2a077410",
          1417 => x"77077872",
          1418 => x"31ff119f",
          1419 => x"2c708106",
          1420 => x"7b720675",
          1421 => x"7131ff1c",
          1422 => x"5c565252",
          1423 => x"55585553",
          1424 => x"74da3872",
          1425 => x"84bb840c",
          1426 => x"883d0d04",
          1427 => x"fa3d0d78",
          1428 => x"9f2c7a9f",
          1429 => x"2c7a9f2c",
          1430 => x"7b327c9f",
          1431 => x"2c7d3273",
          1432 => x"73327174",
          1433 => x"31577275",
          1434 => x"31565956",
          1435 => x"595556fc",
          1436 => x"b43f84bb",
          1437 => x"84087532",
          1438 => x"753184bb",
          1439 => x"840c883d",
          1440 => x"0d04f73d",
          1441 => x"0d7b7d5b",
          1442 => x"5780707b",
          1443 => x"0c770870",
          1444 => x"33565659",
          1445 => x"73a02e09",
          1446 => x"81068f38",
          1447 => x"81157078",
          1448 => x"0c703355",
          1449 => x"5573a02e",
          1450 => x"f33873ad",
          1451 => x"2e80f538",
          1452 => x"73b02e81",
          1453 => x"8338d014",
          1454 => x"58805677",
          1455 => x"892680db",
          1456 => x"388a5880",
          1457 => x"56a07427",
          1458 => x"80c43880",
          1459 => x"e0742789",
          1460 => x"38e01470",
          1461 => x"81ff0655",
          1462 => x"53d01470",
          1463 => x"81ff0651",
          1464 => x"53907327",
          1465 => x"8f38f913",
          1466 => x"7081ff06",
          1467 => x"54548973",
          1468 => x"27818938",
          1469 => x"72782781",
          1470 => x"83387776",
          1471 => x"29138116",
          1472 => x"70790c70",
          1473 => x"33565656",
          1474 => x"73a026ff",
          1475 => x"be387880",
          1476 => x"2e843875",
          1477 => x"3056757a",
          1478 => x"0c815675",
          1479 => x"84bb840c",
          1480 => x"8b3d0d04",
          1481 => x"81701670",
          1482 => x"790c7033",
          1483 => x"56565973",
          1484 => x"b02e0981",
          1485 => x"06feff38",
          1486 => x"81157078",
          1487 => x"0c703355",
          1488 => x"557380e2",
          1489 => x"2ea63890",
          1490 => x"587380f8",
          1491 => x"2ea03881",
          1492 => x"56a07427",
          1493 => x"c638d014",
          1494 => x"53805688",
          1495 => x"58897327",
          1496 => x"fee13875",
          1497 => x"84bb840c",
          1498 => x"8b3d0d04",
          1499 => x"82588115",
          1500 => x"70780c70",
          1501 => x"33555580",
          1502 => x"56feca39",
          1503 => x"800b84bb",
          1504 => x"840c8b3d",
          1505 => x"0d04f73d",
          1506 => x"0d7b7d5b",
          1507 => x"5780707b",
          1508 => x"0c770870",
          1509 => x"33565659",
          1510 => x"73a02e09",
          1511 => x"81068f38",
          1512 => x"81157078",
          1513 => x"0c703355",
          1514 => x"5573a02e",
          1515 => x"f33873ad",
          1516 => x"2e80f538",
          1517 => x"73b02e81",
          1518 => x"8338d014",
          1519 => x"58805677",
          1520 => x"892680db",
          1521 => x"388a5880",
          1522 => x"56a07427",
          1523 => x"80c43880",
          1524 => x"e0742789",
          1525 => x"38e01470",
          1526 => x"81ff0655",
          1527 => x"53d01470",
          1528 => x"81ff0651",
          1529 => x"53907327",
          1530 => x"8f38f913",
          1531 => x"7081ff06",
          1532 => x"54548973",
          1533 => x"27818938",
          1534 => x"72782781",
          1535 => x"83387776",
          1536 => x"29138116",
          1537 => x"70790c70",
          1538 => x"33565656",
          1539 => x"73a026ff",
          1540 => x"be387880",
          1541 => x"2e843875",
          1542 => x"3056757a",
          1543 => x"0c815675",
          1544 => x"84bb840c",
          1545 => x"8b3d0d04",
          1546 => x"81701670",
          1547 => x"790c7033",
          1548 => x"56565973",
          1549 => x"b02e0981",
          1550 => x"06feff38",
          1551 => x"81157078",
          1552 => x"0c703355",
          1553 => x"557380e2",
          1554 => x"2ea63890",
          1555 => x"587380f8",
          1556 => x"2ea03881",
          1557 => x"56a07427",
          1558 => x"c638d014",
          1559 => x"53805688",
          1560 => x"58897327",
          1561 => x"fee13875",
          1562 => x"84bb840c",
          1563 => x"8b3d0d04",
          1564 => x"82588115",
          1565 => x"70780c70",
          1566 => x"33555580",
          1567 => x"56feca39",
          1568 => x"800b84bb",
          1569 => x"840c8b3d",
          1570 => x"0d0480d8",
          1571 => x"aa3f84bb",
          1572 => x"840881ff",
          1573 => x"0684bb84",
          1574 => x"0c04ff3d",
          1575 => x"0d735271",
          1576 => x"93268c38",
          1577 => x"71101083",
          1578 => x"bf940552",
          1579 => x"71080483",
          1580 => x"cfac51ef",
          1581 => x"be3f833d",
          1582 => x"0d0483cf",
          1583 => x"bc51efb3",
          1584 => x"3f833d0d",
          1585 => x"0483cfd4",
          1586 => x"51efa83f",
          1587 => x"833d0d04",
          1588 => x"83cfec51",
          1589 => x"ef9d3f83",
          1590 => x"3d0d0483",
          1591 => x"d08451ef",
          1592 => x"923f833d",
          1593 => x"0d0483d0",
          1594 => x"9451ef87",
          1595 => x"3f833d0d",
          1596 => x"0483d0b4",
          1597 => x"51eefc3f",
          1598 => x"833d0d04",
          1599 => x"83d0c451",
          1600 => x"eef13f83",
          1601 => x"3d0d0483",
          1602 => x"d0ec51ee",
          1603 => x"e63f833d",
          1604 => x"0d0483d1",
          1605 => x"8051eedb",
          1606 => x"3f833d0d",
          1607 => x"0483d19c",
          1608 => x"51eed03f",
          1609 => x"833d0d04",
          1610 => x"83d1b451",
          1611 => x"eec53f83",
          1612 => x"3d0d0483",
          1613 => x"d1cc51ee",
          1614 => x"ba3f833d",
          1615 => x"0d0483d1",
          1616 => x"e451eeaf",
          1617 => x"3f833d0d",
          1618 => x"0483d1f4",
          1619 => x"51eea43f",
          1620 => x"833d0d04",
          1621 => x"83d28851",
          1622 => x"ee993f83",
          1623 => x"3d0d0483",
          1624 => x"d29851ee",
          1625 => x"8e3f833d",
          1626 => x"0d0483d2",
          1627 => x"a851ee83",
          1628 => x"3f833d0d",
          1629 => x"0483d2b8",
          1630 => x"51edf83f",
          1631 => x"833d0d04",
          1632 => x"83d2c851",
          1633 => x"eded3f83",
          1634 => x"3d0d0483",
          1635 => x"d2d451ed",
          1636 => x"e23f833d",
          1637 => x"0d04feec",
          1638 => x"3d0d8197",
          1639 => x"3d080284",
          1640 => x"0584e305",
          1641 => x"335b5880",
          1642 => x"0b81993d",
          1643 => x"08793070",
          1644 => x"7b077325",
          1645 => x"51575759",
          1646 => x"78577587",
          1647 => x"ff268338",
          1648 => x"81577477",
          1649 => x"077081ff",
          1650 => x"06515593",
          1651 => x"577480e2",
          1652 => x"38815377",
          1653 => x"528c3d70",
          1654 => x"52588297",
          1655 => x"993f84bb",
          1656 => x"84085784",
          1657 => x"bb840880",
          1658 => x"2e80d138",
          1659 => x"775182af",
          1660 => x"983f7630",
          1661 => x"70780780",
          1662 => x"257b3070",
          1663 => x"9f2a7206",
          1664 => x"53575758",
          1665 => x"77802eaa",
          1666 => x"3887c098",
          1667 => x"88085574",
          1668 => x"87e72680",
          1669 => x"e3387452",
          1670 => x"7887e829",
          1671 => x"51f5863f",
          1672 => x"84bb8408",
          1673 => x"5483d384",
          1674 => x"53785283",
          1675 => x"d2e051df",
          1676 => x"d73f7684",
          1677 => x"bb840c81",
          1678 => x"963d0d04",
          1679 => x"84bb8408",
          1680 => x"87c09888",
          1681 => x"0c84bb84",
          1682 => x"08598196",
          1683 => x"3dfbd405",
          1684 => x"54848053",
          1685 => x"75527751",
          1686 => x"829fea3f",
          1687 => x"84bb8408",
          1688 => x"5784bb84",
          1689 => x"08ff8538",
          1690 => x"7a557480",
          1691 => x"2efefd38",
          1692 => x"74197517",
          1693 => x"5759d339",
          1694 => x"87e85274",
          1695 => x"51f4a63f",
          1696 => x"84bb8408",
          1697 => x"527851f4",
          1698 => x"9c3f84bb",
          1699 => x"84085483",
          1700 => x"d3845378",
          1701 => x"5283d2e0",
          1702 => x"51deed3f",
          1703 => x"ff9439f8",
          1704 => x"3d0d7c02",
          1705 => x"8405b705",
          1706 => x"335859ff",
          1707 => x"5880537b",
          1708 => x"527a51fd",
          1709 => x"e13f84bb",
          1710 => x"84088b38",
          1711 => x"76802e91",
          1712 => x"3876812e",
          1713 => x"8a387784",
          1714 => x"bb840c8a",
          1715 => x"3d0d0478",
          1716 => x"0484e6e4",
          1717 => x"56615560",
          1718 => x"5484bb84",
          1719 => x"537f527e",
          1720 => x"51782d84",
          1721 => x"bb840884",
          1722 => x"bb840c8a",
          1723 => x"3d0d04f3",
          1724 => x"3d0d7f61",
          1725 => x"63028c05",
          1726 => x"80cf0533",
          1727 => x"73731568",
          1728 => x"415f5c5c",
          1729 => x"5f5d5e78",
          1730 => x"802e8382",
          1731 => x"387a5283",
          1732 => x"d38c51dd",
          1733 => x"f33f83d3",
          1734 => x"9451ddec",
          1735 => x"3f805473",
          1736 => x"7927b238",
          1737 => x"7c902e81",
          1738 => x"ed387ca0",
          1739 => x"2e82a838",
          1740 => x"73185372",
          1741 => x"7a2781a7",
          1742 => x"38723352",
          1743 => x"83d39851",
          1744 => x"ddc63f81",
          1745 => x"1484e6e8",
          1746 => x"085354a0",
          1747 => x"51ec9f3f",
          1748 => x"787426dc",
          1749 => x"3883d3a0",
          1750 => x"51ddad3f",
          1751 => x"80567579",
          1752 => x"2780c038",
          1753 => x"75187033",
          1754 => x"55538055",
          1755 => x"727a2783",
          1756 => x"38815580",
          1757 => x"539f7427",
          1758 => x"83388153",
          1759 => x"74730670",
          1760 => x"81ff0656",
          1761 => x"5774802e",
          1762 => x"883880fe",
          1763 => x"742781ee",
          1764 => x"3884e6e8",
          1765 => x"0852a051",
          1766 => x"ebd43f81",
          1767 => x"16567876",
          1768 => x"26c23883",
          1769 => x"d3a451e9",
          1770 => x"ca3f7818",
          1771 => x"791c5c58",
          1772 => x"80519dc8",
          1773 => x"3f84bb84",
          1774 => x"08982b70",
          1775 => x"982c5854",
          1776 => x"76a02e81",
          1777 => x"ee38769b",
          1778 => x"2e82c338",
          1779 => x"7b1e5776",
          1780 => x"7826feb9",
          1781 => x"38ff0b84",
          1782 => x"bb840c8f",
          1783 => x"3d0d0483",
          1784 => x"d3a851dc",
          1785 => x"a33f8114",
          1786 => x"84e6e808",
          1787 => x"5354a051",
          1788 => x"eafc3f78",
          1789 => x"7426feb8",
          1790 => x"38feda39",
          1791 => x"83d3b851",
          1792 => x"dc863f82",
          1793 => x"1484e6e8",
          1794 => x"085354a0",
          1795 => x"51eadf3f",
          1796 => x"737927fe",
          1797 => x"c0387318",
          1798 => x"53727a27",
          1799 => x"df387222",
          1800 => x"5283d3ac",
          1801 => x"51dbe13f",
          1802 => x"821484e6",
          1803 => x"e8085354",
          1804 => x"a051eaba",
          1805 => x"3f787426",
          1806 => x"dd38fe99",
          1807 => x"3983d3b4",
          1808 => x"51dbc53f",
          1809 => x"841484e6",
          1810 => x"e8085354",
          1811 => x"a051ea9e",
          1812 => x"3f737927",
          1813 => x"fdff3873",
          1814 => x"1853727a",
          1815 => x"27df3872",
          1816 => x"085283d3",
          1817 => x"8c51dba0",
          1818 => x"3f841484",
          1819 => x"e6e80853",
          1820 => x"54a051e9",
          1821 => x"f93f7874",
          1822 => x"26dd38fd",
          1823 => x"d83984e6",
          1824 => x"e8085273",
          1825 => x"51e9e73f",
          1826 => x"811656fe",
          1827 => x"913980d0",
          1828 => x"a63f84bb",
          1829 => x"840881ff",
          1830 => x"06538859",
          1831 => x"72a82efc",
          1832 => x"ec38a059",
          1833 => x"7280d02e",
          1834 => x"098106fc",
          1835 => x"e0389059",
          1836 => x"fcdb3980",
          1837 => x"519bc53f",
          1838 => x"84bb8408",
          1839 => x"982b7098",
          1840 => x"2c70a032",
          1841 => x"7030729b",
          1842 => x"32703070",
          1843 => x"72077375",
          1844 => x"07065155",
          1845 => x"58595758",
          1846 => x"53728025",
          1847 => x"fde83880",
          1848 => x"519b993f",
          1849 => x"84bb8408",
          1850 => x"982b7098",
          1851 => x"2c70a032",
          1852 => x"7030729b",
          1853 => x"32703070",
          1854 => x"72077375",
          1855 => x"07065155",
          1856 => x"58595758",
          1857 => x"53807324",
          1858 => x"ffa938fd",
          1859 => x"b939800b",
          1860 => x"84bb840c",
          1861 => x"8f3d0d04",
          1862 => x"fe3d0d87",
          1863 => x"c0968008",
          1864 => x"53aadd3f",
          1865 => x"81519d8d",
          1866 => x"3f83d4d0",
          1867 => x"519d9e3f",
          1868 => x"80519d81",
          1869 => x"3f72812a",
          1870 => x"70810651",
          1871 => x"527182b7",
          1872 => x"3872822a",
          1873 => x"70810651",
          1874 => x"52718289",
          1875 => x"3872832a",
          1876 => x"70810651",
          1877 => x"527181db",
          1878 => x"3872842a",
          1879 => x"70810651",
          1880 => x"527181ad",
          1881 => x"3872852a",
          1882 => x"70810651",
          1883 => x"527180ff",
          1884 => x"3872862a",
          1885 => x"70810651",
          1886 => x"527180d2",
          1887 => x"3872872a",
          1888 => x"70810651",
          1889 => x"5271a938",
          1890 => x"72882a81",
          1891 => x"06537288",
          1892 => x"38a9f53f",
          1893 => x"843d0d04",
          1894 => x"81519c99",
          1895 => x"3f83d4e8",
          1896 => x"519caa3f",
          1897 => x"80519c8d",
          1898 => x"3fa9dd3f",
          1899 => x"843d0d04",
          1900 => x"81519c81",
          1901 => x"3f83d4fc",
          1902 => x"519c923f",
          1903 => x"80519bf5",
          1904 => x"3f72882a",
          1905 => x"81065372",
          1906 => x"802ec638",
          1907 => x"cb398151",
          1908 => x"9be33f83",
          1909 => x"d590519b",
          1910 => x"f43f8051",
          1911 => x"9bd73f72",
          1912 => x"872a7081",
          1913 => x"06515271",
          1914 => x"802eff9c",
          1915 => x"38c23981",
          1916 => x"519bc23f",
          1917 => x"83d5a451",
          1918 => x"9bd33f80",
          1919 => x"519bb63f",
          1920 => x"72862a70",
          1921 => x"81065152",
          1922 => x"71802efe",
          1923 => x"f038ffbe",
          1924 => x"3981519b",
          1925 => x"a03f83d5",
          1926 => x"b8519bb1",
          1927 => x"3f80519b",
          1928 => x"943f7285",
          1929 => x"2a708106",
          1930 => x"51527180",
          1931 => x"2efec238",
          1932 => x"ffbd3981",
          1933 => x"519afe3f",
          1934 => x"83d5cc51",
          1935 => x"9b8f3f80",
          1936 => x"519af23f",
          1937 => x"72842a70",
          1938 => x"81065152",
          1939 => x"71802efe",
          1940 => x"9438ffbd",
          1941 => x"3981519a",
          1942 => x"dc3f83d5",
          1943 => x"e0519aed",
          1944 => x"3f80519a",
          1945 => x"d03f7283",
          1946 => x"2a708106",
          1947 => x"51527180",
          1948 => x"2efde638",
          1949 => x"ffbd3981",
          1950 => x"519aba3f",
          1951 => x"83d5f051",
          1952 => x"9acb3f80",
          1953 => x"519aae3f",
          1954 => x"72822a70",
          1955 => x"81065152",
          1956 => x"71802efd",
          1957 => x"b838ffbd",
          1958 => x"39ca3d0d",
          1959 => x"80704141",
          1960 => x"ff6184de",
          1961 => x"900c4281",
          1962 => x"52605181",
          1963 => x"b7c93f84",
          1964 => x"bb840881",
          1965 => x"ff069b3d",
          1966 => x"40597861",
          1967 => x"2e84b538",
          1968 => x"83d6c451",
          1969 => x"e3ad3f98",
          1970 => x"3d4383d6",
          1971 => x"fc51d6b8",
          1972 => x"3f7e4880",
          1973 => x"f8538052",
          1974 => x"7e51eba3",
          1975 => x"3f0b0b83",
          1976 => x"eff83370",
          1977 => x"81ff065b",
          1978 => x"5979802e",
          1979 => x"82f13879",
          1980 => x"812e8388",
          1981 => x"387881ff",
          1982 => x"065e7d82",
          1983 => x"2e83c138",
          1984 => x"67705a5a",
          1985 => x"79802e83",
          1986 => x"e0387933",
          1987 => x"5c7ba02e",
          1988 => x"0981068c",
          1989 => x"38811a70",
          1990 => x"335d5a7b",
          1991 => x"a02ef638",
          1992 => x"805c7b9b",
          1993 => x"26be387b",
          1994 => x"902983ef",
          1995 => x"fc057008",
          1996 => x"525be7f4",
          1997 => x"3f84bb84",
          1998 => x"0884bb84",
          1999 => x"08547a53",
          2000 => x"7b08525d",
          2001 => x"e8cf3f84",
          2002 => x"bb84088b",
          2003 => x"38841b33",
          2004 => x"5e7d812e",
          2005 => x"83843881",
          2006 => x"1c7081ff",
          2007 => x"065d5b9b",
          2008 => x"7c27c438",
          2009 => x"9a3d335c",
          2010 => x"7b802efe",
          2011 => x"dd3880f8",
          2012 => x"527e51e9",
          2013 => x"873f84bb",
          2014 => x"84085e84",
          2015 => x"bb840880",
          2016 => x"2e8dce38",
          2017 => x"84bb8408",
          2018 => x"48b83dff",
          2019 => x"80055191",
          2020 => x"a93f84bb",
          2021 => x"84086062",
          2022 => x"065c5c7a",
          2023 => x"802e8184",
          2024 => x"3884bb84",
          2025 => x"0851e780",
          2026 => x"3f84bb84",
          2027 => x"088f2680",
          2028 => x"f338810b",
          2029 => x"a53d5e5b",
          2030 => x"7a822e8d",
          2031 => x"8a387a82",
          2032 => x"248ce738",
          2033 => x"7a812e82",
          2034 => x"e8387b54",
          2035 => x"805383d7",
          2036 => x"80527c51",
          2037 => x"d5d23f83",
          2038 => x"f3c05884",
          2039 => x"bbb4577d",
          2040 => x"56675580",
          2041 => x"5490800a",
          2042 => x"5390800a",
          2043 => x"527c51f5",
          2044 => x"ae3f84bb",
          2045 => x"840884bb",
          2046 => x"84080970",
          2047 => x"30707207",
          2048 => x"8025515b",
          2049 => x"5b42805a",
          2050 => x"7a832683",
          2051 => x"38815a78",
          2052 => x"7a065978",
          2053 => x"802e8d38",
          2054 => x"811b7081",
          2055 => x"ff065c5a",
          2056 => x"7aff9538",
          2057 => x"7f813261",
          2058 => x"8132075d",
          2059 => x"7c81f238",
          2060 => x"61ff2e81",
          2061 => x"ec387d51",
          2062 => x"81969e3f",
          2063 => x"83d6fc51",
          2064 => x"d3c63f7e",
          2065 => x"4880f853",
          2066 => x"80527e51",
          2067 => x"e8b13f0b",
          2068 => x"0b83eff8",
          2069 => x"337081ff",
          2070 => x"065b5979",
          2071 => x"fd913881",
          2072 => x"5383d6a8",
          2073 => x"5284de94",
          2074 => x"51828a8a",
          2075 => x"3f84bb84",
          2076 => x"0880c538",
          2077 => x"810b0b0b",
          2078 => x"83eff834",
          2079 => x"84de9453",
          2080 => x"80f8527e",
          2081 => x"5182f7cc",
          2082 => x"3f84bb84",
          2083 => x"08802ea0",
          2084 => x"3884bb84",
          2085 => x"0851dfdb",
          2086 => x"3f0b0b83",
          2087 => x"eff83370",
          2088 => x"81ff065f",
          2089 => x"597d822e",
          2090 => x"098106fc",
          2091 => x"d3389139",
          2092 => x"84de9451",
          2093 => x"82a1d23f",
          2094 => x"820b0b0b",
          2095 => x"83eff834",
          2096 => x"805583d6",
          2097 => x"b8548053",
          2098 => x"80f8527e",
          2099 => x"51a7d73f",
          2100 => x"67705a5a",
          2101 => x"79fcb338",
          2102 => x"90397c1a",
          2103 => x"630c851b",
          2104 => x"33597881",
          2105 => x"8926fcfc",
          2106 => x"38781010",
          2107 => x"83bfe405",
          2108 => x"5a790804",
          2109 => x"835383d7",
          2110 => x"88527e51",
          2111 => x"e4ec3f60",
          2112 => x"537e5284",
          2113 => x"c8b05182",
          2114 => x"86bd3f84",
          2115 => x"bb840861",
          2116 => x"2e098106",
          2117 => x"fbaa3881",
          2118 => x"709a3d45",
          2119 => x"4141fbaa",
          2120 => x"3983d78c",
          2121 => x"51decc3f",
          2122 => x"7d518194",
          2123 => x"ac3ffe8c",
          2124 => x"3983d79c",
          2125 => x"567b5583",
          2126 => x"d7a05480",
          2127 => x"5383d7a4",
          2128 => x"527c51d2",
          2129 => x"e33ffd8f",
          2130 => x"39818de4",
          2131 => x"3ffafb39",
          2132 => x"9af93ffa",
          2133 => x"f5398152",
          2134 => x"835180c0",
          2135 => x"dc3ffaea",
          2136 => x"39818f8e",
          2137 => x"3ffae339",
          2138 => x"83d7b451",
          2139 => x"de853f80",
          2140 => x"59780483",
          2141 => x"d7c851dd",
          2142 => x"fa3fd0ed",
          2143 => x"3ffacb39",
          2144 => x"b83dff84",
          2145 => x"1153ff80",
          2146 => x"0551ebfa",
          2147 => x"3f84bb84",
          2148 => x"08802efa",
          2149 => x"b5386852",
          2150 => x"83d7e451",
          2151 => x"d0ea3f68",
          2152 => x"5a792d84",
          2153 => x"bb840880",
          2154 => x"2efa9f38",
          2155 => x"84bb8408",
          2156 => x"5283d880",
          2157 => x"51d0d13f",
          2158 => x"fa9039b8",
          2159 => x"3dff8411",
          2160 => x"53ff8005",
          2161 => x"51ebbf3f",
          2162 => x"84bb8408",
          2163 => x"802ef9fa",
          2164 => x"38685283",
          2165 => x"d89c51d0",
          2166 => x"af3f6859",
          2167 => x"7804b83d",
          2168 => x"fef41153",
          2169 => x"ff800551",
          2170 => x"e9983f84",
          2171 => x"bb840880",
          2172 => x"2ef9d738",
          2173 => x"b83dfef0",
          2174 => x"1153ff80",
          2175 => x"0551e982",
          2176 => x"3f84bb84",
          2177 => x"0886d038",
          2178 => x"64597808",
          2179 => x"53785283",
          2180 => x"d8b851cf",
          2181 => x"f33f84e6",
          2182 => x"e4085380",
          2183 => x"f8527e51",
          2184 => x"d0813f7e",
          2185 => x"487e3359",
          2186 => x"78ae2ef9",
          2187 => x"9d38789f",
          2188 => x"2687d338",
          2189 => x"64840570",
          2190 => x"4659cf39",
          2191 => x"b83dfef4",
          2192 => x"1153ff80",
          2193 => x"0551e8ba",
          2194 => x"3f84bb84",
          2195 => x"08802ef8",
          2196 => x"f938b83d",
          2197 => x"fef01153",
          2198 => x"ff800551",
          2199 => x"e8a43f84",
          2200 => x"bb840886",
          2201 => x"b0386459",
          2202 => x"78225378",
          2203 => x"5283d8c8",
          2204 => x"51cf953f",
          2205 => x"84e6e408",
          2206 => x"5380f852",
          2207 => x"7e51cfa3",
          2208 => x"3f7e487e",
          2209 => x"335978ae",
          2210 => x"2ef8bf38",
          2211 => x"789f2687",
          2212 => x"ca386482",
          2213 => x"05704659",
          2214 => x"cf39b83d",
          2215 => x"ff841153",
          2216 => x"ff800551",
          2217 => x"e9e03f84",
          2218 => x"bb840880",
          2219 => x"2ef89b38",
          2220 => x"b83dfefc",
          2221 => x"1153ff80",
          2222 => x"0551e9ca",
          2223 => x"3f84bb84",
          2224 => x"08802ef8",
          2225 => x"8538b83d",
          2226 => x"fef81153",
          2227 => x"ff800551",
          2228 => x"e9b43f84",
          2229 => x"bb840880",
          2230 => x"2ef7ef38",
          2231 => x"83d8d451",
          2232 => x"cea63f68",
          2233 => x"675d5978",
          2234 => x"7c27838d",
          2235 => x"38657033",
          2236 => x"7a335f5c",
          2237 => x"5a7a7d2e",
          2238 => x"95387a55",
          2239 => x"79547833",
          2240 => x"53785283",
          2241 => x"d8e451cd",
          2242 => x"ff3f6666",
          2243 => x"5b5c8119",
          2244 => x"811b4759",
          2245 => x"d239b83d",
          2246 => x"ff841153",
          2247 => x"ff800551",
          2248 => x"e8e43f84",
          2249 => x"bb840880",
          2250 => x"2ef79f38",
          2251 => x"b83dfefc",
          2252 => x"1153ff80",
          2253 => x"0551e8ce",
          2254 => x"3f84bb84",
          2255 => x"08802ef7",
          2256 => x"8938b83d",
          2257 => x"fef81153",
          2258 => x"ff800551",
          2259 => x"e8b83f84",
          2260 => x"bb840880",
          2261 => x"2ef6f338",
          2262 => x"83d98051",
          2263 => x"cdaa3f68",
          2264 => x"5a796727",
          2265 => x"82933865",
          2266 => x"5c797081",
          2267 => x"055b337c",
          2268 => x"34658105",
          2269 => x"46eb39b8",
          2270 => x"3dff8411",
          2271 => x"53ff8005",
          2272 => x"51e8833f",
          2273 => x"84bb8408",
          2274 => x"802ef6be",
          2275 => x"38b83dfe",
          2276 => x"fc1153ff",
          2277 => x"800551e7",
          2278 => x"ed3f84bb",
          2279 => x"8408b138",
          2280 => x"68703354",
          2281 => x"5283d98c",
          2282 => x"51ccdd3f",
          2283 => x"84e6e408",
          2284 => x"5380f852",
          2285 => x"7e51cceb",
          2286 => x"3f7e487e",
          2287 => x"335978ae",
          2288 => x"2ef68738",
          2289 => x"789f2684",
          2290 => x"97386881",
          2291 => x"0549d139",
          2292 => x"68590280",
          2293 => x"db053379",
          2294 => x"34688105",
          2295 => x"49b83dfe",
          2296 => x"fc1153ff",
          2297 => x"800551e7",
          2298 => x"9d3f84bb",
          2299 => x"8408802e",
          2300 => x"f5d83868",
          2301 => x"590280db",
          2302 => x"05337934",
          2303 => x"68810549",
          2304 => x"b83dfefc",
          2305 => x"1153ff80",
          2306 => x"0551e6fa",
          2307 => x"3f84bb84",
          2308 => x"08ffbd38",
          2309 => x"f5b439b8",
          2310 => x"3dff8411",
          2311 => x"53ff8005",
          2312 => x"51e6e33f",
          2313 => x"84bb8408",
          2314 => x"802ef59e",
          2315 => x"38b83dfe",
          2316 => x"fc1153ff",
          2317 => x"800551e6",
          2318 => x"cd3f84bb",
          2319 => x"8408802e",
          2320 => x"f58838b8",
          2321 => x"3dfef811",
          2322 => x"53ff8005",
          2323 => x"51e6b73f",
          2324 => x"84bb8408",
          2325 => x"863884bb",
          2326 => x"84084683",
          2327 => x"d99851cb",
          2328 => x"a73f6867",
          2329 => x"5b59787a",
          2330 => x"278f3865",
          2331 => x"5b7a7970",
          2332 => x"84055b0c",
          2333 => x"797926f5",
          2334 => x"388a51d9",
          2335 => x"e13ff4ca",
          2336 => x"39b83dff",
          2337 => x"80055187",
          2338 => x"b13f84bb",
          2339 => x"8408b93d",
          2340 => x"ff800552",
          2341 => x"5988f33f",
          2342 => x"815384bb",
          2343 => x"84085278",
          2344 => x"51e9f33f",
          2345 => x"84bb8408",
          2346 => x"802ef49e",
          2347 => x"3884bb84",
          2348 => x"0851e7e6",
          2349 => x"3ff49339",
          2350 => x"b83dff84",
          2351 => x"1153ff80",
          2352 => x"0551e5c2",
          2353 => x"3f84bb84",
          2354 => x"08913883",
          2355 => x"f488335a",
          2356 => x"79802e83",
          2357 => x"c03883f3",
          2358 => x"c00849b8",
          2359 => x"3dfefc11",
          2360 => x"53ff8005",
          2361 => x"51e59f3f",
          2362 => x"84bb8408",
          2363 => x"913883f4",
          2364 => x"88335a79",
          2365 => x"802e838a",
          2366 => x"3883f3c4",
          2367 => x"0847b83d",
          2368 => x"fef81153",
          2369 => x"ff800551",
          2370 => x"e4fc3f84",
          2371 => x"bb840880",
          2372 => x"2ea53880",
          2373 => x"665c5c7a",
          2374 => x"882e8338",
          2375 => x"815c7a90",
          2376 => x"32703070",
          2377 => x"72079f2a",
          2378 => x"7e065c5f",
          2379 => x"5d79802e",
          2380 => x"88387aa0",
          2381 => x"2e833888",
          2382 => x"4683d9a8",
          2383 => x"51d6b43f",
          2384 => x"80556854",
          2385 => x"65536652",
          2386 => x"6851eba3",
          2387 => x"3f83d9b4",
          2388 => x"51d6a03f",
          2389 => x"f2f43964",
          2390 => x"64710c59",
          2391 => x"64840545",
          2392 => x"b83dfef0",
          2393 => x"1153ff80",
          2394 => x"0551e296",
          2395 => x"3f84bb84",
          2396 => x"08802ef2",
          2397 => x"d5386464",
          2398 => x"710c5964",
          2399 => x"840545b8",
          2400 => x"3dfef011",
          2401 => x"53ff8005",
          2402 => x"51e1f73f",
          2403 => x"84bb8408",
          2404 => x"c638f2b6",
          2405 => x"39645e02",
          2406 => x"80ce0522",
          2407 => x"7e708205",
          2408 => x"40237d45",
          2409 => x"b83dfef0",
          2410 => x"1153ff80",
          2411 => x"0551e1d2",
          2412 => x"3f84bb84",
          2413 => x"08802ef2",
          2414 => x"9138645e",
          2415 => x"0280ce05",
          2416 => x"227e7082",
          2417 => x"0540237d",
          2418 => x"45b83dfe",
          2419 => x"f01153ff",
          2420 => x"800551e1",
          2421 => x"ad3f84bb",
          2422 => x"8408ffb9",
          2423 => x"38f1eb39",
          2424 => x"b83dfefc",
          2425 => x"1153ff80",
          2426 => x"0551e39a",
          2427 => x"3f84bb84",
          2428 => x"08802e81",
          2429 => x"dc38685c",
          2430 => x"0280db05",
          2431 => x"337c3468",
          2432 => x"810549fb",
          2433 => x"9b39b83d",
          2434 => x"fef01153",
          2435 => x"ff800551",
          2436 => x"e0f03f84",
          2437 => x"bb840880",
          2438 => x"2e819838",
          2439 => x"6464710c",
          2440 => x"5d648405",
          2441 => x"704659f7",
          2442 => x"e1397a83",
          2443 => x"2e098106",
          2444 => x"f398387b",
          2445 => x"5583d7a0",
          2446 => x"54805383",
          2447 => x"d9c0527c",
          2448 => x"51c8e53f",
          2449 => x"f391397b",
          2450 => x"527c51d9",
          2451 => x"fa3ff387",
          2452 => x"3983d9cc",
          2453 => x"51d49c3f",
          2454 => x"f0f039b8",
          2455 => x"3dfef011",
          2456 => x"53ff8005",
          2457 => x"51e09b3f",
          2458 => x"84bb8408",
          2459 => x"802eb838",
          2460 => x"64590280",
          2461 => x"ce052279",
          2462 => x"7082055b",
          2463 => x"237845f7",
          2464 => x"e73983f4",
          2465 => x"89335c7b",
          2466 => x"802e80cf",
          2467 => x"3883f3cc",
          2468 => x"0847fcea",
          2469 => x"3983f489",
          2470 => x"335c7b80",
          2471 => x"2ea13883",
          2472 => x"f3c80849",
          2473 => x"fcb53983",
          2474 => x"d9f851d3",
          2475 => x"c63f6459",
          2476 => x"f7b63983",
          2477 => x"d9f851d3",
          2478 => x"ba3f6459",
          2479 => x"f6cc3983",
          2480 => x"f48a3359",
          2481 => x"78802ea5",
          2482 => x"3883f3d0",
          2483 => x"0849fc8b",
          2484 => x"3983d9f8",
          2485 => x"51d39c3f",
          2486 => x"f9c63983",
          2487 => x"f48a3359",
          2488 => x"78802e9b",
          2489 => x"3883f3d4",
          2490 => x"0847fc92",
          2491 => x"3983f48b",
          2492 => x"335e7d80",
          2493 => x"2e9b3883",
          2494 => x"f3d80849",
          2495 => x"fbdd3983",
          2496 => x"f48b335e",
          2497 => x"7d802e9b",
          2498 => x"3883f3dc",
          2499 => x"0847fbee",
          2500 => x"3983f486",
          2501 => x"335d7c80",
          2502 => x"2e9b3883",
          2503 => x"f3e00849",
          2504 => x"fbb93983",
          2505 => x"f486335d",
          2506 => x"7c802e94",
          2507 => x"3883f3e4",
          2508 => x"0847fbca",
          2509 => x"3983f3f0",
          2510 => x"08fc8005",
          2511 => x"49fb9c39",
          2512 => x"83f3f008",
          2513 => x"880547fb",
          2514 => x"b539f33d",
          2515 => x"0d800b84",
          2516 => x"bbb43487",
          2517 => x"c0948c70",
          2518 => x"08565787",
          2519 => x"84805274",
          2520 => x"51dac23f",
          2521 => x"84bb8408",
          2522 => x"902b7708",
          2523 => x"57558784",
          2524 => x"80527551",
          2525 => x"daaf3f74",
          2526 => x"84bb8408",
          2527 => x"07770c87",
          2528 => x"c0949c70",
          2529 => x"08565787",
          2530 => x"84805274",
          2531 => x"51da963f",
          2532 => x"84bb8408",
          2533 => x"902b7708",
          2534 => x"57558784",
          2535 => x"80527551",
          2536 => x"da833f74",
          2537 => x"84bb8408",
          2538 => x"07770c8c",
          2539 => x"80830b87",
          2540 => x"c094840c",
          2541 => x"8c80830b",
          2542 => x"87c09494",
          2543 => x"0c81beba",
          2544 => x"5c81c9b9",
          2545 => x"5d830284",
          2546 => x"05a10534",
          2547 => x"805e84e6",
          2548 => x"e40b893d",
          2549 => x"7088130c",
          2550 => x"70720c84",
          2551 => x"e6e80c56",
          2552 => x"b8bd3f89",
          2553 => x"9e3f9598",
          2554 => x"3fba9851",
          2555 => x"958d3f83",
          2556 => x"d3c05283",
          2557 => x"d3c451c4",
          2558 => x"8f3f83f3",
          2559 => x"f4702252",
          2560 => x"5594983f",
          2561 => x"83d3cc54",
          2562 => x"83d3d853",
          2563 => x"81153352",
          2564 => x"83d3e051",
          2565 => x"c3f23f8d",
          2566 => x"b23f83d3",
          2567 => x"fc51d0d3",
          2568 => x"3f805283",
          2569 => x"d48051c3",
          2570 => x"df3f9080",
          2571 => x"0a5283d4",
          2572 => x"a851c3d4",
          2573 => x"3fece23f",
          2574 => x"8004fb3d",
          2575 => x"0d777008",
          2576 => x"56568075",
          2577 => x"52537473",
          2578 => x"2e818338",
          2579 => x"74337081",
          2580 => x"ff065252",
          2581 => x"70a02e09",
          2582 => x"81069138",
          2583 => x"81157033",
          2584 => x"7081ff06",
          2585 => x"53535570",
          2586 => x"a02ef138",
          2587 => x"7181ff06",
          2588 => x"5473a22e",
          2589 => x"81823874",
          2590 => x"5272812e",
          2591 => x"80e73880",
          2592 => x"72337081",
          2593 => x"ff065354",
          2594 => x"5470a02e",
          2595 => x"83388154",
          2596 => x"70802e8b",
          2597 => x"3873802e",
          2598 => x"86388112",
          2599 => x"52e13980",
          2600 => x"7381ff06",
          2601 => x"525470a0",
          2602 => x"2e098106",
          2603 => x"83388154",
          2604 => x"70a23270",
          2605 => x"30708025",
          2606 => x"76075252",
          2607 => x"5372802e",
          2608 => x"88388072",
          2609 => x"70810554",
          2610 => x"3471760c",
          2611 => x"74517084",
          2612 => x"bb840c87",
          2613 => x"3d0d0470",
          2614 => x"802ec438",
          2615 => x"73802eff",
          2616 => x"be388112",
          2617 => x"52807233",
          2618 => x"7081ff06",
          2619 => x"53545470",
          2620 => x"a22ee438",
          2621 => x"8154e039",
          2622 => x"81155581",
          2623 => x"75535372",
          2624 => x"812e0981",
          2625 => x"06fef838",
          2626 => x"dc39fc3d",
          2627 => x"0d765372",
          2628 => x"088b3880",
          2629 => x"0b84bb84",
          2630 => x"0c863d0d",
          2631 => x"04863dfc",
          2632 => x"05527251",
          2633 => x"dadc3f84",
          2634 => x"bb840880",
          2635 => x"2ee53874",
          2636 => x"84bb840c",
          2637 => x"863d0d04",
          2638 => x"fc3d0d76",
          2639 => x"821133ff",
          2640 => x"05525381",
          2641 => x"52708b26",
          2642 => x"81983883",
          2643 => x"1333ff05",
          2644 => x"54825273",
          2645 => x"9e26818a",
          2646 => x"38841333",
          2647 => x"51835270",
          2648 => x"972680fe",
          2649 => x"38851333",
          2650 => x"54845273",
          2651 => x"bb2680f2",
          2652 => x"38861333",
          2653 => x"55855274",
          2654 => x"bb2680e6",
          2655 => x"38881322",
          2656 => x"55865274",
          2657 => x"87e72680",
          2658 => x"d9388a13",
          2659 => x"22548752",
          2660 => x"7387e726",
          2661 => x"80cc3881",
          2662 => x"0b87c098",
          2663 => x"9c0c7222",
          2664 => x"87c098bc",
          2665 => x"0c821333",
          2666 => x"87c098b8",
          2667 => x"0c831333",
          2668 => x"87c098b4",
          2669 => x"0c841333",
          2670 => x"87c098b0",
          2671 => x"0c851333",
          2672 => x"87c098ac",
          2673 => x"0c861333",
          2674 => x"87c098a8",
          2675 => x"0c7487c0",
          2676 => x"98a40c73",
          2677 => x"87c098a0",
          2678 => x"0c800b87",
          2679 => x"c0989c0c",
          2680 => x"80527184",
          2681 => x"bb840c86",
          2682 => x"3d0d04f3",
          2683 => x"3d0d7f5b",
          2684 => x"87c0989c",
          2685 => x"5d817d0c",
          2686 => x"87c098bc",
          2687 => x"085e7d7b",
          2688 => x"2387c098",
          2689 => x"b8085c7b",
          2690 => x"821c3487",
          2691 => x"c098b408",
          2692 => x"5a79831c",
          2693 => x"3487c098",
          2694 => x"b0085c7b",
          2695 => x"841c3487",
          2696 => x"c098ac08",
          2697 => x"5a79851c",
          2698 => x"3487c098",
          2699 => x"a8085c7b",
          2700 => x"861c3487",
          2701 => x"c098a408",
          2702 => x"5c7b881c",
          2703 => x"2387c098",
          2704 => x"a0085a79",
          2705 => x"8a1c2380",
          2706 => x"7d0c7983",
          2707 => x"ffff0659",
          2708 => x"7b83ffff",
          2709 => x"0658861b",
          2710 => x"3357851b",
          2711 => x"3356841b",
          2712 => x"3355831b",
          2713 => x"3354821b",
          2714 => x"33537d83",
          2715 => x"ffff0652",
          2716 => x"83d9fc51",
          2717 => x"ffbf913f",
          2718 => x"8f3d0d04",
          2719 => x"fe3d0d02",
          2720 => x"93053353",
          2721 => x"72812ea8",
          2722 => x"38725180",
          2723 => x"e9de3f84",
          2724 => x"bb840898",
          2725 => x"2b70982c",
          2726 => x"515271ff",
          2727 => x"2e098106",
          2728 => x"86387283",
          2729 => x"2ee33871",
          2730 => x"84bb840c",
          2731 => x"843d0d04",
          2732 => x"725180e9",
          2733 => x"b73f84bb",
          2734 => x"8408982b",
          2735 => x"70982c51",
          2736 => x"5271ff2e",
          2737 => x"098106df",
          2738 => x"38725180",
          2739 => x"e99e3f84",
          2740 => x"bb840898",
          2741 => x"2b70982c",
          2742 => x"515271ff",
          2743 => x"2ed238c7",
          2744 => x"39fd3d0d",
          2745 => x"80705452",
          2746 => x"71882b54",
          2747 => x"815180e8",
          2748 => x"fb3f84bb",
          2749 => x"8408982b",
          2750 => x"70982c51",
          2751 => x"5271ff2e",
          2752 => x"eb387372",
          2753 => x"07811454",
          2754 => x"52837325",
          2755 => x"db387184",
          2756 => x"bb840c85",
          2757 => x"3d0d04fc",
          2758 => x"3d0d029b",
          2759 => x"053383f3",
          2760 => x"bc337081",
          2761 => x"ff065355",
          2762 => x"5570802e",
          2763 => x"80f43887",
          2764 => x"c0949408",
          2765 => x"70962a70",
          2766 => x"81065354",
          2767 => x"5270802e",
          2768 => x"8c387191",
          2769 => x"2a708106",
          2770 => x"515170e3",
          2771 => x"38728132",
          2772 => x"81065372",
          2773 => x"802e8a38",
          2774 => x"71932a81",
          2775 => x"065271cf",
          2776 => x"387381ff",
          2777 => x"065187c0",
          2778 => x"94805270",
          2779 => x"802e8638",
          2780 => x"87c09490",
          2781 => x"5274720c",
          2782 => x"7484bb84",
          2783 => x"0c863d0d",
          2784 => x"0471912a",
          2785 => x"70810651",
          2786 => x"51709738",
          2787 => x"72813281",
          2788 => x"06537280",
          2789 => x"2ecb3871",
          2790 => x"932a8106",
          2791 => x"5271802e",
          2792 => x"c03887c0",
          2793 => x"94840870",
          2794 => x"962a7081",
          2795 => x"06535452",
          2796 => x"70cf38d8",
          2797 => x"39ff3d0d",
          2798 => x"028f0533",
          2799 => x"7030709f",
          2800 => x"2a515252",
          2801 => x"7083f3bc",
          2802 => x"34833d0d",
          2803 => x"04fa3d0d",
          2804 => x"78558075",
          2805 => x"33705652",
          2806 => x"5770772e",
          2807 => x"80e73881",
          2808 => x"1583f3bc",
          2809 => x"337081ff",
          2810 => x"06545755",
          2811 => x"71802e80",
          2812 => x"ff3887c0",
          2813 => x"94940870",
          2814 => x"962a7081",
          2815 => x"06535452",
          2816 => x"70802e8c",
          2817 => x"3871912a",
          2818 => x"70810651",
          2819 => x"5170e338",
          2820 => x"72813281",
          2821 => x"06537280",
          2822 => x"2e8a3871",
          2823 => x"932a8106",
          2824 => x"5271cf38",
          2825 => x"7581ff06",
          2826 => x"5187c094",
          2827 => x"80527080",
          2828 => x"2e863887",
          2829 => x"c0949052",
          2830 => x"73720c81",
          2831 => x"17753355",
          2832 => x"5773ff9b",
          2833 => x"387684bb",
          2834 => x"840c883d",
          2835 => x"0d047191",
          2836 => x"2a708106",
          2837 => x"51517098",
          2838 => x"38728132",
          2839 => x"81065372",
          2840 => x"802ec138",
          2841 => x"71932a81",
          2842 => x"06527180",
          2843 => x"2effb538",
          2844 => x"87c09484",
          2845 => x"0870962a",
          2846 => x"70810653",
          2847 => x"545270ce",
          2848 => x"38d739ff",
          2849 => x"3d0d87c0",
          2850 => x"9e800870",
          2851 => x"9c2a8a06",
          2852 => x"52527080",
          2853 => x"2e84ab38",
          2854 => x"87c09ea4",
          2855 => x"0883f3c0",
          2856 => x"0c87c09e",
          2857 => x"a80883f3",
          2858 => x"c40c87c0",
          2859 => x"9e940883",
          2860 => x"f3c80c87",
          2861 => x"c09e9808",
          2862 => x"83f3cc0c",
          2863 => x"87c09e9c",
          2864 => x"0883f3d0",
          2865 => x"0c87c09e",
          2866 => x"a00883f3",
          2867 => x"d40c87c0",
          2868 => x"9eac0883",
          2869 => x"f3d80c87",
          2870 => x"c09eb008",
          2871 => x"83f3dc0c",
          2872 => x"87c09eb4",
          2873 => x"0883f3e0",
          2874 => x"0c87c09e",
          2875 => x"b80883f3",
          2876 => x"e40c87c0",
          2877 => x"9ebc0883",
          2878 => x"f3e80c87",
          2879 => x"c09ec008",
          2880 => x"83f3ec0c",
          2881 => x"87c09ec4",
          2882 => x"0883f3f0",
          2883 => x"0c87c09e",
          2884 => x"80085271",
          2885 => x"83f3f423",
          2886 => x"87c09e84",
          2887 => x"0883f3f8",
          2888 => x"0c87c09e",
          2889 => x"880883f3",
          2890 => x"fc0c87c0",
          2891 => x"9e8c0883",
          2892 => x"f4800c81",
          2893 => x"0b83f484",
          2894 => x"34800b87",
          2895 => x"c09e9008",
          2896 => x"7084800a",
          2897 => x"06515252",
          2898 => x"7082fb38",
          2899 => x"7183f485",
          2900 => x"34800b87",
          2901 => x"c09e9008",
          2902 => x"7088800a",
          2903 => x"06515252",
          2904 => x"70802e83",
          2905 => x"38815271",
          2906 => x"83f48634",
          2907 => x"800b87c0",
          2908 => x"9e900870",
          2909 => x"90800a06",
          2910 => x"51525270",
          2911 => x"802e8338",
          2912 => x"81527183",
          2913 => x"f4873480",
          2914 => x"0b87c09e",
          2915 => x"90087088",
          2916 => x"80800651",
          2917 => x"52527080",
          2918 => x"2e833881",
          2919 => x"527183f4",
          2920 => x"8834800b",
          2921 => x"87c09e90",
          2922 => x"0870a080",
          2923 => x"80065152",
          2924 => x"5270802e",
          2925 => x"83388152",
          2926 => x"7183f489",
          2927 => x"34800b87",
          2928 => x"c09e9008",
          2929 => x"70908080",
          2930 => x"06515252",
          2931 => x"70802e83",
          2932 => x"38815271",
          2933 => x"83f48a34",
          2934 => x"800b87c0",
          2935 => x"9e900870",
          2936 => x"84808006",
          2937 => x"51525270",
          2938 => x"802e8338",
          2939 => x"81527183",
          2940 => x"f48b3480",
          2941 => x"0b87c09e",
          2942 => x"90087082",
          2943 => x"80800651",
          2944 => x"52527080",
          2945 => x"2e833881",
          2946 => x"527183f4",
          2947 => x"8c34800b",
          2948 => x"87c09e90",
          2949 => x"08708180",
          2950 => x"80065152",
          2951 => x"5270802e",
          2952 => x"83388152",
          2953 => x"7183f48d",
          2954 => x"34800b87",
          2955 => x"c09e9008",
          2956 => x"7080c080",
          2957 => x"06515252",
          2958 => x"70802e83",
          2959 => x"38815271",
          2960 => x"83f48e34",
          2961 => x"800b87c0",
          2962 => x"9e900870",
          2963 => x"a0800651",
          2964 => x"52527080",
          2965 => x"2e833881",
          2966 => x"527183f4",
          2967 => x"8f3487c0",
          2968 => x"9e900898",
          2969 => x"8006708a",
          2970 => x"2a535171",
          2971 => x"83f49034",
          2972 => x"800b87c0",
          2973 => x"9e900870",
          2974 => x"84800651",
          2975 => x"52527080",
          2976 => x"2e833881",
          2977 => x"527183f4",
          2978 => x"913487c0",
          2979 => x"9e900883",
          2980 => x"f0067084",
          2981 => x"2a535171",
          2982 => x"83f49234",
          2983 => x"800b87c0",
          2984 => x"9e900870",
          2985 => x"88065152",
          2986 => x"5270802e",
          2987 => x"83388152",
          2988 => x"7183f493",
          2989 => x"3487c09e",
          2990 => x"90088706",
          2991 => x"517083f4",
          2992 => x"9434833d",
          2993 => x"0d048152",
          2994 => x"fd8239fb",
          2995 => x"3d0d83da",
          2996 => x"9451ffb6",
          2997 => x"b33f83f4",
          2998 => x"84335473",
          2999 => x"86a03883",
          3000 => x"daa851c3",
          3001 => x"8e3f83f4",
          3002 => x"86335574",
          3003 => x"85f03883",
          3004 => x"f48b3354",
          3005 => x"7385c738",
          3006 => x"83f48833",
          3007 => x"5675859e",
          3008 => x"3883f489",
          3009 => x"33557484",
          3010 => x"f53883f4",
          3011 => x"8a335473",
          3012 => x"84cc3883",
          3013 => x"f48f3356",
          3014 => x"7584a938",
          3015 => x"83f49333",
          3016 => x"54738486",
          3017 => x"3883f491",
          3018 => x"33557483",
          3019 => x"e33883f4",
          3020 => x"85335675",
          3021 => x"83c53883",
          3022 => x"f4873354",
          3023 => x"7383a738",
          3024 => x"83f48c33",
          3025 => x"55748389",
          3026 => x"3883f48d",
          3027 => x"33567582",
          3028 => x"ea3883f4",
          3029 => x"8e335473",
          3030 => x"81e13883",
          3031 => x"dac051c2",
          3032 => x"923f83f3",
          3033 => x"e8085283",
          3034 => x"dacc51ff",
          3035 => x"b59a3f83",
          3036 => x"f3ec0852",
          3037 => x"83daf451",
          3038 => x"ffb58d3f",
          3039 => x"83f3f008",
          3040 => x"5283db9c",
          3041 => x"51ffb580",
          3042 => x"3f83dbc4",
          3043 => x"51c1e43f",
          3044 => x"83f3f422",
          3045 => x"5283dbcc",
          3046 => x"51ffb4ec",
          3047 => x"3f83f3f8",
          3048 => x"0856bd84",
          3049 => x"c0527551",
          3050 => x"c9fb3f84",
          3051 => x"bb8408bd",
          3052 => x"84c02976",
          3053 => x"71315454",
          3054 => x"84bb8408",
          3055 => x"5283dbf4",
          3056 => x"51ffb4c4",
          3057 => x"3f83f48b",
          3058 => x"335574b9",
          3059 => x"3883f486",
          3060 => x"33557485",
          3061 => x"38873d0d",
          3062 => x"0483f480",
          3063 => x"0856bd84",
          3064 => x"c0527551",
          3065 => x"c9bf3f84",
          3066 => x"bb8408bd",
          3067 => x"84c02976",
          3068 => x"71315454",
          3069 => x"84bb8408",
          3070 => x"5283dca0",
          3071 => x"51ffb488",
          3072 => x"3f873d0d",
          3073 => x"0483f3fc",
          3074 => x"0856bd84",
          3075 => x"c0527551",
          3076 => x"c9933f84",
          3077 => x"bb8408bd",
          3078 => x"84c02976",
          3079 => x"71315454",
          3080 => x"84bb8408",
          3081 => x"5283dccc",
          3082 => x"51ffb3dc",
          3083 => x"3f83f486",
          3084 => x"33557480",
          3085 => x"2eff9e38",
          3086 => x"ff9f3983",
          3087 => x"dcf851c0",
          3088 => x"b23f83da",
          3089 => x"c051c0ab",
          3090 => x"3f83f3e8",
          3091 => x"085283da",
          3092 => x"cc51ffb3",
          3093 => x"b33f83f3",
          3094 => x"ec085283",
          3095 => x"daf451ff",
          3096 => x"b3a63f83",
          3097 => x"f3f00852",
          3098 => x"83db9c51",
          3099 => x"ffb3993f",
          3100 => x"83dbc451",
          3101 => x"ffbffc3f",
          3102 => x"83f3f422",
          3103 => x"5283dbcc",
          3104 => x"51ffb384",
          3105 => x"3f83f3f8",
          3106 => x"0856bd84",
          3107 => x"c0527551",
          3108 => x"c8933f84",
          3109 => x"bb8408bd",
          3110 => x"84c02976",
          3111 => x"71315454",
          3112 => x"84bb8408",
          3113 => x"5283dbf4",
          3114 => x"51ffb2dc",
          3115 => x"3f83f48b",
          3116 => x"33557480",
          3117 => x"2efe9638",
          3118 => x"fecb3983",
          3119 => x"dd8051ff",
          3120 => x"bfb13f83",
          3121 => x"f48e3354",
          3122 => x"73802efd",
          3123 => x"8e38feeb",
          3124 => x"3983dd88",
          3125 => x"51ffbf9b",
          3126 => x"3f83f48d",
          3127 => x"33567580",
          3128 => x"2efcef38",
          3129 => x"d63983dd",
          3130 => x"9451ffbf",
          3131 => x"863f83f4",
          3132 => x"8c335574",
          3133 => x"802efcd1",
          3134 => x"38d73983",
          3135 => x"dda051ff",
          3136 => x"bef13f83",
          3137 => x"f4873354",
          3138 => x"73802efc",
          3139 => x"b338d739",
          3140 => x"83f49233",
          3141 => x"5283ddb4",
          3142 => x"51ffb1ec",
          3143 => x"3f83f485",
          3144 => x"33567580",
          3145 => x"2efc9038",
          3146 => x"d23983f4",
          3147 => x"94335283",
          3148 => x"ddd451ff",
          3149 => x"b1d23f83",
          3150 => x"f4913355",
          3151 => x"74802efb",
          3152 => x"ed38cd39",
          3153 => x"83f49033",
          3154 => x"5283ddf4",
          3155 => x"51ffb1b8",
          3156 => x"3f83f493",
          3157 => x"33547380",
          3158 => x"2efbca38",
          3159 => x"cd3983f3",
          3160 => x"d00883f3",
          3161 => x"d4081154",
          3162 => x"5283de94",
          3163 => x"51ffb198",
          3164 => x"3f83f48f",
          3165 => x"33567580",
          3166 => x"2efba138",
          3167 => x"c73983f3",
          3168 => x"c80883f3",
          3169 => x"cc081154",
          3170 => x"5283deb0",
          3171 => x"51ffb0f8",
          3172 => x"3f83f48a",
          3173 => x"33547380",
          3174 => x"2efaf838",
          3175 => x"c13983f3",
          3176 => x"c00883f3",
          3177 => x"c4081154",
          3178 => x"5283decc",
          3179 => x"51ffb0d8",
          3180 => x"3f83f489",
          3181 => x"33557480",
          3182 => x"2efacf38",
          3183 => x"c13983f3",
          3184 => x"d80883f3",
          3185 => x"dc081154",
          3186 => x"5283dee8",
          3187 => x"51ffb0b8",
          3188 => x"3f83f488",
          3189 => x"33567580",
          3190 => x"2efaa638",
          3191 => x"c13983f3",
          3192 => x"e00883f3",
          3193 => x"e4081154",
          3194 => x"5283df84",
          3195 => x"51ffb098",
          3196 => x"3f83f48b",
          3197 => x"33547380",
          3198 => x"2ef9fd38",
          3199 => x"c13983df",
          3200 => x"a051ffb0",
          3201 => x"833f83da",
          3202 => x"a851ffbc",
          3203 => x"e63f83f4",
          3204 => x"86335574",
          3205 => x"802ef9d7",
          3206 => x"38c439ff",
          3207 => x"3d0d028e",
          3208 => x"05335271",
          3209 => x"85268c38",
          3210 => x"71101083",
          3211 => x"c48c0552",
          3212 => x"71080483",
          3213 => x"dfb451ff",
          3214 => x"afce3f83",
          3215 => x"3d0d0483",
          3216 => x"dfbc51ff",
          3217 => x"afc23f83",
          3218 => x"3d0d0483",
          3219 => x"dfc451ff",
          3220 => x"afb63f83",
          3221 => x"3d0d0483",
          3222 => x"dfcc51ff",
          3223 => x"afaa3f83",
          3224 => x"3d0d0483",
          3225 => x"dfd451ff",
          3226 => x"af9e3f83",
          3227 => x"3d0d0483",
          3228 => x"dfdc51ff",
          3229 => x"af923f83",
          3230 => x"3d0d0471",
          3231 => x"88800c04",
          3232 => x"800b87c0",
          3233 => x"96840c04",
          3234 => x"83f49808",
          3235 => x"87c09684",
          3236 => x"0c04d93d",
          3237 => x"0daa3d08",
          3238 => x"ad3d085a",
          3239 => x"5a817057",
          3240 => x"58805283",
          3241 => x"f4ec0851",
          3242 => x"8287fb3f",
          3243 => x"84bb8408",
          3244 => x"80ed388b",
          3245 => x"3d57ff0b",
          3246 => x"83f4ec08",
          3247 => x"545580f8",
          3248 => x"52765182",
          3249 => x"d38e3f84",
          3250 => x"bb840880",
          3251 => x"2ea43876",
          3252 => x"51c0d53f",
          3253 => x"84bb8408",
          3254 => x"81175755",
          3255 => x"800b84bb",
          3256 => x"8408258e",
          3257 => x"3884bb84",
          3258 => x"08ff0570",
          3259 => x"18555580",
          3260 => x"74347409",
          3261 => x"70307072",
          3262 => x"079f2a51",
          3263 => x"55557876",
          3264 => x"2e853873",
          3265 => x"ffb03883",
          3266 => x"f4ec088c",
          3267 => x"11085351",
          3268 => x"8287933f",
          3269 => x"84bb8408",
          3270 => x"8f387876",
          3271 => x"2e9a3877",
          3272 => x"84bb840c",
          3273 => x"a93d0d04",
          3274 => x"83e3b851",
          3275 => x"ffadd93f",
          3276 => x"78762e09",
          3277 => x"8106e838",
          3278 => x"76527951",
          3279 => x"c0893f79",
          3280 => x"51ffbfe4",
          3281 => x"3fab3d08",
          3282 => x"5684bb84",
          3283 => x"08763476",
          3284 => x"5283e3e4",
          3285 => x"51ffadb0",
          3286 => x"3f800b84",
          3287 => x"bb840ca9",
          3288 => x"3d0d04d8",
          3289 => x"3d0dab3d",
          3290 => x"08ad3d08",
          3291 => x"71725d72",
          3292 => x"3357575a",
          3293 => x"5773a02e",
          3294 => x"81923880",
          3295 => x"0b8d3d59",
          3296 => x"56751010",
          3297 => x"1083f4f8",
          3298 => x"05700852",
          3299 => x"54ffbf98",
          3300 => x"3f84bb84",
          3301 => x"08537952",
          3302 => x"730851ff",
          3303 => x"bff73f84",
          3304 => x"bb840890",
          3305 => x"38841433",
          3306 => x"5473812e",
          3307 => x"81883873",
          3308 => x"822e9938",
          3309 => x"81167081",
          3310 => x"ff065754",
          3311 => x"827627c1",
          3312 => x"38805473",
          3313 => x"84bb840c",
          3314 => x"aa3d0d04",
          3315 => x"811a5aaa",
          3316 => x"3dff8411",
          3317 => x"53ff8005",
          3318 => x"51c7ab3f",
          3319 => x"84bb8408",
          3320 => x"802ed138",
          3321 => x"ff1b5378",
          3322 => x"527651fd",
          3323 => x"a53f84bb",
          3324 => x"840881ff",
          3325 => x"06547380",
          3326 => x"2ec93881",
          3327 => x"167081ff",
          3328 => x"06575482",
          3329 => x"7627fef9",
          3330 => x"38ffb639",
          3331 => x"78337705",
          3332 => x"56767627",
          3333 => x"fee53881",
          3334 => x"15705b70",
          3335 => x"33555573",
          3336 => x"a02e0981",
          3337 => x"06fed438",
          3338 => x"757526eb",
          3339 => x"38800b8d",
          3340 => x"3d5956fe",
          3341 => x"cc397384",
          3342 => x"bb840853",
          3343 => x"83f4ec08",
          3344 => x"52568284",
          3345 => x"e13f84bb",
          3346 => x"840880d0",
          3347 => x"3883f4ec",
          3348 => x"085380f8",
          3349 => x"52775182",
          3350 => x"cffa3f84",
          3351 => x"bb840880",
          3352 => x"2eba3877",
          3353 => x"51ffbdc0",
          3354 => x"3f84bb84",
          3355 => x"0855800b",
          3356 => x"84bb8408",
          3357 => x"259d3884",
          3358 => x"bb8408ff",
          3359 => x"05701958",
          3360 => x"55807734",
          3361 => x"77537552",
          3362 => x"811683e3",
          3363 => x"ac5256ff",
          3364 => x"aaf63f74",
          3365 => x"ff2e0981",
          3366 => x"06ffb238",
          3367 => x"810b84bb",
          3368 => x"840caa3d",
          3369 => x"0d04cd3d",
          3370 => x"0db63d08",
          3371 => x"b83d08ba",
          3372 => x"3d08bc3d",
          3373 => x"08be3d08",
          3374 => x"425b5842",
          3375 => x"5c800bb5",
          3376 => x"3d3483f4",
          3377 => x"f4335d75",
          3378 => x"83f4f034",
          3379 => x"83f4ec08",
          3380 => x"55749e38",
          3381 => x"747681ff",
          3382 => x"06565774",
          3383 => x"802e82ed",
          3384 => x"3877802e",
          3385 => x"91883881",
          3386 => x"7078065a",
          3387 => x"5678908b",
          3388 => x"3877802e",
          3389 => x"90f83894",
          3390 => x"3db53d40",
          3391 => x"408051ea",
          3392 => x"fb3f84bb",
          3393 => x"8408982b",
          3394 => x"70982c5b",
          3395 => x"5779ff2e",
          3396 => x"81d73879",
          3397 => x"81ff0684",
          3398 => x"e2c03370",
          3399 => x"982b7098",
          3400 => x"2c84e2bc",
          3401 => x"3370982b",
          3402 => x"70972c71",
          3403 => x"982c0570",
          3404 => x"101083df",
          3405 => x"e0057008",
          3406 => x"15703351",
          3407 => x"53495d5a",
          3408 => x"525b585c",
          3409 => x"59815774",
          3410 => x"792e80cd",
          3411 => x"38787527",
          3412 => x"81a83875",
          3413 => x"81800a29",
          3414 => x"81ff0a05",
          3415 => x"70982c57",
          3416 => x"42807624",
          3417 => x"81ec3875",
          3418 => x"10167082",
          3419 => x"2b565780",
          3420 => x"0b83dfe4",
          3421 => x"16334357",
          3422 => x"77622591",
          3423 => x"3883dfe0",
          3424 => x"15081870",
          3425 => x"33564278",
          3426 => x"752e81b6",
          3427 => x"3876802e",
          3428 => x"c2387584",
          3429 => x"e2bc3481",
          3430 => x"5776802e",
          3431 => x"81ba3881",
          3432 => x"1b70982b",
          3433 => x"70982c84",
          3434 => x"e2bc3370",
          3435 => x"982b7097",
          3436 => x"2c71982c",
          3437 => x"0570822b",
          3438 => x"83dfe411",
          3439 => x"335f535e",
          3440 => x"5e585d57",
          3441 => x"577a782e",
          3442 => x"81b13876",
          3443 => x"84e2c034",
          3444 => x"8051e9a8",
          3445 => x"3f84bb84",
          3446 => x"08982b70",
          3447 => x"982c5b57",
          3448 => x"79ff2e09",
          3449 => x"8106feab",
          3450 => x"387d802e",
          3451 => x"fe8f387d",
          3452 => x"2dfe8a39",
          3453 => x"815776ff",
          3454 => x"99387581",
          3455 => x"800a2981",
          3456 => x"800a0570",
          3457 => x"982c7081",
          3458 => x"ff065957",
          3459 => x"42769526",
          3460 => x"80c03875",
          3461 => x"10167082",
          3462 => x"2b515580",
          3463 => x"0b83dfe4",
          3464 => x"16334357",
          3465 => x"776225ce",
          3466 => x"3883dfe0",
          3467 => x"15081870",
          3468 => x"33435578",
          3469 => x"622effbc",
          3470 => x"3876802e",
          3471 => x"ffbc38fe",
          3472 => x"d1398157",
          3473 => x"76802efe",
          3474 => x"8a38fec6",
          3475 => x"398157fd",
          3476 => x"90398057",
          3477 => x"76fec838",
          3478 => x"7684e2c0",
          3479 => x"347684e2",
          3480 => x"bc34797f",
          3481 => x"3476600c",
          3482 => x"63557495",
          3483 => x"26fd8e38",
          3484 => x"74101083",
          3485 => x"c4a40557",
          3486 => x"76080483",
          3487 => x"dfe81508",
          3488 => x"600c800b",
          3489 => x"84e2c034",
          3490 => x"800b84e2",
          3491 => x"bc34d939",
          3492 => x"84e2c833",
          3493 => x"5675802e",
          3494 => x"fce33884",
          3495 => x"e6e80852",
          3496 => x"8851ffb5",
          3497 => x"c93f84e2",
          3498 => x"c833ff05",
          3499 => x"5b7a84e2",
          3500 => x"c834fcc9",
          3501 => x"3984e2c8",
          3502 => x"337081ff",
          3503 => x"0684e2c4",
          3504 => x"335a5755",
          3505 => x"757827fc",
          3506 => x"b43884e6",
          3507 => x"e8085281",
          3508 => x"15426184",
          3509 => x"e2c8347b",
          3510 => x"16703352",
          3511 => x"55ffb58e",
          3512 => x"3ffc9a39",
          3513 => x"7c932e90",
          3514 => x"bd387c92",
          3515 => x"2690387c",
          3516 => x"101083f4",
          3517 => x"a0057008",
          3518 => x"5758758f",
          3519 => x"a538800b",
          3520 => x"84e2c434",
          3521 => x"807c3484",
          3522 => x"e2c43384",
          3523 => x"e2c83356",
          3524 => x"5674802e",
          3525 => x"b63884e6",
          3526 => x"e8085288",
          3527 => x"51ffb4ce",
          3528 => x"3f84e6e8",
          3529 => x"0852a051",
          3530 => x"ffb4c33f",
          3531 => x"84e6e808",
          3532 => x"528851ff",
          3533 => x"b4b83f84",
          3534 => x"e2c833ff",
          3535 => x"05597884",
          3536 => x"e2c83478",
          3537 => x"81ff0655",
          3538 => x"74cc387b",
          3539 => x"51ffa5b8",
          3540 => x"3f7584e2",
          3541 => x"c834fba5",
          3542 => x"397c8a38",
          3543 => x"83f4e808",
          3544 => x"56758cf1",
          3545 => x"38ff1d70",
          3546 => x"81ff0658",
          3547 => x"58769226",
          3548 => x"90387c10",
          3549 => x"1083f498",
          3550 => x"05700857",
          3551 => x"55758dbc",
          3552 => x"387c9326",
          3553 => x"faf7387c",
          3554 => x"101083f4",
          3555 => x"9c057008",
          3556 => x"57597580",
          3557 => x"2efae638",
          3558 => x"7551ffb7",
          3559 => x"8b3f84bb",
          3560 => x"840884e2",
          3561 => x"c43484bb",
          3562 => x"840881ff",
          3563 => x"06810553",
          3564 => x"75527b51",
          3565 => x"ffb7b33f",
          3566 => x"84e2c433",
          3567 => x"84e2c833",
          3568 => x"56567480",
          3569 => x"2eff8438",
          3570 => x"84e6e808",
          3571 => x"528851ff",
          3572 => x"b39c3f84",
          3573 => x"e6e80852",
          3574 => x"a051ffb3",
          3575 => x"913f84e6",
          3576 => x"e8085288",
          3577 => x"51ffb386",
          3578 => x"3f84e2c8",
          3579 => x"33ff0555",
          3580 => x"7484e2c8",
          3581 => x"347481ff",
          3582 => x"0655c739",
          3583 => x"84e2c833",
          3584 => x"7081ff06",
          3585 => x"84e2c433",
          3586 => x"5c575575",
          3587 => x"7a27f9ed",
          3588 => x"3884e6e8",
          3589 => x"08528115",
          3590 => x"577684e2",
          3591 => x"c8347b16",
          3592 => x"70335255",
          3593 => x"ffb2c73f",
          3594 => x"84e2c833",
          3595 => x"7081ff06",
          3596 => x"84e2c433",
          3597 => x"5a575575",
          3598 => x"7827f9c1",
          3599 => x"3884e6e8",
          3600 => x"08528115",
          3601 => x"577684e2",
          3602 => x"c8347b16",
          3603 => x"70335255",
          3604 => x"ffb29b3f",
          3605 => x"84e2c833",
          3606 => x"7081ff06",
          3607 => x"84e2c433",
          3608 => x"5a575577",
          3609 => x"7626ffa9",
          3610 => x"38f99239",
          3611 => x"84e2c833",
          3612 => x"84e2c433",
          3613 => x"56567476",
          3614 => x"2ef98238",
          3615 => x"ff155b7a",
          3616 => x"84e2c434",
          3617 => x"75982b70",
          3618 => x"982c7c81",
          3619 => x"ff064457",
          3620 => x"59617624",
          3621 => x"80ef3884",
          3622 => x"e6e80852",
          3623 => x"a051ffb1",
          3624 => x"cd3f84e2",
          3625 => x"c8337098",
          3626 => x"2b70982c",
          3627 => x"84e2c433",
          3628 => x"5a574356",
          3629 => x"747724f8",
          3630 => x"c43884e6",
          3631 => x"e8085288",
          3632 => x"51ffb1aa",
          3633 => x"3f748180",
          3634 => x"0a298180",
          3635 => x"0a057098",
          3636 => x"2c84e2c4",
          3637 => x"335d5659",
          3638 => x"747b24f8",
          3639 => x"a03884e6",
          3640 => x"e8085288",
          3641 => x"51ffb186",
          3642 => x"3f748180",
          3643 => x"0a298180",
          3644 => x"0a057098",
          3645 => x"2c84e2c4",
          3646 => x"335d5659",
          3647 => x"7a7525ff",
          3648 => x"b938f7f9",
          3649 => x"397b1658",
          3650 => x"81183378",
          3651 => x"3484e6e8",
          3652 => x"08527733",
          3653 => x"51ffb0d6",
          3654 => x"3f758180",
          3655 => x"0a298180",
          3656 => x"0a057098",
          3657 => x"2c84e2c4",
          3658 => x"335c5755",
          3659 => x"757a25fe",
          3660 => x"e6387b16",
          3661 => x"58811833",
          3662 => x"783484e6",
          3663 => x"e8085277",
          3664 => x"3351ffb0",
          3665 => x"a93f7581",
          3666 => x"800a2981",
          3667 => x"800a0570",
          3668 => x"982c84e2",
          3669 => x"c4335c57",
          3670 => x"55797624",
          3671 => x"ffa738fe",
          3672 => x"b63984e2",
          3673 => x"c8335574",
          3674 => x"802ef791",
          3675 => x"3884e6e8",
          3676 => x"08528851",
          3677 => x"ffaff73f",
          3678 => x"84e2c833",
          3679 => x"ff055776",
          3680 => x"84e2c834",
          3681 => x"7681ff06",
          3682 => x"55dd3984",
          3683 => x"e2c4337c",
          3684 => x"05418061",
          3685 => x"3484e6e8",
          3686 => x"08528a51",
          3687 => x"ffafcf3f",
          3688 => x"84e2c452",
          3689 => x"7b51f3bb",
          3690 => x"3f84bb84",
          3691 => x"0881ff06",
          3692 => x"58778ada",
          3693 => x"3884e2c4",
          3694 => x"33577680",
          3695 => x"2e80f038",
          3696 => x"83f4f433",
          3697 => x"70101083",
          3698 => x"f49c0570",
          3699 => x"08574156",
          3700 => x"748bc238",
          3701 => x"75822b87",
          3702 => x"fc0683f4",
          3703 => x"9c058118",
          3704 => x"70535759",
          3705 => x"80e8e23f",
          3706 => x"84bb8408",
          3707 => x"790c83f4",
          3708 => x"f4337010",
          3709 => x"1083f49c",
          3710 => x"05700854",
          3711 => x"4383e394",
          3712 => x"525bffa0",
          3713 => x"833f83f4",
          3714 => x"f4337010",
          3715 => x"1083f49c",
          3716 => x"05700857",
          3717 => x"5e5e748b",
          3718 => x"cf3883f4",
          3719 => x"ec085675",
          3720 => x"802e8c38",
          3721 => x"83f4f033",
          3722 => x"5877802e",
          3723 => x"8bde3880",
          3724 => x"0b84e2c8",
          3725 => x"34800b84",
          3726 => x"e2c4347b",
          3727 => x"84bb840c",
          3728 => x"b53d0d04",
          3729 => x"84e2c833",
          3730 => x"5574802e",
          3731 => x"b63884e6",
          3732 => x"e8085288",
          3733 => x"51ffae96",
          3734 => x"3f84e6e8",
          3735 => x"0852a051",
          3736 => x"ffae8b3f",
          3737 => x"84e6e808",
          3738 => x"528851ff",
          3739 => x"ae803f84",
          3740 => x"e2c833ff",
          3741 => x"05426184",
          3742 => x"e2c83461",
          3743 => x"81ff0655",
          3744 => x"74cc3883",
          3745 => x"d38051ff",
          3746 => x"9efe3f80",
          3747 => x"0b84e2c8",
          3748 => x"34800b84",
          3749 => x"e2c434f4",
          3750 => x"e43984e2",
          3751 => x"c8337081",
          3752 => x"ff065c56",
          3753 => x"7a802ef4",
          3754 => x"d43884e2",
          3755 => x"c433ff05",
          3756 => x"5a7984e2",
          3757 => x"c434ff16",
          3758 => x"587784e2",
          3759 => x"c83484e6",
          3760 => x"e8085288",
          3761 => x"51ffada6",
          3762 => x"3f84e2c8",
          3763 => x"3370982b",
          3764 => x"70982c84",
          3765 => x"e2c4335a",
          3766 => x"525a5676",
          3767 => x"762480ef",
          3768 => x"3884e6e8",
          3769 => x"0852a051",
          3770 => x"ffad833f",
          3771 => x"84e2c833",
          3772 => x"70982b70",
          3773 => x"982c84e2",
          3774 => x"c4335c57",
          3775 => x"59567479",
          3776 => x"24f3fa38",
          3777 => x"84e6e808",
          3778 => x"528851ff",
          3779 => x"ace03f74",
          3780 => x"81800a29",
          3781 => x"81800a05",
          3782 => x"70982c84",
          3783 => x"e2c4335c",
          3784 => x"5155747a",
          3785 => x"24f3d638",
          3786 => x"84e6e808",
          3787 => x"528851ff",
          3788 => x"acbc3f74",
          3789 => x"81800a29",
          3790 => x"81800a05",
          3791 => x"70982c84",
          3792 => x"e2c4335c",
          3793 => x"51557975",
          3794 => x"25ffb938",
          3795 => x"f3af397b",
          3796 => x"16578117",
          3797 => x"33773484",
          3798 => x"e6e80852",
          3799 => x"763351ff",
          3800 => x"ac8c3f75",
          3801 => x"81800a29",
          3802 => x"81800a05",
          3803 => x"70982c84",
          3804 => x"e2c43344",
          3805 => x"575b7562",
          3806 => x"25fee638",
          3807 => x"7b165781",
          3808 => x"17337734",
          3809 => x"84e6e808",
          3810 => x"52763351",
          3811 => x"ffabdf3f",
          3812 => x"7581800a",
          3813 => x"2981800a",
          3814 => x"0570982c",
          3815 => x"84e2c433",
          3816 => x"44575b61",
          3817 => x"7624ffa7",
          3818 => x"38feb639",
          3819 => x"837c3480",
          3820 => x"0b811d34",
          3821 => x"84e2c833",
          3822 => x"5574802e",
          3823 => x"b63884e6",
          3824 => x"e8085288",
          3825 => x"51ffaba6",
          3826 => x"3f84e6e8",
          3827 => x"0852a051",
          3828 => x"ffab9b3f",
          3829 => x"84e6e808",
          3830 => x"528851ff",
          3831 => x"ab903f84",
          3832 => x"e2c833ff",
          3833 => x"055d7c84",
          3834 => x"e2c8347c",
          3835 => x"81ff0655",
          3836 => x"74cc3883",
          3837 => x"d38051ff",
          3838 => x"9c8e3f80",
          3839 => x"0b84e2c8",
          3840 => x"34800b84",
          3841 => x"e2c4347b",
          3842 => x"84bb840c",
          3843 => x"b53d0d04",
          3844 => x"84e2c833",
          3845 => x"7081ff06",
          3846 => x"58587661",
          3847 => x"2ef1de38",
          3848 => x"84e2c433",
          3849 => x"55767527",
          3850 => x"ae387498",
          3851 => x"2b70982c",
          3852 => x"57427676",
          3853 => x"24a1387b",
          3854 => x"165b7a33",
          3855 => x"811c3475",
          3856 => x"81800a29",
          3857 => x"81ff0a05",
          3858 => x"70982c84",
          3859 => x"e2c83352",
          3860 => x"57587578",
          3861 => x"25e13881",
          3862 => x"18557484",
          3863 => x"e2c83477",
          3864 => x"81ff067c",
          3865 => x"0559b43d",
          3866 => x"33793484",
          3867 => x"e2c43357",
          3868 => x"7661258b",
          3869 => x"38811756",
          3870 => x"7584e2c4",
          3871 => x"34755784",
          3872 => x"e2c83370",
          3873 => x"81800a29",
          3874 => x"81ff0a05",
          3875 => x"70982c79",
          3876 => x"81ff0645",
          3877 => x"585c5861",
          3878 => x"76248190",
          3879 => x"3877982b",
          3880 => x"70982c78",
          3881 => x"81ff065b",
          3882 => x"575a7579",
          3883 => x"25f0ce38",
          3884 => x"84e6e808",
          3885 => x"528851ff",
          3886 => x"a9b43f75",
          3887 => x"81800a29",
          3888 => x"81800a05",
          3889 => x"70982c84",
          3890 => x"e2c43357",
          3891 => x"57427575",
          3892 => x"25f0aa38",
          3893 => x"84e6e808",
          3894 => x"528851ff",
          3895 => x"a9903f75",
          3896 => x"81800a29",
          3897 => x"81800a05",
          3898 => x"70982c84",
          3899 => x"e2c43357",
          3900 => x"57427476",
          3901 => x"24ffb938",
          3902 => x"f0833984",
          3903 => x"a85180e2",
          3904 => x"c83f84bb",
          3905 => x"840883f4",
          3906 => x"ec0c84bb",
          3907 => x"84085283",
          3908 => x"e2c051ff",
          3909 => x"99f23f83",
          3910 => x"f4ec0855",
          3911 => x"7486a638",
          3912 => x"7583f4f0",
          3913 => x"3477efcf",
          3914 => x"3880c339",
          3915 => x"84e6e808",
          3916 => x"527b1670",
          3917 => x"335258ff",
          3918 => x"a8b43f75",
          3919 => x"81800a29",
          3920 => x"81800a05",
          3921 => x"70982c84",
          3922 => x"e2c43352",
          3923 => x"57577676",
          3924 => x"24da3884",
          3925 => x"e2c83370",
          3926 => x"982b7098",
          3927 => x"2c7981ff",
          3928 => x"065c585b",
          3929 => x"58757925",
          3930 => x"ef9338fe",
          3931 => x"c33983f4",
          3932 => x"ec08802e",
          3933 => x"ef813883",
          3934 => x"f49c5793",
          3935 => x"56760855",
          3936 => x"74bb38ff",
          3937 => x"16841858",
          3938 => x"56758025",
          3939 => x"f038800b",
          3940 => x"83f4f434",
          3941 => x"83f4ec08",
          3942 => x"5574802e",
          3943 => x"eed93874",
          3944 => x"5181e7e5",
          3945 => x"3f83f4ec",
          3946 => x"085180db",
          3947 => x"ac3f800b",
          3948 => x"83f4ec0c",
          3949 => x"943db53d",
          3950 => x"4040eec1",
          3951 => x"39745180",
          3952 => x"db973f80",
          3953 => x"770cff16",
          3954 => x"84185856",
          3955 => x"758025ff",
          3956 => x"ac38ffba",
          3957 => x"397551ff",
          3958 => x"aace3f84",
          3959 => x"bb840884",
          3960 => x"e2c43484",
          3961 => x"bb840881",
          3962 => x"ff068105",
          3963 => x"5375527b",
          3964 => x"51ffaaf6",
          3965 => x"3f930b84",
          3966 => x"e2c43384",
          3967 => x"e2c83357",
          3968 => x"575d7480",
          3969 => x"2ef2c438",
          3970 => x"84e6e808",
          3971 => x"528851ff",
          3972 => x"a6dc3f84",
          3973 => x"e6e80852",
          3974 => x"a051ffa6",
          3975 => x"d13f84e6",
          3976 => x"e8085288",
          3977 => x"51ffa6c6",
          3978 => x"3f84e2c8",
          3979 => x"33ff0559",
          3980 => x"7884e2c8",
          3981 => x"347881ff",
          3982 => x"0655c739",
          3983 => x"7551ffa9",
          3984 => x"e73f84bb",
          3985 => x"840884e2",
          3986 => x"c43484bb",
          3987 => x"840881ff",
          3988 => x"06810553",
          3989 => x"75527b51",
          3990 => x"ffaa8f3f",
          3991 => x"7684e2c4",
          3992 => x"3384e2c8",
          3993 => x"3357575d",
          3994 => x"74802ef1",
          3995 => x"de3884e6",
          3996 => x"e8085288",
          3997 => x"51ffa5f6",
          3998 => x"3f84e6e8",
          3999 => x"0852a051",
          4000 => x"ffa5eb3f",
          4001 => x"84e6e808",
          4002 => x"528851ff",
          4003 => x"a5e03f84",
          4004 => x"e2c833ff",
          4005 => x"05577684",
          4006 => x"e2c83476",
          4007 => x"81ff0655",
          4008 => x"c7397551",
          4009 => x"ffa9813f",
          4010 => x"84bb8408",
          4011 => x"84e2c434",
          4012 => x"84bb8408",
          4013 => x"81ff0681",
          4014 => x"05537552",
          4015 => x"7b51ffa9",
          4016 => x"a93f811d",
          4017 => x"7081ff06",
          4018 => x"84e2c433",
          4019 => x"84e2c833",
          4020 => x"58525e56",
          4021 => x"74802ef0",
          4022 => x"f23884e6",
          4023 => x"e8085288",
          4024 => x"51ffa58a",
          4025 => x"3f84e6e8",
          4026 => x"0852a051",
          4027 => x"ffa4ff3f",
          4028 => x"84e6e808",
          4029 => x"528851ff",
          4030 => x"a4f43f84",
          4031 => x"e2c833ff",
          4032 => x"055b7a84",
          4033 => x"e2c8347a",
          4034 => x"81ff0655",
          4035 => x"c739807c",
          4036 => x"34800b84",
          4037 => x"e2c83480",
          4038 => x"0b84e2c4",
          4039 => x"347b84bb",
          4040 => x"840cb53d",
          4041 => x"0d0483f4",
          4042 => x"9c085675",
          4043 => x"802eefce",
          4044 => x"387551ff",
          4045 => x"a7f23f84",
          4046 => x"bb840884",
          4047 => x"e2c43484",
          4048 => x"bb840881",
          4049 => x"ff068105",
          4050 => x"5375527b",
          4051 => x"51ffa89a",
          4052 => x"3f84e2c4",
          4053 => x"3384e2c8",
          4054 => x"33565674",
          4055 => x"802eefeb",
          4056 => x"3884e6e8",
          4057 => x"08528851",
          4058 => x"ffa4833f",
          4059 => x"84e6e808",
          4060 => x"52a051ff",
          4061 => x"a3f83f84",
          4062 => x"e6e80852",
          4063 => x"8851ffa3",
          4064 => x"ed3f84e2",
          4065 => x"c833ff05",
          4066 => x"597884e2",
          4067 => x"c8347881",
          4068 => x"ff0655c7",
          4069 => x"39745180",
          4070 => x"d7bf3f83",
          4071 => x"f4f43370",
          4072 => x"822b87fc",
          4073 => x"0683f49c",
          4074 => x"05811970",
          4075 => x"54525a56",
          4076 => x"80dd963f",
          4077 => x"84bb8408",
          4078 => x"790c83f4",
          4079 => x"f4337010",
          4080 => x"1083f49c",
          4081 => x"05700854",
          4082 => x"4383e394",
          4083 => x"525bff94",
          4084 => x"b73f83f4",
          4085 => x"f4337010",
          4086 => x"1083f49c",
          4087 => x"05700857",
          4088 => x"5e5e7480",
          4089 => x"2ef4b338",
          4090 => x"75537b52",
          4091 => x"7451ffa6",
          4092 => x"f93f83f4",
          4093 => x"f4338105",
          4094 => x"7081ff06",
          4095 => x"56569375",
          4096 => x"27839f38",
          4097 => x"7783f4f4",
          4098 => x"34f48f39",
          4099 => x"b53dfef8",
          4100 => x"05547653",
          4101 => x"7b527551",
          4102 => x"81d98a3f",
          4103 => x"83f4ec08",
          4104 => x"528a5182",
          4105 => x"b9fc3f83",
          4106 => x"f4ec0851",
          4107 => x"81de893f",
          4108 => x"800b84e2",
          4109 => x"c834800b",
          4110 => x"84e2c434",
          4111 => x"7b84bb84",
          4112 => x"0cb53d0d",
          4113 => x"04935377",
          4114 => x"52745181",
          4115 => x"caa83f84",
          4116 => x"bb840882",
          4117 => x"d53884bb",
          4118 => x"8408973d",
          4119 => x"5c5d83f4",
          4120 => x"ec085380",
          4121 => x"f8527a51",
          4122 => x"82b7e93f",
          4123 => x"84bb8408",
          4124 => x"5a84bb84",
          4125 => x"087b2e09",
          4126 => x"8106e8f5",
          4127 => x"3884bb84",
          4128 => x"0851ffa5",
          4129 => x"a33f84bb",
          4130 => x"84085780",
          4131 => x"0b84bb84",
          4132 => x"082580fb",
          4133 => x"3884bb84",
          4134 => x"08ff0570",
          4135 => x"1b575780",
          4136 => x"76347681",
          4137 => x"ff0683f4",
          4138 => x"f4337010",
          4139 => x"1083f49c",
          4140 => x"05700858",
          4141 => x"41575974",
          4142 => x"818a3875",
          4143 => x"822b87fc",
          4144 => x"0683f49c",
          4145 => x"05811a70",
          4146 => x"53575f80",
          4147 => x"dafb3f84",
          4148 => x"bb84087f",
          4149 => x"0c83f4f4",
          4150 => x"33701010",
          4151 => x"83f49c05",
          4152 => x"70085456",
          4153 => x"83e39452",
          4154 => x"59ff929c",
          4155 => x"3f83f4f4",
          4156 => x"33701010",
          4157 => x"83f49c05",
          4158 => x"70085741",
          4159 => x"4274a038",
          4160 => x"811d7081",
          4161 => x"ff065e56",
          4162 => x"937d2783",
          4163 => x"38805d76",
          4164 => x"ff2e0981",
          4165 => x"06fec738",
          4166 => x"77e7dc38",
          4167 => x"f8d03975",
          4168 => x"53795274",
          4169 => x"51ffa4c2",
          4170 => x"3f83f4f4",
          4171 => x"33810570",
          4172 => x"81ff065b",
          4173 => x"56937a27",
          4174 => x"80e03880",
          4175 => x"0b83f4f4",
          4176 => x"34ffbd39",
          4177 => x"745180d4",
          4178 => x"903f83f4",
          4179 => x"f4337082",
          4180 => x"2b87fc06",
          4181 => x"83f49c05",
          4182 => x"811b7054",
          4183 => x"52405680",
          4184 => x"d9e73f84",
          4185 => x"bb84087f",
          4186 => x"0c83f4f4",
          4187 => x"33701010",
          4188 => x"83f49c05",
          4189 => x"70085456",
          4190 => x"83e39452",
          4191 => x"59ff9188",
          4192 => x"3f83f4f4",
          4193 => x"33701010",
          4194 => x"83f49c05",
          4195 => x"70085741",
          4196 => x"4274802e",
          4197 => x"feea38ff",
          4198 => x"86397583",
          4199 => x"f4f434fe",
          4200 => x"df397583",
          4201 => x"f4f434f0",
          4202 => x"f13983e2",
          4203 => x"d451ff9d",
          4204 => x"c23f77e6",
          4205 => x"c238f7b6",
          4206 => x"39f23d0d",
          4207 => x"0280c305",
          4208 => x"33028405",
          4209 => x"80c70533",
          4210 => x"5b537283",
          4211 => x"26818d38",
          4212 => x"72812e81",
          4213 => x"8b388173",
          4214 => x"25839e38",
          4215 => x"72822e82",
          4216 => x"a83886c7",
          4217 => x"a0805986",
          4218 => x"c7b08070",
          4219 => x"5e578056",
          4220 => x"9fa05879",
          4221 => x"762e9038",
          4222 => x"7583fab4",
          4223 => x"347583fa",
          4224 => x"b5347583",
          4225 => x"fab22383",
          4226 => x"fab03370",
          4227 => x"982b7190",
          4228 => x"2b077188",
          4229 => x"2b077107",
          4230 => x"7a7f5656",
          4231 => x"565b7877",
          4232 => x"27943880",
          4233 => x"74708405",
          4234 => x"560c7473",
          4235 => x"70840555",
          4236 => x"0c767426",
          4237 => x"ee387578",
          4238 => x"27a23883",
          4239 => x"fab03384",
          4240 => x"99d61779",
          4241 => x"78315555",
          4242 => x"55a00be0",
          4243 => x"e0153474",
          4244 => x"74708105",
          4245 => x"5634ff13",
          4246 => x"5372ee38",
          4247 => x"903d0d04",
          4248 => x"86c7a080",
          4249 => x"0b83fab4",
          4250 => x"33701010",
          4251 => x"1183fab5",
          4252 => x"33719029",
          4253 => x"1174055b",
          4254 => x"41584059",
          4255 => x"86c7b080",
          4256 => x"0b84b8f8",
          4257 => x"337081ff",
          4258 => x"0684b8f7",
          4259 => x"337081ff",
          4260 => x"0683fab2",
          4261 => x"227083ff",
          4262 => x"ff067075",
          4263 => x"295d595d",
          4264 => x"585e575b",
          4265 => x"5d737326",
          4266 => x"87387274",
          4267 => x"31752956",
          4268 => x"7981ff06",
          4269 => x"7e81ff06",
          4270 => x"7c81ff06",
          4271 => x"7a83ffff",
          4272 => x"066281ff",
          4273 => x"06707529",
          4274 => x"145d4257",
          4275 => x"575b5c74",
          4276 => x"74268f38",
          4277 => x"83fab433",
          4278 => x"74763105",
          4279 => x"707d291b",
          4280 => x"595f7683",
          4281 => x"065c7b80",
          4282 => x"2efe9c38",
          4283 => x"787d5553",
          4284 => x"727726fe",
          4285 => x"c1388073",
          4286 => x"70810555",
          4287 => x"3483fab0",
          4288 => x"33747081",
          4289 => x"055634e8",
          4290 => x"3986c7a0",
          4291 => x"805986c7",
          4292 => x"b0807084",
          4293 => x"b8f83370",
          4294 => x"81ff0684",
          4295 => x"b8f73370",
          4296 => x"81ff0683",
          4297 => x"fab22270",
          4298 => x"74295d5b",
          4299 => x"5d575e56",
          4300 => x"5e577478",
          4301 => x"2781df38",
          4302 => x"7381ff06",
          4303 => x"7381ff06",
          4304 => x"71712918",
          4305 => x"5a545479",
          4306 => x"802efdbb",
          4307 => x"38800b83",
          4308 => x"fab43480",
          4309 => x"0b83fab5",
          4310 => x"3483fab0",
          4311 => x"3370982b",
          4312 => x"71902b07",
          4313 => x"71882b07",
          4314 => x"71077a7f",
          4315 => x"5656565b",
          4316 => x"767926fd",
          4317 => x"ae38fdbe",
          4318 => x"3972fce6",
          4319 => x"3883fab4",
          4320 => x"337081ff",
          4321 => x"06701010",
          4322 => x"1183fab5",
          4323 => x"33719029",
          4324 => x"1186c7a0",
          4325 => x"80115e57",
          4326 => x"5b56565f",
          4327 => x"86c7b080",
          4328 => x"701484b8",
          4329 => x"f8337081",
          4330 => x"ff0684b8",
          4331 => x"f7337081",
          4332 => x"ff0683fa",
          4333 => x"b2227083",
          4334 => x"ffff067c",
          4335 => x"75296005",
          4336 => x"5e5a415f",
          4337 => x"585f405e",
          4338 => x"57797326",
          4339 => x"8b38727a",
          4340 => x"3115707d",
          4341 => x"29195753",
          4342 => x"7d81ff06",
          4343 => x"7481ff06",
          4344 => x"7171297d",
          4345 => x"83ffff06",
          4346 => x"6281ff06",
          4347 => x"70752958",
          4348 => x"5f5b5c5d",
          4349 => x"557b7826",
          4350 => x"85387775",
          4351 => x"29537973",
          4352 => x"31167983",
          4353 => x"065b5879",
          4354 => x"fde23876",
          4355 => x"83065c7b",
          4356 => x"fdda38fb",
          4357 => x"f2397478",
          4358 => x"317b2956",
          4359 => x"fe9a39fb",
          4360 => x"3d0d878e",
          4361 => x"808c53ff",
          4362 => x"8a733487",
          4363 => x"73348573",
          4364 => x"34817334",
          4365 => x"878e809c",
          4366 => x"5580f475",
          4367 => x"34ffb075",
          4368 => x"34878e80",
          4369 => x"98568076",
          4370 => x"34807634",
          4371 => x"878e8094",
          4372 => x"548a7434",
          4373 => x"807434ff",
          4374 => x"80753481",
          4375 => x"528351fa",
          4376 => x"d83f86c0",
          4377 => x"87e07008",
          4378 => x"545481f8",
          4379 => x"5686c081",
          4380 => x"f8737706",
          4381 => x"84075455",
          4382 => x"72753473",
          4383 => x"087080ff",
          4384 => x"0680c007",
          4385 => x"51537275",
          4386 => x"3486c087",
          4387 => x"cc087077",
          4388 => x"06810751",
          4389 => x"537286c0",
          4390 => x"81f33473",
          4391 => x"0881f706",
          4392 => x"88075372",
          4393 => x"753480d0",
          4394 => x"0b84b8f8",
          4395 => x"34800b84",
          4396 => x"bb840c87",
          4397 => x"3d0d0484",
          4398 => x"b8f83384",
          4399 => x"bb840c04",
          4400 => x"f73d0d02",
          4401 => x"af053302",
          4402 => x"8405b305",
          4403 => x"3384b8f7",
          4404 => x"335b5956",
          4405 => x"81537579",
          4406 => x"2682da38",
          4407 => x"84b8f833",
          4408 => x"83fab533",
          4409 => x"83fab433",
          4410 => x"72712912",
          4411 => x"86c7a080",
          4412 => x"1183fab2",
          4413 => x"225f5157",
          4414 => x"59717c29",
          4415 => x"057083ff",
          4416 => x"ff0683f9",
          4417 => x"8a335357",
          4418 => x"58537281",
          4419 => x"2e83c438",
          4420 => x"83fab222",
          4421 => x"76055574",
          4422 => x"83fab223",
          4423 => x"83fab433",
          4424 => x"76057081",
          4425 => x"ff067a81",
          4426 => x"ff06555b",
          4427 => x"55727a26",
          4428 => x"828c38ff",
          4429 => x"19537283",
          4430 => x"fab43483",
          4431 => x"fab22270",
          4432 => x"83ffff06",
          4433 => x"84b8f633",
          4434 => x"5c555779",
          4435 => x"74268289",
          4436 => x"3884b8f8",
          4437 => x"33767129",
          4438 => x"54588054",
          4439 => x"729f9f26",
          4440 => x"ac388499",
          4441 => x"d6701454",
          4442 => x"55e0e013",
          4443 => x"33e0e016",
          4444 => x"34727081",
          4445 => x"05543375",
          4446 => x"70810557",
          4447 => x"34811454",
          4448 => x"84b8f573",
          4449 => x"27e33873",
          4450 => x"9f9f26a1",
          4451 => x"3883fab0",
          4452 => x"338499d6",
          4453 => x"155455a0",
          4454 => x"0be0e014",
          4455 => x"34747370",
          4456 => x"81055534",
          4457 => x"8114549f",
          4458 => x"9f7427eb",
          4459 => x"3884b8f6",
          4460 => x"33ff0556",
          4461 => x"7583fab2",
          4462 => x"23755778",
          4463 => x"81ff0677",
          4464 => x"83ffff06",
          4465 => x"54547373",
          4466 => x"2681fd38",
          4467 => x"72743181",
          4468 => x"0584b8f8",
          4469 => x"33717129",
          4470 => x"58555775",
          4471 => x"5586c7a0",
          4472 => x"805886c7",
          4473 => x"b0807981",
          4474 => x"ff067581",
          4475 => x"ff067171",
          4476 => x"29195c5c",
          4477 => x"54577579",
          4478 => x"27b93884",
          4479 => x"99d61654",
          4480 => x"e0e01433",
          4481 => x"5384b980",
          4482 => x"13337870",
          4483 => x"81055a34",
          4484 => x"73708105",
          4485 => x"55337770",
          4486 => x"81055934",
          4487 => x"811584b8",
          4488 => x"f83384b8",
          4489 => x"f7337171",
          4490 => x"2919565c",
          4491 => x"5a557275",
          4492 => x"26ce3880",
          4493 => x"537284bb",
          4494 => x"840c8b3d",
          4495 => x"0d047483",
          4496 => x"fab43483",
          4497 => x"fab22270",
          4498 => x"83ffff06",
          4499 => x"84b8f633",
          4500 => x"5c555773",
          4501 => x"7a27fdf9",
          4502 => x"3877802e",
          4503 => x"fedd3878",
          4504 => x"81ff06ff",
          4505 => x"0583fab4",
          4506 => x"33565372",
          4507 => x"752e0981",
          4508 => x"06fec838",
          4509 => x"73763181",
          4510 => x"0584b8f8",
          4511 => x"33717129",
          4512 => x"78722911",
          4513 => x"56525954",
          4514 => x"737327fe",
          4515 => x"ae3883fa",
          4516 => x"b0338499",
          4517 => x"d6157476",
          4518 => x"31555656",
          4519 => x"a00be0e0",
          4520 => x"16347575",
          4521 => x"70810557",
          4522 => x"34ff1353",
          4523 => x"72802efe",
          4524 => x"8a38a00b",
          4525 => x"e0e01634",
          4526 => x"75757081",
          4527 => x"055734ff",
          4528 => x"135372d8",
          4529 => x"38fdf439",
          4530 => x"800b84b8",
          4531 => x"f8335556",
          4532 => x"fe893983",
          4533 => x"fab61533",
          4534 => x"5984b980",
          4535 => x"19337434",
          4536 => x"84b8f733",
          4537 => x"59fca939",
          4538 => x"fc3d0d76",
          4539 => x"0284059f",
          4540 => x"05335351",
          4541 => x"7086269b",
          4542 => x"38701010",
          4543 => x"83c4fc05",
          4544 => x"51700804",
          4545 => x"84b8f833",
          4546 => x"51717127",
          4547 => x"86387183",
          4548 => x"fab53480",
          4549 => x"0b84bb84",
          4550 => x"0c863d0d",
          4551 => x"04800b83",
          4552 => x"fab53483",
          4553 => x"fab43370",
          4554 => x"81ff0654",
          4555 => x"5272802e",
          4556 => x"e238ff12",
          4557 => x"517083fa",
          4558 => x"b434800b",
          4559 => x"84bb840c",
          4560 => x"863d0d04",
          4561 => x"83fab433",
          4562 => x"70733170",
          4563 => x"09709f2c",
          4564 => x"72065455",
          4565 => x"53547083",
          4566 => x"fab434de",
          4567 => x"3983fab4",
          4568 => x"33720584",
          4569 => x"b8f733ff",
          4570 => x"11555651",
          4571 => x"70752583",
          4572 => x"38705372",
          4573 => x"83fab434",
          4574 => x"800b84bb",
          4575 => x"840c863d",
          4576 => x"0d0483fa",
          4577 => x"b5337073",
          4578 => x"31700970",
          4579 => x"9f2c7206",
          4580 => x"54565355",
          4581 => x"7083fab5",
          4582 => x"34800b84",
          4583 => x"bb840c86",
          4584 => x"3d0d0483",
          4585 => x"fab53372",
          4586 => x"0584b8f8",
          4587 => x"33ff1155",
          4588 => x"55517074",
          4589 => x"25833870",
          4590 => x"537283fa",
          4591 => x"b534800b",
          4592 => x"84bb840c",
          4593 => x"863d0d04",
          4594 => x"800b83fa",
          4595 => x"b53483fa",
          4596 => x"b43384b8",
          4597 => x"f733ff05",
          4598 => x"56527175",
          4599 => x"25feb438",
          4600 => x"81125170",
          4601 => x"83fab434",
          4602 => x"fed039ff",
          4603 => x"3d0d028f",
          4604 => x"05335170",
          4605 => x"b126b338",
          4606 => x"70101083",
          4607 => x"c5980551",
          4608 => x"70080483",
          4609 => x"fab03370",
          4610 => x"80f00671",
          4611 => x"842b80f0",
          4612 => x"06707284",
          4613 => x"2a075152",
          4614 => x"53517180",
          4615 => x"f02e0981",
          4616 => x"069c3880",
          4617 => x"f20b83fa",
          4618 => x"b034800b",
          4619 => x"84bb840c",
          4620 => x"833d0d04",
          4621 => x"83fab033",
          4622 => x"819f0690",
          4623 => x"07517083",
          4624 => x"fab03480",
          4625 => x"0b84bb84",
          4626 => x"0c833d0d",
          4627 => x"0483fab0",
          4628 => x"3380f007",
          4629 => x"517083fa",
          4630 => x"b034e839",
          4631 => x"83fab033",
          4632 => x"81fe0686",
          4633 => x"07517083",
          4634 => x"fab034d7",
          4635 => x"3980f10b",
          4636 => x"83fab034",
          4637 => x"800b84bb",
          4638 => x"840c833d",
          4639 => x"0d0483fa",
          4640 => x"b03381fc",
          4641 => x"06840751",
          4642 => x"7083fab0",
          4643 => x"34ffb439",
          4644 => x"83fab033",
          4645 => x"87075170",
          4646 => x"83fab034",
          4647 => x"ffa53983",
          4648 => x"fab03381",
          4649 => x"fd068507",
          4650 => x"517083fa",
          4651 => x"b034ff93",
          4652 => x"3983fab0",
          4653 => x"3381fb06",
          4654 => x"83075170",
          4655 => x"83fab034",
          4656 => x"ff813983",
          4657 => x"fab03381",
          4658 => x"f9068107",
          4659 => x"517083fa",
          4660 => x"b034feef",
          4661 => x"3983fab0",
          4662 => x"3381f806",
          4663 => x"517083fa",
          4664 => x"b034fedf",
          4665 => x"3983fab0",
          4666 => x"3381df06",
          4667 => x"80d00751",
          4668 => x"7083fab0",
          4669 => x"34fecc39",
          4670 => x"83fab033",
          4671 => x"81bf06b0",
          4672 => x"07517083",
          4673 => x"fab034fe",
          4674 => x"ba3983fa",
          4675 => x"b03381ef",
          4676 => x"0680e007",
          4677 => x"517083fa",
          4678 => x"b034fea7",
          4679 => x"3983fab0",
          4680 => x"3381cf06",
          4681 => x"80c00751",
          4682 => x"7083fab0",
          4683 => x"34fe9439",
          4684 => x"83fab033",
          4685 => x"81af06a0",
          4686 => x"07517083",
          4687 => x"fab034fe",
          4688 => x"823983fa",
          4689 => x"b033818f",
          4690 => x"06517083",
          4691 => x"fab034fd",
          4692 => x"f23983fa",
          4693 => x"b03381fa",
          4694 => x"06820751",
          4695 => x"7083fab0",
          4696 => x"34fde039",
          4697 => x"f33d0d02",
          4698 => x"bf053302",
          4699 => x"840580c3",
          4700 => x"053383fa",
          4701 => x"b43383fa",
          4702 => x"b33383fa",
          4703 => x"b53384b8",
          4704 => x"fa334341",
          4705 => x"5f5d5b59",
          4706 => x"78822e82",
          4707 => x"a1387882",
          4708 => x"24a53878",
          4709 => x"812e8182",
          4710 => x"387d84b8",
          4711 => x"fa34800b",
          4712 => x"84b8fc34",
          4713 => x"7a83fab4",
          4714 => x"347b83fa",
          4715 => x"b2237c83",
          4716 => x"fab5348f",
          4717 => x"3d0d0478",
          4718 => x"832e0981",
          4719 => x"06db3880",
          4720 => x"0b84b8fa",
          4721 => x"34810b84",
          4722 => x"b8fc3482",
          4723 => x"0b83fab4",
          4724 => x"34a80b83",
          4725 => x"fab53482",
          4726 => x"0b83fab2",
          4727 => x"23795884",
          4728 => x"b8f83357",
          4729 => x"84b8f733",
          4730 => x"5684b8f6",
          4731 => x"33557b54",
          4732 => x"7c537a52",
          4733 => x"83e4f851",
          4734 => x"ff808d3f",
          4735 => x"7d84b8fa",
          4736 => x"34800b84",
          4737 => x"b8fc347a",
          4738 => x"83fab434",
          4739 => x"7b83fab2",
          4740 => x"237c83fa",
          4741 => x"b5348f3d",
          4742 => x"0d04800b",
          4743 => x"84b8fa34",
          4744 => x"810b84b8",
          4745 => x"fc34800b",
          4746 => x"83fab434",
          4747 => x"a80b83fa",
          4748 => x"b534800b",
          4749 => x"83fab223",
          4750 => x"84ba8733",
          4751 => x"5884ba86",
          4752 => x"335784ba",
          4753 => x"85335679",
          4754 => x"557b547c",
          4755 => x"537a5283",
          4756 => x"e59451fe",
          4757 => x"ffb23f80",
          4758 => x"0b84ba85",
          4759 => x"335a5a79",
          4760 => x"7927a538",
          4761 => x"791084ba",
          4762 => x"d8057022",
          4763 => x"535983e5",
          4764 => x"ac51feff",
          4765 => x"933f811a",
          4766 => x"7081ff06",
          4767 => x"84ba8533",
          4768 => x"525b5978",
          4769 => x"7a26dd38",
          4770 => x"83d3b451",
          4771 => x"fefef93f",
          4772 => x"7d84b8fa",
          4773 => x"34800b84",
          4774 => x"b8fc347a",
          4775 => x"83fab434",
          4776 => x"7b83fab2",
          4777 => x"237c83fa",
          4778 => x"b5348f3d",
          4779 => x"0d04800b",
          4780 => x"84b8fa34",
          4781 => x"810b84b8",
          4782 => x"fc34810b",
          4783 => x"83fab434",
          4784 => x"a80b83fa",
          4785 => x"b534810b",
          4786 => x"83fab223",
          4787 => x"83f8e851",
          4788 => x"ff90d53f",
          4789 => x"84bb8408",
          4790 => x"5283e5b0",
          4791 => x"51fefea8",
          4792 => x"3f805983",
          4793 => x"f8e851ff",
          4794 => x"90be3f78",
          4795 => x"84bb8408",
          4796 => x"27fda638",
          4797 => x"83f8e819",
          4798 => x"335283e5",
          4799 => x"b851fefe",
          4800 => x"873f8119",
          4801 => x"7081ff06",
          4802 => x"5a5ad839",
          4803 => x"f93d0d7a",
          4804 => x"028405a7",
          4805 => x"053384b8",
          4806 => x"f83383fa",
          4807 => x"b53383fa",
          4808 => x"b4337271",
          4809 => x"291286c7",
          4810 => x"a0801183",
          4811 => x"fab22253",
          4812 => x"51595c71",
          4813 => x"7c290570",
          4814 => x"83ffff06",
          4815 => x"83f98a33",
          4816 => x"52595155",
          4817 => x"57577281",
          4818 => x"2e81e938",
          4819 => x"75892e81",
          4820 => x"f9387589",
          4821 => x"2481b938",
          4822 => x"75812e83",
          4823 => x"85387588",
          4824 => x"2e82d538",
          4825 => x"84b8f833",
          4826 => x"83fab433",
          4827 => x"83fab533",
          4828 => x"72722905",
          4829 => x"55565484",
          4830 => x"b9801633",
          4831 => x"86c7a080",
          4832 => x"143484b8",
          4833 => x"f83383fa",
          4834 => x"b53383fa",
          4835 => x"b2227271",
          4836 => x"29125a5a",
          4837 => x"56537583",
          4838 => x"fab61834",
          4839 => x"83fab433",
          4840 => x"73712916",
          4841 => x"585483fa",
          4842 => x"b03386c7",
          4843 => x"b0801834",
          4844 => x"84b8f833",
          4845 => x"7081ff06",
          4846 => x"83fab222",
          4847 => x"83fab533",
          4848 => x"72722911",
          4849 => x"575b5755",
          4850 => x"5783fab0",
          4851 => x"338499d6",
          4852 => x"14348118",
          4853 => x"7081ff06",
          4854 => x"59557378",
          4855 => x"26819938",
          4856 => x"84b8f933",
          4857 => x"587781ea",
          4858 => x"38ff1753",
          4859 => x"7283fab5",
          4860 => x"3484b8fb",
          4861 => x"33537280",
          4862 => x"2e8c3884",
          4863 => x"b8fc3357",
          4864 => x"76802e80",
          4865 => x"fb38800b",
          4866 => x"84bb840c",
          4867 => x"893d0d04",
          4868 => x"758d2e97",
          4869 => x"38758d24",
          4870 => x"80f73875",
          4871 => x"8a2e0981",
          4872 => x"06fec138",
          4873 => x"81528151",
          4874 => x"f1963f80",
          4875 => x"0b83fab5",
          4876 => x"34ffbe39",
          4877 => x"83fab615",
          4878 => x"335384b9",
          4879 => x"80133374",
          4880 => x"3475892e",
          4881 => x"098106fe",
          4882 => x"89388053",
          4883 => x"7652a051",
          4884 => x"fdba3f81",
          4885 => x"137081ff",
          4886 => x"06545472",
          4887 => x"8326ff91",
          4888 => x"387652a0",
          4889 => x"51fda53f",
          4890 => x"81137081",
          4891 => x"ff065454",
          4892 => x"837327d8",
          4893 => x"38fefa39",
          4894 => x"7483fab5",
          4895 => x"34fef239",
          4896 => x"75528351",
          4897 => x"f9de3f80",
          4898 => x"0b84bb84",
          4899 => x"0c893d0d",
          4900 => x"047580ff",
          4901 => x"2e098106",
          4902 => x"fdca3883",
          4903 => x"fab53370",
          4904 => x"81ff0655",
          4905 => x"ff055373",
          4906 => x"83387353",
          4907 => x"7283fab5",
          4908 => x"347652a0",
          4909 => x"51fcd53f",
          4910 => x"83fab533",
          4911 => x"7081ff06",
          4912 => x"55ff0553",
          4913 => x"73fea538",
          4914 => x"73537283",
          4915 => x"fab534fe",
          4916 => x"a039800b",
          4917 => x"83fab534",
          4918 => x"81528151",
          4919 => x"efe23ffe",
          4920 => x"90398052",
          4921 => x"7551efd8",
          4922 => x"3ffe8639",
          4923 => x"e63d0d02",
          4924 => x"80f30533",
          4925 => x"84ba8008",
          4926 => x"57597581",
          4927 => x"2e81b838",
          4928 => x"75822e83",
          4929 => x"8238788a",
          4930 => x"2e84b538",
          4931 => x"788a2482",
          4932 => x"d1387888",
          4933 => x"2e84b938",
          4934 => x"78892e88",
          4935 => x"8f3884b8",
          4936 => x"f83383fa",
          4937 => x"b43383fa",
          4938 => x"b5337272",
          4939 => x"2905585e",
          4940 => x"5c84b980",
          4941 => x"193386c7",
          4942 => x"a0801734",
          4943 => x"84b8f833",
          4944 => x"83fab533",
          4945 => x"83fab222",
          4946 => x"72712912",
          4947 => x"5a5a4240",
          4948 => x"7883fab6",
          4949 => x"183483fa",
          4950 => x"b4336071",
          4951 => x"29620540",
          4952 => x"5a83fab0",
          4953 => x"337f86c7",
          4954 => x"b0800534",
          4955 => x"84b8f833",
          4956 => x"7081ff06",
          4957 => x"83fab222",
          4958 => x"83fab533",
          4959 => x"72722911",
          4960 => x"42405d58",
          4961 => x"5983fab0",
          4962 => x"338499d6",
          4963 => x"1f34811d",
          4964 => x"7081ff06",
          4965 => x"42587661",
          4966 => x"2681b838",
          4967 => x"84b8f933",
          4968 => x"5a7986f1",
          4969 => x"38ff1956",
          4970 => x"7583fab5",
          4971 => x"34800b84",
          4972 => x"bb840c9c",
          4973 => x"3d0d0478",
          4974 => x"b72e848a",
          4975 => x"38b77925",
          4976 => x"81fd3878",
          4977 => x"b82e9bb3",
          4978 => x"387880db",
          4979 => x"2e89cc38",
          4980 => x"800b84ba",
          4981 => x"800c84b8",
          4982 => x"f83383fa",
          4983 => x"b43383fa",
          4984 => x"b5337272",
          4985 => x"29055e40",
          4986 => x"4084b980",
          4987 => x"193386c7",
          4988 => x"a0801d34",
          4989 => x"84b8f833",
          4990 => x"83fab533",
          4991 => x"83fab222",
          4992 => x"72712912",
          4993 => x"415f5956",
          4994 => x"7883fab6",
          4995 => x"1f3483fa",
          4996 => x"b4337671",
          4997 => x"29195b57",
          4998 => x"83fab033",
          4999 => x"86c7b080",
          5000 => x"1b3484b8",
          5001 => x"f8337081",
          5002 => x"ff0683fa",
          5003 => x"b22283fa",
          5004 => x"b5337272",
          5005 => x"29114442",
          5006 => x"43585983",
          5007 => x"fab03360",
          5008 => x"8499d605",
          5009 => x"34811f58",
          5010 => x"7781ff06",
          5011 => x"41607727",
          5012 => x"feca3877",
          5013 => x"83fab534",
          5014 => x"800b84bb",
          5015 => x"840c9c3d",
          5016 => x"0d04789b",
          5017 => x"2e82b738",
          5018 => x"789b2483",
          5019 => x"8138788d",
          5020 => x"2e098106",
          5021 => x"fda83880",
          5022 => x"0b83fab5",
          5023 => x"34800b84",
          5024 => x"bb840c9c",
          5025 => x"3d0d0478",
          5026 => x"9b2e82aa",
          5027 => x"38d01956",
          5028 => x"75892684",
          5029 => x"d03884ba",
          5030 => x"84338111",
          5031 => x"59577784",
          5032 => x"ba843478",
          5033 => x"84ba8818",
          5034 => x"347781ff",
          5035 => x"0659800b",
          5036 => x"84ba881a",
          5037 => x"34800b84",
          5038 => x"bb840c9c",
          5039 => x"3d0d0478",
          5040 => x"9b2efde9",
          5041 => x"38800b84",
          5042 => x"ba800c84",
          5043 => x"b8f83383",
          5044 => x"fab43383",
          5045 => x"fab53372",
          5046 => x"7229055e",
          5047 => x"404084b9",
          5048 => x"80193386",
          5049 => x"c7a0801d",
          5050 => x"3484b8f8",
          5051 => x"3383fab5",
          5052 => x"3383fab2",
          5053 => x"22727129",
          5054 => x"12415f59",
          5055 => x"567883fa",
          5056 => x"b61f3483",
          5057 => x"fab43376",
          5058 => x"7129195b",
          5059 => x"5783fab0",
          5060 => x"3386c7b0",
          5061 => x"801b3484",
          5062 => x"b8f83370",
          5063 => x"81ff0683",
          5064 => x"fab22283",
          5065 => x"fab53372",
          5066 => x"72291144",
          5067 => x"42435859",
          5068 => x"83fab033",
          5069 => x"608499d6",
          5070 => x"0534811f",
          5071 => x"58fe8939",
          5072 => x"81528151",
          5073 => x"eafa3f80",
          5074 => x"0b83fab5",
          5075 => x"34feae39",
          5076 => x"84b8f833",
          5077 => x"83fab533",
          5078 => x"7081ff06",
          5079 => x"83fab433",
          5080 => x"73712912",
          5081 => x"86c7a080",
          5082 => x"0583fab2",
          5083 => x"2240515d",
          5084 => x"727e2905",
          5085 => x"7083ffff",
          5086 => x"0683f98a",
          5087 => x"335a5159",
          5088 => x"5a5c7581",
          5089 => x"2e86a438",
          5090 => x"7881ff06",
          5091 => x"ff1a5757",
          5092 => x"76fc9538",
          5093 => x"76567583",
          5094 => x"fab534fc",
          5095 => x"9039800b",
          5096 => x"84ba8434",
          5097 => x"800b84ba",
          5098 => x"8534800b",
          5099 => x"84ba8634",
          5100 => x"800b84ba",
          5101 => x"8734810b",
          5102 => x"84ba800c",
          5103 => x"800b84bb",
          5104 => x"840c9c3d",
          5105 => x"0d0483fa",
          5106 => x"b43384ba",
          5107 => x"ec3483fa",
          5108 => x"b53384ba",
          5109 => x"ed3483fa",
          5110 => x"b33384ba",
          5111 => x"ee34800b",
          5112 => x"84ba800c",
          5113 => x"800b84bb",
          5114 => x"840c9c3d",
          5115 => x"0d047880",
          5116 => x"ff2e0981",
          5117 => x"06faa738",
          5118 => x"83fab433",
          5119 => x"84b8f833",
          5120 => x"7081ff06",
          5121 => x"83fab533",
          5122 => x"7081ff06",
          5123 => x"72752911",
          5124 => x"86c7a080",
          5125 => x"0583fab2",
          5126 => x"225c4072",
          5127 => x"7b290570",
          5128 => x"83ffff06",
          5129 => x"83f98a33",
          5130 => x"445c435c",
          5131 => x"425b5c7d",
          5132 => x"812e85fe",
          5133 => x"387881ff",
          5134 => x"06ff1a58",
          5135 => x"56758338",
          5136 => x"75577683",
          5137 => x"fab5347b",
          5138 => x"81ff067a",
          5139 => x"81ff0678",
          5140 => x"81ff0672",
          5141 => x"7229055f",
          5142 => x"405b84b9",
          5143 => x"a03386c7",
          5144 => x"a0801e34",
          5145 => x"84b8f833",
          5146 => x"83fab533",
          5147 => x"83fab222",
          5148 => x"72712912",
          5149 => x"5a5e4240",
          5150 => x"a00b83fa",
          5151 => x"b6183483",
          5152 => x"fab43360",
          5153 => x"71296205",
          5154 => x"5a5683fa",
          5155 => x"b03386c7",
          5156 => x"b0801a34",
          5157 => x"84b8f833",
          5158 => x"7081ff06",
          5159 => x"83fab222",
          5160 => x"83fab533",
          5161 => x"72722911",
          5162 => x"435d5a5e",
          5163 => x"5983fab0",
          5164 => x"337f8499",
          5165 => x"d6053481",
          5166 => x"1a7081ff",
          5167 => x"065c587c",
          5168 => x"7b2695ea",
          5169 => x"3884b8f9",
          5170 => x"335a7996",
          5171 => x"d038ff19",
          5172 => x"587783fa",
          5173 => x"b53483fa",
          5174 => x"b5337081",
          5175 => x"ff0658ff",
          5176 => x"0556fdac",
          5177 => x"3978bb2e",
          5178 => x"95d83878",
          5179 => x"bd2e83d7",
          5180 => x"3878bf2e",
          5181 => x"95a83884",
          5182 => x"ba84335f",
          5183 => x"7e83f938",
          5184 => x"ffbf1956",
          5185 => x"75b42684",
          5186 => x"c8387510",
          5187 => x"1083c6e0",
          5188 => x"05587708",
          5189 => x"04800b83",
          5190 => x"fab53480",
          5191 => x"528151e7",
          5192 => x"9f3f800b",
          5193 => x"84bb840c",
          5194 => x"9c3d0d04",
          5195 => x"83fab433",
          5196 => x"84b8f833",
          5197 => x"7081ff06",
          5198 => x"83fab533",
          5199 => x"7081ff06",
          5200 => x"72752911",
          5201 => x"86c7a080",
          5202 => x"0583fab2",
          5203 => x"225c4172",
          5204 => x"7b290570",
          5205 => x"83ffff06",
          5206 => x"83f98a33",
          5207 => x"4653455c",
          5208 => x"595b5b7f",
          5209 => x"812e82ef",
          5210 => x"38805c7a",
          5211 => x"81ff067a",
          5212 => x"81ff067a",
          5213 => x"81ff0672",
          5214 => x"7229055c",
          5215 => x"584084b9",
          5216 => x"a03386c7",
          5217 => x"a0801b34",
          5218 => x"84b8f833",
          5219 => x"83fab533",
          5220 => x"83fab222",
          5221 => x"72712912",
          5222 => x"5e415e56",
          5223 => x"a00b83fa",
          5224 => x"b61c3483",
          5225 => x"fab43376",
          5226 => x"71291e5a",
          5227 => x"5e83fab0",
          5228 => x"3386c7b0",
          5229 => x"801a3484",
          5230 => x"b8f83370",
          5231 => x"81ff0683",
          5232 => x"fab22283",
          5233 => x"fab53372",
          5234 => x"7229115b",
          5235 => x"445a4059",
          5236 => x"83fab033",
          5237 => x"8499d618",
          5238 => x"34608105",
          5239 => x"7081ff06",
          5240 => x"5b587e7a",
          5241 => x"2681ac38",
          5242 => x"84b8f933",
          5243 => x"587792fb",
          5244 => x"38ff1956",
          5245 => x"7583fab5",
          5246 => x"34811c70",
          5247 => x"81ff065d",
          5248 => x"597b8326",
          5249 => x"f7a73883",
          5250 => x"fab43384",
          5251 => x"b8f83383",
          5252 => x"fab53372",
          5253 => x"81ff0672",
          5254 => x"81ff0672",
          5255 => x"81ff0672",
          5256 => x"72290554",
          5257 => x"5b435b5b",
          5258 => x"5b84b9a0",
          5259 => x"3386c7a0",
          5260 => x"801b3484",
          5261 => x"b8f83383",
          5262 => x"fab53383",
          5263 => x"fab22272",
          5264 => x"7129125e",
          5265 => x"415e56a0",
          5266 => x"0b83fab6",
          5267 => x"1c3483fa",
          5268 => x"b4337671",
          5269 => x"291e5a5e",
          5270 => x"83fab033",
          5271 => x"86c7b080",
          5272 => x"1a3484b8",
          5273 => x"f8337081",
          5274 => x"ff0683fa",
          5275 => x"b22283fa",
          5276 => x"b5337272",
          5277 => x"29115b44",
          5278 => x"5a405983",
          5279 => x"fab03384",
          5280 => x"99d61834",
          5281 => x"60810570",
          5282 => x"81ff065b",
          5283 => x"58797f27",
          5284 => x"fed63877",
          5285 => x"83fab534",
          5286 => x"fedf3982",
          5287 => x"0b84ba80",
          5288 => x"0c800b84",
          5289 => x"bb840c9c",
          5290 => x"3d0d0483",
          5291 => x"fab61733",
          5292 => x"5984b980",
          5293 => x"19337a34",
          5294 => x"83fab533",
          5295 => x"7081ff06",
          5296 => x"58ff0556",
          5297 => x"f9ca3981",
          5298 => x"0b84ba86",
          5299 => x"34800b84",
          5300 => x"bb840c9c",
          5301 => x"3d0d0483",
          5302 => x"fab61733",
          5303 => x"5b84b980",
          5304 => x"1b337c34",
          5305 => x"83fab433",
          5306 => x"84b8f833",
          5307 => x"83fab533",
          5308 => x"5b5b5b80",
          5309 => x"5cfcf439",
          5310 => x"84ba8842",
          5311 => x"9c3ddc11",
          5312 => x"53d80551",
          5313 => x"ff88ff3f",
          5314 => x"84bb8408",
          5315 => x"802efbf0",
          5316 => x"3884ba85",
          5317 => x"33811157",
          5318 => x"5a7584ba",
          5319 => x"85347910",
          5320 => x"83fe0641",
          5321 => x"0280ca05",
          5322 => x"226184ba",
          5323 => x"d80523fb",
          5324 => x"cf3983fa",
          5325 => x"b617335c",
          5326 => x"84b9801c",
          5327 => x"337b3483",
          5328 => x"fab43384",
          5329 => x"b8f83383",
          5330 => x"fab5335b",
          5331 => x"5b5cf9e5",
          5332 => x"3984b8f8",
          5333 => x"3383fab4",
          5334 => x"3383fab5",
          5335 => x"33727229",
          5336 => x"05415d5b",
          5337 => x"84b98019",
          5338 => x"337f86c7",
          5339 => x"a0800534",
          5340 => x"84b8f833",
          5341 => x"83fab533",
          5342 => x"83fab222",
          5343 => x"72712912",
          5344 => x"5a435b56",
          5345 => x"7883fab6",
          5346 => x"183483fa",
          5347 => x"b4337671",
          5348 => x"291b415e",
          5349 => x"83fab033",
          5350 => x"6086c7b0",
          5351 => x"80053484",
          5352 => x"b8f83370",
          5353 => x"81ff0683",
          5354 => x"fab22283",
          5355 => x"fab53372",
          5356 => x"72291141",
          5357 => x"5f5a425a",
          5358 => x"83fab033",
          5359 => x"8499d61e",
          5360 => x"34811c70",
          5361 => x"81ff065c",
          5362 => x"58607b26",
          5363 => x"90a23884",
          5364 => x"b8f93358",
          5365 => x"7790e238",
          5366 => x"ff1a5675",
          5367 => x"83fab534",
          5368 => x"800b84ba",
          5369 => x"800c84b8",
          5370 => x"fb33407f",
          5371 => x"802ef3bd",
          5372 => x"3884b8fc",
          5373 => x"335675f3",
          5374 => x"b4387852",
          5375 => x"8151eae4",
          5376 => x"3f800b84",
          5377 => x"bb840c9c",
          5378 => x"3d0d0484",
          5379 => x"baec3383",
          5380 => x"fab43484",
          5381 => x"baed3383",
          5382 => x"fab53484",
          5383 => x"baee3357",
          5384 => x"7683fab2",
          5385 => x"23ffb939",
          5386 => x"83fab433",
          5387 => x"84baec34",
          5388 => x"83fab533",
          5389 => x"84baed34",
          5390 => x"83fab333",
          5391 => x"84baee34",
          5392 => x"ff9e3984",
          5393 => x"ba85335b",
          5394 => x"7a802eff",
          5395 => x"933884ba",
          5396 => x"d8225d7c",
          5397 => x"862e0981",
          5398 => x"06ff8538",
          5399 => x"83fab533",
          5400 => x"81055583",
          5401 => x"fab43381",
          5402 => x"05549b53",
          5403 => x"83e5c052",
          5404 => x"943d7052",
          5405 => x"57feecb0",
          5406 => x"3f7651fe",
          5407 => x"fdaa3f84",
          5408 => x"bb840881",
          5409 => x"ff0683f9",
          5410 => x"88335776",
          5411 => x"054160a0",
          5412 => x"24fecd38",
          5413 => x"765283f8",
          5414 => x"e851fefb",
          5415 => x"f53ffec0",
          5416 => x"39800b84",
          5417 => x"ba85335b",
          5418 => x"587981ff",
          5419 => x"065b777b",
          5420 => x"27fead38",
          5421 => x"771084ba",
          5422 => x"d8058111",
          5423 => x"33574175",
          5424 => x"b1268aa5",
          5425 => x"38751010",
          5426 => x"83c8b405",
          5427 => x"5f7e0804",
          5428 => x"84ba8533",
          5429 => x"5e7d802e",
          5430 => x"8fa43883",
          5431 => x"fab43384",
          5432 => x"bad93371",
          5433 => x"71317009",
          5434 => x"709f2c72",
          5435 => x"065a4259",
          5436 => x"5e5c7583",
          5437 => x"fab434fd",
          5438 => x"e73984ba",
          5439 => x"85335675",
          5440 => x"802e8ee7",
          5441 => x"3884bad9",
          5442 => x"33ff0570",
          5443 => x"81ff0684",
          5444 => x"b8f8335d",
          5445 => x"575f757b",
          5446 => x"27fdc538",
          5447 => x"7583fab5",
          5448 => x"34fdbd39",
          5449 => x"800b83fa",
          5450 => x"b53483fa",
          5451 => x"b4337081",
          5452 => x"ff065d57",
          5453 => x"7b802efd",
          5454 => x"a738ff17",
          5455 => x"567583fa",
          5456 => x"b434fd9c",
          5457 => x"39800b83",
          5458 => x"fab53483",
          5459 => x"fab43384",
          5460 => x"b8f733ff",
          5461 => x"05575776",
          5462 => x"7625fd84",
          5463 => x"38811756",
          5464 => x"7583fab4",
          5465 => x"34fcf939",
          5466 => x"84ba8533",
          5467 => x"407f802e",
          5468 => x"8de03883",
          5469 => x"fab53384",
          5470 => x"bad93371",
          5471 => x"71317009",
          5472 => x"709f2c72",
          5473 => x"065a4159",
          5474 => x"425a7583",
          5475 => x"fab534fc",
          5476 => x"cf3984ba",
          5477 => x"85335b7a",
          5478 => x"802efcc4",
          5479 => x"3884bad8",
          5480 => x"22416099",
          5481 => x"2e098106",
          5482 => x"fcb63884",
          5483 => x"b8f83383",
          5484 => x"fab53383",
          5485 => x"fab43372",
          5486 => x"71291286",
          5487 => x"c7a08011",
          5488 => x"83fab222",
          5489 => x"43515a58",
          5490 => x"71602905",
          5491 => x"7083ffff",
          5492 => x"0683f988",
          5493 => x"0887fffe",
          5494 => x"8006425a",
          5495 => x"5d5d7e84",
          5496 => x"82802e92",
          5497 => x"bf38800b",
          5498 => x"83f98934",
          5499 => x"fbf23984",
          5500 => x"ba85335a",
          5501 => x"79802efb",
          5502 => x"e73884ba",
          5503 => x"d8225877",
          5504 => x"992e0981",
          5505 => x"06fbd938",
          5506 => x"810b83f9",
          5507 => x"8934fbd0",
          5508 => x"3984ba85",
          5509 => x"33567580",
          5510 => x"2e90be38",
          5511 => x"84bad933",
          5512 => x"83fab533",
          5513 => x"5d7c0584",
          5514 => x"b8f833ff",
          5515 => x"11595e56",
          5516 => x"757d2583",
          5517 => x"38755776",
          5518 => x"83fab534",
          5519 => x"fba23984",
          5520 => x"ba853357",
          5521 => x"76802e8c",
          5522 => x"c83884ba",
          5523 => x"d93383fa",
          5524 => x"b4334261",
          5525 => x"0584b8f7",
          5526 => x"33ff1159",
          5527 => x"41567560",
          5528 => x"25833875",
          5529 => x"577683fa",
          5530 => x"b434faf4",
          5531 => x"3983e5cc",
          5532 => x"51fee794",
          5533 => x"3f800b84",
          5534 => x"ba853357",
          5535 => x"57767627",
          5536 => x"8bc73876",
          5537 => x"1084bad8",
          5538 => x"05702253",
          5539 => x"5a83e5ac",
          5540 => x"51fee6f4",
          5541 => x"3f811770",
          5542 => x"81ff0684",
          5543 => x"ba853358",
          5544 => x"5858da39",
          5545 => x"820b84ba",
          5546 => x"85335f57",
          5547 => x"7d802e8d",
          5548 => x"3884bad8",
          5549 => x"22567583",
          5550 => x"26833875",
          5551 => x"57815276",
          5552 => x"81ff0651",
          5553 => x"d5f33ffa",
          5554 => x"973984ba",
          5555 => x"85335781",
          5556 => x"77278eb7",
          5557 => x"3884badb",
          5558 => x"33ff0570",
          5559 => x"81ff0684",
          5560 => x"bad933ff",
          5561 => x"057081ff",
          5562 => x"0684b8f7",
          5563 => x"337081ff",
          5564 => x"06ff1140",
          5565 => x"43525b59",
          5566 => x"5c5c777e",
          5567 => x"27833877",
          5568 => x"5a7983fa",
          5569 => x"b2237681",
          5570 => x"ff06ff18",
          5571 => x"585f777f",
          5572 => x"27833877",
          5573 => x"577683fa",
          5574 => x"b43484b8",
          5575 => x"f833ff11",
          5576 => x"57407a60",
          5577 => x"27f9b438",
          5578 => x"7a567583",
          5579 => x"fab534f9",
          5580 => x"af3984ba",
          5581 => x"85335f7e",
          5582 => x"802e8aef",
          5583 => x"3884bad9",
          5584 => x"3384b8f7",
          5585 => x"33405b7a",
          5586 => x"7f26f994",
          5587 => x"3883fab4",
          5588 => x"3384b8f8",
          5589 => x"337081ff",
          5590 => x"0683fab5",
          5591 => x"33717429",
          5592 => x"1186c7a0",
          5593 => x"800583fa",
          5594 => x"b2225f40",
          5595 => x"717e2905",
          5596 => x"7083ffff",
          5597 => x"0683f98a",
          5598 => x"33465259",
          5599 => x"595f5d60",
          5600 => x"812e84f0",
          5601 => x"387983ff",
          5602 => x"ff06707c",
          5603 => x"315d5780",
          5604 => x"7c248efe",
          5605 => x"3884b8f7",
          5606 => x"33567676",
          5607 => x"278ed638",
          5608 => x"ff165675",
          5609 => x"83fab223",
          5610 => x"7c81ff06",
          5611 => x"707c3141",
          5612 => x"57806024",
          5613 => x"8ee53884",
          5614 => x"b8f73356",
          5615 => x"7676278d",
          5616 => x"ee38ff16",
          5617 => x"567583fa",
          5618 => x"b4347e81",
          5619 => x"ff0683fa",
          5620 => x"b2225757",
          5621 => x"805a7676",
          5622 => x"26903875",
          5623 => x"77318105",
          5624 => x"7e81ff06",
          5625 => x"7171295c",
          5626 => x"5e5b7958",
          5627 => x"86c7a080",
          5628 => x"5b86c7b0",
          5629 => x"807f81ff",
          5630 => x"067f81ff",
          5631 => x"06717129",
          5632 => x"1d425842",
          5633 => x"5c797f27",
          5634 => x"f7d63884",
          5635 => x"99d61a57",
          5636 => x"e0e01733",
          5637 => x"5f84b980",
          5638 => x"1f337b70",
          5639 => x"81055d34",
          5640 => x"76708105",
          5641 => x"58337c70",
          5642 => x"81055e34",
          5643 => x"811884b8",
          5644 => x"f83384b8",
          5645 => x"f7337171",
          5646 => x"291d4340",
          5647 => x"5e587760",
          5648 => x"27f79d38",
          5649 => x"e0e01733",
          5650 => x"5f84b980",
          5651 => x"1f337b70",
          5652 => x"81055d34",
          5653 => x"76708105",
          5654 => x"58337c70",
          5655 => x"81055e34",
          5656 => x"811884b8",
          5657 => x"f83384b8",
          5658 => x"f7337171",
          5659 => x"291d4340",
          5660 => x"5e587f78",
          5661 => x"26ff9938",
          5662 => x"f6e63984",
          5663 => x"ba853356",
          5664 => x"75802e87",
          5665 => x"e0388052",
          5666 => x"84bad933",
          5667 => x"51d8b13f",
          5668 => x"f6ce3980",
          5669 => x"0b84b8f8",
          5670 => x"33ff1184",
          5671 => x"ba85335d",
          5672 => x"59405879",
          5673 => x"782e9438",
          5674 => x"84bad822",
          5675 => x"5675782e",
          5676 => x"0981068b",
          5677 => x"be3883fa",
          5678 => x"b5335876",
          5679 => x"81ff0683",
          5680 => x"fab43379",
          5681 => x"435c5c76",
          5682 => x"ff2e81ed",
          5683 => x"3884b8f7",
          5684 => x"33407a60",
          5685 => x"26f68938",
          5686 => x"7e81ff06",
          5687 => x"56607626",
          5688 => x"f5fe387b",
          5689 => x"7626617d",
          5690 => x"27075776",
          5691 => x"f5f2387a",
          5692 => x"10101b70",
          5693 => x"90296205",
          5694 => x"86c7a080",
          5695 => x"11701f5d",
          5696 => x"5a86c7b0",
          5697 => x"80057983",
          5698 => x"0658515d",
          5699 => x"758bac38",
          5700 => x"79830657",
          5701 => x"768ba438",
          5702 => x"83fab033",
          5703 => x"70982b71",
          5704 => x"902b0771",
          5705 => x"882b0771",
          5706 => x"07797f59",
          5707 => x"525f5777",
          5708 => x"7a279e38",
          5709 => x"80777084",
          5710 => x"05590c7d",
          5711 => x"76708405",
          5712 => x"580c7977",
          5713 => x"26ee3884",
          5714 => x"b8f83384",
          5715 => x"b8f73341",
          5716 => x"5f7e81ff",
          5717 => x"066081ff",
          5718 => x"0683fab2",
          5719 => x"227d7329",
          5720 => x"64055959",
          5721 => x"595a7777",
          5722 => x"268c3876",
          5723 => x"78311b70",
          5724 => x"7b296205",
          5725 => x"57407576",
          5726 => x"1d575776",
          5727 => x"7626f4e0",
          5728 => x"3883fab0",
          5729 => x"338499d6",
          5730 => x"18595aa0",
          5731 => x"0be0e019",
          5732 => x"34797870",
          5733 => x"81055a34",
          5734 => x"81175776",
          5735 => x"7626f4c0",
          5736 => x"38a00be0",
          5737 => x"e0193479",
          5738 => x"78708105",
          5739 => x"5a348117",
          5740 => x"57757727",
          5741 => x"d638f4a8",
          5742 => x"39ff1f70",
          5743 => x"81ff065d",
          5744 => x"58fe8a39",
          5745 => x"83fab033",
          5746 => x"7080f006",
          5747 => x"71842b80",
          5748 => x"f0067184",
          5749 => x"2a07585d",
          5750 => x"577b80f0",
          5751 => x"2e098106",
          5752 => x"be3880f2",
          5753 => x"0b83fab0",
          5754 => x"34811870",
          5755 => x"81ff0659",
          5756 => x"56f5b639",
          5757 => x"83fab617",
          5758 => x"335e84b9",
          5759 => x"801e337c",
          5760 => x"3483fab4",
          5761 => x"3384b8f8",
          5762 => x"3383fab2",
          5763 => x"2284b8f7",
          5764 => x"33425c5f",
          5765 => x"5dfaee39",
          5766 => x"83fab033",
          5767 => x"87075675",
          5768 => x"83fab034",
          5769 => x"81187081",
          5770 => x"ff065956",
          5771 => x"f4fb3983",
          5772 => x"fab03381",
          5773 => x"fd068507",
          5774 => x"567583fa",
          5775 => x"b034e539",
          5776 => x"83fab033",
          5777 => x"81fb0683",
          5778 => x"07567583",
          5779 => x"fab034d4",
          5780 => x"3983fab0",
          5781 => x"3381f906",
          5782 => x"81075675",
          5783 => x"83fab034",
          5784 => x"c33983fa",
          5785 => x"b033819f",
          5786 => x"06900756",
          5787 => x"7583fab0",
          5788 => x"34ffb139",
          5789 => x"80f10b83",
          5790 => x"fab03481",
          5791 => x"187081ff",
          5792 => x"065956f4",
          5793 => x"a43983fa",
          5794 => x"b033818f",
          5795 => x"06567583",
          5796 => x"fab034ff",
          5797 => x"8f3983fa",
          5798 => x"b033819f",
          5799 => x"06900756",
          5800 => x"7583fab0",
          5801 => x"34fefd39",
          5802 => x"83fab033",
          5803 => x"81ef0680",
          5804 => x"e0075675",
          5805 => x"83fab034",
          5806 => x"feea3983",
          5807 => x"fab03381",
          5808 => x"cf0680c0",
          5809 => x"07567583",
          5810 => x"fab034fe",
          5811 => x"d73983fa",
          5812 => x"b03381af",
          5813 => x"06a00756",
          5814 => x"7583fab0",
          5815 => x"34fec539",
          5816 => x"83fab033",
          5817 => x"81fe0686",
          5818 => x"07567583",
          5819 => x"fab034fe",
          5820 => x"b33983fa",
          5821 => x"b03381fc",
          5822 => x"06840756",
          5823 => x"7583fab0",
          5824 => x"34fea139",
          5825 => x"83fab033",
          5826 => x"81fa0682",
          5827 => x"07567583",
          5828 => x"fab034fe",
          5829 => x"8f3983fa",
          5830 => x"b03381f8",
          5831 => x"06567583",
          5832 => x"fab034fd",
          5833 => x"ff3983fa",
          5834 => x"b03380f0",
          5835 => x"07567583",
          5836 => x"fab034fd",
          5837 => x"ef3983fa",
          5838 => x"b03380f0",
          5839 => x"07567583",
          5840 => x"fab034fd",
          5841 => x"df3983fa",
          5842 => x"b03381df",
          5843 => x"0680d007",
          5844 => x"567583fa",
          5845 => x"b034fdcc",
          5846 => x"3983fab0",
          5847 => x"3381bf06",
          5848 => x"b0075675",
          5849 => x"83fab034",
          5850 => x"fdba3980",
          5851 => x"0b83fab5",
          5852 => x"34805281",
          5853 => x"51d2c93f",
          5854 => x"ecff3984",
          5855 => x"baec3383",
          5856 => x"fab43484",
          5857 => x"baed3383",
          5858 => x"fab53484",
          5859 => x"baee3359",
          5860 => x"7883fab2",
          5861 => x"23800b84",
          5862 => x"ba800ce8",
          5863 => x"c739810b",
          5864 => x"84ba8734",
          5865 => x"800b84bb",
          5866 => x"840c9c3d",
          5867 => x"0d047783",
          5868 => x"fab53483",
          5869 => x"fab53370",
          5870 => x"81ff0658",
          5871 => x"ff0556e7",
          5872 => x"cf3984ba",
          5873 => x"88429c3d",
          5874 => x"dc1153d8",
          5875 => x"0551fef7",
          5876 => x"b53f84bb",
          5877 => x"8408a138",
          5878 => x"84bb8408",
          5879 => x"84ba800c",
          5880 => x"800b84ba",
          5881 => x"8434800b",
          5882 => x"84bb840c",
          5883 => x"9c3d0d04",
          5884 => x"7783fab5",
          5885 => x"34efe939",
          5886 => x"84ba8533",
          5887 => x"81115c5c",
          5888 => x"7a84ba85",
          5889 => x"347b1083",
          5890 => x"fe065d02",
          5891 => x"80ca0522",
          5892 => x"84bad81e",
          5893 => x"23800b84",
          5894 => x"ba8434ca",
          5895 => x"39800b83",
          5896 => x"fab53480",
          5897 => x"528151d1",
          5898 => x"973f83fa",
          5899 => x"b5337081",
          5900 => x"ff0658ff",
          5901 => x"0556e6d8",
          5902 => x"39800b83",
          5903 => x"fab53480",
          5904 => x"528151d0",
          5905 => x"fb3fef98",
          5906 => x"398a51fe",
          5907 => x"ea903fef",
          5908 => x"8f3983fa",
          5909 => x"b533ff05",
          5910 => x"7009709f",
          5911 => x"2c720658",
          5912 => x"5f57f2a6",
          5913 => x"39755281",
          5914 => x"51d93984",
          5915 => x"b8f83340",
          5916 => x"756027ee",
          5917 => x"eb387583",
          5918 => x"fab534ee",
          5919 => x"e33983fa",
          5920 => x"b433ff05",
          5921 => x"7009709f",
          5922 => x"2c720658",
          5923 => x"4057f0e2",
          5924 => x"3983fab4",
          5925 => x"33810584",
          5926 => x"b8f733ff",
          5927 => x"11595956",
          5928 => x"757825f3",
          5929 => x"c0387557",
          5930 => x"f3bb3984",
          5931 => x"b8f73370",
          5932 => x"81ff0658",
          5933 => x"5c817726",
          5934 => x"eea63883",
          5935 => x"fab43384",
          5936 => x"b8f83370",
          5937 => x"81ff0683",
          5938 => x"fab53371",
          5939 => x"74291186",
          5940 => x"c7a08005",
          5941 => x"83fab222",
          5942 => x"5f5f717e",
          5943 => x"29057083",
          5944 => x"ffff0683",
          5945 => x"f98a335d",
          5946 => x"5b44425f",
          5947 => x"5d77812e",
          5948 => x"81f53879",
          5949 => x"83ffff06",
          5950 => x"ff115c57",
          5951 => x"807b2484",
          5952 => x"893884b8",
          5953 => x"f7335676",
          5954 => x"76278398",
          5955 => x"38ff1656",
          5956 => x"7583fab2",
          5957 => x"237c81ff",
          5958 => x"06ff1157",
          5959 => x"57807624",
          5960 => x"83df3884",
          5961 => x"b8f73356",
          5962 => x"76762782",
          5963 => x"ec38ff16",
          5964 => x"567583fa",
          5965 => x"b4347b81",
          5966 => x"ff0683fa",
          5967 => x"b2225757",
          5968 => x"805a7676",
          5969 => x"26903875",
          5970 => x"77318105",
          5971 => x"7e81ff06",
          5972 => x"7171295c",
          5973 => x"5e5f7958",
          5974 => x"86c7a080",
          5975 => x"5b86c7b0",
          5976 => x"807c81ff",
          5977 => x"067f81ff",
          5978 => x"06717129",
          5979 => x"1d414242",
          5980 => x"5d797e27",
          5981 => x"ecea3884",
          5982 => x"99d61a57",
          5983 => x"e0e01733",
          5984 => x"5e84b980",
          5985 => x"1e337b70",
          5986 => x"81055d34",
          5987 => x"76708105",
          5988 => x"58337d70",
          5989 => x"81055f34",
          5990 => x"811884b8",
          5991 => x"f83384b8",
          5992 => x"f7337171",
          5993 => x"291d5941",
          5994 => x"5d587776",
          5995 => x"27ecb138",
          5996 => x"e0e01733",
          5997 => x"5e84b980",
          5998 => x"1e337b70",
          5999 => x"81055d34",
          6000 => x"76708105",
          6001 => x"58337d70",
          6002 => x"81055f34",
          6003 => x"811884b8",
          6004 => x"f83384b8",
          6005 => x"f7337171",
          6006 => x"291d5941",
          6007 => x"5d587578",
          6008 => x"26ff9938",
          6009 => x"ebfa3983",
          6010 => x"fab61733",
          6011 => x"5c84b980",
          6012 => x"1c337b34",
          6013 => x"83fab433",
          6014 => x"84b8f833",
          6015 => x"83fab222",
          6016 => x"84b8f733",
          6017 => x"5f5c5f5d",
          6018 => x"fde93976",
          6019 => x"ebd23884",
          6020 => x"b8f73370",
          6021 => x"81ff06ff",
          6022 => x"115c4258",
          6023 => x"76612783",
          6024 => x"38765a79",
          6025 => x"83fab223",
          6026 => x"7781ff06",
          6027 => x"ff19585a",
          6028 => x"807a2783",
          6029 => x"38805776",
          6030 => x"83fab434",
          6031 => x"84b8f833",
          6032 => x"7081ff06",
          6033 => x"ff125259",
          6034 => x"56807827",
          6035 => x"eb8d3880",
          6036 => x"567583fa",
          6037 => x"b534eb88",
          6038 => x"3983fab5",
          6039 => x"33810584",
          6040 => x"b8f833ff",
          6041 => x"11594056",
          6042 => x"757f25ef",
          6043 => x"ca387557",
          6044 => x"efc53975",
          6045 => x"812e0981",
          6046 => x"06f4c038",
          6047 => x"83fab533",
          6048 => x"7081ff06",
          6049 => x"83fab433",
          6050 => x"7a445d5d",
          6051 => x"5776ff2e",
          6052 => x"098106f4",
          6053 => x"b838f6a1",
          6054 => x"39ff1d56",
          6055 => x"7583fab4",
          6056 => x"34fd9339",
          6057 => x"ff1a5675",
          6058 => x"83fab223",
          6059 => x"fce7397c",
          6060 => x"7b315675",
          6061 => x"83fab434",
          6062 => x"f2903977",
          6063 => x"7d585677",
          6064 => x"7a26f58d",
          6065 => x"38807670",
          6066 => x"81055834",
          6067 => x"83fab033",
          6068 => x"77708105",
          6069 => x"5934757a",
          6070 => x"26f4ec38",
          6071 => x"80767081",
          6072 => x"05583483",
          6073 => x"fab03377",
          6074 => x"70810559",
          6075 => x"34797627",
          6076 => x"d438f4d3",
          6077 => x"39797b31",
          6078 => x"567583fa",
          6079 => x"b223f1a8",
          6080 => x"39800b83",
          6081 => x"fab434fc",
          6082 => x"ad397e83",
          6083 => x"fab223fc",
          6084 => x"8439800b",
          6085 => x"83fab223",
          6086 => x"f18e3980",
          6087 => x"0b83fab4",
          6088 => x"34f1a739",
          6089 => x"83fab618",
          6090 => x"335a84b9",
          6091 => x"801a3377",
          6092 => x"34800b83",
          6093 => x"f98934e9",
          6094 => x"a739fd3d",
          6095 => x"0d029705",
          6096 => x"3384b8fa",
          6097 => x"33545472",
          6098 => x"802e9038",
          6099 => x"7351db9c",
          6100 => x"3f800b84",
          6101 => x"bb840c85",
          6102 => x"3d0d0476",
          6103 => x"527351d7",
          6104 => x"ab3f800b",
          6105 => x"84bb840c",
          6106 => x"853d0d04",
          6107 => x"f33d0d02",
          6108 => x"bf05335c",
          6109 => x"ff0b83f9",
          6110 => x"88337081",
          6111 => x"ff0683f8",
          6112 => x"e8113358",
          6113 => x"55555974",
          6114 => x"802e80d6",
          6115 => x"38811456",
          6116 => x"7583f988",
          6117 => x"34745978",
          6118 => x"84bb840c",
          6119 => x"8f3d0d04",
          6120 => x"83f8e408",
          6121 => x"54825373",
          6122 => x"802e9138",
          6123 => x"73733270",
          6124 => x"30710770",
          6125 => x"09709f2a",
          6126 => x"565d5e58",
          6127 => x"7283f8e4",
          6128 => x"0cff5980",
          6129 => x"547b812e",
          6130 => x"09810683",
          6131 => x"387b547b",
          6132 => x"83327030",
          6133 => x"70802576",
          6134 => x"075c5c5d",
          6135 => x"79802e85",
          6136 => x"c43884b8",
          6137 => x"f83383fa",
          6138 => x"b53383fa",
          6139 => x"b4337271",
          6140 => x"291286c7",
          6141 => x"a0800583",
          6142 => x"fab2225b",
          6143 => x"595d7179",
          6144 => x"29057083",
          6145 => x"ffff0683",
          6146 => x"f9893358",
          6147 => x"59555874",
          6148 => x"812e838c",
          6149 => x"3881f054",
          6150 => x"73878e80",
          6151 => x"8034800b",
          6152 => x"87c09888",
          6153 => x"0c87c098",
          6154 => x"88085675",
          6155 => x"802ef638",
          6156 => x"878e8084",
          6157 => x"08577683",
          6158 => x"f6b41534",
          6159 => x"81147081",
          6160 => x"ff065555",
          6161 => x"81f97427",
          6162 => x"cf388054",
          6163 => x"83f8a414",
          6164 => x"337081ff",
          6165 => x"0683f8ae",
          6166 => x"16335854",
          6167 => x"5572762e",
          6168 => x"85c13872",
          6169 => x"81ff2e86",
          6170 => x"b4387483",
          6171 => x"f8b81534",
          6172 => x"7581ff06",
          6173 => x"5a7981ff",
          6174 => x"2e85cd38",
          6175 => x"7583f8c2",
          6176 => x"153483f8",
          6177 => x"a4143383",
          6178 => x"f8ae1534",
          6179 => x"81147081",
          6180 => x"ff06555e",
          6181 => x"897427ff",
          6182 => x"b33883f8",
          6183 => x"ac337098",
          6184 => x"2b708025",
          6185 => x"58565475",
          6186 => x"83f8dc34",
          6187 => x"7381ff06",
          6188 => x"70862a81",
          6189 => x"32708106",
          6190 => x"51545872",
          6191 => x"802e85e7",
          6192 => x"38810b83",
          6193 => x"f8dd3473",
          6194 => x"09810653",
          6195 => x"72802e85",
          6196 => x"e438810b",
          6197 => x"83f8de34",
          6198 => x"800b83f8",
          6199 => x"dd3383f8",
          6200 => x"e40883f8",
          6201 => x"de337083",
          6202 => x"f8e03383",
          6203 => x"f8df335d",
          6204 => x"5d425e5c",
          6205 => x"5e5683f8",
          6206 => x"b8163355",
          6207 => x"7481ff2e",
          6208 => x"8d3883f8",
          6209 => x"cc163354",
          6210 => x"73802e82",
          6211 => x"823883f8",
          6212 => x"c2163353",
          6213 => x"7281ff2e",
          6214 => x"8b3883f8",
          6215 => x"cc163354",
          6216 => x"7381ec38",
          6217 => x"7481ff06",
          6218 => x"547381ff",
          6219 => x"2e8d3883",
          6220 => x"f8cc1633",
          6221 => x"5372812e",
          6222 => x"81da3874",
          6223 => x"81ff0653",
          6224 => x"7281ff2e",
          6225 => x"848c3883",
          6226 => x"f8cc1633",
          6227 => x"54817427",
          6228 => x"84803883",
          6229 => x"f8d80887",
          6230 => x"e80587c0",
          6231 => x"989c0854",
          6232 => x"54737327",
          6233 => x"83ec3881",
          6234 => x"0b87c098",
          6235 => x"9c0883f8",
          6236 => x"d80c5881",
          6237 => x"167081ff",
          6238 => x"06575489",
          6239 => x"7627fef6",
          6240 => x"387683f8",
          6241 => x"df347783",
          6242 => x"f8e034fe",
          6243 => x"9e195372",
          6244 => x"9c26828b",
          6245 => x"38721010",
          6246 => x"83c9fc05",
          6247 => x"5a790804",
          6248 => x"83f98c08",
          6249 => x"5473802e",
          6250 => x"913883f4",
          6251 => x"1487c098",
          6252 => x"9c085e5e",
          6253 => x"7d7d27fc",
          6254 => x"dc38800b",
          6255 => x"83f98a33",
          6256 => x"54547281",
          6257 => x"2e833874",
          6258 => x"547383f9",
          6259 => x"8a3487c0",
          6260 => x"989c0883",
          6261 => x"f98c0c73",
          6262 => x"81ff0658",
          6263 => x"77812e94",
          6264 => x"3883fab6",
          6265 => x"17335484",
          6266 => x"b9801433",
          6267 => x"763481f0",
          6268 => x"54fca539",
          6269 => x"83f8e408",
          6270 => x"5372802e",
          6271 => x"829c3872",
          6272 => x"812e83f4",
          6273 => x"3880c376",
          6274 => x"3481f054",
          6275 => x"fc8a3980",
          6276 => x"58fee039",
          6277 => x"80745657",
          6278 => x"83597c81",
          6279 => x"2e9b3879",
          6280 => x"772e0981",
          6281 => x"0683b438",
          6282 => x"7d812e80",
          6283 => x"ed387981",
          6284 => x"2e80d738",
          6285 => x"7981ff06",
          6286 => x"59877727",
          6287 => x"75982b54",
          6288 => x"54728025",
          6289 => x"a1387380",
          6290 => x"2e9c3881",
          6291 => x"177081ff",
          6292 => x"06761081",
          6293 => x"fe068772",
          6294 => x"2771982b",
          6295 => x"57535758",
          6296 => x"54807324",
          6297 => x"e1387810",
          6298 => x"10107910",
          6299 => x"05761183",
          6300 => x"2b780583",
          6301 => x"f5940570",
          6302 => x"335b5654",
          6303 => x"7887c098",
          6304 => x"9c0883f8",
          6305 => x"d80c57fd",
          6306 => x"ea398059",
          6307 => x"7d812eff",
          6308 => x"a8387981",
          6309 => x"ff0659ff",
          6310 => x"a0398259",
          6311 => x"ff9b3978",
          6312 => x"ff2efa9f",
          6313 => x"38800b84",
          6314 => x"b8fa3354",
          6315 => x"5472812e",
          6316 => x"83e8387b",
          6317 => x"82327030",
          6318 => x"70802576",
          6319 => x"07405956",
          6320 => x"7d8a387b",
          6321 => x"832e0981",
          6322 => x"06f9cc38",
          6323 => x"78ff2ef9",
          6324 => x"c6388053",
          6325 => x"72101010",
          6326 => x"83f99005",
          6327 => x"70335d54",
          6328 => x"787c2e83",
          6329 => x"ba388113",
          6330 => x"7081ff06",
          6331 => x"54579373",
          6332 => x"27e23884",
          6333 => x"b8fb3353",
          6334 => x"72802ef9",
          6335 => x"9a3884b8",
          6336 => x"fc335574",
          6337 => x"f9913878",
          6338 => x"81ff0652",
          6339 => x"8251ccd4",
          6340 => x"3f7884bb",
          6341 => x"840c8f3d",
          6342 => x"0d04be76",
          6343 => x"3481f054",
          6344 => x"f9f63972",
          6345 => x"81ff2e92",
          6346 => x"3883f8cc",
          6347 => x"14338105",
          6348 => x"5b7a83f8",
          6349 => x"cc1534fa",
          6350 => x"c939800b",
          6351 => x"83f8cc15",
          6352 => x"34ff0b83",
          6353 => x"f8b81534",
          6354 => x"ff0b83f8",
          6355 => x"c21534fa",
          6356 => x"b1397481",
          6357 => x"ff065372",
          6358 => x"81ff2efc",
          6359 => x"963883f8",
          6360 => x"cc163355",
          6361 => x"817527fc",
          6362 => x"8a387781",
          6363 => x"ff065473",
          6364 => x"812e0981",
          6365 => x"06fbfc38",
          6366 => x"83f8d808",
          6367 => x"81fa0587",
          6368 => x"c0989c08",
          6369 => x"54557473",
          6370 => x"27fbe838",
          6371 => x"87c0989c",
          6372 => x"0883f8d8",
          6373 => x"0c7681ff",
          6374 => x"0659fbd7",
          6375 => x"39ff0b83",
          6376 => x"f8b81534",
          6377 => x"f9ca3972",
          6378 => x"83f8dd34",
          6379 => x"73098106",
          6380 => x"5372fa9e",
          6381 => x"387283f8",
          6382 => x"de34800b",
          6383 => x"83f8dd33",
          6384 => x"83f8e408",
          6385 => x"83f8de33",
          6386 => x"7083f8e0",
          6387 => x"3383f8df",
          6388 => x"335d5d42",
          6389 => x"5e5c5e56",
          6390 => x"fa9c3979",
          6391 => x"822e0981",
          6392 => x"06fccb38",
          6393 => x"7a597a81",
          6394 => x"2efcce38",
          6395 => x"79812e09",
          6396 => x"8106fcc0",
          6397 => x"38fd9339",
          6398 => x"ef763481",
          6399 => x"f054f898",
          6400 => x"39800b84",
          6401 => x"b8fb3357",
          6402 => x"54758338",
          6403 => x"81547384",
          6404 => x"b8fb34ff",
          6405 => x"59f7ac39",
          6406 => x"800b84b8",
          6407 => x"fa335854",
          6408 => x"76833881",
          6409 => x"547384b8",
          6410 => x"fa34ff59",
          6411 => x"f7953981",
          6412 => x"5383f8e4",
          6413 => x"08842ef7",
          6414 => x"8338840b",
          6415 => x"83f8e40c",
          6416 => x"f6ff3984",
          6417 => x"b8f73370",
          6418 => x"81ff06ff",
          6419 => x"11575a54",
          6420 => x"80792783",
          6421 => x"38805574",
          6422 => x"83fab223",
          6423 => x"7381ff06",
          6424 => x"ff155553",
          6425 => x"80732783",
          6426 => x"38805473",
          6427 => x"83fab434",
          6428 => x"84b8f833",
          6429 => x"7081ff06",
          6430 => x"56ff0553",
          6431 => x"80752783",
          6432 => x"38805372",
          6433 => x"83fab534",
          6434 => x"ff59f6b7",
          6435 => x"39815283",
          6436 => x"51ffbaa5",
          6437 => x"3fff59f6",
          6438 => x"aa397254",
          6439 => x"fc953984",
          6440 => x"14085283",
          6441 => x"f8e851fe",
          6442 => x"dd9d3f81",
          6443 => x"0b83f988",
          6444 => x"3483f8e8",
          6445 => x"3359fcbb",
          6446 => x"39803d0d",
          6447 => x"8151f5ac",
          6448 => x"3f823d0d",
          6449 => x"04fa3d0d",
          6450 => x"800b83f5",
          6451 => x"90085357",
          6452 => x"02a30533",
          6453 => x"82133483",
          6454 => x"f5900851",
          6455 => x"80e07134",
          6456 => x"850b83f5",
          6457 => x"90085556",
          6458 => x"fe0b8115",
          6459 => x"34800b87",
          6460 => x"9080e834",
          6461 => x"87c0989c",
          6462 => x"0883f590",
          6463 => x"085580ce",
          6464 => x"90055387",
          6465 => x"c0989c08",
          6466 => x"5287c098",
          6467 => x"9c085170",
          6468 => x"722ef638",
          6469 => x"81143387",
          6470 => x"c0989c08",
          6471 => x"56527473",
          6472 => x"27873871",
          6473 => x"81fe2edb",
          6474 => x"3887c098",
          6475 => x"a40851ff",
          6476 => x"55707327",
          6477 => x"80c83871",
          6478 => x"5571ff2e",
          6479 => x"80c03887",
          6480 => x"c0989c08",
          6481 => x"80ce9005",
          6482 => x"5387c098",
          6483 => x"9c085287",
          6484 => x"c0989c08",
          6485 => x"5574722e",
          6486 => x"f6388114",
          6487 => x"3387c098",
          6488 => x"9c085252",
          6489 => x"70732787",
          6490 => x"387181ff",
          6491 => x"2edb3887",
          6492 => x"c098a408",
          6493 => x"55727526",
          6494 => x"8338ff52",
          6495 => x"7155ff16",
          6496 => x"7081ff06",
          6497 => x"57537580",
          6498 => x"2e983874",
          6499 => x"81ff0652",
          6500 => x"71fed538",
          6501 => x"74ff2e8a",
          6502 => x"387684bb",
          6503 => x"840c883d",
          6504 => x"0d04810b",
          6505 => x"84bb840c",
          6506 => x"883d0d04",
          6507 => x"fa3d0d79",
          6508 => x"028405a3",
          6509 => x"05335652",
          6510 => x"800b83f5",
          6511 => x"90087388",
          6512 => x"2b87fc80",
          6513 => x"80067075",
          6514 => x"982a0751",
          6515 => x"55555771",
          6516 => x"83153472",
          6517 => x"902a5170",
          6518 => x"84153471",
          6519 => x"902a5675",
          6520 => x"85153472",
          6521 => x"86153483",
          6522 => x"f5900852",
          6523 => x"74821334",
          6524 => x"83f59008",
          6525 => x"5180e171",
          6526 => x"34850b83",
          6527 => x"f5900855",
          6528 => x"56fe0b81",
          6529 => x"1534800b",
          6530 => x"879080e8",
          6531 => x"3487c098",
          6532 => x"9c0883f5",
          6533 => x"90085580",
          6534 => x"ce900553",
          6535 => x"87c0989c",
          6536 => x"085287c0",
          6537 => x"989c0851",
          6538 => x"70722ef6",
          6539 => x"38811433",
          6540 => x"87c0989c",
          6541 => x"08565274",
          6542 => x"73278738",
          6543 => x"7181fe2e",
          6544 => x"db3887c0",
          6545 => x"98a40851",
          6546 => x"ff557073",
          6547 => x"2780c838",
          6548 => x"715571ff",
          6549 => x"2e80c038",
          6550 => x"87c0989c",
          6551 => x"0880ce90",
          6552 => x"055387c0",
          6553 => x"989c0852",
          6554 => x"87c0989c",
          6555 => x"08557472",
          6556 => x"2ef63881",
          6557 => x"143387c0",
          6558 => x"989c0852",
          6559 => x"52707327",
          6560 => x"87387181",
          6561 => x"ff2edb38",
          6562 => x"87c098a4",
          6563 => x"08557275",
          6564 => x"268338ff",
          6565 => x"527155ff",
          6566 => x"167081ff",
          6567 => x"06575375",
          6568 => x"802e80c7",
          6569 => x"387481ff",
          6570 => x"065271fe",
          6571 => x"d4387451",
          6572 => x"7081ff06",
          6573 => x"5675aa38",
          6574 => x"80c6147b",
          6575 => x"84801155",
          6576 => x"52527073",
          6577 => x"27923871",
          6578 => x"70810553",
          6579 => x"33717081",
          6580 => x"05533472",
          6581 => x"7126f038",
          6582 => x"7684bb84",
          6583 => x"0c883d0d",
          6584 => x"04810b84",
          6585 => x"bb840c88",
          6586 => x"3d0d04ff",
          6587 => x"51c239fa",
          6588 => x"3d0d7902",
          6589 => x"8405a305",
          6590 => x"33565680",
          6591 => x"0b83f590",
          6592 => x"0877882b",
          6593 => x"87fc8080",
          6594 => x"06707998",
          6595 => x"2a075155",
          6596 => x"55577583",
          6597 => x"15347290",
          6598 => x"2a517084",
          6599 => x"15347590",
          6600 => x"2a527185",
          6601 => x"15347286",
          6602 => x"15347a83",
          6603 => x"f5900880",
          6604 => x"c6118480",
          6605 => x"13565455",
          6606 => x"51707327",
          6607 => x"97387070",
          6608 => x"81055233",
          6609 => x"72708105",
          6610 => x"54347271",
          6611 => x"26f03883",
          6612 => x"f5900854",
          6613 => x"74821534",
          6614 => x"83f59008",
          6615 => x"5580e275",
          6616 => x"34850b83",
          6617 => x"f5900855",
          6618 => x"56fe0b81",
          6619 => x"1534800b",
          6620 => x"879080e8",
          6621 => x"3487c098",
          6622 => x"9c0883f5",
          6623 => x"90085580",
          6624 => x"ce900553",
          6625 => x"87c0989c",
          6626 => x"085287c0",
          6627 => x"989c0851",
          6628 => x"70722ef6",
          6629 => x"38811433",
          6630 => x"87c0989c",
          6631 => x"08565274",
          6632 => x"73278738",
          6633 => x"7181fe2e",
          6634 => x"db3887c0",
          6635 => x"98a40851",
          6636 => x"ff557073",
          6637 => x"2780c838",
          6638 => x"715571ff",
          6639 => x"2e80c038",
          6640 => x"87c0989c",
          6641 => x"0880ce90",
          6642 => x"055387c0",
          6643 => x"989c0852",
          6644 => x"87c0989c",
          6645 => x"08557472",
          6646 => x"2ef63881",
          6647 => x"143387c0",
          6648 => x"989c0852",
          6649 => x"52707327",
          6650 => x"87387181",
          6651 => x"ff2edb38",
          6652 => x"87c098a4",
          6653 => x"08557275",
          6654 => x"268338ff",
          6655 => x"527155ff",
          6656 => x"167081ff",
          6657 => x"06575375",
          6658 => x"802ea138",
          6659 => x"7481ff06",
          6660 => x"5271fed5",
          6661 => x"38745170",
          6662 => x"81ff0654",
          6663 => x"73802e83",
          6664 => x"38815776",
          6665 => x"84bb840c",
          6666 => x"883d0d04",
          6667 => x"ff51e839",
          6668 => x"fb3d0d83",
          6669 => x"f5900851",
          6670 => x"80d07134",
          6671 => x"850b83f5",
          6672 => x"90085656",
          6673 => x"fe0b8116",
          6674 => x"34800b87",
          6675 => x"9080e834",
          6676 => x"87c0989c",
          6677 => x"0883f590",
          6678 => x"085680ce",
          6679 => x"90055487",
          6680 => x"c0989c08",
          6681 => x"5287c098",
          6682 => x"9c085372",
          6683 => x"722ef638",
          6684 => x"81153387",
          6685 => x"c0989c08",
          6686 => x"52527074",
          6687 => x"27873871",
          6688 => x"81fe2edb",
          6689 => x"3887c098",
          6690 => x"a40851ff",
          6691 => x"53707427",
          6692 => x"80c83871",
          6693 => x"5371ff2e",
          6694 => x"80c03887",
          6695 => x"c0989c08",
          6696 => x"80ce9005",
          6697 => x"5387c098",
          6698 => x"9c085287",
          6699 => x"c0989c08",
          6700 => x"5170722e",
          6701 => x"f6388115",
          6702 => x"3387c098",
          6703 => x"9c085552",
          6704 => x"73732787",
          6705 => x"387181ff",
          6706 => x"2edb3887",
          6707 => x"c098a408",
          6708 => x"51727126",
          6709 => x"8338ff52",
          6710 => x"7153ff16",
          6711 => x"7081ff06",
          6712 => x"57527580",
          6713 => x"2e8a3872",
          6714 => x"81ff0654",
          6715 => x"73fed538",
          6716 => x"ff39803d",
          6717 => x"0d83e688",
          6718 => x"51fecef7",
          6719 => x"3f823d0d",
          6720 => x"04f93d0d",
          6721 => x"84baf408",
          6722 => x"7a713183",
          6723 => x"2a7083ff",
          6724 => x"ff067083",
          6725 => x"2b731170",
          6726 => x"33811233",
          6727 => x"718b2b71",
          6728 => x"832b0777",
          6729 => x"11703381",
          6730 => x"12337198",
          6731 => x"2b71902b",
          6732 => x"075c5441",
          6733 => x"53535d57",
          6734 => x"59525657",
          6735 => x"53807124",
          6736 => x"81af3872",
          6737 => x"16821133",
          6738 => x"83123371",
          6739 => x"8b2b7183",
          6740 => x"2b077605",
          6741 => x"70338112",
          6742 => x"3371982b",
          6743 => x"71902b07",
          6744 => x"57535c52",
          6745 => x"59565280",
          6746 => x"7124839e",
          6747 => x"38841333",
          6748 => x"85143371",
          6749 => x"8b2b7183",
          6750 => x"2b077505",
          6751 => x"76882a52",
          6752 => x"54565774",
          6753 => x"86133473",
          6754 => x"81ff0654",
          6755 => x"73871334",
          6756 => x"84baf408",
          6757 => x"70178412",
          6758 => x"33851333",
          6759 => x"71882b07",
          6760 => x"70882a5c",
          6761 => x"55595451",
          6762 => x"77841434",
          6763 => x"71851434",
          6764 => x"84baf408",
          6765 => x"1652800b",
          6766 => x"86133480",
          6767 => x"0b871334",
          6768 => x"84baf408",
          6769 => x"53748414",
          6770 => x"34738514",
          6771 => x"3484baf4",
          6772 => x"08167033",
          6773 => x"81123371",
          6774 => x"882b0782",
          6775 => x"80800770",
          6776 => x"882a5858",
          6777 => x"52527472",
          6778 => x"34758113",
          6779 => x"34893d0d",
          6780 => x"04861233",
          6781 => x"87133371",
          6782 => x"8b2b7183",
          6783 => x"2b077511",
          6784 => x"84163385",
          6785 => x"17337188",
          6786 => x"2b077088",
          6787 => x"2a585854",
          6788 => x"51535858",
          6789 => x"71841234",
          6790 => x"72851234",
          6791 => x"84baf408",
          6792 => x"70168411",
          6793 => x"33851233",
          6794 => x"718b2b71",
          6795 => x"832b0756",
          6796 => x"5a5a5272",
          6797 => x"05861233",
          6798 => x"87133371",
          6799 => x"882b0770",
          6800 => x"882a5255",
          6801 => x"59527786",
          6802 => x"13347287",
          6803 => x"133484ba",
          6804 => x"f4081570",
          6805 => x"33811233",
          6806 => x"71882b07",
          6807 => x"81ffff06",
          6808 => x"70882a5a",
          6809 => x"5a545276",
          6810 => x"72347781",
          6811 => x"133484ba",
          6812 => x"f4087017",
          6813 => x"70338112",
          6814 => x"33718b2b",
          6815 => x"71832b07",
          6816 => x"74057033",
          6817 => x"81123371",
          6818 => x"882b0770",
          6819 => x"832b8fff",
          6820 => x"f8067705",
          6821 => x"7b882a54",
          6822 => x"5253545c",
          6823 => x"5a575452",
          6824 => x"77821434",
          6825 => x"73831434",
          6826 => x"84baf408",
          6827 => x"70177033",
          6828 => x"81123371",
          6829 => x"8b2b7183",
          6830 => x"2b077405",
          6831 => x"70338112",
          6832 => x"3371882b",
          6833 => x"0781ffff",
          6834 => x"0670882a",
          6835 => x"5f525355",
          6836 => x"5a575452",
          6837 => x"77733470",
          6838 => x"81143484",
          6839 => x"baf40870",
          6840 => x"17821133",
          6841 => x"83123371",
          6842 => x"8b2b7183",
          6843 => x"2b077405",
          6844 => x"70338112",
          6845 => x"3371982b",
          6846 => x"71902b07",
          6847 => x"58535d52",
          6848 => x"5a575353",
          6849 => x"708025fc",
          6850 => x"e4387133",
          6851 => x"81133371",
          6852 => x"882b0782",
          6853 => x"80800770",
          6854 => x"882a5959",
          6855 => x"54767534",
          6856 => x"77811634",
          6857 => x"84baf408",
          6858 => x"70177033",
          6859 => x"81123371",
          6860 => x"8b2b7183",
          6861 => x"2b077405",
          6862 => x"82143383",
          6863 => x"15337188",
          6864 => x"2b077088",
          6865 => x"2a575c5c",
          6866 => x"52585652",
          6867 => x"53728215",
          6868 => x"34758315",
          6869 => x"34893d0d",
          6870 => x"04f93d0d",
          6871 => x"7984baf4",
          6872 => x"08585876",
          6873 => x"802e8f38",
          6874 => x"77802e86",
          6875 => x"387751fb",
          6876 => x"903f893d",
          6877 => x"0d0484ff",
          6878 => x"f40b84ba",
          6879 => x"f40ca080",
          6880 => x"0b84baf0",
          6881 => x"23828080",
          6882 => x"53765284",
          6883 => x"fff451fe",
          6884 => x"d1ed3f84",
          6885 => x"baf40855",
          6886 => x"76753481",
          6887 => x"0b811634",
          6888 => x"84baf408",
          6889 => x"54768415",
          6890 => x"34810b85",
          6891 => x"153484ba",
          6892 => x"f4085676",
          6893 => x"86173481",
          6894 => x"0b871734",
          6895 => x"84baf408",
          6896 => x"84baf022",
          6897 => x"ff05fe80",
          6898 => x"80077083",
          6899 => x"ffff0670",
          6900 => x"882a5851",
          6901 => x"55567488",
          6902 => x"17347389",
          6903 => x"173484ba",
          6904 => x"f0227010",
          6905 => x"101084ba",
          6906 => x"f40805f8",
          6907 => x"05555576",
          6908 => x"82153481",
          6909 => x"0b831534",
          6910 => x"feee39f7",
          6911 => x"3d0d7b52",
          6912 => x"80538151",
          6913 => x"8472278e",
          6914 => x"38fb1283",
          6915 => x"2a820570",
          6916 => x"83ffff06",
          6917 => x"51517083",
          6918 => x"ffff0684",
          6919 => x"baf40884",
          6920 => x"11338512",
          6921 => x"3371882b",
          6922 => x"07705259",
          6923 => x"5a585581",
          6924 => x"ffff5475",
          6925 => x"802e80cc",
          6926 => x"38751010",
          6927 => x"10177033",
          6928 => x"81123371",
          6929 => x"882b0770",
          6930 => x"81ffff06",
          6931 => x"79317083",
          6932 => x"ffff0670",
          6933 => x"7a275653",
          6934 => x"5c5c5452",
          6935 => x"7274278a",
          6936 => x"3870802e",
          6937 => x"85387573",
          6938 => x"55588412",
          6939 => x"33851333",
          6940 => x"71882b07",
          6941 => x"575a75c1",
          6942 => x"387381ff",
          6943 => x"ff2e8538",
          6944 => x"77745456",
          6945 => x"8076832b",
          6946 => x"78117033",
          6947 => x"81123371",
          6948 => x"882b0770",
          6949 => x"81ffff06",
          6950 => x"56565d56",
          6951 => x"59597079",
          6952 => x"2e833881",
          6953 => x"59805174",
          6954 => x"7326828d",
          6955 => x"38785178",
          6956 => x"802e8285",
          6957 => x"3872752e",
          6958 => x"82883874",
          6959 => x"1670832b",
          6960 => x"78117482",
          6961 => x"80800770",
          6962 => x"882a5b5c",
          6963 => x"56565a76",
          6964 => x"74347881",
          6965 => x"153484ba",
          6966 => x"f4081576",
          6967 => x"882a5353",
          6968 => x"71821434",
          6969 => x"75831434",
          6970 => x"84baf408",
          6971 => x"70197033",
          6972 => x"81123371",
          6973 => x"882b0770",
          6974 => x"832b8fff",
          6975 => x"f8067405",
          6976 => x"7e83ffff",
          6977 => x"0670882a",
          6978 => x"5c585357",
          6979 => x"59525275",
          6980 => x"82123472",
          6981 => x"81ff0653",
          6982 => x"72831234",
          6983 => x"84baf408",
          6984 => x"18547574",
          6985 => x"34728115",
          6986 => x"3484baf4",
          6987 => x"08701986",
          6988 => x"11338712",
          6989 => x"33718b2b",
          6990 => x"71832b07",
          6991 => x"7405585c",
          6992 => x"5c535775",
          6993 => x"84153472",
          6994 => x"85153484",
          6995 => x"baf40870",
          6996 => x"16557805",
          6997 => x"86113387",
          6998 => x"12337188",
          6999 => x"2b077088",
          7000 => x"2a545458",
          7001 => x"59708615",
          7002 => x"34718715",
          7003 => x"3484baf4",
          7004 => x"08701984",
          7005 => x"11338512",
          7006 => x"33718b2b",
          7007 => x"71832b07",
          7008 => x"7405585a",
          7009 => x"5c5a5275",
          7010 => x"86153472",
          7011 => x"87153484",
          7012 => x"baf40870",
          7013 => x"16557805",
          7014 => x"84113385",
          7015 => x"12337188",
          7016 => x"2b077088",
          7017 => x"2a545c57",
          7018 => x"59708415",
          7019 => x"34798515",
          7020 => x"3484baf4",
          7021 => x"08188405",
          7022 => x"517084bb",
          7023 => x"840c8b3d",
          7024 => x"0d048614",
          7025 => x"33871533",
          7026 => x"718b2b71",
          7027 => x"832b0779",
          7028 => x"05841733",
          7029 => x"85183371",
          7030 => x"882b0770",
          7031 => x"882a5a5b",
          7032 => x"59535452",
          7033 => x"74841234",
          7034 => x"76851234",
          7035 => x"84baf408",
          7036 => x"70198411",
          7037 => x"33851233",
          7038 => x"718b2b71",
          7039 => x"832b0774",
          7040 => x"05861433",
          7041 => x"87153371",
          7042 => x"882b0770",
          7043 => x"882a585d",
          7044 => x"5f52565b",
          7045 => x"57527086",
          7046 => x"1a347687",
          7047 => x"1a3484ba",
          7048 => x"f4081870",
          7049 => x"33811233",
          7050 => x"71882b07",
          7051 => x"81ffff06",
          7052 => x"70882a59",
          7053 => x"57545775",
          7054 => x"77347481",
          7055 => x"183484ba",
          7056 => x"f4081884",
          7057 => x"0551fef1",
          7058 => x"39f93d0d",
          7059 => x"7984baf4",
          7060 => x"08585876",
          7061 => x"802ea038",
          7062 => x"7754778a",
          7063 => x"387384bb",
          7064 => x"840c893d",
          7065 => x"0d047751",
          7066 => x"fb913f84",
          7067 => x"bb840884",
          7068 => x"bb840c89",
          7069 => x"3d0d0484",
          7070 => x"fff40b84",
          7071 => x"baf40ca0",
          7072 => x"800b84ba",
          7073 => x"f0238280",
          7074 => x"80537652",
          7075 => x"84fff451",
          7076 => x"fecbec3f",
          7077 => x"84baf408",
          7078 => x"55767534",
          7079 => x"810b8116",
          7080 => x"3484baf4",
          7081 => x"08547684",
          7082 => x"1534810b",
          7083 => x"85153484",
          7084 => x"baf40856",
          7085 => x"76861734",
          7086 => x"810b8717",
          7087 => x"3484baf4",
          7088 => x"0884baf0",
          7089 => x"22ff05fe",
          7090 => x"80800770",
          7091 => x"83ffff06",
          7092 => x"70882a58",
          7093 => x"51555674",
          7094 => x"88173473",
          7095 => x"89173484",
          7096 => x"baf02270",
          7097 => x"10101084",
          7098 => x"baf40805",
          7099 => x"f8055555",
          7100 => x"76821534",
          7101 => x"810b8315",
          7102 => x"34775477",
          7103 => x"802efedd",
          7104 => x"38fee339",
          7105 => x"ed3d0d65",
          7106 => x"67415f80",
          7107 => x"7084baf4",
          7108 => x"08594541",
          7109 => x"76612e84",
          7110 => x"aa387e80",
          7111 => x"2e85af38",
          7112 => x"7f802e88",
          7113 => x"d7388154",
          7114 => x"8460278f",
          7115 => x"387ffb05",
          7116 => x"832a8205",
          7117 => x"7083ffff",
          7118 => x"06555873",
          7119 => x"83ffff06",
          7120 => x"7f783183",
          7121 => x"2a7083ff",
          7122 => x"ff067083",
          7123 => x"2b7a1170",
          7124 => x"33811233",
          7125 => x"71882b07",
          7126 => x"70753170",
          7127 => x"83ffff06",
          7128 => x"70101010",
          7129 => x"fc057383",
          7130 => x"2b611170",
          7131 => x"33811233",
          7132 => x"71882b07",
          7133 => x"70902b70",
          7134 => x"902c5342",
          7135 => x"45464453",
          7136 => x"5443445c",
          7137 => x"4859525e",
          7138 => x"5f42807a",
          7139 => x"2485fd38",
          7140 => x"82153383",
          7141 => x"16337188",
          7142 => x"2b077010",
          7143 => x"10101970",
          7144 => x"33811233",
          7145 => x"71982b71",
          7146 => x"902b0753",
          7147 => x"5c535656",
          7148 => x"56807424",
          7149 => x"85c9387a",
          7150 => x"622782f6",
          7151 => x"38631b58",
          7152 => x"77622e87",
          7153 => x"a2386080",
          7154 => x"2e85f938",
          7155 => x"601b5877",
          7156 => x"622587be",
          7157 => x"38631859",
          7158 => x"61792492",
          7159 => x"f738761e",
          7160 => x"70338112",
          7161 => x"33718b2b",
          7162 => x"71832b07",
          7163 => x"7a117033",
          7164 => x"81123371",
          7165 => x"982b7190",
          7166 => x"2b074743",
          7167 => x"59525357",
          7168 => x"5b588060",
          7169 => x"248cba38",
          7170 => x"761e8211",
          7171 => x"33831233",
          7172 => x"718b2b71",
          7173 => x"832b077a",
          7174 => x"11861133",
          7175 => x"87123371",
          7176 => x"8b2b7183",
          7177 => x"2b077e05",
          7178 => x"84143385",
          7179 => x"15337188",
          7180 => x"2b077088",
          7181 => x"2a595748",
          7182 => x"525b4158",
          7183 => x"535c5956",
          7184 => x"77841d34",
          7185 => x"79851d34",
          7186 => x"84baf408",
          7187 => x"70178411",
          7188 => x"33851233",
          7189 => x"718b2b71",
          7190 => x"832b0774",
          7191 => x"05861433",
          7192 => x"87153371",
          7193 => x"882b0770",
          7194 => x"882a5f42",
          7195 => x"5e524057",
          7196 => x"41577786",
          7197 => x"16347b87",
          7198 => x"163484ba",
          7199 => x"f4081670",
          7200 => x"33811233",
          7201 => x"71882b07",
          7202 => x"81ffff06",
          7203 => x"70882a5a",
          7204 => x"5c5e5976",
          7205 => x"79347981",
          7206 => x"1a3484ba",
          7207 => x"f408701f",
          7208 => x"82113383",
          7209 => x"1233718b",
          7210 => x"2b71832b",
          7211 => x"07740573",
          7212 => x"33811533",
          7213 => x"71882b07",
          7214 => x"70882a41",
          7215 => x"5c455d5f",
          7216 => x"5a555579",
          7217 => x"79347581",
          7218 => x"1a3484ba",
          7219 => x"f408701f",
          7220 => x"70338112",
          7221 => x"33718b2b",
          7222 => x"71832b07",
          7223 => x"74058214",
          7224 => x"33831533",
          7225 => x"71882b07",
          7226 => x"70882a41",
          7227 => x"5c455d5f",
          7228 => x"5a555579",
          7229 => x"821a3475",
          7230 => x"831a3484",
          7231 => x"baf40870",
          7232 => x"1f821133",
          7233 => x"83123371",
          7234 => x"882b0766",
          7235 => x"57625670",
          7236 => x"832b4252",
          7237 => x"5a5d7e05",
          7238 => x"840551fe",
          7239 => x"c3a43f84",
          7240 => x"baf4081e",
          7241 => x"84056165",
          7242 => x"051c7083",
          7243 => x"ffff065d",
          7244 => x"445f7a62",
          7245 => x"2681b638",
          7246 => x"7e547384",
          7247 => x"bb840c95",
          7248 => x"3d0d0484",
          7249 => x"fff40b84",
          7250 => x"baf40ca0",
          7251 => x"800b84ba",
          7252 => x"f0238280",
          7253 => x"80536052",
          7254 => x"84fff451",
          7255 => x"fec6a03f",
          7256 => x"84baf408",
          7257 => x"5e607e34",
          7258 => x"810b811f",
          7259 => x"3484baf4",
          7260 => x"085d6084",
          7261 => x"1e34810b",
          7262 => x"851e3484",
          7263 => x"baf4085c",
          7264 => x"60861d34",
          7265 => x"810b871d",
          7266 => x"3484baf4",
          7267 => x"0884baf0",
          7268 => x"22ff05fe",
          7269 => x"80800770",
          7270 => x"83ffff06",
          7271 => x"70882a5c",
          7272 => x"5a5b5778",
          7273 => x"88183477",
          7274 => x"89183484",
          7275 => x"baf02270",
          7276 => x"10101084",
          7277 => x"baf40805",
          7278 => x"f8055556",
          7279 => x"60821534",
          7280 => x"810b8315",
          7281 => x"3484baf4",
          7282 => x"08577efa",
          7283 => x"d3387680",
          7284 => x"2e828c38",
          7285 => x"7e547f80",
          7286 => x"2efedf38",
          7287 => x"7f51f49b",
          7288 => x"3f84bb84",
          7289 => x"0884bb84",
          7290 => x"0c953d0d",
          7291 => x"04611c84",
          7292 => x"baf40871",
          7293 => x"832b7111",
          7294 => x"5e447f05",
          7295 => x"70338112",
          7296 => x"3371882b",
          7297 => x"0781ffff",
          7298 => x"0670882a",
          7299 => x"48445b5e",
          7300 => x"40637b34",
          7301 => x"60811c34",
          7302 => x"6184baf4",
          7303 => x"08057c88",
          7304 => x"2a575875",
          7305 => x"8219347b",
          7306 => x"83193484",
          7307 => x"baf40870",
          7308 => x"1f703381",
          7309 => x"12337188",
          7310 => x"2b077083",
          7311 => x"2b8ffff8",
          7312 => x"06740564",
          7313 => x"83ffff06",
          7314 => x"70882a4a",
          7315 => x"5c47575e",
          7316 => x"5b5d6363",
          7317 => x"82053476",
          7318 => x"81ff0641",
          7319 => x"60638305",
          7320 => x"3484baf4",
          7321 => x"081e5b63",
          7322 => x"7b346081",
          7323 => x"1c346184",
          7324 => x"baf40805",
          7325 => x"840551ed",
          7326 => x"883f7e54",
          7327 => x"fdbc397b",
          7328 => x"75317083",
          7329 => x"ffff0642",
          7330 => x"54faac39",
          7331 => x"7781ffff",
          7332 => x"06763170",
          7333 => x"83ffff06",
          7334 => x"82173383",
          7335 => x"18337188",
          7336 => x"2b077010",
          7337 => x"10101b70",
          7338 => x"33811233",
          7339 => x"71982b71",
          7340 => x"902b0753",
          7341 => x"5e535458",
          7342 => x"58455473",
          7343 => x"8025f9f7",
          7344 => x"38ffbc39",
          7345 => x"617824fa",
          7346 => x"8338807a",
          7347 => x"248b8f38",
          7348 => x"7783ffff",
          7349 => x"065b617b",
          7350 => x"27fcdd38",
          7351 => x"fe8f3984",
          7352 => x"fff40b84",
          7353 => x"baf40ca0",
          7354 => x"800b84ba",
          7355 => x"f0238280",
          7356 => x"80537e52",
          7357 => x"84fff451",
          7358 => x"fec3843f",
          7359 => x"84baf408",
          7360 => x"5a7e7a34",
          7361 => x"810b811b",
          7362 => x"3484baf4",
          7363 => x"08597e84",
          7364 => x"1a34810b",
          7365 => x"851a3484",
          7366 => x"baf40858",
          7367 => x"7e861934",
          7368 => x"810b8719",
          7369 => x"3484baf4",
          7370 => x"0884baf0",
          7371 => x"22ff05fe",
          7372 => x"80800770",
          7373 => x"83ffff06",
          7374 => x"70882a58",
          7375 => x"56574474",
          7376 => x"64880534",
          7377 => x"73648905",
          7378 => x"3484baf0",
          7379 => x"22701010",
          7380 => x"1084baf4",
          7381 => x"0805f805",
          7382 => x"42437e61",
          7383 => x"82053481",
          7384 => x"61830534",
          7385 => x"fcee3980",
          7386 => x"7a2483de",
          7387 => x"386183ff",
          7388 => x"ff065b61",
          7389 => x"7b27fbc0",
          7390 => x"38fcf239",
          7391 => x"76802e82",
          7392 => x"bd387e51",
          7393 => x"eafb3f7f",
          7394 => x"547384bb",
          7395 => x"840c953d",
          7396 => x"0d04761e",
          7397 => x"82113383",
          7398 => x"1233718b",
          7399 => x"2b71832b",
          7400 => x"077a1186",
          7401 => x"11338712",
          7402 => x"33718b2b",
          7403 => x"71832b07",
          7404 => x"7e058414",
          7405 => x"33851533",
          7406 => x"71882b07",
          7407 => x"70882a43",
          7408 => x"4445565b",
          7409 => x"4658535c",
          7410 => x"45567864",
          7411 => x"8405347a",
          7412 => x"64850534",
          7413 => x"84baf408",
          7414 => x"70178411",
          7415 => x"33851233",
          7416 => x"718b2b71",
          7417 => x"832b0774",
          7418 => x"05861433",
          7419 => x"87153371",
          7420 => x"882b0770",
          7421 => x"882a5b41",
          7422 => x"42485d59",
          7423 => x"5d417364",
          7424 => x"8605347a",
          7425 => x"64870534",
          7426 => x"84baf408",
          7427 => x"16703381",
          7428 => x"12337188",
          7429 => x"2b0781ff",
          7430 => x"ff067088",
          7431 => x"2a5f5c5a",
          7432 => x"5d7b7d34",
          7433 => x"79811e34",
          7434 => x"84baf408",
          7435 => x"701f8211",
          7436 => x"33831233",
          7437 => x"718b2b71",
          7438 => x"832b0774",
          7439 => x"05733381",
          7440 => x"15337188",
          7441 => x"2b077088",
          7442 => x"2a5e5c5e",
          7443 => x"40435745",
          7444 => x"54767c34",
          7445 => x"75811d34",
          7446 => x"84baf408",
          7447 => x"701f7033",
          7448 => x"81123371",
          7449 => x"8b2b7183",
          7450 => x"2b077405",
          7451 => x"82143383",
          7452 => x"15337188",
          7453 => x"2b077088",
          7454 => x"2a404740",
          7455 => x"5b405c55",
          7456 => x"55788218",
          7457 => x"34608318",
          7458 => x"3484baf4",
          7459 => x"08701f82",
          7460 => x"11338312",
          7461 => x"3371882b",
          7462 => x"07665762",
          7463 => x"5670832b",
          7464 => x"4252585d",
          7465 => x"7e058405",
          7466 => x"51febc96",
          7467 => x"3f84baf4",
          7468 => x"081e8405",
          7469 => x"7883ffff",
          7470 => x"065c5ffc",
          7471 => x"993984ff",
          7472 => x"f40b84ba",
          7473 => x"f40ca080",
          7474 => x"0b84baf0",
          7475 => x"23828080",
          7476 => x"537f5284",
          7477 => x"fff451fe",
          7478 => x"bfa53f84",
          7479 => x"baf40856",
          7480 => x"7f763481",
          7481 => x"0b811734",
          7482 => x"84baf408",
          7483 => x"557f8416",
          7484 => x"34810b85",
          7485 => x"163484ba",
          7486 => x"f408547f",
          7487 => x"86153481",
          7488 => x"0b871534",
          7489 => x"84baf408",
          7490 => x"84baf022",
          7491 => x"ff05fe80",
          7492 => x"80077083",
          7493 => x"ffff0670",
          7494 => x"882a4543",
          7495 => x"445e6188",
          7496 => x"1f346089",
          7497 => x"1f3484ba",
          7498 => x"f0227010",
          7499 => x"101084ba",
          7500 => x"f40805f8",
          7501 => x"055c5d7f",
          7502 => x"821c3481",
          7503 => x"0b831c34",
          7504 => x"7e51e7bd",
          7505 => x"3f7f54fc",
          7506 => x"c0398619",
          7507 => x"33871a33",
          7508 => x"718b2b71",
          7509 => x"832b0779",
          7510 => x"05841c33",
          7511 => x"851d3371",
          7512 => x"882b0770",
          7513 => x"882a5c48",
          7514 => x"5e435955",
          7515 => x"76618405",
          7516 => x"34636185",
          7517 => x"053484ba",
          7518 => x"f408701e",
          7519 => x"84113385",
          7520 => x"1233718b",
          7521 => x"2b71832b",
          7522 => x"07740586",
          7523 => x"14338715",
          7524 => x"3371882b",
          7525 => x"0770882a",
          7526 => x"415f4848",
          7527 => x"59565940",
          7528 => x"79648605",
          7529 => x"34786487",
          7530 => x"053484ba",
          7531 => x"f4081d70",
          7532 => x"33811233",
          7533 => x"71882b07",
          7534 => x"81ffff06",
          7535 => x"70882a59",
          7536 => x"42585875",
          7537 => x"78347f81",
          7538 => x"193484ba",
          7539 => x"f408701f",
          7540 => x"70338112",
          7541 => x"33718b2b",
          7542 => x"71832b07",
          7543 => x"74057033",
          7544 => x"81123371",
          7545 => x"882b0770",
          7546 => x"832b8fff",
          7547 => x"f8067705",
          7548 => x"63882a48",
          7549 => x"5d5d5a5d",
          7550 => x"405d4441",
          7551 => x"7f821734",
          7552 => x"7b831734",
          7553 => x"84baf408",
          7554 => x"701f7033",
          7555 => x"81123371",
          7556 => x"8b2b7183",
          7557 => x"2b077405",
          7558 => x"70338112",
          7559 => x"3371882b",
          7560 => x"0781ffff",
          7561 => x"0670882a",
          7562 => x"485d5e5e",
          7563 => x"465a415b",
          7564 => x"60603476",
          7565 => x"60810534",
          7566 => x"6183ffff",
          7567 => x"065bfab3",
          7568 => x"39861533",
          7569 => x"87163371",
          7570 => x"8b2b7183",
          7571 => x"2b077905",
          7572 => x"84183385",
          7573 => x"19337188",
          7574 => x"2b077088",
          7575 => x"2a5e5e5a",
          7576 => x"52415d78",
          7577 => x"841e3479",
          7578 => x"851e3484",
          7579 => x"baf40870",
          7580 => x"19841133",
          7581 => x"85123371",
          7582 => x"8b2b7183",
          7583 => x"2b077405",
          7584 => x"86143387",
          7585 => x"15337188",
          7586 => x"2b077088",
          7587 => x"2a44565e",
          7588 => x"525a4255",
          7589 => x"567c6086",
          7590 => x"05347560",
          7591 => x"87053484",
          7592 => x"baf40818",
          7593 => x"70338112",
          7594 => x"3371882b",
          7595 => x"0781ffff",
          7596 => x"0670882a",
          7597 => x"5b5b5855",
          7598 => x"77753478",
          7599 => x"81163484",
          7600 => x"baf40870",
          7601 => x"1f703381",
          7602 => x"1233718b",
          7603 => x"2b71832b",
          7604 => x"07740570",
          7605 => x"33811233",
          7606 => x"71882b07",
          7607 => x"70832b8f",
          7608 => x"fff80677",
          7609 => x"0563882a",
          7610 => x"56545f5f",
          7611 => x"5859425e",
          7612 => x"557f8217",
          7613 => x"347b8317",
          7614 => x"3484baf4",
          7615 => x"08701f70",
          7616 => x"33811233",
          7617 => x"718b2b71",
          7618 => x"832b0774",
          7619 => x"05703381",
          7620 => x"12337188",
          7621 => x"2b0781ff",
          7622 => x"ff067088",
          7623 => x"2a5d545e",
          7624 => x"585b595d",
          7625 => x"55757c34",
          7626 => x"76811d34",
          7627 => x"84baf408",
          7628 => x"701f8211",
          7629 => x"33831233",
          7630 => x"718b2b71",
          7631 => x"832b0774",
          7632 => x"11861133",
          7633 => x"87123371",
          7634 => x"8b2b7183",
          7635 => x"2b077805",
          7636 => x"84143385",
          7637 => x"15337188",
          7638 => x"2b077088",
          7639 => x"2a595749",
          7640 => x"525c4259",
          7641 => x"535d5a57",
          7642 => x"5777841d",
          7643 => x"3479851d",
          7644 => x"3484baf4",
          7645 => x"08701784",
          7646 => x"11338512",
          7647 => x"33718b2b",
          7648 => x"71832b07",
          7649 => x"74058614",
          7650 => x"33871533",
          7651 => x"71882b07",
          7652 => x"70882a5f",
          7653 => x"425e5240",
          7654 => x"57415777",
          7655 => x"8616347b",
          7656 => x"87163484",
          7657 => x"baf40816",
          7658 => x"70338112",
          7659 => x"3371882b",
          7660 => x"0781ffff",
          7661 => x"0670882a",
          7662 => x"5a5c5e59",
          7663 => x"76793479",
          7664 => x"811a3484",
          7665 => x"baf40870",
          7666 => x"1f821133",
          7667 => x"83123371",
          7668 => x"8b2b7183",
          7669 => x"2b077405",
          7670 => x"73338115",
          7671 => x"3371882b",
          7672 => x"0770882a",
          7673 => x"415c455d",
          7674 => x"5f5a5555",
          7675 => x"79793475",
          7676 => x"811a3484",
          7677 => x"baf40870",
          7678 => x"1f703381",
          7679 => x"1233718b",
          7680 => x"2b71832b",
          7681 => x"07740582",
          7682 => x"14338315",
          7683 => x"3371882b",
          7684 => x"0770882a",
          7685 => x"415c455d",
          7686 => x"5f5a5555",
          7687 => x"79821a34",
          7688 => x"75831a34",
          7689 => x"84baf408",
          7690 => x"701f8211",
          7691 => x"33831233",
          7692 => x"71882b07",
          7693 => x"66576256",
          7694 => x"70832b42",
          7695 => x"525a5d7e",
          7696 => x"05840551",
          7697 => x"feb4fb3f",
          7698 => x"84baf408",
          7699 => x"1e840561",
          7700 => x"65051c70",
          7701 => x"83ffff06",
          7702 => x"5d445ff1",
          7703 => x"d5398619",
          7704 => x"33871a33",
          7705 => x"718b2b71",
          7706 => x"832b0779",
          7707 => x"05841c33",
          7708 => x"851d3371",
          7709 => x"882b0770",
          7710 => x"882a4048",
          7711 => x"5d434155",
          7712 => x"7a618405",
          7713 => x"34636185",
          7714 => x"053484ba",
          7715 => x"f408701e",
          7716 => x"84113385",
          7717 => x"1233718b",
          7718 => x"2b71832b",
          7719 => x"07740586",
          7720 => x"14338715",
          7721 => x"3371882b",
          7722 => x"0770882a",
          7723 => x"5b415f48",
          7724 => x"5c594156",
          7725 => x"73648605",
          7726 => x"347a6487",
          7727 => x"053484ba",
          7728 => x"f4081d70",
          7729 => x"33811233",
          7730 => x"71882b07",
          7731 => x"81ffff06",
          7732 => x"70882a5c",
          7733 => x"5f425578",
          7734 => x"75347c81",
          7735 => x"163484ba",
          7736 => x"f408701f",
          7737 => x"70338112",
          7738 => x"33718b2b",
          7739 => x"71832b07",
          7740 => x"74057033",
          7741 => x"81123371",
          7742 => x"882b0770",
          7743 => x"832b8fff",
          7744 => x"f8067705",
          7745 => x"63882a5d",
          7746 => x"445c4958",
          7747 => x"5e455840",
          7748 => x"74821e34",
          7749 => x"7b831e34",
          7750 => x"84baf408",
          7751 => x"701f7033",
          7752 => x"81123371",
          7753 => x"8b2b7183",
          7754 => x"2b077405",
          7755 => x"70338112",
          7756 => x"3371882b",
          7757 => x"0781ffff",
          7758 => x"0670882a",
          7759 => x"475f4958",
          7760 => x"46595e5b",
          7761 => x"7f7d3478",
          7762 => x"811e3477",
          7763 => x"83ffff06",
          7764 => x"5bf38339",
          7765 => x"7e605254",
          7766 => x"e5a13f84",
          7767 => x"bb84085f",
          7768 => x"84bb8408",
          7769 => x"802e9338",
          7770 => x"62537352",
          7771 => x"84bb8408",
          7772 => x"51feb3f6",
          7773 => x"3f7351df",
          7774 => x"883f615b",
          7775 => x"617b27ef",
          7776 => x"b738f0e9",
          7777 => x"39f93d0d",
          7778 => x"7a7a2984",
          7779 => x"baf40858",
          7780 => x"5876802e",
          7781 => x"b7387754",
          7782 => x"778a3873",
          7783 => x"84bb840c",
          7784 => x"893d0d04",
          7785 => x"7751e4d3",
          7786 => x"3f84bb84",
          7787 => x"085484bb",
          7788 => x"8408802e",
          7789 => x"e6387753",
          7790 => x"805284bb",
          7791 => x"840851fe",
          7792 => x"b5bd3f73",
          7793 => x"84bb840c",
          7794 => x"893d0d04",
          7795 => x"84fff40b",
          7796 => x"84baf40c",
          7797 => x"a0800b84",
          7798 => x"baf02382",
          7799 => x"80805376",
          7800 => x"5284fff4",
          7801 => x"51feb597",
          7802 => x"3f84baf4",
          7803 => x"08557675",
          7804 => x"34810b81",
          7805 => x"163484ba",
          7806 => x"f4085476",
          7807 => x"84153481",
          7808 => x"0b851534",
          7809 => x"84baf408",
          7810 => x"56768617",
          7811 => x"34810b87",
          7812 => x"173484ba",
          7813 => x"f40884ba",
          7814 => x"f022ff05",
          7815 => x"fe808007",
          7816 => x"7083ffff",
          7817 => x"0670882a",
          7818 => x"58515556",
          7819 => x"74881734",
          7820 => x"73891734",
          7821 => x"84baf022",
          7822 => x"70101010",
          7823 => x"84baf408",
          7824 => x"05f80555",
          7825 => x"55768215",
          7826 => x"34810b83",
          7827 => x"15347754",
          7828 => x"77802efe",
          7829 => x"c638fecc",
          7830 => x"39ff3d0d",
          7831 => x"028f0533",
          7832 => x"51815270",
          7833 => x"72268738",
          7834 => x"84bb8011",
          7835 => x"33527184",
          7836 => x"bb840c83",
          7837 => x"3d0d04fe",
          7838 => x"3d0d0293",
          7839 => x"05335283",
          7840 => x"53718126",
          7841 => x"9d387151",
          7842 => x"d4bb3f84",
          7843 => x"bb840881",
          7844 => x"ff065372",
          7845 => x"87387284",
          7846 => x"bb801334",
          7847 => x"84bb8012",
          7848 => x"33537284",
          7849 => x"bb840c84",
          7850 => x"3d0d04f7",
          7851 => x"3d0d7c7e",
          7852 => x"60028c05",
          7853 => x"af05335a",
          7854 => x"5c575981",
          7855 => x"54767426",
          7856 => x"873884bb",
          7857 => x"80173354",
          7858 => x"73810654",
          7859 => x"835573bd",
          7860 => x"38735885",
          7861 => x"0b87c098",
          7862 => x"8c0c7853",
          7863 => x"75527651",
          7864 => x"d5ca3f84",
          7865 => x"bb840881",
          7866 => x"ff065574",
          7867 => x"802ea738",
          7868 => x"87c0988c",
          7869 => x"085473e2",
          7870 => x"38797826",
          7871 => x"d63874fc",
          7872 => x"80800654",
          7873 => x"73802e83",
          7874 => x"38815473",
          7875 => x"557484bb",
          7876 => x"840c8b3d",
          7877 => x"0d048480",
          7878 => x"16811970",
          7879 => x"81ff065a",
          7880 => x"55567978",
          7881 => x"26ffac38",
          7882 => x"d539f73d",
          7883 => x"0d7c7e60",
          7884 => x"028c05af",
          7885 => x"05335a5c",
          7886 => x"57598154",
          7887 => x"76742687",
          7888 => x"3884bb80",
          7889 => x"17335473",
          7890 => x"81065483",
          7891 => x"5573bd38",
          7892 => x"7358850b",
          7893 => x"87c0988c",
          7894 => x"0c785375",
          7895 => x"527651d7",
          7896 => x"8e3f84bb",
          7897 => x"840881ff",
          7898 => x"06557480",
          7899 => x"2ea73887",
          7900 => x"c0988c08",
          7901 => x"5473e238",
          7902 => x"797826d6",
          7903 => x"3874fc80",
          7904 => x"80065473",
          7905 => x"802e8338",
          7906 => x"81547355",
          7907 => x"7484bb84",
          7908 => x"0c8b3d0d",
          7909 => x"04848016",
          7910 => x"81197081",
          7911 => x"ff065a55",
          7912 => x"56797826",
          7913 => x"ffac38d5",
          7914 => x"39fc3d0d",
          7915 => x"78028405",
          7916 => x"9b053302",
          7917 => x"88059f05",
          7918 => x"33535355",
          7919 => x"81537173",
          7920 => x"26873884",
          7921 => x"bb801233",
          7922 => x"53728106",
          7923 => x"54835373",
          7924 => x"9b38850b",
          7925 => x"87c0988c",
          7926 => x"0c815370",
          7927 => x"732e9638",
          7928 => x"727125ad",
          7929 => x"3870832e",
          7930 => x"9a388453",
          7931 => x"7284bb84",
          7932 => x"0c863d0d",
          7933 => x"0488800a",
          7934 => x"750c7384",
          7935 => x"bb840c86",
          7936 => x"3d0d0481",
          7937 => x"80750c80",
          7938 => x"0b84bb84",
          7939 => x"0c863d0d",
          7940 => x"0471842b",
          7941 => x"87c0928c",
          7942 => x"11535470",
          7943 => x"cd387108",
          7944 => x"70812a81",
          7945 => x"06515170",
          7946 => x"802e8a38",
          7947 => x"87c0988c",
          7948 => x"085574ea",
          7949 => x"3887c098",
          7950 => x"8c085170",
          7951 => x"ca388172",
          7952 => x"0c87c092",
          7953 => x"8c145271",
          7954 => x"08820654",
          7955 => x"73802eff",
          7956 => x"9b387108",
          7957 => x"82065473",
          7958 => x"ee38ff90",
          7959 => x"39f63d0d",
          7960 => x"7c58800b",
          7961 => x"83193371",
          7962 => x"5b565774",
          7963 => x"772e0981",
          7964 => x"06a83877",
          7965 => x"33567583",
          7966 => x"2e818738",
          7967 => x"80538052",
          7968 => x"81183351",
          7969 => x"fea33f84",
          7970 => x"bb840880",
          7971 => x"2e833881",
          7972 => x"597884bb",
          7973 => x"840c8c3d",
          7974 => x"0d048154",
          7975 => x"b4180853",
          7976 => x"b8187053",
          7977 => x"81193352",
          7978 => x"5afcff3f",
          7979 => x"815984bb",
          7980 => x"8408772e",
          7981 => x"098106d9",
          7982 => x"3884bb84",
          7983 => x"08831934",
          7984 => x"b4180870",
          7985 => x"a81a0831",
          7986 => x"a01a0884",
          7987 => x"bb84085c",
          7988 => x"58565b74",
          7989 => x"7627ff9b",
          7990 => x"38821833",
          7991 => x"5574822e",
          7992 => x"098106ff",
          7993 => x"8e388154",
          7994 => x"751b5379",
          7995 => x"52811833",
          7996 => x"51fcb73f",
          7997 => x"76783357",
          7998 => x"5975832e",
          7999 => x"098106fe",
          8000 => x"fb388418",
          8001 => x"33577681",
          8002 => x"2e098106",
          8003 => x"feee38b8",
          8004 => x"185a8480",
          8005 => x"7a565780",
          8006 => x"75708105",
          8007 => x"5734ff17",
          8008 => x"5776f438",
          8009 => x"80d50b84",
          8010 => x"b61934ff",
          8011 => x"aa0b84b7",
          8012 => x"193480d2",
          8013 => x"7a3480d2",
          8014 => x"0bb91934",
          8015 => x"80e10bba",
          8016 => x"193480c1",
          8017 => x"0bbb1934",
          8018 => x"80f20b84",
          8019 => x"9c193480",
          8020 => x"f20b849d",
          8021 => x"193480c1",
          8022 => x"0b849e19",
          8023 => x"3480e10b",
          8024 => x"849f1934",
          8025 => x"94180855",
          8026 => x"7484a019",
          8027 => x"3474882a",
          8028 => x"5b7a84a1",
          8029 => x"19347490",
          8030 => x"2a567584",
          8031 => x"a2193474",
          8032 => x"982a5b7a",
          8033 => x"84a31934",
          8034 => x"9018085b",
          8035 => x"7a84a419",
          8036 => x"347a882a",
          8037 => x"557484a5",
          8038 => x"19347a90",
          8039 => x"2a567584",
          8040 => x"a619347a",
          8041 => x"982a5574",
          8042 => x"84a71934",
          8043 => x"a4180881",
          8044 => x"0570b41a",
          8045 => x"0c5b8154",
          8046 => x"7a537952",
          8047 => x"81183351",
          8048 => x"fae83f76",
          8049 => x"84193480",
          8050 => x"53805281",
          8051 => x"183351fb",
          8052 => x"d83f84bb",
          8053 => x"8408802e",
          8054 => x"fdb738fd",
          8055 => x"b239f33d",
          8056 => x"0d606070",
          8057 => x"08595656",
          8058 => x"81762788",
          8059 => x"389c1708",
          8060 => x"76268c38",
          8061 => x"81587784",
          8062 => x"bb840c8f",
          8063 => x"3d0d04ff",
          8064 => x"77335658",
          8065 => x"74822e81",
          8066 => x"cc387482",
          8067 => x"2482a538",
          8068 => x"74812e09",
          8069 => x"8106dd38",
          8070 => x"75812a16",
          8071 => x"70892aa8",
          8072 => x"1908055a",
          8073 => x"5a805bb4",
          8074 => x"1708792e",
          8075 => x"b0388317",
          8076 => x"335c7b7b",
          8077 => x"2e098106",
          8078 => x"83de3881",
          8079 => x"547853b8",
          8080 => x"17528117",
          8081 => x"3351f8e3",
          8082 => x"3f84bb84",
          8083 => x"08802e85",
          8084 => x"38ff5981",
          8085 => x"5b78b418",
          8086 => x"0c7aff9a",
          8087 => x"387983ff",
          8088 => x"0617b811",
          8089 => x"33811c70",
          8090 => x"892aa81b",
          8091 => x"0805535d",
          8092 => x"5d59b417",
          8093 => x"08792eb5",
          8094 => x"38800b83",
          8095 => x"1833715c",
          8096 => x"565d747d",
          8097 => x"2e098106",
          8098 => x"84b53881",
          8099 => x"547853b8",
          8100 => x"17528117",
          8101 => x"3351f893",
          8102 => x"3f84bb84",
          8103 => x"08802e85",
          8104 => x"38ff5981",
          8105 => x"5a78b418",
          8106 => x"0c79feca",
          8107 => x"387a83ff",
          8108 => x"0617b811",
          8109 => x"3370882b",
          8110 => x"7e077881",
          8111 => x"0671842a",
          8112 => x"535d5959",
          8113 => x"5d79feae",
          8114 => x"38769fff",
          8115 => x"0684bb84",
          8116 => x"0c8f3d0d",
          8117 => x"0475882a",
          8118 => x"a8180805",
          8119 => x"59b41708",
          8120 => x"792eb538",
          8121 => x"800b8318",
          8122 => x"33715c5d",
          8123 => x"5b7b7b2e",
          8124 => x"09810681",
          8125 => x"c2388154",
          8126 => x"7853b817",
          8127 => x"52811733",
          8128 => x"51f7a83f",
          8129 => x"84bb8408",
          8130 => x"802e8538",
          8131 => x"ff59815a",
          8132 => x"78b4180c",
          8133 => x"79fddf38",
          8134 => x"751083fe",
          8135 => x"067705b8",
          8136 => x"05811133",
          8137 => x"71337188",
          8138 => x"2b0784bb",
          8139 => x"840c575b",
          8140 => x"8f3d0d04",
          8141 => x"74832e09",
          8142 => x"8106fdb8",
          8143 => x"3875872a",
          8144 => x"a8180805",
          8145 => x"59b41708",
          8146 => x"792eb538",
          8147 => x"800b8318",
          8148 => x"33715c5e",
          8149 => x"5b7c7b2e",
          8150 => x"09810682",
          8151 => x"81388154",
          8152 => x"7853b817",
          8153 => x"52811733",
          8154 => x"51f6c03f",
          8155 => x"84bb8408",
          8156 => x"802e8538",
          8157 => x"ff59815a",
          8158 => x"78b4180c",
          8159 => x"79fcf738",
          8160 => x"75822b83",
          8161 => x"fc067705",
          8162 => x"b8058311",
          8163 => x"33821233",
          8164 => x"71902b71",
          8165 => x"882b0781",
          8166 => x"14337072",
          8167 => x"07882b75",
          8168 => x"337180ff",
          8169 => x"fffe8006",
          8170 => x"0784bb84",
          8171 => x"0c415c5e",
          8172 => x"595a568f",
          8173 => x"3d0d0481",
          8174 => x"54b41708",
          8175 => x"53b81770",
          8176 => x"53811833",
          8177 => x"525cf6e2",
          8178 => x"3f815a84",
          8179 => x"bb84087b",
          8180 => x"2e098106",
          8181 => x"febe3884",
          8182 => x"bb840883",
          8183 => x"1834b417",
          8184 => x"08a81808",
          8185 => x"3184bb84",
          8186 => x"085b5e7d",
          8187 => x"a0180827",
          8188 => x"fe843882",
          8189 => x"17335574",
          8190 => x"822e0981",
          8191 => x"06fdf738",
          8192 => x"8154b417",
          8193 => x"08a01808",
          8194 => x"05537b52",
          8195 => x"81173351",
          8196 => x"f6983f7a",
          8197 => x"5afddf39",
          8198 => x"8154b417",
          8199 => x"0853b817",
          8200 => x"70538118",
          8201 => x"33525cf6",
          8202 => x"813f84bb",
          8203 => x"84087b2e",
          8204 => x"09810682",
          8205 => x"813884bb",
          8206 => x"84088318",
          8207 => x"34b41708",
          8208 => x"a8180831",
          8209 => x"5d7ca018",
          8210 => x"08278b38",
          8211 => x"8217335e",
          8212 => x"7d822e81",
          8213 => x"cb3884bb",
          8214 => x"84085bfb",
          8215 => x"de398154",
          8216 => x"b4170853",
          8217 => x"b8177053",
          8218 => x"81183352",
          8219 => x"5cf5bb3f",
          8220 => x"815a84bb",
          8221 => x"84087b2e",
          8222 => x"098106fd",
          8223 => x"ff3884bb",
          8224 => x"84088318",
          8225 => x"34b41708",
          8226 => x"a8180831",
          8227 => x"84bb8408",
          8228 => x"5b5e7da0",
          8229 => x"180827fd",
          8230 => x"c5388217",
          8231 => x"33557482",
          8232 => x"2e098106",
          8233 => x"fdb83881",
          8234 => x"54b41708",
          8235 => x"a0180805",
          8236 => x"537b5281",
          8237 => x"173351f4",
          8238 => x"f13f7a5a",
          8239 => x"fda03981",
          8240 => x"54b41708",
          8241 => x"53b81770",
          8242 => x"53811833",
          8243 => x"525ef4da",
          8244 => x"3f815a84",
          8245 => x"bb84087d",
          8246 => x"2e098106",
          8247 => x"fbcb3884",
          8248 => x"bb840883",
          8249 => x"1834b417",
          8250 => x"08a81808",
          8251 => x"3184bb84",
          8252 => x"085b5574",
          8253 => x"a0180827",
          8254 => x"fb913882",
          8255 => x"17335574",
          8256 => x"822e0981",
          8257 => x"06fb8438",
          8258 => x"8154b417",
          8259 => x"08a01808",
          8260 => x"05537d52",
          8261 => x"81173351",
          8262 => x"f4903f7c",
          8263 => x"5afaec39",
          8264 => x"8154b417",
          8265 => x"08a01808",
          8266 => x"05537b52",
          8267 => x"81173351",
          8268 => x"f3f83ffa",
          8269 => x"8639815b",
          8270 => x"7af9bb38",
          8271 => x"fa9f39f2",
          8272 => x"3d0d6062",
          8273 => x"645d5759",
          8274 => x"82588176",
          8275 => x"279c3875",
          8276 => x"9c1a0827",
          8277 => x"95387833",
          8278 => x"5574782e",
          8279 => x"96387478",
          8280 => x"24818038",
          8281 => x"74812e82",
          8282 => x"8a387784",
          8283 => x"bb840c90",
          8284 => x"3d0d0475",
          8285 => x"882aa81a",
          8286 => x"08055880",
          8287 => x"0bb41a08",
          8288 => x"585c7678",
          8289 => x"2e86b638",
          8290 => x"8319337c",
          8291 => x"5b5d7c7c",
          8292 => x"2e098106",
          8293 => x"83fa3881",
          8294 => x"547753b8",
          8295 => x"19528119",
          8296 => x"3351f287",
          8297 => x"3f84bb84",
          8298 => x"08802e85",
          8299 => x"38ff5881",
          8300 => x"5a77b41a",
          8301 => x"0c795879",
          8302 => x"ffb03875",
          8303 => x"1083fe06",
          8304 => x"79057b83",
          8305 => x"ffff0658",
          8306 => x"5e76b81f",
          8307 => x"3476882a",
          8308 => x"5a79b91f",
          8309 => x"34810b83",
          8310 => x"1a347784",
          8311 => x"bb840c90",
          8312 => x"3d0d0474",
          8313 => x"832e0981",
          8314 => x"06feff38",
          8315 => x"75872aa8",
          8316 => x"1a080558",
          8317 => x"800bb41a",
          8318 => x"08585c76",
          8319 => x"782e85e1",
          8320 => x"38831933",
          8321 => x"7c5b5d7c",
          8322 => x"7c2e0981",
          8323 => x"0684bd38",
          8324 => x"81547753",
          8325 => x"b8195281",
          8326 => x"193351f1",
          8327 => x"8e3f84bb",
          8328 => x"8408802e",
          8329 => x"8538ff58",
          8330 => x"815a77b4",
          8331 => x"1a0c7958",
          8332 => x"79feb738",
          8333 => x"75822b83",
          8334 => x"fc067905",
          8335 => x"b8118311",
          8336 => x"3370982b",
          8337 => x"8f0a067e",
          8338 => x"f00a0607",
          8339 => x"41575e5c",
          8340 => x"7d7d347d",
          8341 => x"882a5675",
          8342 => x"b91d347d",
          8343 => x"902a5a79",
          8344 => x"ba1d347d",
          8345 => x"982a5b7a",
          8346 => x"bb1d3481",
          8347 => x"0b831a34",
          8348 => x"fee83975",
          8349 => x"812a1670",
          8350 => x"892aa81b",
          8351 => x"0805b41b",
          8352 => x"0859595a",
          8353 => x"76782eb7",
          8354 => x"38800b83",
          8355 => x"1a33715e",
          8356 => x"565d747d",
          8357 => x"2e098106",
          8358 => x"82d43881",
          8359 => x"547753b8",
          8360 => x"19528119",
          8361 => x"3351f083",
          8362 => x"3f84bb84",
          8363 => x"08802e85",
          8364 => x"38ff5881",
          8365 => x"5c77b41a",
          8366 => x"0c7b587b",
          8367 => x"fdac3879",
          8368 => x"83ff0619",
          8369 => x"b805811b",
          8370 => x"7781065f",
          8371 => x"5f577a55",
          8372 => x"7c802e8f",
          8373 => x"387a842b",
          8374 => x"9ff00677",
          8375 => x"338f0671",
          8376 => x"07565a74",
          8377 => x"7734810b",
          8378 => x"831a347d",
          8379 => x"892aa81a",
          8380 => x"08055680",
          8381 => x"0bb41a08",
          8382 => x"565f7476",
          8383 => x"2e83dd38",
          8384 => x"81547453",
          8385 => x"b8197053",
          8386 => x"811a3352",
          8387 => x"57f09b3f",
          8388 => x"815884bb",
          8389 => x"84087f2e",
          8390 => x"09810680",
          8391 => x"c73884bb",
          8392 => x"8408831a",
          8393 => x"34b41908",
          8394 => x"70a81b08",
          8395 => x"31a01b08",
          8396 => x"84bb8408",
          8397 => x"5b5c565c",
          8398 => x"747a278b",
          8399 => x"38821933",
          8400 => x"5574822e",
          8401 => x"82e43881",
          8402 => x"54755376",
          8403 => x"52811933",
          8404 => x"51eed83f",
          8405 => x"84bb8408",
          8406 => x"802e8538",
          8407 => x"ff568158",
          8408 => x"75b41a0c",
          8409 => x"77fc8338",
          8410 => x"7d83ff06",
          8411 => x"19b8057b",
          8412 => x"842a5656",
          8413 => x"7c8f387a",
          8414 => x"882a7633",
          8415 => x"81f00671",
          8416 => x"8f060756",
          8417 => x"5c747634",
          8418 => x"810b831a",
          8419 => x"34fccb39",
          8420 => x"81547653",
          8421 => x"b8197053",
          8422 => x"811a3352",
          8423 => x"5def8b3f",
          8424 => x"815a84bb",
          8425 => x"84087c2e",
          8426 => x"098106fc",
          8427 => x"883884bb",
          8428 => x"8408831a",
          8429 => x"34b41908",
          8430 => x"70a81b08",
          8431 => x"31a01b08",
          8432 => x"84bb8408",
          8433 => x"5d59405e",
          8434 => x"7e7727fb",
          8435 => x"ca388219",
          8436 => x"33557482",
          8437 => x"2e098106",
          8438 => x"fbbd3881",
          8439 => x"54761e53",
          8440 => x"7c528119",
          8441 => x"3351eec2",
          8442 => x"3f7b5afb",
          8443 => x"aa398154",
          8444 => x"7653b819",
          8445 => x"7053811a",
          8446 => x"335257ee",
          8447 => x"ad3f815c",
          8448 => x"84bb8408",
          8449 => x"7d2e0981",
          8450 => x"06fdae38",
          8451 => x"84bb8408",
          8452 => x"831a34b4",
          8453 => x"190870a8",
          8454 => x"1b0831a0",
          8455 => x"1b0884bb",
          8456 => x"84085f40",
          8457 => x"565f747e",
          8458 => x"27fcf038",
          8459 => x"82193355",
          8460 => x"74822e09",
          8461 => x"8106fce3",
          8462 => x"3881547d",
          8463 => x"1f537652",
          8464 => x"81193351",
          8465 => x"ede43f7c",
          8466 => x"5cfcd039",
          8467 => x"81547653",
          8468 => x"b8197053",
          8469 => x"811a3352",
          8470 => x"57edcf3f",
          8471 => x"815a84bb",
          8472 => x"84087c2e",
          8473 => x"098106fb",
          8474 => x"c53884bb",
          8475 => x"8408831a",
          8476 => x"34b41908",
          8477 => x"70a81b08",
          8478 => x"31a01b08",
          8479 => x"84bb8408",
          8480 => x"5d5f405e",
          8481 => x"7e7d27fb",
          8482 => x"87388219",
          8483 => x"33557482",
          8484 => x"2e098106",
          8485 => x"fafa3881",
          8486 => x"547c1e53",
          8487 => x"76528119",
          8488 => x"3351ed86",
          8489 => x"3f7b5afa",
          8490 => x"e7398154",
          8491 => x"791c5376",
          8492 => x"52811933",
          8493 => x"51ecf33f",
          8494 => x"7e58fd8b",
          8495 => x"397b7610",
          8496 => x"83fe067a",
          8497 => x"057c83ff",
          8498 => x"ff06595f",
          8499 => x"5876b81f",
          8500 => x"3476882a",
          8501 => x"5a79b91f",
          8502 => x"34f9fa39",
          8503 => x"7e58fd88",
          8504 => x"397b7682",
          8505 => x"2b83fc06",
          8506 => x"7a05b811",
          8507 => x"83113370",
          8508 => x"982b8f0a",
          8509 => x"067ff00a",
          8510 => x"06074258",
          8511 => x"5f5d587d",
          8512 => x"7d347d88",
          8513 => x"2a5675b9",
          8514 => x"1d347d90",
          8515 => x"2a5a79ba",
          8516 => x"1d347d98",
          8517 => x"2a5b7abb",
          8518 => x"1d34facf",
          8519 => x"39f63d0d",
          8520 => x"7c7e7108",
          8521 => x"5b5c5a7a",
          8522 => x"818a3890",
          8523 => x"19085776",
          8524 => x"802e80f4",
          8525 => x"38769c1a",
          8526 => x"082780ec",
          8527 => x"38941908",
          8528 => x"70565473",
          8529 => x"802e80d7",
          8530 => x"38767b2e",
          8531 => x"81933876",
          8532 => x"56811656",
          8533 => x"9c190876",
          8534 => x"26893882",
          8535 => x"56757726",
          8536 => x"82b23875",
          8537 => x"527951f0",
          8538 => x"f53f84bb",
          8539 => x"8408802e",
          8540 => x"81d03880",
          8541 => x"5884bb84",
          8542 => x"08812eb1",
          8543 => x"3884bb84",
          8544 => x"08097030",
          8545 => x"70720780",
          8546 => x"25707b07",
          8547 => x"51515555",
          8548 => x"7382aa38",
          8549 => x"75772e09",
          8550 => x"8106ffb5",
          8551 => x"38735574",
          8552 => x"84bb840c",
          8553 => x"8c3d0d04",
          8554 => x"8157ff91",
          8555 => x"3984bb84",
          8556 => x"0858ca39",
          8557 => x"7a527951",
          8558 => x"f0a43f81",
          8559 => x"557484bb",
          8560 => x"840827db",
          8561 => x"3884bb84",
          8562 => x"085584bb",
          8563 => x"8408ff2e",
          8564 => x"ce389c19",
          8565 => x"0884bb84",
          8566 => x"0826c438",
          8567 => x"7a57fedd",
          8568 => x"39811b56",
          8569 => x"9c190876",
          8570 => x"26833882",
          8571 => x"56755279",
          8572 => x"51efeb3f",
          8573 => x"805884bb",
          8574 => x"8408812e",
          8575 => x"81a03884",
          8576 => x"bb840809",
          8577 => x"70307072",
          8578 => x"07802570",
          8579 => x"7b0784bb",
          8580 => x"84085451",
          8581 => x"51555573",
          8582 => x"ff853884",
          8583 => x"bb840880",
          8584 => x"2e9a3890",
          8585 => x"19085481",
          8586 => x"7427fea3",
          8587 => x"38739c1a",
          8588 => x"0827fe9b",
          8589 => x"38737057",
          8590 => x"57fe9639",
          8591 => x"75802efe",
          8592 => x"8e38ff53",
          8593 => x"75527851",
          8594 => x"f5f53f84",
          8595 => x"bb840884",
          8596 => x"bb840830",
          8597 => x"7084bb84",
          8598 => x"08078025",
          8599 => x"5658557a",
          8600 => x"80c43874",
          8601 => x"80e33875",
          8602 => x"901a0c9c",
          8603 => x"1908fe05",
          8604 => x"941a0856",
          8605 => x"58747826",
          8606 => x"8638ff15",
          8607 => x"941a0c84",
          8608 => x"19338107",
          8609 => x"5a79841a",
          8610 => x"34755574",
          8611 => x"84bb840c",
          8612 => x"8c3d0d04",
          8613 => x"800b84bb",
          8614 => x"840c8c3d",
          8615 => x"0d0484bb",
          8616 => x"840858fe",
          8617 => x"da397380",
          8618 => x"2effb838",
          8619 => x"75537a52",
          8620 => x"7851f58b",
          8621 => x"3f84bb84",
          8622 => x"0855ffa7",
          8623 => x"3984bb84",
          8624 => x"0884bb84",
          8625 => x"0c8c3d0d",
          8626 => x"04ff5674",
          8627 => x"812effb9",
          8628 => x"388155ff",
          8629 => x"b639f83d",
          8630 => x"0d7a7c71",
          8631 => x"08595558",
          8632 => x"73f0800a",
          8633 => x"2680df38",
          8634 => x"739f0653",
          8635 => x"7280d738",
          8636 => x"7390190c",
          8637 => x"88180855",
          8638 => x"7480df38",
          8639 => x"76335675",
          8640 => x"822680cc",
          8641 => x"3873852a",
          8642 => x"53820b88",
          8643 => x"18225a56",
          8644 => x"727927a9",
          8645 => x"38ac1708",
          8646 => x"98190c74",
          8647 => x"94190c98",
          8648 => x"18085382",
          8649 => x"5672802e",
          8650 => x"94387389",
          8651 => x"2a139819",
          8652 => x"0c7383ff",
          8653 => x"0617b805",
          8654 => x"9c190c80",
          8655 => x"567584bb",
          8656 => x"840c8a3d",
          8657 => x"0d04820b",
          8658 => x"84bb840c",
          8659 => x"8a3d0d04",
          8660 => x"ac170855",
          8661 => x"74802eff",
          8662 => x"ac388a17",
          8663 => x"2270892b",
          8664 => x"57597376",
          8665 => x"27a5389c",
          8666 => x"170853fe",
          8667 => x"15fe1454",
          8668 => x"56805975",
          8669 => x"73278d38",
          8670 => x"8a172276",
          8671 => x"7129b019",
          8672 => x"08055a53",
          8673 => x"7898190c",
          8674 => x"ff913974",
          8675 => x"527751ec",
          8676 => x"cd3f84bb",
          8677 => x"84085584",
          8678 => x"bb8408ff",
          8679 => x"2ea43881",
          8680 => x"0b84bb84",
          8681 => x"0827ff9e",
          8682 => x"389c1708",
          8683 => x"5384bb84",
          8684 => x"087327ff",
          8685 => x"91387376",
          8686 => x"31547376",
          8687 => x"27cd38ff",
          8688 => x"aa39810b",
          8689 => x"84bb840c",
          8690 => x"8a3d0d04",
          8691 => x"f33d0d7f",
          8692 => x"70089012",
          8693 => x"08a0055c",
          8694 => x"5a57f080",
          8695 => x"0a7a2786",
          8696 => x"38800b98",
          8697 => x"180c9817",
          8698 => x"08558456",
          8699 => x"74802eb2",
          8700 => x"387983ff",
          8701 => x"065b7a9d",
          8702 => x"38811594",
          8703 => x"18085758",
          8704 => x"75a93879",
          8705 => x"852a881a",
          8706 => x"22575574",
          8707 => x"762781f5",
          8708 => x"38779818",
          8709 => x"0c799018",
          8710 => x"0c781bb8",
          8711 => x"059c180c",
          8712 => x"80567584",
          8713 => x"bb840c8f",
          8714 => x"3d0d0477",
          8715 => x"98180c8a",
          8716 => x"1922ff05",
          8717 => x"7a892a06",
          8718 => x"5c7bda38",
          8719 => x"75527651",
          8720 => x"eb9c3f84",
          8721 => x"bb84085d",
          8722 => x"8256810b",
          8723 => x"84bb8408",
          8724 => x"27d03881",
          8725 => x"5684bb84",
          8726 => x"08ff2ec6",
          8727 => x"389c1908",
          8728 => x"84bb8408",
          8729 => x"26829138",
          8730 => x"60802e81",
          8731 => x"98389417",
          8732 => x"08527651",
          8733 => x"f9a73f84",
          8734 => x"bb84085d",
          8735 => x"875684bb",
          8736 => x"8408802e",
          8737 => x"ff9c3882",
          8738 => x"5684bb84",
          8739 => x"08812eff",
          8740 => x"91388156",
          8741 => x"84bb8408",
          8742 => x"ff2eff86",
          8743 => x"3884bb84",
          8744 => x"08831a33",
          8745 => x"5f587d80",
          8746 => x"ea38fe18",
          8747 => x"9c1a08fe",
          8748 => x"05595680",
          8749 => x"5c757827",
          8750 => x"8d388a19",
          8751 => x"22767129",
          8752 => x"b01b0805",
          8753 => x"5d5e7bb4",
          8754 => x"1a0cb819",
          8755 => x"58848078",
          8756 => x"57558076",
          8757 => x"70810558",
          8758 => x"34ff1555",
          8759 => x"74f43874",
          8760 => x"568a1922",
          8761 => x"55757527",
          8762 => x"81803881",
          8763 => x"54751c53",
          8764 => x"77528119",
          8765 => x"3351e4b2",
          8766 => x"3f84bb84",
          8767 => x"0880e738",
          8768 => x"811656dd",
          8769 => x"397a9818",
          8770 => x"0c840b84",
          8771 => x"bb840c8f",
          8772 => x"3d0d0475",
          8773 => x"54b41908",
          8774 => x"53b81970",
          8775 => x"53811a33",
          8776 => x"5256e486",
          8777 => x"3f84bb84",
          8778 => x"0880f338",
          8779 => x"84bb8408",
          8780 => x"831a34b4",
          8781 => x"1908a81a",
          8782 => x"08315574",
          8783 => x"a01a0827",
          8784 => x"fee83882",
          8785 => x"19335c7b",
          8786 => x"822e0981",
          8787 => x"06fedb38",
          8788 => x"8154b419",
          8789 => x"08a01a08",
          8790 => x"05537552",
          8791 => x"81193351",
          8792 => x"e3c83ffe",
          8793 => x"c5398a19",
          8794 => x"22557483",
          8795 => x"ffff0655",
          8796 => x"74762e09",
          8797 => x"8106a738",
          8798 => x"7c94180c",
          8799 => x"fe1d9c1a",
          8800 => x"08fe055e",
          8801 => x"56805875",
          8802 => x"7d27fd85",
          8803 => x"388a1922",
          8804 => x"767129b0",
          8805 => x"1b080598",
          8806 => x"190c5cfc",
          8807 => x"f839810b",
          8808 => x"84bb840c",
          8809 => x"8f3d0d04",
          8810 => x"ee3d0d64",
          8811 => x"66415c84",
          8812 => x"7c085a5b",
          8813 => x"81ff7098",
          8814 => x"1e08585e",
          8815 => x"5e75802e",
          8816 => x"82d238b8",
          8817 => x"195f755a",
          8818 => x"8058b419",
          8819 => x"08762e82",
          8820 => x"d1388319",
          8821 => x"33785855",
          8822 => x"74782e09",
          8823 => x"81068194",
          8824 => x"38815475",
          8825 => x"53b81952",
          8826 => x"81193351",
          8827 => x"e1bd3f84",
          8828 => x"bb840880",
          8829 => x"2e8538ff",
          8830 => x"5a815779",
          8831 => x"b41a0c76",
          8832 => x"5b768290",
          8833 => x"389c1c08",
          8834 => x"70335858",
          8835 => x"76802e82",
          8836 => x"81388b18",
          8837 => x"33bf0670",
          8838 => x"81ff065b",
          8839 => x"4160861d",
          8840 => x"347681e5",
          8841 => x"32703078",
          8842 => x"ae327030",
          8843 => x"72802571",
          8844 => x"80250754",
          8845 => x"45455755",
          8846 => x"74933874",
          8847 => x"7adf0643",
          8848 => x"5661882e",
          8849 => x"81bf3875",
          8850 => x"602e8186",
          8851 => x"3881ff5d",
          8852 => x"80527b51",
          8853 => x"faf63f84",
          8854 => x"bb84085b",
          8855 => x"84bb8408",
          8856 => x"81b23898",
          8857 => x"1c085675",
          8858 => x"fedc387a",
          8859 => x"84bb840c",
          8860 => x"943d0d04",
          8861 => x"8154b419",
          8862 => x"08537e52",
          8863 => x"81193351",
          8864 => x"e1a83f81",
          8865 => x"5784bb84",
          8866 => x"08782e09",
          8867 => x"8106feef",
          8868 => x"3884bb84",
          8869 => x"08831a34",
          8870 => x"b41908a8",
          8871 => x"1a083184",
          8872 => x"bb840858",
          8873 => x"5b7aa01a",
          8874 => x"0827feb5",
          8875 => x"38821933",
          8876 => x"4160822e",
          8877 => x"098106fe",
          8878 => x"a8388154",
          8879 => x"b41908a0",
          8880 => x"1a080553",
          8881 => x"7e528119",
          8882 => x"3351e0de",
          8883 => x"3f7757fe",
          8884 => x"9039798f",
          8885 => x"2e098106",
          8886 => x"81e73876",
          8887 => x"862a8106",
          8888 => x"5b7a802e",
          8889 => x"93388d18",
          8890 => x"337781bf",
          8891 => x"0670901f",
          8892 => x"087fac05",
          8893 => x"0c595e5e",
          8894 => x"767d2eab",
          8895 => x"3881ff55",
          8896 => x"745dfecc",
          8897 => x"39815675",
          8898 => x"602e0981",
          8899 => x"06febe38",
          8900 => x"c139845b",
          8901 => x"800b981d",
          8902 => x"0c7a84bb",
          8903 => x"840c943d",
          8904 => x"0d04775b",
          8905 => x"fddf398d",
          8906 => x"1833577d",
          8907 => x"772e0981",
          8908 => x"06cb388c",
          8909 => x"19089b19",
          8910 => x"339a1a33",
          8911 => x"71882b07",
          8912 => x"58564175",
          8913 => x"ffb73877",
          8914 => x"337081bf",
          8915 => x"068d29f3",
          8916 => x"05515a81",
          8917 => x"76585b83",
          8918 => x"e7841733",
          8919 => x"78058111",
          8920 => x"33713371",
          8921 => x"882b0752",
          8922 => x"44567a80",
          8923 => x"2e80c538",
          8924 => x"7981fe26",
          8925 => x"ff873879",
          8926 => x"10610576",
          8927 => x"5c427562",
          8928 => x"23811a5a",
          8929 => x"8117578c",
          8930 => x"7727cc38",
          8931 => x"77337086",
          8932 => x"2a810659",
          8933 => x"5777802e",
          8934 => x"90387981",
          8935 => x"fe26fedd",
          8936 => x"38791061",
          8937 => x"05438063",
          8938 => x"23ff1d70",
          8939 => x"81ff065e",
          8940 => x"41fd9d39",
          8941 => x"7583ffff",
          8942 => x"2eca3881",
          8943 => x"ff55fec0",
          8944 => x"397ca838",
          8945 => x"7c558b57",
          8946 => x"74812a75",
          8947 => x"81802905",
          8948 => x"78708105",
          8949 => x"5a33407f",
          8950 => x"057081ff",
          8951 => x"06ff1959",
          8952 => x"565976e4",
          8953 => x"38747e2e",
          8954 => x"fd8138ff",
          8955 => x"0bac1d0c",
          8956 => x"7a84bb84",
          8957 => x"0c943d0d",
          8958 => x"04ef3d0d",
          8959 => x"6370085c",
          8960 => x"5c80527b",
          8961 => x"51f5cf3f",
          8962 => x"84bb8408",
          8963 => x"5a84bb84",
          8964 => x"08828038",
          8965 => x"81ff7040",
          8966 => x"5dff0bac",
          8967 => x"1d0cb81b",
          8968 => x"5e981c08",
          8969 => x"568058b4",
          8970 => x"1b08762e",
          8971 => x"82cc3883",
          8972 => x"1b337858",
          8973 => x"5574782e",
          8974 => x"09810681",
          8975 => x"df388154",
          8976 => x"7553b81b",
          8977 => x"52811b33",
          8978 => x"51dce03f",
          8979 => x"84bb8408",
          8980 => x"802e8538",
          8981 => x"ff568157",
          8982 => x"75b41c0c",
          8983 => x"765a7681",
          8984 => x"b2389c1c",
          8985 => x"08703358",
          8986 => x"5976802e",
          8987 => x"8499388b",
          8988 => x"1933bf06",
          8989 => x"7081ff06",
          8990 => x"57587786",
          8991 => x"1d347681",
          8992 => x"e52e80f2",
          8993 => x"3875832a",
          8994 => x"81065575",
          8995 => x"8f2e81ef",
          8996 => x"387480e2",
          8997 => x"38758f2e",
          8998 => x"81e5387c",
          8999 => x"aa38787d",
          9000 => x"56588b57",
          9001 => x"74812a75",
          9002 => x"81802905",
          9003 => x"78708105",
          9004 => x"5a335776",
          9005 => x"057081ff",
          9006 => x"06ff1959",
          9007 => x"565d76e4",
          9008 => x"38747f2e",
          9009 => x"80cd38ab",
          9010 => x"1c338106",
          9011 => x"5776a738",
          9012 => x"8b0ba01d",
          9013 => x"59577870",
          9014 => x"81055a33",
          9015 => x"78708105",
          9016 => x"5a337171",
          9017 => x"31ff1a5a",
          9018 => x"58424076",
          9019 => x"802e81dc",
          9020 => x"3875802e",
          9021 => x"e13881ff",
          9022 => x"5dff0bac",
          9023 => x"1d0c8052",
          9024 => x"7b51f5c8",
          9025 => x"3f84bb84",
          9026 => x"085a84bb",
          9027 => x"8408802e",
          9028 => x"fe8f3879",
          9029 => x"84bb840c",
          9030 => x"933d0d04",
          9031 => x"8154b41b",
          9032 => x"08537d52",
          9033 => x"811b3351",
          9034 => x"dc803f81",
          9035 => x"5784bb84",
          9036 => x"08782e09",
          9037 => x"8106fea4",
          9038 => x"3884bb84",
          9039 => x"08831c34",
          9040 => x"b41b08a8",
          9041 => x"1c083184",
          9042 => x"bb840858",
          9043 => x"5978a01c",
          9044 => x"0827fdea",
          9045 => x"38821b33",
          9046 => x"5a79822e",
          9047 => x"098106fd",
          9048 => x"dd388154",
          9049 => x"b41b08a0",
          9050 => x"1c080553",
          9051 => x"7d52811b",
          9052 => x"3351dbb6",
          9053 => x"3f7757fd",
          9054 => x"c539775a",
          9055 => x"fde439ab",
          9056 => x"1c337086",
          9057 => x"2a810642",
          9058 => x"5560fef2",
          9059 => x"3876862a",
          9060 => x"81065a79",
          9061 => x"802e9338",
          9062 => x"8d193377",
          9063 => x"81bf0670",
          9064 => x"901f087f",
          9065 => x"ac050c59",
          9066 => x"5e5f767d",
          9067 => x"2eaf3881",
          9068 => x"ff55745d",
          9069 => x"80527b51",
          9070 => x"f4923f84",
          9071 => x"bb84085a",
          9072 => x"84bb8408",
          9073 => x"802efcd9",
          9074 => x"38fec839",
          9075 => x"75802efe",
          9076 => x"c23881ff",
          9077 => x"5dff0bac",
          9078 => x"1d0cfea2",
          9079 => x"398d1933",
          9080 => x"577e772e",
          9081 => x"098106c7",
          9082 => x"388c1b08",
          9083 => x"9b1a339a",
          9084 => x"1b337188",
          9085 => x"2b075942",
          9086 => x"4076ffb3",
          9087 => x"38783370",
          9088 => x"bf068d29",
          9089 => x"f3055b55",
          9090 => x"81775956",
          9091 => x"83e78418",
          9092 => x"33790581",
          9093 => x"11337133",
          9094 => x"71882b07",
          9095 => x"52425775",
          9096 => x"802e80ed",
          9097 => x"387981fe",
          9098 => x"26ff8438",
          9099 => x"765181a0",
          9100 => x"d13f84bb",
          9101 => x"84087a10",
          9102 => x"61057022",
          9103 => x"5343811b",
          9104 => x"5b5681a0",
          9105 => x"bd3f7584",
          9106 => x"bb84082e",
          9107 => x"098106fe",
          9108 => x"de387656",
          9109 => x"8118588c",
          9110 => x"7827ffb0",
          9111 => x"38783370",
          9112 => x"862a8106",
          9113 => x"56597580",
          9114 => x"2e923874",
          9115 => x"802e8d38",
          9116 => x"79106005",
          9117 => x"70224141",
          9118 => x"7ffeb438",
          9119 => x"ff1d7081",
          9120 => x"ff065e5a",
          9121 => x"feae3984",
          9122 => x"0b84bb84",
          9123 => x"0c933d0d",
          9124 => x"047683ff",
          9125 => x"ff2effbc",
          9126 => x"3881ff55",
          9127 => x"fe9439ea",
          9128 => x"3d0d6870",
          9129 => x"0870ab13",
          9130 => x"3381a006",
          9131 => x"585a5d5e",
          9132 => x"86567485",
          9133 => x"b538748c",
          9134 => x"1d087022",
          9135 => x"57575d74",
          9136 => x"802e8e38",
          9137 => x"811d7010",
          9138 => x"17702251",
          9139 => x"565d74f4",
          9140 => x"38953da0",
          9141 => x"1f5b408c",
          9142 => x"607b5858",
          9143 => x"55757081",
          9144 => x"05573377",
          9145 => x"70810559",
          9146 => x"34ff1555",
          9147 => x"74ef3802",
          9148 => x"80db0533",
          9149 => x"70810658",
          9150 => x"5676802e",
          9151 => x"82aa3880",
          9152 => x"c00bab1f",
          9153 => x"34810b94",
          9154 => x"3d405b8c",
          9155 => x"1c087b58",
          9156 => x"598b7a61",
          9157 => x"5a575577",
          9158 => x"70810559",
          9159 => x"33767081",
          9160 => x"055834ff",
          9161 => x"155574ef",
          9162 => x"38857b27",
          9163 => x"80c2387a",
          9164 => x"79225657",
          9165 => x"74802eb8",
          9166 => x"3874821a",
          9167 => x"5a568f58",
          9168 => x"75810677",
          9169 => x"10077681",
          9170 => x"2a7083ff",
          9171 => x"ff067290",
          9172 => x"2a810644",
          9173 => x"58565760",
          9174 => x"802e8738",
          9175 => x"7684a0a1",
          9176 => x"3257ff18",
          9177 => x"58778025",
          9178 => x"d7387822",
          9179 => x"5574ca38",
          9180 => x"87028405",
          9181 => x"80cf0557",
          9182 => x"5876b007",
          9183 => x"bf0655b9",
          9184 => x"75278438",
          9185 => x"87155574",
          9186 => x"7634ff16",
          9187 => x"ff197884",
          9188 => x"2a595956",
          9189 => x"76e33877",
          9190 => x"1f5980fe",
          9191 => x"7934767a",
          9192 => x"58568078",
          9193 => x"27a03879",
          9194 => x"335574a0",
          9195 => x"2e983881",
          9196 => x"16567578",
          9197 => x"2788a238",
          9198 => x"751a7033",
          9199 => x"565774a0",
          9200 => x"2e098106",
          9201 => x"ea388116",
          9202 => x"56a05577",
          9203 => x"87268e38",
          9204 => x"983d7805",
          9205 => x"ec058119",
          9206 => x"71335759",
          9207 => x"41747734",
          9208 => x"87762787",
          9209 => x"f4387d51",
          9210 => x"f88f3f84",
          9211 => x"bb84088b",
          9212 => x"38811b5b",
          9213 => x"80e37b27",
          9214 => x"fe913887",
          9215 => x"567a80e4",
          9216 => x"2e82e738",
          9217 => x"84bb8408",
          9218 => x"5684bb84",
          9219 => x"08842e09",
          9220 => x"810682d6",
          9221 => x"380280db",
          9222 => x"0533ab1f",
          9223 => x"347d0802",
          9224 => x"840580db",
          9225 => x"05335758",
          9226 => x"75812a81",
          9227 => x"065f815b",
          9228 => x"7e802e90",
          9229 => x"388d528c",
          9230 => x"1d51fe88",
          9231 => x"e83f84bb",
          9232 => x"84081b5b",
          9233 => x"80527d51",
          9234 => x"ed8c3f84",
          9235 => x"bb840856",
          9236 => x"84bb8408",
          9237 => x"81823884",
          9238 => x"bb8408b8",
          9239 => x"195e5998",
          9240 => x"1e085680",
          9241 => x"57b41808",
          9242 => x"762e85f3",
          9243 => x"38831833",
          9244 => x"407f772e",
          9245 => x"09810682",
          9246 => x"a3388154",
          9247 => x"7553b818",
          9248 => x"52811833",
          9249 => x"51d4a43f",
          9250 => x"84bb8408",
          9251 => x"802e8538",
          9252 => x"ff568157",
          9253 => x"75b4190c",
          9254 => x"765676bc",
          9255 => x"389c1e08",
          9256 => x"70335642",
          9257 => x"7481e52e",
          9258 => x"81c93874",
          9259 => x"30708025",
          9260 => x"7807565f",
          9261 => x"74802e81",
          9262 => x"c9388119",
          9263 => x"59787b2e",
          9264 => x"86893881",
          9265 => x"527d51ee",
          9266 => x"833f84bb",
          9267 => x"84085684",
          9268 => x"bb840880",
          9269 => x"2eff8838",
          9270 => x"87587584",
          9271 => x"2e818938",
          9272 => x"75587581",
          9273 => x"8338ff1b",
          9274 => x"407f81f3",
          9275 => x"38981e08",
          9276 => x"57b41c08",
          9277 => x"772eaf38",
          9278 => x"831c3378",
          9279 => x"57407f84",
          9280 => x"82388154",
          9281 => x"7653b81c",
          9282 => x"52811c33",
          9283 => x"51d39c3f",
          9284 => x"84bb8408",
          9285 => x"802e8538",
          9286 => x"ff578156",
          9287 => x"76b41d0c",
          9288 => x"75587580",
          9289 => x"c338a00b",
          9290 => x"9c1f0857",
          9291 => x"55807670",
          9292 => x"81055834",
          9293 => x"ff155574",
          9294 => x"f4388b0b",
          9295 => x"9c1f087b",
          9296 => x"58585575",
          9297 => x"70810557",
          9298 => x"33777081",
          9299 => x"055934ff",
          9300 => x"155574ef",
          9301 => x"389c1e08",
          9302 => x"ab1f3398",
          9303 => x"065e5a7c",
          9304 => x"8c1b3481",
          9305 => x"0b831d34",
          9306 => x"77567584",
          9307 => x"bb840c98",
          9308 => x"3d0d0481",
          9309 => x"75307080",
          9310 => x"25720757",
          9311 => x"405774fe",
          9312 => x"b9387459",
          9313 => x"81527d51",
          9314 => x"ecc23f84",
          9315 => x"bb840856",
          9316 => x"84bb8408",
          9317 => x"802efdc7",
          9318 => x"38febd39",
          9319 => x"8154b418",
          9320 => x"08537c52",
          9321 => x"81183351",
          9322 => x"d3803f84",
          9323 => x"bb840877",
          9324 => x"2e098106",
          9325 => x"83bf3884",
          9326 => x"bb840883",
          9327 => x"1934b418",
          9328 => x"08a81908",
          9329 => x"315574a0",
          9330 => x"1908278b",
          9331 => x"38821833",
          9332 => x"4160822e",
          9333 => x"84ac3884",
          9334 => x"bb840857",
          9335 => x"fd9c397f",
          9336 => x"852b901f",
          9337 => x"08713153",
          9338 => x"587d51e9",
          9339 => x"e93f84bb",
          9340 => x"84085884",
          9341 => x"bb8408fe",
          9342 => x"ef387984",
          9343 => x"bb840856",
          9344 => x"588b5774",
          9345 => x"812a7581",
          9346 => x"80290578",
          9347 => x"7081055a",
          9348 => x"33577605",
          9349 => x"7081ff06",
          9350 => x"ff195956",
          9351 => x"5d76e438",
          9352 => x"7481ff06",
          9353 => x"b81d4341",
          9354 => x"981e0857",
          9355 => x"8056b41c",
          9356 => x"08772eb2",
          9357 => x"38831c33",
          9358 => x"5b7a762e",
          9359 => x"09810682",
          9360 => x"c9388154",
          9361 => x"7653b81c",
          9362 => x"52811c33",
          9363 => x"51d0dc3f",
          9364 => x"84bb8408",
          9365 => x"802e8538",
          9366 => x"ff578156",
          9367 => x"76b41d0c",
          9368 => x"755875fe",
          9369 => x"83388c1c",
          9370 => x"089c1f08",
          9371 => x"6181ff06",
          9372 => x"5f5c5f60",
          9373 => x"8d1c348f",
          9374 => x"0b8b1c34",
          9375 => x"758c1c34",
          9376 => x"759a1c34",
          9377 => x"759b1c34",
          9378 => x"7c8d29f3",
          9379 => x"0576775a",
          9380 => x"58597683",
          9381 => x"ffff2e8b",
          9382 => x"3878101f",
          9383 => x"7022811b",
          9384 => x"5b585683",
          9385 => x"e7841833",
          9386 => x"7b055576",
          9387 => x"75708105",
          9388 => x"57347688",
          9389 => x"2a567575",
          9390 => x"34768538",
          9391 => x"83ffff57",
          9392 => x"8118588c",
          9393 => x"7827cb38",
          9394 => x"7683ffff",
          9395 => x"2e81b338",
          9396 => x"78101f70",
          9397 => x"22585876",
          9398 => x"802e81a6",
          9399 => x"387c7b34",
          9400 => x"810b831d",
          9401 => x"3480527d",
          9402 => x"51e9e13f",
          9403 => x"84bb8408",
          9404 => x"5884bb84",
          9405 => x"08fcf138",
          9406 => x"7fff0540",
          9407 => x"7ffea938",
          9408 => x"fbeb3981",
          9409 => x"54b41c08",
          9410 => x"53b81c70",
          9411 => x"53811d33",
          9412 => x"5259d096",
          9413 => x"3f815684",
          9414 => x"bb8408fc",
          9415 => x"833884bb",
          9416 => x"8408831d",
          9417 => x"34b41c08",
          9418 => x"a81d0831",
          9419 => x"84bb8408",
          9420 => x"574160a0",
          9421 => x"1d0827fb",
          9422 => x"c938821c",
          9423 => x"33426182",
          9424 => x"2e098106",
          9425 => x"fbbc3881",
          9426 => x"54b41c08",
          9427 => x"a01d0805",
          9428 => x"53785281",
          9429 => x"1c3351cf",
          9430 => x"d13f7756",
          9431 => x"fba43976",
          9432 => x"9c1f0870",
          9433 => x"33574356",
          9434 => x"7481e52e",
          9435 => x"098106fa",
          9436 => x"ba38fbff",
          9437 => x"39817057",
          9438 => x"5776802e",
          9439 => x"fa9f38fa",
          9440 => x"d7397c80",
          9441 => x"c0075dfe",
          9442 => x"d4398154",
          9443 => x"b41c0853",
          9444 => x"6152811c",
          9445 => x"3351cf92",
          9446 => x"3f84bb84",
          9447 => x"08762e09",
          9448 => x"8106bc38",
          9449 => x"84bb8408",
          9450 => x"831d34b4",
          9451 => x"1c08a81d",
          9452 => x"08315574",
          9453 => x"a01d0827",
          9454 => x"8a38821c",
          9455 => x"335f7e82",
          9456 => x"2eaa3884",
          9457 => x"bb840856",
          9458 => x"fcf83975",
          9459 => x"ff1c4158",
          9460 => x"7f802efa",
          9461 => x"9838fc87",
          9462 => x"39751a57",
          9463 => x"f7e83981",
          9464 => x"70595675",
          9465 => x"802efcfe",
          9466 => x"38fafd39",
          9467 => x"8154b41c",
          9468 => x"08a01d08",
          9469 => x"05536152",
          9470 => x"811c3351",
          9471 => x"ceac3ffc",
          9472 => x"c1398154",
          9473 => x"b41808a0",
          9474 => x"19080553",
          9475 => x"7c528118",
          9476 => x"3351ce96",
          9477 => x"3ff8e339",
          9478 => x"f33d0d7f",
          9479 => x"61710840",
          9480 => x"5e5c800b",
          9481 => x"961e3498",
          9482 => x"1c08802e",
          9483 => x"82b538ac",
          9484 => x"1c08ff2e",
          9485 => x"80d93880",
          9486 => x"7071608c",
          9487 => x"05087022",
          9488 => x"57585b5c",
          9489 => x"5872782e",
          9490 => x"bc387754",
          9491 => x"74147022",
          9492 => x"811b5b55",
          9493 => x"567a8295",
          9494 => x"3880d080",
          9495 => x"147083ff",
          9496 => x"ff06585a",
          9497 => x"768fff26",
          9498 => x"82833873",
          9499 => x"791a7611",
          9500 => x"70225d58",
          9501 => x"555b79d4",
          9502 => x"387a3070",
          9503 => x"80257030",
          9504 => x"7a065a5c",
          9505 => x"5e7c1894",
          9506 => x"0557800b",
          9507 => x"82183480",
          9508 => x"70891f59",
          9509 => x"57589c1c",
          9510 => x"08167033",
          9511 => x"81185856",
          9512 => x"5374a02e",
          9513 => x"b2387485",
          9514 => x"2e81bc38",
          9515 => x"75893270",
          9516 => x"30707207",
          9517 => x"8025555b",
          9518 => x"54778b26",
          9519 => x"90387280",
          9520 => x"2e8b38ae",
          9521 => x"77708105",
          9522 => x"59348118",
          9523 => x"58747770",
          9524 => x"81055934",
          9525 => x"8118588a",
          9526 => x"7627ffba",
          9527 => x"387c1888",
          9528 => x"0555800b",
          9529 => x"81163496",
          9530 => x"1d335372",
          9531 => x"a5387781",
          9532 => x"f338bf0b",
          9533 => x"961e3481",
          9534 => x"577c1794",
          9535 => x"0556800b",
          9536 => x"8217349c",
          9537 => x"1c088c11",
          9538 => x"33555373",
          9539 => x"89387389",
          9540 => x"1e349c1c",
          9541 => x"08538b13",
          9542 => x"33881e34",
          9543 => x"9c1c089c",
          9544 => x"11831133",
          9545 => x"82123371",
          9546 => x"902b7188",
          9547 => x"2b078114",
          9548 => x"33707207",
          9549 => x"882b7533",
          9550 => x"7107640c",
          9551 => x"59971633",
          9552 => x"96173371",
          9553 => x"882b075f",
          9554 => x"415b405a",
          9555 => x"565b5577",
          9556 => x"861e2399",
          9557 => x"15339816",
          9558 => x"3371882b",
          9559 => x"075d547b",
          9560 => x"841e238f",
          9561 => x"3d0d0481",
          9562 => x"e555fec0",
          9563 => x"39771d96",
          9564 => x"1181ff7a",
          9565 => x"31585b57",
          9566 => x"83b5527a",
          9567 => x"902b7407",
          9568 => x"518190d0",
          9569 => x"3f84bb84",
          9570 => x"0883ffff",
          9571 => x"065581ff",
          9572 => x"7527ad38",
          9573 => x"81762781",
          9574 => x"b3387488",
          9575 => x"2a54737a",
          9576 => x"34749718",
          9577 => x"34827805",
          9578 => x"58800b8c",
          9579 => x"1f08565b",
          9580 => x"78197511",
          9581 => x"70225c57",
          9582 => x"5479fd90",
          9583 => x"38fdba39",
          9584 => x"74307630",
          9585 => x"70780780",
          9586 => x"25728025",
          9587 => x"07585557",
          9588 => x"7580f938",
          9589 => x"747a3481",
          9590 => x"78055880",
          9591 => x"0b8c1f08",
          9592 => x"565bcd39",
          9593 => x"7273891f",
          9594 => x"335a5757",
          9595 => x"77802efe",
          9596 => x"88387c96",
          9597 => x"1e7e5759",
          9598 => x"54891433",
          9599 => x"ffbf115a",
          9600 => x"54789926",
          9601 => x"a4389c1c",
          9602 => x"088c1133",
          9603 => x"545b8876",
          9604 => x"27b43872",
          9605 => x"842a5372",
          9606 => x"81065e7d",
          9607 => x"802e8a38",
          9608 => x"a0147083",
          9609 => x"ffff0655",
          9610 => x"53737870",
          9611 => x"81055a34",
          9612 => x"81168116",
          9613 => x"81197189",
          9614 => x"13335e57",
          9615 => x"59565679",
          9616 => x"ffb738fd",
          9617 => x"b4397283",
          9618 => x"2a53cc39",
          9619 => x"807b3070",
          9620 => x"80257030",
          9621 => x"7306535d",
          9622 => x"5f58fca9",
          9623 => x"39ef3d0d",
          9624 => x"63700870",
          9625 => x"42575c80",
          9626 => x"65703357",
          9627 => x"555374af",
          9628 => x"2e833881",
          9629 => x"537480dc",
          9630 => x"2e81df38",
          9631 => x"72802e81",
          9632 => x"d9389816",
          9633 => x"08881d0c",
          9634 => x"7333963d",
          9635 => x"943d4142",
          9636 => x"559f7527",
          9637 => x"82a73873",
          9638 => x"428c1608",
          9639 => x"58805761",
          9640 => x"70708105",
          9641 => x"52335553",
          9642 => x"7381df38",
          9643 => x"727f0c73",
          9644 => x"ff2e81ec",
          9645 => x"3883ffff",
          9646 => x"74278b38",
          9647 => x"76101856",
          9648 => x"80762381",
          9649 => x"17577383",
          9650 => x"ffff0670",
          9651 => x"af327030",
          9652 => x"9f732771",
          9653 => x"80250757",
          9654 => x"5b5b5573",
          9655 => x"82903874",
          9656 => x"80dc2e82",
          9657 => x"89387480",
          9658 => x"ff26b238",
          9659 => x"83e6a00b",
          9660 => x"83e6a033",
          9661 => x"7081ff06",
          9662 => x"56545673",
          9663 => x"802e81ab",
          9664 => x"3873752e",
          9665 => x"8f388116",
          9666 => x"70337081",
          9667 => x"ff065654",
          9668 => x"5673ee38",
          9669 => x"7281ff06",
          9670 => x"5b7a8184",
          9671 => x"387681fe",
          9672 => x"2680fd38",
          9673 => x"7610185d",
          9674 => x"747d2381",
          9675 => x"17627070",
          9676 => x"81055233",
          9677 => x"56545773",
          9678 => x"802efef0",
          9679 => x"3880cb39",
          9680 => x"817380dc",
          9681 => x"32703070",
          9682 => x"80257307",
          9683 => x"51555855",
          9684 => x"72802ea1",
          9685 => x"38811470",
          9686 => x"46548074",
          9687 => x"33545572",
          9688 => x"af2edd38",
          9689 => x"7280dc32",
          9690 => x"70307080",
          9691 => x"25770751",
          9692 => x"545772e1",
          9693 => x"3872881d",
          9694 => x"0c733396",
          9695 => x"3d943d41",
          9696 => x"4255749f",
          9697 => x"26fe9038",
          9698 => x"b43983b5",
          9699 => x"52735181",
          9700 => x"8dae3f84",
          9701 => x"bb840883",
          9702 => x"ffff0654",
          9703 => x"73fe8d38",
          9704 => x"86547384",
          9705 => x"bb840c93",
          9706 => x"3d0d0483",
          9707 => x"e6a03370",
          9708 => x"81ff065c",
          9709 => x"537a802e",
          9710 => x"fee338e4",
          9711 => x"39ff800b",
          9712 => x"ab1d3480",
          9713 => x"527b51de",
          9714 => x"8d3f84bb",
          9715 => x"840884bb",
          9716 => x"840c933d",
          9717 => x"0d048173",
          9718 => x"80dc3270",
          9719 => x"30708025",
          9720 => x"73074155",
          9721 => x"5a567d80",
          9722 => x"2ea13881",
          9723 => x"14428062",
          9724 => x"70335555",
          9725 => x"5672af2e",
          9726 => x"dd387280",
          9727 => x"dc327030",
          9728 => x"70802578",
          9729 => x"07405459",
          9730 => x"7de13873",
          9731 => x"610c9f75",
          9732 => x"27822b5a",
          9733 => x"76812e84",
          9734 => x"f8387682",
          9735 => x"2e83d138",
          9736 => x"76175976",
          9737 => x"802ea738",
          9738 => x"76177811",
          9739 => x"fe057022",
          9740 => x"70a03270",
          9741 => x"30709f2a",
          9742 => x"5242565f",
          9743 => x"56597cae",
          9744 => x"2e843872",
          9745 => x"8938ff17",
          9746 => x"5776dd38",
          9747 => x"76597719",
          9748 => x"56807623",
          9749 => x"76802efe",
          9750 => x"c7388078",
          9751 => x"227083ff",
          9752 => x"ff067258",
          9753 => x"5d55567a",
          9754 => x"a02e82e6",
          9755 => x"387383ff",
          9756 => x"ff065372",
          9757 => x"ae2e82f1",
          9758 => x"3876802e",
          9759 => x"aa387719",
          9760 => x"fe057022",
          9761 => x"5a5478ae",
          9762 => x"2e9d3876",
          9763 => x"1018fe05",
          9764 => x"54ff1757",
          9765 => x"76802e8f",
          9766 => x"38fe1470",
          9767 => x"225e547c",
          9768 => x"ae2e0981",
          9769 => x"06eb388b",
          9770 => x"0ba01d55",
          9771 => x"53a07470",
          9772 => x"81055634",
          9773 => x"ff135372",
          9774 => x"f4387273",
          9775 => x"5c5e8878",
          9776 => x"16702281",
          9777 => x"19595754",
          9778 => x"5d74802e",
          9779 => x"80ed3874",
          9780 => x"a02e83d0",
          9781 => x"3874ae32",
          9782 => x"70307080",
          9783 => x"25555a54",
          9784 => x"75772e85",
          9785 => x"ce387283",
          9786 => x"bb387259",
          9787 => x"7c7b2683",
          9788 => x"38815975",
          9789 => x"77327030",
          9790 => x"70720780",
          9791 => x"25707c07",
          9792 => x"51515454",
          9793 => x"72802e83",
          9794 => x"e0387c8b",
          9795 => x"2e868338",
          9796 => x"75772e8a",
          9797 => x"38798307",
          9798 => x"5a757726",
          9799 => x"9e387656",
          9800 => x"885b8b7e",
          9801 => x"822b81fc",
          9802 => x"06771857",
          9803 => x"5f5d7715",
          9804 => x"70228118",
          9805 => x"58565374",
          9806 => x"ff9538a0",
          9807 => x"1c335776",
          9808 => x"81e52e83",
          9809 => x"84387c88",
          9810 => x"2e82e338",
          9811 => x"7d8c0658",
          9812 => x"778c2e82",
          9813 => x"ed387d83",
          9814 => x"06557483",
          9815 => x"2e82e338",
          9816 => x"79812a81",
          9817 => x"0656759d",
          9818 => x"387d8106",
          9819 => x"5d7c802e",
          9820 => x"85387990",
          9821 => x"075a7d82",
          9822 => x"2a81065e",
          9823 => x"7d802e85",
          9824 => x"38798807",
          9825 => x"5a79ab1d",
          9826 => x"347b51e4",
          9827 => x"ec3f84bb",
          9828 => x"8408ab1d",
          9829 => x"33565484",
          9830 => x"bb840880",
          9831 => x"2e81ac38",
          9832 => x"84bb8408",
          9833 => x"842e0981",
          9834 => x"06fbf738",
          9835 => x"74852a81",
          9836 => x"065a7980",
          9837 => x"2e84f038",
          9838 => x"74822a81",
          9839 => x"06597882",
          9840 => x"98387b08",
          9841 => x"65555673",
          9842 => x"428c1608",
          9843 => x"588057f9",
          9844 => x"ce398116",
          9845 => x"70117911",
          9846 => x"70224040",
          9847 => x"56567ca0",
          9848 => x"2ef03875",
          9849 => x"802efd85",
          9850 => x"38798307",
          9851 => x"5afd8a39",
          9852 => x"82182256",
          9853 => x"75ae2e09",
          9854 => x"8106fcac",
          9855 => x"38772254",
          9856 => x"73ae2e09",
          9857 => x"8106fca0",
          9858 => x"38761018",
          9859 => x"5b807b23",
          9860 => x"800ba01d",
          9861 => x"5653ae54",
          9862 => x"76732683",
          9863 => x"38a05473",
          9864 => x"75708105",
          9865 => x"57348113",
          9866 => x"538a7327",
          9867 => x"e93879a0",
          9868 => x"075877ab",
          9869 => x"1d347b51",
          9870 => x"e3bf3f84",
          9871 => x"bb8408ab",
          9872 => x"1d335654",
          9873 => x"84bb8408",
          9874 => x"fed63874",
          9875 => x"822a8106",
          9876 => x"5877face",
          9877 => x"38861c33",
          9878 => x"70842a81",
          9879 => x"06565d74",
          9880 => x"802e83cd",
          9881 => x"38901c08",
          9882 => x"83ff0660",
          9883 => x"0580d311",
          9884 => x"3380d212",
          9885 => x"3371882b",
          9886 => x"07623341",
          9887 => x"5754547d",
          9888 => x"832e82d8",
          9889 => x"3874881d",
          9890 => x"0c7b0865",
          9891 => x"5556feb7",
          9892 => x"39772255",
          9893 => x"74ae2efe",
          9894 => x"f0387617",
          9895 => x"5976fb88",
          9896 => x"38fbab39",
          9897 => x"79830776",
          9898 => x"17565afd",
          9899 => x"81397d82",
          9900 => x"2b81fc06",
          9901 => x"708c0659",
          9902 => x"5e778c2e",
          9903 => x"098106fd",
          9904 => x"95387982",
          9905 => x"075afd98",
          9906 => x"39850ba0",
          9907 => x"1d347c88",
          9908 => x"2e098106",
          9909 => x"fcf638d6",
          9910 => x"39ff800b",
          9911 => x"ab1d3480",
          9912 => x"0b84bb84",
          9913 => x"0c933d0d",
          9914 => x"047480ff",
          9915 => x"269d3881",
          9916 => x"ff752780",
          9917 => x"c938ff1d",
          9918 => x"59787b26",
          9919 => x"81f73879",
          9920 => x"83077d77",
          9921 => x"18575c5a",
          9922 => x"fca43979",
          9923 => x"82075a83",
          9924 => x"b5527451",
          9925 => x"8185bd3f",
          9926 => x"84bb8408",
          9927 => x"83ffff06",
          9928 => x"70872a81",
          9929 => x"065a5578",
          9930 => x"802ec438",
          9931 => x"7480ff06",
          9932 => x"83e79411",
          9933 => x"33565474",
          9934 => x"81ff26ff",
          9935 => x"b9387480",
          9936 => x"2e818538",
          9937 => x"83e6ac0b",
          9938 => x"83e6ac33",
          9939 => x"7081ff06",
          9940 => x"56545973",
          9941 => x"802e80e0",
          9942 => x"3873752e",
          9943 => x"8f388119",
          9944 => x"70337081",
          9945 => x"ff065654",
          9946 => x"5973ee38",
          9947 => x"7281ff06",
          9948 => x"597880d4",
          9949 => x"38ffbf15",
          9950 => x"54739926",
          9951 => x"8a387d82",
          9952 => x"077081ff",
          9953 => x"065f53ff",
          9954 => x"9f155978",
          9955 => x"99269338",
          9956 => x"7d810770",
          9957 => x"81ff06e0",
          9958 => x"177083ff",
          9959 => x"ff065856",
          9960 => x"5f537b1b",
          9961 => x"a0055974",
          9962 => x"7934811b",
          9963 => x"5b751655",
          9964 => x"fafc3980",
          9965 => x"53fab339",
          9966 => x"83e6ac33",
          9967 => x"7081ff06",
          9968 => x"5a537880",
          9969 => x"2effae38",
          9970 => x"80df7a83",
          9971 => x"077d1da0",
          9972 => x"055b5b55",
          9973 => x"74793481",
          9974 => x"1b5bd239",
          9975 => x"80cd1433",
          9976 => x"80cc1533",
          9977 => x"71982b71",
          9978 => x"902b0777",
          9979 => x"07881f0c",
          9980 => x"5a57fd95",
          9981 => x"397b1ba0",
          9982 => x"0575882a",
          9983 => x"54547274",
          9984 => x"34811b7c",
          9985 => x"11a0055a",
          9986 => x"5b747934",
          9987 => x"811b5bff",
          9988 => x"9c397983",
          9989 => x"07a01d33",
          9990 => x"585a7681",
          9991 => x"e52e0981",
          9992 => x"06faa338",
          9993 => x"fda33974",
          9994 => x"822a8106",
          9995 => x"5c7bf6f2",
          9996 => x"38850b84",
          9997 => x"bb840c93",
          9998 => x"3d0d04eb",
          9999 => x"3d0d6769",
         10000 => x"02880580",
         10001 => x"e7053342",
         10002 => x"425e8061",
         10003 => x"0cff7e08",
         10004 => x"70595b42",
         10005 => x"79802e85",
         10006 => x"d7387970",
         10007 => x"81055b33",
         10008 => x"709f2656",
         10009 => x"5675ba2e",
         10010 => x"85d03874",
         10011 => x"ed3875ba",
         10012 => x"2e85c738",
         10013 => x"84e2e033",
         10014 => x"56807624",
         10015 => x"85b23875",
         10016 => x"101084e2",
         10017 => x"cc057008",
         10018 => x"585a8c58",
         10019 => x"76802e85",
         10020 => x"96387661",
         10021 => x"0c7f81fe",
         10022 => x"0677335d",
         10023 => x"597b802e",
         10024 => x"9b388117",
         10025 => x"3351ffbb",
         10026 => x"b03f84bb",
         10027 => x"840881ff",
         10028 => x"06708106",
         10029 => x"5e587c80",
         10030 => x"2e869638",
         10031 => x"80773475",
         10032 => x"165d84ba",
         10033 => x"f81d3381",
         10034 => x"18348152",
         10035 => x"81173351",
         10036 => x"ffbba43f",
         10037 => x"84bb8408",
         10038 => x"81ff0670",
         10039 => x"81064156",
         10040 => x"83587f84",
         10041 => x"c2387880",
         10042 => x"2e8d3875",
         10043 => x"822a8106",
         10044 => x"418a5860",
         10045 => x"84b13880",
         10046 => x"5b7a8318",
         10047 => x"34ff0bb4",
         10048 => x"180c7a7b",
         10049 => x"5a558154",
         10050 => x"7a53b817",
         10051 => x"70538118",
         10052 => x"335258ff",
         10053 => x"bb953f84",
         10054 => x"bb84087b",
         10055 => x"2e8538ff",
         10056 => x"55815974",
         10057 => x"b4180c84",
         10058 => x"56789938",
         10059 => x"84b71733",
         10060 => x"84b61833",
         10061 => x"71882b07",
         10062 => x"56568356",
         10063 => x"7482d4d5",
         10064 => x"2e85a538",
         10065 => x"7581268b",
         10066 => x"3884baf9",
         10067 => x"1d334261",
         10068 => x"85bf3881",
         10069 => x"5875842e",
         10070 => x"83cd388d",
         10071 => x"58758126",
         10072 => x"83c53880",
         10073 => x"c4173380",
         10074 => x"c3183371",
         10075 => x"882b075e",
         10076 => x"597c8480",
         10077 => x"2e098106",
         10078 => x"83ad3880",
         10079 => x"cf173380",
         10080 => x"ce183371",
         10081 => x"882b0757",
         10082 => x"5a75a438",
         10083 => x"80dc1783",
         10084 => x"11338212",
         10085 => x"3371902b",
         10086 => x"71882b07",
         10087 => x"81143370",
         10088 => x"7207882b",
         10089 => x"75337107",
         10090 => x"565a4543",
         10091 => x"5e5f5675",
         10092 => x"a0180c80",
         10093 => x"c8173382",
         10094 => x"183480c8",
         10095 => x"1733ff11",
         10096 => x"7081ff06",
         10097 => x"5f40598d",
         10098 => x"587c8126",
         10099 => x"82d93878",
         10100 => x"81ff0676",
         10101 => x"712980c5",
         10102 => x"19335a5f",
         10103 => x"5a778a18",
         10104 => x"23775977",
         10105 => x"802e87c4",
         10106 => x"38ff1878",
         10107 => x"06426187",
         10108 => x"bb3880ca",
         10109 => x"173380c9",
         10110 => x"18337188",
         10111 => x"2b075640",
         10112 => x"74881823",
         10113 => x"74758f06",
         10114 => x"5e5a8d58",
         10115 => x"7c829838",
         10116 => x"80cc1733",
         10117 => x"80cb1833",
         10118 => x"71882b07",
         10119 => x"565c74a4",
         10120 => x"3880d817",
         10121 => x"83113382",
         10122 => x"12337190",
         10123 => x"2b71882b",
         10124 => x"07811433",
         10125 => x"70720788",
         10126 => x"2b753371",
         10127 => x"0753445a",
         10128 => x"58424242",
         10129 => x"80c71733",
         10130 => x"80c61833",
         10131 => x"71882b07",
         10132 => x"5d588d58",
         10133 => x"7b802e81",
         10134 => x"ce387d1c",
         10135 => x"7a842a05",
         10136 => x"5a797526",
         10137 => x"81c13878",
         10138 => x"52747a31",
         10139 => x"51fdecb5",
         10140 => x"3f84bb84",
         10141 => x"085684bb",
         10142 => x"8408802e",
         10143 => x"81a93884",
         10144 => x"bb840880",
         10145 => x"fffffff5",
         10146 => x"26833883",
         10147 => x"5d7583ff",
         10148 => x"f5268338",
         10149 => x"825d759f",
         10150 => x"f52685eb",
         10151 => x"38815d82",
         10152 => x"16709c19",
         10153 => x"0c7ba419",
         10154 => x"0c7b1d70",
         10155 => x"a81a0c7b",
         10156 => x"1db01a0c",
         10157 => x"57597c83",
         10158 => x"2e8a8738",
         10159 => x"8817225c",
         10160 => x"8d587b80",
         10161 => x"2e80e038",
         10162 => x"7d16ac18",
         10163 => x"0c781955",
         10164 => x"7c822e8d",
         10165 => x"38781019",
         10166 => x"70812a7a",
         10167 => x"81060556",
         10168 => x"5a83ff15",
         10169 => x"892a598d",
         10170 => x"5878a018",
         10171 => x"0826b838",
         10172 => x"ff0b9418",
         10173 => x"0cff0b90",
         10174 => x"180cff80",
         10175 => x"0b841834",
         10176 => x"7c832e86",
         10177 => x"96387c77",
         10178 => x"3484e2dc",
         10179 => x"2281055d",
         10180 => x"7c84e2dc",
         10181 => x"237c8618",
         10182 => x"2384e2e4",
         10183 => x"0b8c180c",
         10184 => x"800b9818",
         10185 => x"0c805877",
         10186 => x"84bb840c",
         10187 => x"973d0d04",
         10188 => x"8b0b84bb",
         10189 => x"840c973d",
         10190 => x"0d047633",
         10191 => x"d0117081",
         10192 => x"ff065757",
         10193 => x"58748926",
         10194 => x"91388217",
         10195 => x"7881ff06",
         10196 => x"d0055d59",
         10197 => x"787a2e87",
         10198 => x"fe38807e",
         10199 => x"0883e6f4",
         10200 => x"5f405c7c",
         10201 => x"087f5a5b",
         10202 => x"7a708105",
         10203 => x"5c337970",
         10204 => x"81055b33",
         10205 => x"ff9f125a",
         10206 => x"58567799",
         10207 => x"268938e0",
         10208 => x"167081ff",
         10209 => x"065755ff",
         10210 => x"9f175877",
         10211 => x"99268938",
         10212 => x"e0177081",
         10213 => x"ff065855",
         10214 => x"7530709f",
         10215 => x"2a595575",
         10216 => x"772e0981",
         10217 => x"06853877",
         10218 => x"ffbe3878",
         10219 => x"7a327030",
         10220 => x"7072079f",
         10221 => x"2a7a075d",
         10222 => x"58557a80",
         10223 => x"2e879838",
         10224 => x"811c841e",
         10225 => x"5e5c837c",
         10226 => x"25ff9838",
         10227 => x"6156f9a9",
         10228 => x"3978802e",
         10229 => x"fecf3877",
         10230 => x"822a8106",
         10231 => x"5e8a587d",
         10232 => x"fec53880",
         10233 => x"58fec039",
         10234 => x"7a783357",
         10235 => x"597581e9",
         10236 => x"2e098106",
         10237 => x"83388159",
         10238 => x"7581eb32",
         10239 => x"70307080",
         10240 => x"257b075a",
         10241 => x"5b5c7783",
         10242 => x"ad387581",
         10243 => x"e82e83a6",
         10244 => x"38933d77",
         10245 => x"575a8359",
         10246 => x"83fa1633",
         10247 => x"70595b7a",
         10248 => x"802ea538",
         10249 => x"84811633",
         10250 => x"84801733",
         10251 => x"71902b71",
         10252 => x"882b0783",
         10253 => x"ff193370",
         10254 => x"7207882b",
         10255 => x"83fe1b33",
         10256 => x"71075259",
         10257 => x"5b404040",
         10258 => x"777a7084",
         10259 => x"055c0cff",
         10260 => x"19901757",
         10261 => x"59788025",
         10262 => x"ffbe3884",
         10263 => x"baf91d33",
         10264 => x"7030709f",
         10265 => x"2a727131",
         10266 => x"9b3d7110",
         10267 => x"1005f005",
         10268 => x"84b61c44",
         10269 => x"5d52435b",
         10270 => x"4278085b",
         10271 => x"83567a80",
         10272 => x"2e80fb38",
         10273 => x"800b8318",
         10274 => x"34ff0bb4",
         10275 => x"180c7a55",
         10276 => x"80567aff",
         10277 => x"2ea53881",
         10278 => x"547a53b8",
         10279 => x"17528117",
         10280 => x"3351ffb4",
         10281 => x"863f84bb",
         10282 => x"8408762e",
         10283 => x"8538ff55",
         10284 => x"815674b4",
         10285 => x"180c8458",
         10286 => x"75bf3881",
         10287 => x"1f337f33",
         10288 => x"71882b07",
         10289 => x"5d5e8358",
         10290 => x"7b82d4d5",
         10291 => x"2e098106",
         10292 => x"a838800b",
         10293 => x"b8183357",
         10294 => x"587581e9",
         10295 => x"2e82b738",
         10296 => x"7581eb32",
         10297 => x"70307080",
         10298 => x"257a0742",
         10299 => x"42427fbc",
         10300 => x"387581e8",
         10301 => x"2eb63882",
         10302 => x"587781ff",
         10303 => x"0656800b",
         10304 => x"84baf91e",
         10305 => x"335d587b",
         10306 => x"782e0981",
         10307 => x"06833881",
         10308 => x"58817627",
         10309 => x"f8bd3877",
         10310 => x"802ef8b7",
         10311 => x"38811a84",
         10312 => x"1a5a5a83",
         10313 => x"7a27fed1",
         10314 => x"38f8a839",
         10315 => x"830b80ee",
         10316 => x"1883e6b4",
         10317 => x"405d587b",
         10318 => x"7081055d",
         10319 => x"337e7081",
         10320 => x"05403371",
         10321 => x"7131ff1b",
         10322 => x"5b525656",
         10323 => x"77802e80",
         10324 => x"c5387580",
         10325 => x"2ee13885",
         10326 => x"0b818a18",
         10327 => x"83e6b840",
         10328 => x"5d587b70",
         10329 => x"81055d33",
         10330 => x"7e708105",
         10331 => x"40337171",
         10332 => x"31ff1b5b",
         10333 => x"58424077",
         10334 => x"802e858e",
         10335 => x"3875802e",
         10336 => x"e1388258",
         10337 => x"fef3398d",
         10338 => x"587cfa93",
         10339 => x"387784bb",
         10340 => x"840c973d",
         10341 => x"0d047558",
         10342 => x"75802efe",
         10343 => x"dc38850b",
         10344 => x"818a1883",
         10345 => x"e6b8405d",
         10346 => x"58ffb739",
         10347 => x"8d0b84bb",
         10348 => x"840c973d",
         10349 => x"0d04830b",
         10350 => x"80ee1883",
         10351 => x"e6b45c5a",
         10352 => x"58787081",
         10353 => x"055a337a",
         10354 => x"7081055c",
         10355 => x"33717131",
         10356 => x"ff1b5b57",
         10357 => x"5f5f7780",
         10358 => x"2e83d138",
         10359 => x"74802ee1",
         10360 => x"38850b81",
         10361 => x"8a1883e6",
         10362 => x"b85c5a58",
         10363 => x"78708105",
         10364 => x"5a337a70",
         10365 => x"81055c33",
         10366 => x"717131ff",
         10367 => x"1b5b5842",
         10368 => x"4077802e",
         10369 => x"84913875",
         10370 => x"802ee138",
         10371 => x"933d7757",
         10372 => x"5a8359fc",
         10373 => x"83398158",
         10374 => x"fdc63980",
         10375 => x"e9173380",
         10376 => x"e8183371",
         10377 => x"882b0757",
         10378 => x"5575812e",
         10379 => x"098106f9",
         10380 => x"d538811b",
         10381 => x"58805ab4",
         10382 => x"1708782e",
         10383 => x"b1388317",
         10384 => x"335b7a7a",
         10385 => x"2e098106",
         10386 => x"829b3881",
         10387 => x"547753b8",
         10388 => x"17528117",
         10389 => x"3351ffb0",
         10390 => x"d23f84bb",
         10391 => x"8408802e",
         10392 => x"8538ff58",
         10393 => x"815a77b4",
         10394 => x"180c79f9",
         10395 => x"99387984",
         10396 => x"183484b7",
         10397 => x"173384b6",
         10398 => x"18337188",
         10399 => x"2b07575e",
         10400 => x"7582d4d5",
         10401 => x"2e098106",
         10402 => x"f8fc38b8",
         10403 => x"17831133",
         10404 => x"82123371",
         10405 => x"902b7188",
         10406 => x"2b078114",
         10407 => x"33707207",
         10408 => x"882b7533",
         10409 => x"71075e41",
         10410 => x"5945425c",
         10411 => x"5977848b",
         10412 => x"85a4d22e",
         10413 => x"098106f8",
         10414 => x"cd38849c",
         10415 => x"17831133",
         10416 => x"82123371",
         10417 => x"902b7188",
         10418 => x"2b078114",
         10419 => x"33707207",
         10420 => x"882b7533",
         10421 => x"71074744",
         10422 => x"405b5c5a",
         10423 => x"5e60868a",
         10424 => x"85e4f22e",
         10425 => x"098106f8",
         10426 => x"9d3884a0",
         10427 => x"17831133",
         10428 => x"82123371",
         10429 => x"902b7188",
         10430 => x"2b078114",
         10431 => x"33707207",
         10432 => x"882b7533",
         10433 => x"7107941e",
         10434 => x"0c5d84a4",
         10435 => x"1c831133",
         10436 => x"82123371",
         10437 => x"902b7188",
         10438 => x"2b078114",
         10439 => x"33707207",
         10440 => x"882b7533",
         10441 => x"71076290",
         10442 => x"050c5944",
         10443 => x"49465c45",
         10444 => x"40455b56",
         10445 => x"5a7c7734",
         10446 => x"84e2dc22",
         10447 => x"81055d7c",
         10448 => x"84e2dc23",
         10449 => x"7c861823",
         10450 => x"84e2e40b",
         10451 => x"8c180c80",
         10452 => x"0b98180c",
         10453 => x"f7cf397b",
         10454 => x"8324f8f0",
         10455 => x"387b7a7f",
         10456 => x"0c56f295",
         10457 => x"397554b4",
         10458 => x"170853b8",
         10459 => x"17705381",
         10460 => x"18335259",
         10461 => x"ffafb33f",
         10462 => x"84bb8408",
         10463 => x"7a2e0981",
         10464 => x"0681a438",
         10465 => x"84bb8408",
         10466 => x"831834b4",
         10467 => x"1708a818",
         10468 => x"0831407f",
         10469 => x"a0180827",
         10470 => x"8b388217",
         10471 => x"33416082",
         10472 => x"2e818d38",
         10473 => x"84bb8408",
         10474 => x"5afda039",
         10475 => x"74567480",
         10476 => x"2ef39138",
         10477 => x"850b818a",
         10478 => x"1883e6b8",
         10479 => x"5c5a58fc",
         10480 => x"ab3980e3",
         10481 => x"173380e2",
         10482 => x"18337188",
         10483 => x"2b075f5a",
         10484 => x"8d587df6",
         10485 => x"d2388817",
         10486 => x"224261f6",
         10487 => x"ca3880e4",
         10488 => x"17831133",
         10489 => x"82123371",
         10490 => x"902b7188",
         10491 => x"2b078114",
         10492 => x"33707207",
         10493 => x"882b7533",
         10494 => x"7107ac1e",
         10495 => x"0c5a7d82",
         10496 => x"2b5a4344",
         10497 => x"405940f5",
         10498 => x"d8397558",
         10499 => x"75802ef9",
         10500 => x"e8388258",
         10501 => x"f9e33975",
         10502 => x"802ef2a8",
         10503 => x"38933d77",
         10504 => x"575a8359",
         10505 => x"f7f23975",
         10506 => x"5a79f5da",
         10507 => x"38fcbf39",
         10508 => x"7554b417",
         10509 => x"08a01808",
         10510 => x"05537852",
         10511 => x"81173351",
         10512 => x"ffade73f",
         10513 => x"fc8539f0",
         10514 => x"3d0d0280",
         10515 => x"d3053364",
         10516 => x"7043933d",
         10517 => x"41575dff",
         10518 => x"765a4075",
         10519 => x"802e80e9",
         10520 => x"38787081",
         10521 => x"055a3370",
         10522 => x"9f265555",
         10523 => x"74ba2e80",
         10524 => x"e23873ed",
         10525 => x"3874ba2e",
         10526 => x"80d93884",
         10527 => x"e2e03354",
         10528 => x"80742480",
         10529 => x"c4387310",
         10530 => x"1084e2cc",
         10531 => x"05700855",
         10532 => x"5573802e",
         10533 => x"84388074",
         10534 => x"34625473",
         10535 => x"802e8638",
         10536 => x"80743462",
         10537 => x"5473750c",
         10538 => x"7c547c80",
         10539 => x"2e923880",
         10540 => x"53933d70",
         10541 => x"53840551",
         10542 => x"ef813f84",
         10543 => x"bb840854",
         10544 => x"7384bb84",
         10545 => x"0c923d0d",
         10546 => x"048b0b84",
         10547 => x"bb840c92",
         10548 => x"3d0d0475",
         10549 => x"33d01170",
         10550 => x"81ff0656",
         10551 => x"56577389",
         10552 => x"26913882",
         10553 => x"167781ff",
         10554 => x"06d0055c",
         10555 => x"5877792e",
         10556 => x"80f73880",
         10557 => x"7f0883e6",
         10558 => x"f45e5f5b",
         10559 => x"7b087e59",
         10560 => x"5a797081",
         10561 => x"055b3378",
         10562 => x"7081055a",
         10563 => x"33ff9f12",
         10564 => x"59575576",
         10565 => x"99268938",
         10566 => x"e0157081",
         10567 => x"ff065654",
         10568 => x"ff9f1657",
         10569 => x"76992689",
         10570 => x"38e01670",
         10571 => x"81ff0657",
         10572 => x"54743070",
         10573 => x"9f2a5854",
         10574 => x"74762e09",
         10575 => x"81068538",
         10576 => x"76ffbe38",
         10577 => x"77793270",
         10578 => x"30707207",
         10579 => x"9f2a7907",
         10580 => x"5c575479",
         10581 => x"802e9238",
         10582 => x"811b841d",
         10583 => x"5d5b837b",
         10584 => x"25ff9938",
         10585 => x"7f54fe98",
         10586 => x"397a8324",
         10587 => x"f7387a79",
         10588 => x"600c54fe",
         10589 => x"8b39e63d",
         10590 => x"0d6c0284",
         10591 => x"0580fb05",
         10592 => x"33565a89",
         10593 => x"5679802e",
         10594 => x"a63874bf",
         10595 => x"0670549d",
         10596 => x"3dcc0553",
         10597 => x"9e3d8405",
         10598 => x"5259ed9f",
         10599 => x"3f84bb84",
         10600 => x"085784bb",
         10601 => x"8408802e",
         10602 => x"8f38807a",
         10603 => x"0c765675",
         10604 => x"84bb840c",
         10605 => x"9c3d0d04",
         10606 => x"7e406d52",
         10607 => x"903d7052",
         10608 => x"5ce19a3f",
         10609 => x"84bb8408",
         10610 => x"5784bb84",
         10611 => x"08802e81",
         10612 => x"ba38789c",
         10613 => x"065d7c80",
         10614 => x"2e81ca38",
         10615 => x"76802e83",
         10616 => x"e0387684",
         10617 => x"2e84f238",
         10618 => x"78880759",
         10619 => x"76ffbb38",
         10620 => x"78832a81",
         10621 => x"06587780",
         10622 => x"2e81d138",
         10623 => x"669b1133",
         10624 => x"9a123371",
         10625 => x"882b0761",
         10626 => x"70334258",
         10627 => x"5d5e567d",
         10628 => x"832e8697",
         10629 => x"38800b8e",
         10630 => x"1734800b",
         10631 => x"8f1734a1",
         10632 => x"0b901734",
         10633 => x"80cc0b91",
         10634 => x"17346656",
         10635 => x"a00b8b17",
         10636 => x"347e6757",
         10637 => x"5e800b9a",
         10638 => x"1734800b",
         10639 => x"9b17347d",
         10640 => x"335d7c83",
         10641 => x"2e85d738",
         10642 => x"6658800b",
         10643 => x"9c193480",
         10644 => x"0b9d1934",
         10645 => x"800b9e19",
         10646 => x"34800b9f",
         10647 => x"19347e55",
         10648 => x"810b8316",
         10649 => x"347a802e",
         10650 => x"80e2387e",
         10651 => x"b411087c",
         10652 => x"7e085957",
         10653 => x"5f57817b",
         10654 => x"2789389c",
         10655 => x"16087b26",
         10656 => x"83ec3882",
         10657 => x"57807a0c",
         10658 => x"fea33902",
         10659 => x"80e70533",
         10660 => x"70982b5c",
         10661 => x"587a8025",
         10662 => x"feb83886",
         10663 => x"799c065e",
         10664 => x"577cfeb8",
         10665 => x"3876fe82",
         10666 => x"380280c2",
         10667 => x"05337084",
         10668 => x"2a81065d",
         10669 => x"567b82b0",
         10670 => x"3878812a",
         10671 => x"81065d7c",
         10672 => x"802e8938",
         10673 => x"75810658",
         10674 => x"77829538",
         10675 => x"78832a81",
         10676 => x"06567580",
         10677 => x"2e863878",
         10678 => x"80c00759",
         10679 => x"7eb41108",
         10680 => x"a01c0c67",
         10681 => x"a41c0c67",
         10682 => x"9b11339a",
         10683 => x"12337188",
         10684 => x"2b077333",
         10685 => x"405b4057",
         10686 => x"5b7b832e",
         10687 => x"81fb3877",
         10688 => x"881b0c9c",
         10689 => x"16831133",
         10690 => x"82123371",
         10691 => x"902b7188",
         10692 => x"2b078114",
         10693 => x"33707207",
         10694 => x"882b7533",
         10695 => x"7107608c",
         10696 => x"050c437f",
         10697 => x"7f0c4158",
         10698 => x"5e595686",
         10699 => x"1b22841b",
         10700 => x"2378901b",
         10701 => x"34800b91",
         10702 => x"1b34800b",
         10703 => x"9c1b0c80",
         10704 => x"0b941b0c",
         10705 => x"a81a5c84",
         10706 => x"807c5755",
         10707 => x"80767081",
         10708 => x"055834ff",
         10709 => x"155574f4",
         10710 => x"3878852a",
         10711 => x"81065978",
         10712 => x"802efcc9",
         10713 => x"388c1a08",
         10714 => x"5574802e",
         10715 => x"fcbf3874",
         10716 => x"941b0c8a",
         10717 => x"1b227089",
         10718 => x"2b881c08",
         10719 => x"77595a5a",
         10720 => x"5b763070",
         10721 => x"78078025",
         10722 => x"51557876",
         10723 => x"2783e738",
         10724 => x"81707606",
         10725 => x"5e5b7c80",
         10726 => x"2e83db38",
         10727 => x"77527951",
         10728 => x"ffacbb3f",
         10729 => x"84bb8408",
         10730 => x"5884bb84",
         10731 => x"08812683",
         10732 => x"38825784",
         10733 => x"bb8408ff",
         10734 => x"2eb63875",
         10735 => x"793156c1",
         10736 => x"390280c2",
         10737 => x"05339106",
         10738 => x"5e7d9538",
         10739 => x"78822a81",
         10740 => x"06557480",
         10741 => x"2efc9938",
         10742 => x"8857807a",
         10743 => x"0cfbce39",
         10744 => x"8757807a",
         10745 => x"0cfbc639",
         10746 => x"8457807a",
         10747 => x"0cfbbe39",
         10748 => x"7a767a31",
         10749 => x"5757ff89",
         10750 => x"39951633",
         10751 => x"94173371",
         10752 => x"982b7190",
         10753 => x"2b077a07",
         10754 => x"881d0c9c",
         10755 => x"18831133",
         10756 => x"82123371",
         10757 => x"902b7188",
         10758 => x"2b078114",
         10759 => x"33707207",
         10760 => x"882b7533",
         10761 => x"7107628c",
         10762 => x"050c4561",
         10763 => x"610c555a",
         10764 => x"545b585e",
         10765 => x"5c861b22",
         10766 => x"841b2378",
         10767 => x"901b3480",
         10768 => x"0b911b34",
         10769 => x"800b9c1b",
         10770 => x"0c800b94",
         10771 => x"1b0ca81a",
         10772 => x"5c84807c",
         10773 => x"5755fdf4",
         10774 => x"397b51cc",
         10775 => x"c23f84bb",
         10776 => x"84087988",
         10777 => x"075a5776",
         10778 => x"fac038fb",
         10779 => x"83397452",
         10780 => x"7b51ffaa",
         10781 => x"e93f84bb",
         10782 => x"84085d84",
         10783 => x"bb840880",
         10784 => x"2e80cb38",
         10785 => x"84bb8408",
         10786 => x"812efbf7",
         10787 => x"3884bb84",
         10788 => x"08ff2e82",
         10789 => x"b7388053",
         10790 => x"74527551",
         10791 => x"ffb1a03f",
         10792 => x"84bb8408",
         10793 => x"838f389c",
         10794 => x"1608fe11",
         10795 => x"94180859",
         10796 => x"56587675",
         10797 => x"27903881",
         10798 => x"1794170c",
         10799 => x"84163381",
         10800 => x"07557484",
         10801 => x"17347c55",
         10802 => x"777d26ff",
         10803 => x"a138807f",
         10804 => x"7f725f59",
         10805 => x"575db416",
         10806 => x"087e2eaf",
         10807 => x"38831633",
         10808 => x"58777d2e",
         10809 => x"09810681",
         10810 => x"eb388154",
         10811 => x"7d53b816",
         10812 => x"52811633",
         10813 => x"51ffa3b3",
         10814 => x"3f84bb84",
         10815 => x"08802e85",
         10816 => x"38ff5781",
         10817 => x"5c76b417",
         10818 => x"0c7e567b",
         10819 => x"ff1c9018",
         10820 => x"0c577b80",
         10821 => x"2efbb538",
         10822 => x"807a0cf9",
         10823 => x"9039800b",
         10824 => x"94173480",
         10825 => x"0b951734",
         10826 => x"fa9e3995",
         10827 => x"16339417",
         10828 => x"3371982b",
         10829 => x"71902b07",
         10830 => x"7d075d56",
         10831 => x"58800b8e",
         10832 => x"1734800b",
         10833 => x"8f1734a1",
         10834 => x"0b901734",
         10835 => x"80cc0b91",
         10836 => x"17346656",
         10837 => x"a00b8b17",
         10838 => x"347e6757",
         10839 => x"5e800b9a",
         10840 => x"1734800b",
         10841 => x"9b17347d",
         10842 => x"335d7c83",
         10843 => x"2e098106",
         10844 => x"f9d638ff",
         10845 => x"a9397798",
         10846 => x"1b0c76f8",
         10847 => x"ad387583",
         10848 => x"ff065978",
         10849 => x"802ef8a5",
         10850 => x"387efe19",
         10851 => x"9c1208fe",
         10852 => x"05405959",
         10853 => x"777e27f9",
         10854 => x"ea388a19",
         10855 => x"22787129",
         10856 => x"b01b0805",
         10857 => x"565b7480",
         10858 => x"2ef9d838",
         10859 => x"75892a15",
         10860 => x"709c1c0c",
         10861 => x"58815477",
         10862 => x"537b5281",
         10863 => x"193351ff",
         10864 => x"a1e93f84",
         10865 => x"bb840880",
         10866 => x"2ef7e238",
         10867 => x"8157807a",
         10868 => x"0cf7da39",
         10869 => x"8154b416",
         10870 => x"0853b816",
         10871 => x"70538117",
         10872 => x"335258ff",
         10873 => x"a2c43f84",
         10874 => x"bb84087d",
         10875 => x"2e098106",
         10876 => x"80ce3884",
         10877 => x"bb840883",
         10878 => x"1734b416",
         10879 => x"08a81708",
         10880 => x"3184bb84",
         10881 => x"085d5574",
         10882 => x"a0170827",
         10883 => x"fddc3882",
         10884 => x"16335574",
         10885 => x"822e0981",
         10886 => x"06fdcf38",
         10887 => x"8154b416",
         10888 => x"08a01708",
         10889 => x"05537752",
         10890 => x"81163351",
         10891 => x"ffa1fb3f",
         10892 => x"7c5cfdb6",
         10893 => x"3984bb84",
         10894 => x"0857807a",
         10895 => x"0cf6ee39",
         10896 => x"815cfdc5",
         10897 => x"39f23d0d",
         10898 => x"60636564",
         10899 => x"40405b59",
         10900 => x"807e0c89",
         10901 => x"5778802e",
         10902 => x"9f387808",
         10903 => x"5675802e",
         10904 => x"97387533",
         10905 => x"5574802e",
         10906 => x"8f388616",
         10907 => x"22841a22",
         10908 => x"595b7a78",
         10909 => x"2e83b438",
         10910 => x"8055745f",
         10911 => x"76557681",
         10912 => x"e7389119",
         10913 => x"33557481",
         10914 => x"df389019",
         10915 => x"33810657",
         10916 => x"87567680",
         10917 => x"2e81c838",
         10918 => x"9419088c",
         10919 => x"1a087131",
         10920 => x"56567975",
         10921 => x"2681ca38",
         10922 => x"79802e81",
         10923 => x"b0387583",
         10924 => x"ff065c7b",
         10925 => x"8299387e",
         10926 => x"8a1122ff",
         10927 => x"0577892a",
         10928 => x"065d587b",
         10929 => x"9b387582",
         10930 => x"d0388819",
         10931 => x"08558175",
         10932 => x"2783c338",
         10933 => x"74ff2e83",
         10934 => x"ae387498",
         10935 => x"1a0c7e58",
         10936 => x"981908fe",
         10937 => x"059c1908",
         10938 => x"fe055c57",
         10939 => x"767b2783",
         10940 => x"a5388a18",
         10941 => x"22707829",
         10942 => x"b01a0805",
         10943 => x"56567480",
         10944 => x"2e839338",
         10945 => x"7b157a89",
         10946 => x"2a5c577a",
         10947 => x"802e80e6",
         10948 => x"387a1c55",
         10949 => x"75752785",
         10950 => x"38757c31",
         10951 => x"5b7a5476",
         10952 => x"537c5281",
         10953 => x"183351ff",
         10954 => x"9f813f84",
         10955 => x"bb840882",
         10956 => x"d6389019",
         10957 => x"3370982b",
         10958 => x"59568078",
         10959 => x"24828738",
         10960 => x"7a892b57",
         10961 => x"7977317e",
         10962 => x"08187f0c",
         10963 => x"771e941b",
         10964 => x"08197059",
         10965 => x"941c0c5e",
         10966 => x"5a79fed2",
         10967 => x"38805675",
         10968 => x"84bb840c",
         10969 => x"903d0d04",
         10970 => x"7484bb84",
         10971 => x"0c903d0d",
         10972 => x"04745afe",
         10973 => x"b3399c19",
         10974 => x"08567577",
         10975 => x"2e80c838",
         10976 => x"90193370",
         10977 => x"982ba81b",
         10978 => x"525d5b7b",
         10979 => x"8025a338",
         10980 => x"81547553",
         10981 => x"7a528118",
         10982 => x"3351ff9f",
         10983 => x"8d3f84bb",
         10984 => x"840881e3",
         10985 => x"38901933",
         10986 => x"80ff0655",
         10987 => x"74901a34",
         10988 => x"7e588154",
         10989 => x"76537a52",
         10990 => x"81183351",
         10991 => x"ff9dec3f",
         10992 => x"84bb8408",
         10993 => x"81c13876",
         10994 => x"9c1a0c94",
         10995 => x"19085675",
         10996 => x"83ff0684",
         10997 => x"80713158",
         10998 => x"55797727",
         10999 => x"83387957",
         11000 => x"767d7a17",
         11001 => x"a8055759",
         11002 => x"5676802e",
         11003 => x"fed63874",
         11004 => x"70810556",
         11005 => x"33787081",
         11006 => x"055a34ff",
         11007 => x"16567580",
         11008 => x"2efec138",
         11009 => x"74708105",
         11010 => x"56337870",
         11011 => x"81055a34",
         11012 => x"ff165675",
         11013 => x"da38feac",
         11014 => x"39981908",
         11015 => x"527851ff",
         11016 => x"a3bc3f84",
         11017 => x"bb840855",
         11018 => x"fda43981",
         11019 => x"163351ff",
         11020 => x"9ca73f84",
         11021 => x"bb840881",
         11022 => x"065574fc",
         11023 => x"bb387479",
         11024 => x"085657fc",
         11025 => x"b5399c19",
         11026 => x"08773156",
         11027 => x"757b27fd",
         11028 => x"ef388480",
         11029 => x"7671291e",
         11030 => x"a81b5858",
         11031 => x"55757081",
         11032 => x"05573377",
         11033 => x"70810559",
         11034 => x"34ff1555",
         11035 => x"74802efd",
         11036 => x"cf387570",
         11037 => x"81055733",
         11038 => x"77708105",
         11039 => x"5934ff15",
         11040 => x"5574da38",
         11041 => x"fdba3981",
         11042 => x"0b911a34",
         11043 => x"810b84bb",
         11044 => x"840c903d",
         11045 => x"0d04820b",
         11046 => x"911a3482",
         11047 => x"0b84bb84",
         11048 => x"0c903d0d",
         11049 => x"04f13d0d",
         11050 => x"61646665",
         11051 => x"41415c59",
         11052 => x"807f0c89",
         11053 => x"5778802e",
         11054 => x"9f387808",
         11055 => x"5675802e",
         11056 => x"97387533",
         11057 => x"5574802e",
         11058 => x"8f388616",
         11059 => x"22841a22",
         11060 => x"595a7978",
         11061 => x"2e84a838",
         11062 => x"80557440",
         11063 => x"76557682",
         11064 => x"cc389119",
         11065 => x"33557482",
         11066 => x"c4389019",
         11067 => x"3370812a",
         11068 => x"81065858",
         11069 => x"87567680",
         11070 => x"2e82a938",
         11071 => x"9419087b",
         11072 => x"115d577b",
         11073 => x"77278438",
         11074 => x"76095b7a",
         11075 => x"802e8289",
         11076 => x"387683ff",
         11077 => x"065d7c82",
         11078 => x"cd387f8a",
         11079 => x"1122ff05",
         11080 => x"78892a06",
         11081 => x"5e587caa",
         11082 => x"387682f9",
         11083 => x"38881908",
         11084 => x"5574802e",
         11085 => x"838c3874",
         11086 => x"812e83ed",
         11087 => x"3874ff2e",
         11088 => x"83d83874",
         11089 => x"981a0c88",
         11090 => x"19088538",
         11091 => x"74881a0c",
         11092 => x"7f589019",
         11093 => x"3370982b",
         11094 => x"5b57807a",
         11095 => x"2482f938",
         11096 => x"981908fe",
         11097 => x"059c1908",
         11098 => x"fe055d57",
         11099 => x"767c2783",
         11100 => x"b8388a18",
         11101 => x"22707829",
         11102 => x"b01a0805",
         11103 => x"56567480",
         11104 => x"2e83a638",
         11105 => x"7c157b89",
         11106 => x"2a5b5c79",
         11107 => x"802e81a6",
         11108 => x"38791d55",
         11109 => x"75752785",
         11110 => x"38757d31",
         11111 => x"5a79547b",
         11112 => x"537d5281",
         11113 => x"183351ff",
         11114 => x"9b803f84",
         11115 => x"bb840882",
         11116 => x"e9389c19",
         11117 => x"087c3156",
         11118 => x"757a27ab",
         11119 => x"3884800b",
         11120 => x"a81a7772",
         11121 => x"29600558",
         11122 => x"58557570",
         11123 => x"81055733",
         11124 => x"77708105",
         11125 => x"5934ff15",
         11126 => x"5574ef38",
         11127 => x"90193380",
         11128 => x"ff065d7c",
         11129 => x"901a3479",
         11130 => x"892b587a",
         11131 => x"78317f08",
         11132 => x"19600c78",
         11133 => x"1f941b08",
         11134 => x"1a707194",
         11135 => x"1e0c8c1d",
         11136 => x"08595a58",
         11137 => x"5f5b7476",
         11138 => x"27833875",
         11139 => x"55748c1a",
         11140 => x"0c7afdfd",
         11141 => x"38901933",
         11142 => x"587780c0",
         11143 => x"075b7a90",
         11144 => x"1a348056",
         11145 => x"7584bb84",
         11146 => x"0c913d0d",
         11147 => x"047484bb",
         11148 => x"840c913d",
         11149 => x"0d049c19",
         11150 => x"087c2ea2",
         11151 => x"38941908",
         11152 => x"57768c1a",
         11153 => x"08279b38",
         11154 => x"81547b53",
         11155 => x"a8195281",
         11156 => x"183351ff",
         11157 => x"98d53f84",
         11158 => x"bb840881",
         11159 => x"bd389419",
         11160 => x"08577b9c",
         11161 => x"1a0c7683",
         11162 => x"ff068480",
         11163 => x"71315955",
         11164 => x"7a782783",
         11165 => x"387a5877",
         11166 => x"7916a805",
         11167 => x"7f595656",
         11168 => x"77802e93",
         11169 => x"38767081",
         11170 => x"05583375",
         11171 => x"70810557",
         11172 => x"34ff1656",
         11173 => x"75ef3890",
         11174 => x"1933ff80",
         11175 => x"075a7990",
         11176 => x"1a34fec7",
         11177 => x"39981908",
         11178 => x"527851ff",
         11179 => x"acef3f84",
         11180 => x"bb840855",
         11181 => x"84bb8408",
         11182 => x"fcfd3890",
         11183 => x"193358fe",
         11184 => x"d8397652",
         11185 => x"7851ffac",
         11186 => x"d43f84bb",
         11187 => x"84085584",
         11188 => x"bb8408fc",
         11189 => x"e238e439",
         11190 => x"81549c19",
         11191 => x"0853a819",
         11192 => x"52811833",
         11193 => x"51ff98c2",
         11194 => x"3f84bb84",
         11195 => x"08ac3890",
         11196 => x"193380ff",
         11197 => x"06567590",
         11198 => x"1a347f58",
         11199 => x"fce23981",
         11200 => x"163351ff",
         11201 => x"96d33f84",
         11202 => x"bb840881",
         11203 => x"065574fb",
         11204 => x"c7387479",
         11205 => x"085657fb",
         11206 => x"c139810b",
         11207 => x"911a3481",
         11208 => x"0b84bb84",
         11209 => x"0c913d0d",
         11210 => x"04820b91",
         11211 => x"1a34820b",
         11212 => x"84bb840c",
         11213 => x"913d0d04",
         11214 => x"f53d0d7d",
         11215 => x"58895777",
         11216 => x"802e9f38",
         11217 => x"77085675",
         11218 => x"802e9738",
         11219 => x"75335574",
         11220 => x"802e8f38",
         11221 => x"86162284",
         11222 => x"19225a5a",
         11223 => x"79792e83",
         11224 => x"d2388055",
         11225 => x"745c7656",
         11226 => x"7681ee38",
         11227 => x"90183370",
         11228 => x"862a8106",
         11229 => x"5c577a80",
         11230 => x"2e81de38",
         11231 => x"76982b56",
         11232 => x"80762483",
         11233 => x"c9387ba0",
         11234 => x"19085856",
         11235 => x"b4160877",
         11236 => x"2eb83880",
         11237 => x"0b831733",
         11238 => x"715b5c5a",
         11239 => x"7a7a2e09",
         11240 => x"810681c0",
         11241 => x"38815476",
         11242 => x"53b81652",
         11243 => x"81163351",
         11244 => x"ff95f83f",
         11245 => x"84bb8408",
         11246 => x"802e8538",
         11247 => x"ff578159",
         11248 => x"76b4170c",
         11249 => x"78567881",
         11250 => x"9038a418",
         11251 => x"088b1133",
         11252 => x"a0075657",
         11253 => x"748b1834",
         11254 => x"77088819",
         11255 => x"087083ff",
         11256 => x"ff065d5a",
         11257 => x"567a9a18",
         11258 => x"347a882a",
         11259 => x"5a799b18",
         11260 => x"349c1776",
         11261 => x"3396195c",
         11262 => x"565b7483",
         11263 => x"2e81c838",
         11264 => x"8c180855",
         11265 => x"747b3474",
         11266 => x"882a5b7a",
         11267 => x"9d183474",
         11268 => x"902a5675",
         11269 => x"9e183474",
         11270 => x"982a5978",
         11271 => x"9f183480",
         11272 => x"7a34800b",
         11273 => x"971834a1",
         11274 => x"0b981834",
         11275 => x"80cc0b99",
         11276 => x"1834800b",
         11277 => x"92183480",
         11278 => x"0b931834",
         11279 => x"7b5b810b",
         11280 => x"831c347b",
         11281 => x"51ff9895",
         11282 => x"3f84bb84",
         11283 => x"08901933",
         11284 => x"81bf065b",
         11285 => x"56799019",
         11286 => x"34755574",
         11287 => x"84bb840c",
         11288 => x"8d3d0d04",
         11289 => x"8154b416",
         11290 => x"0853b816",
         11291 => x"70538117",
         11292 => x"33525bff",
         11293 => x"95b43f81",
         11294 => x"5984bb84",
         11295 => x"087a2e09",
         11296 => x"8106fec0",
         11297 => x"3884bb84",
         11298 => x"08831734",
         11299 => x"b41608a8",
         11300 => x"17083184",
         11301 => x"bb84085a",
         11302 => x"5574a017",
         11303 => x"0827fe85",
         11304 => x"38821633",
         11305 => x"5574822e",
         11306 => x"098106fd",
         11307 => x"f8388154",
         11308 => x"b41608a0",
         11309 => x"17080553",
         11310 => x"7a528116",
         11311 => x"3351ff94",
         11312 => x"e93f7959",
         11313 => x"fddf3978",
         11314 => x"902a5574",
         11315 => x"94183474",
         11316 => x"882a5675",
         11317 => x"9518348c",
         11318 => x"18085574",
         11319 => x"7b347488",
         11320 => x"2a5b7a9d",
         11321 => x"18347490",
         11322 => x"2a56759e",
         11323 => x"18347498",
         11324 => x"2a59789f",
         11325 => x"1834807a",
         11326 => x"34800b97",
         11327 => x"1834a10b",
         11328 => x"98183480",
         11329 => x"cc0b9918",
         11330 => x"34800b92",
         11331 => x"1834800b",
         11332 => x"9318347b",
         11333 => x"5b810b83",
         11334 => x"1c347b51",
         11335 => x"ff96be3f",
         11336 => x"84bb8408",
         11337 => x"90193381",
         11338 => x"bf065b56",
         11339 => x"79901934",
         11340 => x"fea73981",
         11341 => x"163351ff",
         11342 => x"929f3f84",
         11343 => x"bb840881",
         11344 => x"065574fc",
         11345 => x"9d387478",
         11346 => x"085657fc",
         11347 => x"97398154",
         11348 => x"9c180853",
         11349 => x"a818527b",
         11350 => x"81113352",
         11351 => x"57ff93ca",
         11352 => x"3f815584",
         11353 => x"bb8408fd",
         11354 => x"f2389018",
         11355 => x"3380ff06",
         11356 => x"59789019",
         11357 => x"347ba019",
         11358 => x"085856b4",
         11359 => x"1608772e",
         11360 => x"098106fc",
         11361 => x"8e38fcc2",
         11362 => x"39f93d0d",
         11363 => x"79705255",
         11364 => x"fba63f84",
         11365 => x"bb840854",
         11366 => x"84bb8408",
         11367 => x"b1388956",
         11368 => x"74802e9e",
         11369 => x"38740853",
         11370 => x"72802e96",
         11371 => x"38723352",
         11372 => x"71802e8e",
         11373 => x"38861322",
         11374 => x"84162258",
         11375 => x"5271772e",
         11376 => x"96388052",
         11377 => x"71587554",
         11378 => x"75843875",
         11379 => x"750c7384",
         11380 => x"bb840c89",
         11381 => x"3d0d0481",
         11382 => x"133351ff",
         11383 => x"90fb3f84",
         11384 => x"bb840881",
         11385 => x"065372da",
         11386 => x"38737508",
         11387 => x"5356d539",
         11388 => x"f63d0dff",
         11389 => x"7d705b57",
         11390 => x"5b75802e",
         11391 => x"b2387570",
         11392 => x"81055733",
         11393 => x"709f2652",
         11394 => x"5271ba2e",
         11395 => x"ac3870ee",
         11396 => x"3871ba2e",
         11397 => x"a43884e2",
         11398 => x"e0335180",
         11399 => x"71249038",
         11400 => x"7084e2e0",
         11401 => x"34800b84",
         11402 => x"bb840c8c",
         11403 => x"3d0d048b",
         11404 => x"0b84bb84",
         11405 => x"0c8c3d0d",
         11406 => x"047833d0",
         11407 => x"117081ff",
         11408 => x"06535353",
         11409 => x"70892691",
         11410 => x"38821973",
         11411 => x"81ff06d0",
         11412 => x"05595473",
         11413 => x"762e80f5",
         11414 => x"38800b83",
         11415 => x"e6f45b58",
         11416 => x"79087956",
         11417 => x"57767081",
         11418 => x"05583375",
         11419 => x"70810557",
         11420 => x"33ff9f12",
         11421 => x"53545270",
         11422 => x"99268938",
         11423 => x"e0127081",
         11424 => x"ff065354",
         11425 => x"ff9f1351",
         11426 => x"70992689",
         11427 => x"38e01370",
         11428 => x"81ff0654",
         11429 => x"54713070",
         11430 => x"9f2a5551",
         11431 => x"71732e09",
         11432 => x"81068538",
         11433 => x"73ffbe38",
         11434 => x"74763270",
         11435 => x"30707207",
         11436 => x"9f2a7607",
         11437 => x"59525276",
         11438 => x"802e9238",
         11439 => x"8118841b",
         11440 => x"5b588378",
         11441 => x"25ff9938",
         11442 => x"7a51fecf",
         11443 => x"39778324",
         11444 => x"f7387776",
         11445 => x"5e51fec3",
         11446 => x"39ea3d0d",
         11447 => x"8053983d",
         11448 => x"cc055299",
         11449 => x"3d51d2d3",
         11450 => x"3f84bb84",
         11451 => x"085584bb",
         11452 => x"8408802e",
         11453 => x"8a387484",
         11454 => x"bb840c98",
         11455 => x"3d0d047a",
         11456 => x"5c685298",
         11457 => x"3dd00551",
         11458 => x"c6d33f84",
         11459 => x"bb840855",
         11460 => x"84bb8408",
         11461 => x"80c63802",
         11462 => x"80d70533",
         11463 => x"70982b58",
         11464 => x"5a807724",
         11465 => x"80e23802",
         11466 => x"b2053370",
         11467 => x"842a8106",
         11468 => x"57597580",
         11469 => x"2eb2387a",
         11470 => x"639b1133",
         11471 => x"9a123371",
         11472 => x"882b0773",
         11473 => x"335e5a5b",
         11474 => x"57587983",
         11475 => x"2ea43876",
         11476 => x"98190c74",
         11477 => x"84bb840c",
         11478 => x"983d0d04",
         11479 => x"84bb8408",
         11480 => x"842e0981",
         11481 => x"06ff8f38",
         11482 => x"850b84bb",
         11483 => x"840c983d",
         11484 => x"0d049516",
         11485 => x"33941733",
         11486 => x"71982b71",
         11487 => x"902b0779",
         11488 => x"07981b0c",
         11489 => x"5b54cc39",
         11490 => x"7a7e9812",
         11491 => x"0c587484",
         11492 => x"bb840c98",
         11493 => x"3d0d04ff",
         11494 => x"9e3d0d80",
         11495 => x"e63d0880",
         11496 => x"e63d085d",
         11497 => x"40807c34",
         11498 => x"805380e4",
         11499 => x"3dfdb405",
         11500 => x"5280e53d",
         11501 => x"51d1843f",
         11502 => x"84bb8408",
         11503 => x"5984bb84",
         11504 => x"0883c838",
         11505 => x"6080d93d",
         11506 => x"0c7f6198",
         11507 => x"110880dd",
         11508 => x"3d0c5880",
         11509 => x"db3d085b",
         11510 => x"5879802e",
         11511 => x"82cc3880",
         11512 => x"d83d983d",
         11513 => x"405ba052",
         11514 => x"7a51ffa5",
         11515 => x"e93f84bb",
         11516 => x"84085984",
         11517 => x"bb840883",
         11518 => x"92386080",
         11519 => x"df3d0858",
         11520 => x"56b41608",
         11521 => x"772eb138",
         11522 => x"84bb8408",
         11523 => x"8317335f",
         11524 => x"5d7d83c7",
         11525 => x"38815476",
         11526 => x"53b81652",
         11527 => x"81163351",
         11528 => x"ff8d883f",
         11529 => x"84bb8408",
         11530 => x"802e8538",
         11531 => x"ff578159",
         11532 => x"76b4170c",
         11533 => x"7882d438",
         11534 => x"80df3d08",
         11535 => x"9b11339a",
         11536 => x"12337188",
         11537 => x"2b076370",
         11538 => x"335d4059",
         11539 => x"56567883",
         11540 => x"2e82da38",
         11541 => x"7680db3d",
         11542 => x"0c80527a",
         11543 => x"51ffa4f6",
         11544 => x"3f84bb84",
         11545 => x"085984bb",
         11546 => x"8408829f",
         11547 => x"3880527a",
         11548 => x"51ffaab4",
         11549 => x"3f84bb84",
         11550 => x"085984bb",
         11551 => x"8408bb38",
         11552 => x"80df3d08",
         11553 => x"9b11339a",
         11554 => x"12337188",
         11555 => x"2b076370",
         11556 => x"33425859",
         11557 => x"5e567d83",
         11558 => x"2e81fd38",
         11559 => x"767a2ea4",
         11560 => x"3884bb84",
         11561 => x"08527a51",
         11562 => x"ffa6a13f",
         11563 => x"84bb8408",
         11564 => x"5984bb84",
         11565 => x"08802eff",
         11566 => x"b4387884",
         11567 => x"2e83d838",
         11568 => x"7881c838",
         11569 => x"80e43dfd",
         11570 => x"b805527a",
         11571 => x"51ffbec8",
         11572 => x"3f787f82",
         11573 => x"05335b57",
         11574 => x"79802e90",
         11575 => x"38821f56",
         11576 => x"81178117",
         11577 => x"70335f57",
         11578 => x"577cf538",
         11579 => x"81175675",
         11580 => x"78268195",
         11581 => x"3876802e",
         11582 => x"9c387e17",
         11583 => x"820556ff",
         11584 => x"1880e63d",
         11585 => x"0811ff19",
         11586 => x"ff195959",
         11587 => x"56587533",
         11588 => x"753476eb",
         11589 => x"38ff1880",
         11590 => x"e63d0811",
         11591 => x"5f58af7e",
         11592 => x"3480da3d",
         11593 => x"085a79fd",
         11594 => x"bd387760",
         11595 => x"2e828a38",
         11596 => x"800b84e2",
         11597 => x"e0337010",
         11598 => x"1083e6f4",
         11599 => x"05700870",
         11600 => x"33435959",
         11601 => x"5e5a7e7a",
         11602 => x"2e8d3881",
         11603 => x"1a701770",
         11604 => x"33575f5a",
         11605 => x"74f53882",
         11606 => x"1a5b7a78",
         11607 => x"26ab3880",
         11608 => x"57767a27",
         11609 => x"94387616",
         11610 => x"5f7e337c",
         11611 => x"7081055e",
         11612 => x"34811757",
         11613 => x"797726ee",
         11614 => x"38ba7c70",
         11615 => x"81055e34",
         11616 => x"76ff2e09",
         11617 => x"810681df",
         11618 => x"38915980",
         11619 => x"7c347884",
         11620 => x"bb840c80",
         11621 => x"e43d0d04",
         11622 => x"95163394",
         11623 => x"17337198",
         11624 => x"2b71902b",
         11625 => x"07790759",
         11626 => x"565efdf0",
         11627 => x"39951633",
         11628 => x"94173371",
         11629 => x"982b7190",
         11630 => x"2b077907",
         11631 => x"80dd3d0c",
         11632 => x"5a5d8052",
         11633 => x"7a51ffa2",
         11634 => x"8d3f84bb",
         11635 => x"84085984",
         11636 => x"bb840880",
         11637 => x"2efd9638",
         11638 => x"ffb13981",
         11639 => x"54b41608",
         11640 => x"53b81670",
         11641 => x"53811733",
         11642 => x"525eff8a",
         11643 => x"bd3f8159",
         11644 => x"84bb8408",
         11645 => x"fcbe3884",
         11646 => x"bb840883",
         11647 => x"1734b416",
         11648 => x"08a81708",
         11649 => x"3184bb84",
         11650 => x"085a5574",
         11651 => x"a0170827",
         11652 => x"fc833882",
         11653 => x"16335574",
         11654 => x"822e0981",
         11655 => x"06fbf638",
         11656 => x"8154b416",
         11657 => x"08a01708",
         11658 => x"05537d52",
         11659 => x"81163351",
         11660 => x"ff89f73f",
         11661 => x"7c59fbdd",
         11662 => x"39ff1880",
         11663 => x"e63d0811",
         11664 => x"5c58af7b",
         11665 => x"34800b84",
         11666 => x"e2e03370",
         11667 => x"101083e6",
         11668 => x"f4057008",
         11669 => x"70334359",
         11670 => x"595e5a7e",
         11671 => x"7a2e0981",
         11672 => x"06fde838",
         11673 => x"fdf13980",
         11674 => x"e53d0818",
         11675 => x"8119595a",
         11676 => x"79337c70",
         11677 => x"81055e34",
         11678 => x"776027fe",
         11679 => x"8e3880e5",
         11680 => x"3d081881",
         11681 => x"19595a79",
         11682 => x"337c7081",
         11683 => x"055e347f",
         11684 => x"7826d438",
         11685 => x"fdf53982",
         11686 => x"59807c34",
         11687 => x"7884bb84",
         11688 => x"0c80e43d",
         11689 => x"0d04f53d",
         11690 => x"0d7d7f5a",
         11691 => x"57895876",
         11692 => x"802e9f38",
         11693 => x"76085675",
         11694 => x"802e9738",
         11695 => x"75335574",
         11696 => x"802e8f38",
         11697 => x"86162284",
         11698 => x"18225b5b",
         11699 => x"7a7a2e83",
         11700 => x"ee388055",
         11701 => x"745c7755",
         11702 => x"7782fb38",
         11703 => x"91173355",
         11704 => x"7482f338",
         11705 => x"8c170858",
         11706 => x"78782682",
         11707 => x"f2389417",
         11708 => x"0856805a",
         11709 => x"787a2e83",
         11710 => x"85387b8a",
         11711 => x"11227089",
         11712 => x"2b525c58",
         11713 => x"757a2e82",
         11714 => x"fc387752",
         11715 => x"ff1951fd",
         11716 => x"bb933f84",
         11717 => x"bb8408ff",
         11718 => x"17795470",
         11719 => x"535755fd",
         11720 => x"bb833f84",
         11721 => x"bb840875",
         11722 => x"2682da38",
         11723 => x"77307606",
         11724 => x"7094190c",
         11725 => x"79713198",
         11726 => x"1908585a",
         11727 => x"5b75802e",
         11728 => x"81923877",
         11729 => x"792780d3",
         11730 => x"38787831",
         11731 => x"94180819",
         11732 => x"94190c90",
         11733 => x"18337081",
         11734 => x"2a810651",
         11735 => x"5c597a80",
         11736 => x"2e82cc38",
         11737 => x"75527651",
         11738 => x"ff9bb23f",
         11739 => x"84bb8408",
         11740 => x"5684bb84",
         11741 => x"08802e9e",
         11742 => x"3875ff2e",
         11743 => x"81d13881",
         11744 => x"76278382",
         11745 => x"387b5575",
         11746 => x"9c160827",
         11747 => x"82f83875",
         11748 => x"98180cff",
         11749 => x"ae3984bb",
         11750 => x"84085994",
         11751 => x"17081994",
         11752 => x"180c7883",
         11753 => x"ff065877",
         11754 => x"802ea938",
         11755 => x"7bfe179c",
         11756 => x"1208fe05",
         11757 => x"5c575875",
         11758 => x"7a2782ca",
         11759 => x"388a1822",
         11760 => x"767129b0",
         11761 => x"1a08057a",
         11762 => x"892a115c",
         11763 => x"5c557a80",
         11764 => x"2e82b338",
         11765 => x"8c170858",
         11766 => x"94170856",
         11767 => x"77762790",
         11768 => x"38758c18",
         11769 => x"0c901733",
         11770 => x"80c00759",
         11771 => x"78901834",
         11772 => x"7583ff06",
         11773 => x"5b7a802e",
         11774 => x"81ab389c",
         11775 => x"17085675",
         11776 => x"7a2e81a1",
         11777 => x"38901733",
         11778 => x"70982ba8",
         11779 => x"195a5659",
         11780 => x"748025a2",
         11781 => x"38815475",
         11782 => x"5377527b",
         11783 => x"81113352",
         11784 => x"56ff8686",
         11785 => x"3f84bb84",
         11786 => x"08a53890",
         11787 => x"173380ff",
         11788 => x"06557490",
         11789 => x"18348154",
         11790 => x"79537752",
         11791 => x"7b811133",
         11792 => x"5258ff84",
         11793 => x"e63f84bb",
         11794 => x"8408802e",
         11795 => x"80d33881",
         11796 => x"0b911834",
         11797 => x"81557484",
         11798 => x"bb840c8d",
         11799 => x"3d0d0490",
         11800 => x"17337081",
         11801 => x"2a810657",
         11802 => x"5a75fd82",
         11803 => x"38779418",
         11804 => x"08575980",
         11805 => x"5a787a2e",
         11806 => x"098106fc",
         11807 => x"fd387994",
         11808 => x"180cfed4",
         11809 => x"39800b94",
         11810 => x"180c8817",
         11811 => x"08567580",
         11812 => x"2e80c738",
         11813 => x"7598180c",
         11814 => x"75802efe",
         11815 => x"b738fda3",
         11816 => x"39799c18",
         11817 => x"0c800b84",
         11818 => x"bb840c8d",
         11819 => x"3d0d0475",
         11820 => x"527651ff",
         11821 => x"8aa83f84",
         11822 => x"bb840856",
         11823 => x"fdbb3981",
         11824 => x"163351ff",
         11825 => x"83933f84",
         11826 => x"bb840881",
         11827 => x"065574fc",
         11828 => x"81387477",
         11829 => x"085658fb",
         11830 => x"fb397552",
         11831 => x"7651ff98",
         11832 => x"bc3f84bb",
         11833 => x"84085684",
         11834 => x"bb840881",
         11835 => x"2e983884",
         11836 => x"bb8408ff",
         11837 => x"2efed838",
         11838 => x"84bb8408",
         11839 => x"88180c75",
         11840 => x"98180cff",
         11841 => x"9339820b",
         11842 => x"91183482",
         11843 => x"0b84bb84",
         11844 => x"0c8d3d0d",
         11845 => x"04f63d0d",
         11846 => x"7c568954",
         11847 => x"75802ea2",
         11848 => x"3880538c",
         11849 => x"3dfc0552",
         11850 => x"8d3d8405",
         11851 => x"51c68c3f",
         11852 => x"84bb8408",
         11853 => x"5584bb84",
         11854 => x"08802e8f",
         11855 => x"3880760c",
         11856 => x"74547384",
         11857 => x"bb840c8c",
         11858 => x"3d0d047a",
         11859 => x"760c7d52",
         11860 => x"7551ffba",
         11861 => x"883f84bb",
         11862 => x"84085584",
         11863 => x"bb840880",
         11864 => x"d138ab16",
         11865 => x"3370982b",
         11866 => x"59598078",
         11867 => x"24af3886",
         11868 => x"16337084",
         11869 => x"2a81065b",
         11870 => x"5479802e",
         11871 => x"80c5389c",
         11872 => x"16089b11",
         11873 => x"339a1233",
         11874 => x"71882b07",
         11875 => x"7d70335d",
         11876 => x"5d5a5557",
         11877 => x"78832eb3",
         11878 => x"38778817",
         11879 => x"0c7a5886",
         11880 => x"18228417",
         11881 => x"23745275",
         11882 => x"51ff9aaa",
         11883 => x"3f84bb84",
         11884 => x"08557484",
         11885 => x"2e8d3874",
         11886 => x"802eff84",
         11887 => x"3880760c",
         11888 => x"fefe3985",
         11889 => x"5580760c",
         11890 => x"fef63995",
         11891 => x"17339418",
         11892 => x"3371982b",
         11893 => x"71902b07",
         11894 => x"7a078819",
         11895 => x"0c5a5aff",
         11896 => x"bc39fa3d",
         11897 => x"0d785589",
         11898 => x"5474802e",
         11899 => x"9e387408",
         11900 => x"5372802e",
         11901 => x"96387233",
         11902 => x"5271802e",
         11903 => x"8e388613",
         11904 => x"22841622",
         11905 => x"57527176",
         11906 => x"2e943880",
         11907 => x"52715773",
         11908 => x"84387375",
         11909 => x"0c7384bb",
         11910 => x"840c883d",
         11911 => x"0d048113",
         11912 => x"3351ff80",
         11913 => x"b43f84bb",
         11914 => x"84088106",
         11915 => x"5271dc38",
         11916 => x"71750853",
         11917 => x"54d739f8",
         11918 => x"3d0d7a7c",
         11919 => x"58558956",
         11920 => x"74802e9f",
         11921 => x"38740854",
         11922 => x"73802e97",
         11923 => x"38733353",
         11924 => x"72802e8f",
         11925 => x"38861422",
         11926 => x"84162259",
         11927 => x"5372782e",
         11928 => x"81973880",
         11929 => x"53725975",
         11930 => x"537580c7",
         11931 => x"3876802e",
         11932 => x"80f33875",
         11933 => x"527451ff",
         11934 => x"9eae3f84",
         11935 => x"bb840853",
         11936 => x"84bb8408",
         11937 => x"842eb538",
         11938 => x"84bb8408",
         11939 => x"a6387652",
         11940 => x"7451ffb3",
         11941 => x"833f7252",
         11942 => x"7451ff9a",
         11943 => x"af3f84bb",
         11944 => x"84088432",
         11945 => x"70307072",
         11946 => x"079f2c84",
         11947 => x"bb840806",
         11948 => x"55575472",
         11949 => x"84bb840c",
         11950 => x"8a3d0d04",
         11951 => x"75775375",
         11952 => x"5253ffb2",
         11953 => x"d33f7252",
         11954 => x"7451ff99",
         11955 => x"ff3f84bb",
         11956 => x"84088432",
         11957 => x"70307072",
         11958 => x"079f2c84",
         11959 => x"bb840806",
         11960 => x"555754cf",
         11961 => x"39755274",
         11962 => x"51ff97ea",
         11963 => x"3f84bb84",
         11964 => x"0884bb84",
         11965 => x"0c8a3d0d",
         11966 => x"04811433",
         11967 => x"51fefed9",
         11968 => x"3f84bb84",
         11969 => x"08810653",
         11970 => x"72fed838",
         11971 => x"72750854",
         11972 => x"56fed239",
         11973 => x"ed3d0d66",
         11974 => x"57805389",
         11975 => x"3d705397",
         11976 => x"3d5256c2",
         11977 => x"963f84bb",
         11978 => x"84085584",
         11979 => x"bb840880",
         11980 => x"2e8a3874",
         11981 => x"84bb840c",
         11982 => x"953d0d04",
         11983 => x"65527551",
         11984 => x"ffb69a3f",
         11985 => x"84bb8408",
         11986 => x"5584bb84",
         11987 => x"08e53802",
         11988 => x"80cb0533",
         11989 => x"70982b55",
         11990 => x"58807424",
         11991 => x"97387680",
         11992 => x"2ed13876",
         11993 => x"527551ff",
         11994 => x"b1ae3f74",
         11995 => x"84bb840c",
         11996 => x"953d0d04",
         11997 => x"860b84bb",
         11998 => x"840c953d",
         11999 => x"0d04ed3d",
         12000 => x"0d666856",
         12001 => x"5f805395",
         12002 => x"3dec0552",
         12003 => x"963d51c1",
         12004 => x"aa3f84bb",
         12005 => x"84085a84",
         12006 => x"bb84089a",
         12007 => x"387f750c",
         12008 => x"74089c11",
         12009 => x"08fe1194",
         12010 => x"13085957",
         12011 => x"59577575",
         12012 => x"268d3875",
         12013 => x"7f0c7984",
         12014 => x"bb840c95",
         12015 => x"3d0d0484",
         12016 => x"bb840877",
         12017 => x"335a5b78",
         12018 => x"812e8293",
         12019 => x"3877a818",
         12020 => x"0884bb84",
         12021 => x"085a5d59",
         12022 => x"7780c138",
         12023 => x"7b811d71",
         12024 => x"5c5d56b4",
         12025 => x"1708762e",
         12026 => x"82ef3883",
         12027 => x"1733785f",
         12028 => x"5d7c818d",
         12029 => x"38815475",
         12030 => x"53b81752",
         12031 => x"81173351",
         12032 => x"fefda83f",
         12033 => x"84bb8408",
         12034 => x"802e8538",
         12035 => x"ff5a815e",
         12036 => x"79b4180c",
         12037 => x"7f7e5b57",
         12038 => x"7d80cc38",
         12039 => x"76335e7d",
         12040 => x"822e828d",
         12041 => x"387717b8",
         12042 => x"05831133",
         12043 => x"82123371",
         12044 => x"902b7188",
         12045 => x"2b078114",
         12046 => x"33707207",
         12047 => x"882b7533",
         12048 => x"7180ffff",
         12049 => x"fe800607",
         12050 => x"70307080",
         12051 => x"25630560",
         12052 => x"840583ff",
         12053 => x"0662ff05",
         12054 => x"43414353",
         12055 => x"54525358",
         12056 => x"405e5678",
         12057 => x"fef2387a",
         12058 => x"7f0c7a94",
         12059 => x"180c8417",
         12060 => x"33810758",
         12061 => x"77841834",
         12062 => x"7984bb84",
         12063 => x"0c953d0d",
         12064 => x"048154b4",
         12065 => x"170853b8",
         12066 => x"17705381",
         12067 => x"1833525d",
         12068 => x"fefd973f",
         12069 => x"815e84bb",
         12070 => x"8408fef8",
         12071 => x"3884bb84",
         12072 => x"08831834",
         12073 => x"b41708a8",
         12074 => x"18083184",
         12075 => x"bb84085f",
         12076 => x"5574a018",
         12077 => x"0827febd",
         12078 => x"38821733",
         12079 => x"5574822e",
         12080 => x"098106fe",
         12081 => x"b0388154",
         12082 => x"b41708a0",
         12083 => x"18080553",
         12084 => x"7c528117",
         12085 => x"3351fefc",
         12086 => x"d13f775e",
         12087 => x"fe973982",
         12088 => x"7742923d",
         12089 => x"59567552",
         12090 => x"7751ff81",
         12091 => x"f13f84bb",
         12092 => x"8408ff2e",
         12093 => x"80e83884",
         12094 => x"bb840881",
         12095 => x"2e80f738",
         12096 => x"84bb8408",
         12097 => x"307084bb",
         12098 => x"84080780",
         12099 => x"257c0581",
         12100 => x"18625a58",
         12101 => x"5c5c9c17",
         12102 => x"087626ca",
         12103 => x"387a7f0c",
         12104 => x"7a94180c",
         12105 => x"84173381",
         12106 => x"07587784",
         12107 => x"1834fec8",
         12108 => x"397717b8",
         12109 => x"05811133",
         12110 => x"71337188",
         12111 => x"2b077030",
         12112 => x"7080251f",
         12113 => x"821d83ff",
         12114 => x"06ff1f5f",
         12115 => x"5d5f595f",
         12116 => x"5f5578fd",
         12117 => x"8338fe8f",
         12118 => x"39775afd",
         12119 => x"bf398160",
         12120 => x"585a7a7f",
         12121 => x"0c7a9418",
         12122 => x"0c841733",
         12123 => x"81075877",
         12124 => x"841834fe",
         12125 => x"83398260",
         12126 => x"585ae739",
         12127 => x"f63d0d7c",
         12128 => x"58895777",
         12129 => x"802e9f38",
         12130 => x"77085675",
         12131 => x"802e9738",
         12132 => x"75335574",
         12133 => x"802e8f38",
         12134 => x"86162284",
         12135 => x"19225a5a",
         12136 => x"79792e82",
         12137 => x"81388055",
         12138 => x"745b7681",
         12139 => x"83389118",
         12140 => x"33577680",
         12141 => x"fb389018",
         12142 => x"3370812a",
         12143 => x"81065659",
         12144 => x"87567480",
         12145 => x"2e80eb38",
         12146 => x"94180855",
         12147 => x"748c1908",
         12148 => x"2780dd38",
         12149 => x"7481fb38",
         12150 => x"88180878",
         12151 => x"08585581",
         12152 => x"75278938",
         12153 => x"9c170875",
         12154 => x"2680d838",
         12155 => x"8257800b",
         12156 => x"88190c94",
         12157 => x"18088c19",
         12158 => x"0c7880c0",
         12159 => x"07557490",
         12160 => x"193476a8",
         12161 => x"3874982b",
         12162 => x"5a798025",
         12163 => x"a3388154",
         12164 => x"9c180853",
         12165 => x"a818527a",
         12166 => x"81113352",
         12167 => x"59fefa8a",
         12168 => x"3f84bb84",
         12169 => x"08802e83",
         12170 => x"90388157",
         12171 => x"76911934",
         12172 => x"76567584",
         12173 => x"bb840c8c",
         12174 => x"3d0d0479",
         12175 => x"55797927",
         12176 => x"80ff3874",
         12177 => x"527751fe",
         12178 => x"ff943f84",
         12179 => x"bb84085a",
         12180 => x"84bb8408",
         12181 => x"802e80e9",
         12182 => x"3884bb84",
         12183 => x"08812e82",
         12184 => x"e83884bb",
         12185 => x"8408ff2e",
         12186 => x"82f53880",
         12187 => x"53745276",
         12188 => x"51ff85cb",
         12189 => x"3f84bb84",
         12190 => x"0882d838",
         12191 => x"9c1708fe",
         12192 => x"11941908",
         12193 => x"58565975",
         12194 => x"7527ffaf",
         12195 => x"38811694",
         12196 => x"180c8417",
         12197 => x"33810755",
         12198 => x"74841834",
         12199 => x"7955787a",
         12200 => x"26ffa038",
         12201 => x"9c398116",
         12202 => x"3351fef7",
         12203 => x"ac3f84bb",
         12204 => x"84088106",
         12205 => x"5574fdee",
         12206 => x"38747808",
         12207 => x"5657fde8",
         12208 => x"39800b90",
         12209 => x"19335a55",
         12210 => x"7457800b",
         12211 => x"88190cfe",
         12212 => x"a2399818",
         12213 => x"08527751",
         12214 => x"fefe833f",
         12215 => x"84bb8408",
         12216 => x"ff2e81c2",
         12217 => x"3884bb84",
         12218 => x"08812e81",
         12219 => x"be387681",
         12220 => x"ae387a59",
         12221 => x"84bb8408",
         12222 => x"9c1a0827",
         12223 => x"81a13884",
         12224 => x"bb840898",
         12225 => x"19087908",
         12226 => x"59575581",
         12227 => x"0b84bb84",
         12228 => x"082781a1",
         12229 => x"3884bb84",
         12230 => x"089c1808",
         12231 => x"27819638",
         12232 => x"75802e97",
         12233 => x"38ff5375",
         12234 => x"527651ff",
         12235 => x"84913f84",
         12236 => x"bb840856",
         12237 => x"84bb8408",
         12238 => x"80e33874",
         12239 => x"527751fe",
         12240 => x"fd9c3f84",
         12241 => x"bb84085a",
         12242 => x"84bb8408",
         12243 => x"802e80cb",
         12244 => x"3884bb84",
         12245 => x"08812e80",
         12246 => x"dc3884bb",
         12247 => x"8408ff2e",
         12248 => x"818f3880",
         12249 => x"53745276",
         12250 => x"51ff83d3",
         12251 => x"3f84bb84",
         12252 => x"0880f638",
         12253 => x"9c1708fe",
         12254 => x"11941908",
         12255 => x"58565975",
         12256 => x"75279038",
         12257 => x"81169418",
         12258 => x"0c841733",
         12259 => x"81075574",
         12260 => x"84183479",
         12261 => x"55787a26",
         12262 => x"ffa13880",
         12263 => x"56755790",
         12264 => x"183359fc",
         12265 => x"ce398157",
         12266 => x"febb3982",
         12267 => x"0b901933",
         12268 => x"5a57fcbf",
         12269 => x"398257e7",
         12270 => x"39901833",
         12271 => x"80ff0655",
         12272 => x"74901934",
         12273 => x"7656fcea",
         12274 => x"39820b90",
         12275 => x"19335a55",
         12276 => x"fdf63984",
         12277 => x"bb840890",
         12278 => x"19335a55",
         12279 => x"fdea3981",
         12280 => x"0b901933",
         12281 => x"5a55fde0",
         12282 => x"3984bb84",
         12283 => x"0857ffaf",
         12284 => x"398157ff",
         12285 => x"aa39db3d",
         12286 => x"0d8253a7",
         12287 => x"3dff9c05",
         12288 => x"52a83d51",
         12289 => x"ffb8b43f",
         12290 => x"84bb8408",
         12291 => x"5684bb84",
         12292 => x"08802e8a",
         12293 => x"387584bb",
         12294 => x"840ca73d",
         12295 => x"0d047d4b",
         12296 => x"a83d0852",
         12297 => x"9b3d7052",
         12298 => x"59ffacb1",
         12299 => x"3f84bb84",
         12300 => x"085684bb",
         12301 => x"8408de38",
         12302 => x"02819305",
         12303 => x"3370852a",
         12304 => x"81065957",
         12305 => x"865677cd",
         12306 => x"3876982b",
         12307 => x"5b807b24",
         12308 => x"c4380280",
         12309 => x"ee053370",
         12310 => x"81065d57",
         12311 => x"87567bff",
         12312 => x"b4387da3",
         12313 => x"3d089b11",
         12314 => x"339a1233",
         12315 => x"71882b07",
         12316 => x"7333415e",
         12317 => x"5c57587c",
         12318 => x"832e80d5",
         12319 => x"3876842a",
         12320 => x"81065776",
         12321 => x"802e80ed",
         12322 => x"38875698",
         12323 => x"18087b2e",
         12324 => x"ff833877",
         12325 => x"5f7a4184",
         12326 => x"bb840852",
         12327 => x"8f3d7052",
         12328 => x"55ff8cb2",
         12329 => x"3f84bb84",
         12330 => x"085684bb",
         12331 => x"8408fee5",
         12332 => x"3884bb84",
         12333 => x"08527451",
         12334 => x"ff91ed3f",
         12335 => x"84bb8408",
         12336 => x"5684bb84",
         12337 => x"08a03887",
         12338 => x"0b84bb84",
         12339 => x"0ca73d0d",
         12340 => x"04951633",
         12341 => x"94173371",
         12342 => x"982b7190",
         12343 => x"2b077d07",
         12344 => x"5d5d5dff",
         12345 => x"983984bb",
         12346 => x"8408842e",
         12347 => x"883884bb",
         12348 => x"8408fea1",
         12349 => x"3878086f",
         12350 => x"a83d0857",
         12351 => x"5d5774ff",
         12352 => x"2e80d338",
         12353 => x"74527851",
         12354 => x"ff8bcb3f",
         12355 => x"84bb8408",
         12356 => x"5684bb84",
         12357 => x"08802ebe",
         12358 => x"38753070",
         12359 => x"77078025",
         12360 => x"565a7a80",
         12361 => x"2e9a3874",
         12362 => x"802e9538",
         12363 => x"7a790858",
         12364 => x"55817b27",
         12365 => x"89389c17",
         12366 => x"087b2681",
         12367 => x"fd388256",
         12368 => x"75fdd238",
         12369 => x"7d51fef6",
         12370 => x"943f84bb",
         12371 => x"840884bb",
         12372 => x"840ca73d",
         12373 => x"0d04b817",
         12374 => x"5d981908",
         12375 => x"56805ab4",
         12376 => x"1708762e",
         12377 => x"82b93883",
         12378 => x"17337a59",
         12379 => x"55747a2e",
         12380 => x"09810680",
         12381 => x"dd388154",
         12382 => x"7553b817",
         12383 => x"52811733",
         12384 => x"51fef2a7",
         12385 => x"3f84bb84",
         12386 => x"08802e85",
         12387 => x"38ff5681",
         12388 => x"5875b418",
         12389 => x"0c775677",
         12390 => x"ab389c19",
         12391 => x"0858e578",
         12392 => x"34810b83",
         12393 => x"18349019",
         12394 => x"087c27fe",
         12395 => x"ec388052",
         12396 => x"7851ff8c",
         12397 => x"973f84bb",
         12398 => x"84085684",
         12399 => x"bb840880",
         12400 => x"2eff9638",
         12401 => x"75842e09",
         12402 => x"8106fecd",
         12403 => x"388256fe",
         12404 => x"c8398154",
         12405 => x"b4170853",
         12406 => x"7c528117",
         12407 => x"3351fef2",
         12408 => x"c93f8158",
         12409 => x"84bb8408",
         12410 => x"7a2e0981",
         12411 => x"06ffa638",
         12412 => x"84bb8408",
         12413 => x"831834b4",
         12414 => x"1708a818",
         12415 => x"083184bb",
         12416 => x"84085955",
         12417 => x"74a01808",
         12418 => x"27feeb38",
         12419 => x"82173355",
         12420 => x"74822e09",
         12421 => x"8106fede",
         12422 => x"388154b4",
         12423 => x"1708a018",
         12424 => x"0805537c",
         12425 => x"52811733",
         12426 => x"51fef1fe",
         12427 => x"3f7958fe",
         12428 => x"c5397955",
         12429 => x"79782780",
         12430 => x"e1387452",
         12431 => x"7851fef7",
         12432 => x"9d3f84bb",
         12433 => x"84085a84",
         12434 => x"bb840880",
         12435 => x"2e80cb38",
         12436 => x"84bb8408",
         12437 => x"812efde6",
         12438 => x"3884bb84",
         12439 => x"08ff2e80",
         12440 => x"cb388053",
         12441 => x"74527651",
         12442 => x"fefdd43f",
         12443 => x"84bb8408",
         12444 => x"b3389c17",
         12445 => x"08fe1194",
         12446 => x"1908585c",
         12447 => x"58757b27",
         12448 => x"ffb03881",
         12449 => x"1694180c",
         12450 => x"84173381",
         12451 => x"075c7b84",
         12452 => x"18347955",
         12453 => x"777a26ff",
         12454 => x"a1388056",
         12455 => x"fda23979",
         12456 => x"56fdf739",
         12457 => x"84bb8408",
         12458 => x"56fd9539",
         12459 => x"8156fd90",
         12460 => x"39e33d0d",
         12461 => x"82539f3d",
         12462 => x"ffbc0552",
         12463 => x"a03d51ff",
         12464 => x"b2f93f84",
         12465 => x"bb840856",
         12466 => x"84bb8408",
         12467 => x"802e8a38",
         12468 => x"7584bb84",
         12469 => x"0c9f3d0d",
         12470 => x"047d436f",
         12471 => x"52933d70",
         12472 => x"525affa6",
         12473 => x"f83f84bb",
         12474 => x"84085684",
         12475 => x"bb84088b",
         12476 => x"38880b84",
         12477 => x"bb840c9f",
         12478 => x"3d0d0484",
         12479 => x"bb840884",
         12480 => x"2e098106",
         12481 => x"cb380280",
         12482 => x"f3053370",
         12483 => x"852a8106",
         12484 => x"56588656",
         12485 => x"74ffb938",
         12486 => x"7d5f7452",
         12487 => x"8f3d7052",
         12488 => x"5dff83f9",
         12489 => x"3f84bb84",
         12490 => x"0875575c",
         12491 => x"84bb8408",
         12492 => x"83388756",
         12493 => x"84bb8408",
         12494 => x"812e80f9",
         12495 => x"3884bb84",
         12496 => x"08ff2e81",
         12497 => x"cb387581",
         12498 => x"c9387d84",
         12499 => x"bb840883",
         12500 => x"12335d5a",
         12501 => x"577a80e2",
         12502 => x"38fe199c",
         12503 => x"1808fe05",
         12504 => x"5a56805b",
         12505 => x"7579278d",
         12506 => x"388a1722",
         12507 => x"767129b0",
         12508 => x"1908055c",
         12509 => x"587ab418",
         12510 => x"0cb81759",
         12511 => x"84807957",
         12512 => x"55807670",
         12513 => x"81055834",
         12514 => x"ff155574",
         12515 => x"f4387458",
         12516 => x"8a172255",
         12517 => x"77752781",
         12518 => x"f9388154",
         12519 => x"771b5378",
         12520 => x"52811733",
         12521 => x"51feef82",
         12522 => x"3f84bb84",
         12523 => x"0881df38",
         12524 => x"811858dc",
         12525 => x"398256ff",
         12526 => x"84398154",
         12527 => x"b4170853",
         12528 => x"b8177053",
         12529 => x"81183352",
         12530 => x"58feeede",
         12531 => x"3f815684",
         12532 => x"bb8408be",
         12533 => x"3884bb84",
         12534 => x"08831834",
         12535 => x"b41708a8",
         12536 => x"18083155",
         12537 => x"74a01808",
         12538 => x"27feee38",
         12539 => x"8217335b",
         12540 => x"7a822e09",
         12541 => x"8106fee1",
         12542 => x"387554b4",
         12543 => x"1708a018",
         12544 => x"08055377",
         12545 => x"52811733",
         12546 => x"51feee9e",
         12547 => x"3ffeca39",
         12548 => x"81567b7d",
         12549 => x"08585581",
         12550 => x"7c27fdb4",
         12551 => x"387b9c18",
         12552 => x"0827fdac",
         12553 => x"3874527c",
         12554 => x"51fef3b2",
         12555 => x"3f84bb84",
         12556 => x"085a84bb",
         12557 => x"8408802e",
         12558 => x"fd963884",
         12559 => x"bb840881",
         12560 => x"2efd8d38",
         12561 => x"84bb8408",
         12562 => x"ff2efd84",
         12563 => x"38805374",
         12564 => x"527651fe",
         12565 => x"f9e93f84",
         12566 => x"bb8408fc",
         12567 => x"f3389c17",
         12568 => x"08fe1194",
         12569 => x"19085a5c",
         12570 => x"59777b27",
         12571 => x"90388118",
         12572 => x"94180c84",
         12573 => x"17338107",
         12574 => x"5c7b8418",
         12575 => x"34795578",
         12576 => x"7a26ffa1",
         12577 => x"387584bb",
         12578 => x"840c9f3d",
         12579 => x"0d048a17",
         12580 => x"22557483",
         12581 => x"ffff0657",
         12582 => x"81567678",
         12583 => x"2e098106",
         12584 => x"fef0388b",
         12585 => x"0bb81f56",
         12586 => x"56a07570",
         12587 => x"81055734",
         12588 => x"ff165675",
         12589 => x"f4387d57",
         12590 => x"ae0bb818",
         12591 => x"347d5890",
         12592 => x"0b80c319",
         12593 => x"347d5975",
         12594 => x"80ce1a34",
         12595 => x"7580cf1a",
         12596 => x"34a10b80",
         12597 => x"d01a3480",
         12598 => x"cc0b80d1",
         12599 => x"1a347d7c",
         12600 => x"83ffff06",
         12601 => x"59567780",
         12602 => x"d2173477",
         12603 => x"882a5b7a",
         12604 => x"80d31734",
         12605 => x"75335574",
         12606 => x"832e81cc",
         12607 => x"387d59a0",
         12608 => x"0b80d81a",
         12609 => x"b81b5758",
         12610 => x"56747081",
         12611 => x"05563377",
         12612 => x"70810559",
         12613 => x"34ff1656",
         12614 => x"75ef387d",
         12615 => x"56ae0b80",
         12616 => x"d9173464",
         12617 => x"7e7183ff",
         12618 => x"ff065b57",
         12619 => x"577880f2",
         12620 => x"17347888",
         12621 => x"2a5b7a80",
         12622 => x"f3173475",
         12623 => x"33557483",
         12624 => x"2e80f038",
         12625 => x"7d5b810b",
         12626 => x"831c3479",
         12627 => x"51ff92cf",
         12628 => x"3f84bb84",
         12629 => x"085684bb",
         12630 => x"8408fdb6",
         12631 => x"38695684",
         12632 => x"bb840896",
         12633 => x"173484bb",
         12634 => x"84089717",
         12635 => x"34a10b98",
         12636 => x"173480cc",
         12637 => x"0b991734",
         12638 => x"7d6a585d",
         12639 => x"779a1834",
         12640 => x"77882a59",
         12641 => x"789b1834",
         12642 => x"7c335a79",
         12643 => x"832e80d9",
         12644 => x"38695590",
         12645 => x"0b8b1634",
         12646 => x"7d57810b",
         12647 => x"8318347d",
         12648 => x"51feedb9",
         12649 => x"3f84bb84",
         12650 => x"08567584",
         12651 => x"bb840c9f",
         12652 => x"3d0d0476",
         12653 => x"902a5574",
         12654 => x"80ec1734",
         12655 => x"74882a57",
         12656 => x"7680ed17",
         12657 => x"34fefd39",
         12658 => x"7b902a5b",
         12659 => x"7a80cc17",
         12660 => x"347a882a",
         12661 => x"557480cd",
         12662 => x"17347d59",
         12663 => x"a00b80d8",
         12664 => x"1ab81b57",
         12665 => x"5856fea1",
         12666 => x"397b902a",
         12667 => x"58779418",
         12668 => x"3477882a",
         12669 => x"5c7b9518",
         12670 => x"34695590",
         12671 => x"0b8b1634",
         12672 => x"7d57810b",
         12673 => x"8318347d",
         12674 => x"51feecd1",
         12675 => x"3f84bb84",
         12676 => x"0856ff96",
         12677 => x"39d13d0d",
         12678 => x"b33db43d",
         12679 => x"0870595b",
         12680 => x"5f79802e",
         12681 => x"9b387970",
         12682 => x"81055b33",
         12683 => x"709f2656",
         12684 => x"5675ba2e",
         12685 => x"81b83874",
         12686 => x"ed3875ba",
         12687 => x"2e81af38",
         12688 => x"8253b13d",
         12689 => x"fefc0552",
         12690 => x"b23d51ff",
         12691 => x"abed3f84",
         12692 => x"bb840856",
         12693 => x"84bb8408",
         12694 => x"802e8a38",
         12695 => x"7584bb84",
         12696 => x"0cb13d0d",
         12697 => x"047fa63d",
         12698 => x"0cb23d08",
         12699 => x"52a53d70",
         12700 => x"5259ff9f",
         12701 => x"e83f84bb",
         12702 => x"84085684",
         12703 => x"bb8408dc",
         12704 => x"380281bb",
         12705 => x"053381a0",
         12706 => x"065d8656",
         12707 => x"7cce38a0",
         12708 => x"0b923dae",
         12709 => x"3d085858",
         12710 => x"55757081",
         12711 => x"05573377",
         12712 => x"70810559",
         12713 => x"34ff1555",
         12714 => x"74ef3899",
         12715 => x"3d58b078",
         12716 => x"7a585855",
         12717 => x"75708105",
         12718 => x"57337770",
         12719 => x"81055934",
         12720 => x"ff155574",
         12721 => x"ef38b33d",
         12722 => x"08527751",
         12723 => x"ff9f8e3f",
         12724 => x"84bb8408",
         12725 => x"5684bb84",
         12726 => x"0885d838",
         12727 => x"6aa83d08",
         12728 => x"2e81cb38",
         12729 => x"880b84bb",
         12730 => x"840cb13d",
         12731 => x"0d047633",
         12732 => x"d0117081",
         12733 => x"ff065757",
         12734 => x"58748926",
         12735 => x"91388217",
         12736 => x"7881ff06",
         12737 => x"d0055d59",
         12738 => x"787a2e80",
         12739 => x"fa38807f",
         12740 => x"0883e6f4",
         12741 => x"7008725d",
         12742 => x"5e5f5f5c",
         12743 => x"7a708105",
         12744 => x"5c337970",
         12745 => x"81055b33",
         12746 => x"ff9f125a",
         12747 => x"58567799",
         12748 => x"268938e0",
         12749 => x"167081ff",
         12750 => x"065755ff",
         12751 => x"9f175877",
         12752 => x"99268938",
         12753 => x"e0177081",
         12754 => x"ff065855",
         12755 => x"7530709f",
         12756 => x"2a595575",
         12757 => x"772e0981",
         12758 => x"06853877",
         12759 => x"ffbe3878",
         12760 => x"7a327030",
         12761 => x"7072079f",
         12762 => x"2a7a075d",
         12763 => x"58557a80",
         12764 => x"2e953881",
         12765 => x"1c841e5e",
         12766 => x"5c7b8324",
         12767 => x"fdc2387c",
         12768 => x"087e5a5b",
         12769 => x"ff96397b",
         12770 => x"8324fdb4",
         12771 => x"38797f0c",
         12772 => x"8253b13d",
         12773 => x"fefc0552",
         12774 => x"b23d51ff",
         12775 => x"a99d3f84",
         12776 => x"bb840856",
         12777 => x"84bb8408",
         12778 => x"fdb238fd",
         12779 => x"b8396caa",
         12780 => x"3d082e09",
         12781 => x"8106feac",
         12782 => x"387751ff",
         12783 => x"8de13f84",
         12784 => x"bb840856",
         12785 => x"84bb8408",
         12786 => x"fd92386f",
         12787 => x"58930b8d",
         12788 => x"19028805",
         12789 => x"80cd0558",
         12790 => x"565a7570",
         12791 => x"81055733",
         12792 => x"75708105",
         12793 => x"5734ff1a",
         12794 => x"5a79ef38",
         12795 => x"0280cb05",
         12796 => x"338b1934",
         12797 => x"8b183370",
         12798 => x"842a8106",
         12799 => x"40567e89",
         12800 => x"3875a007",
         12801 => x"57768b19",
         12802 => x"347f5d81",
         12803 => x"0b831e34",
         12804 => x"8b183370",
         12805 => x"842a8106",
         12806 => x"575c7580",
         12807 => x"2e81c538",
         12808 => x"a73d086b",
         12809 => x"2e81bd38",
         12810 => x"7f9b1933",
         12811 => x"9a1a3371",
         12812 => x"882b0772",
         12813 => x"3341585c",
         12814 => x"577d832e",
         12815 => x"82e038fe",
         12816 => x"169c1808",
         12817 => x"fe055e56",
         12818 => x"757d2782",
         12819 => x"c7388a17",
         12820 => x"22767129",
         12821 => x"b0190805",
         12822 => x"575e7580",
         12823 => x"2e82b538",
         12824 => x"757a5d58",
         12825 => x"b4170876",
         12826 => x"2eaa3883",
         12827 => x"17335f7e",
         12828 => x"83bc3881",
         12829 => x"547553b8",
         12830 => x"17528117",
         12831 => x"3351fee4",
         12832 => x"aa3f84bb",
         12833 => x"8408802e",
         12834 => x"8538ff58",
         12835 => x"815c77b4",
         12836 => x"180c7f57",
         12837 => x"7b80d818",
         12838 => x"56567bfb",
         12839 => x"bf388115",
         12840 => x"335a79ae",
         12841 => x"2e098106",
         12842 => x"bb386a70",
         12843 => x"83ffff06",
         12844 => x"5d567b80",
         12845 => x"f218347b",
         12846 => x"882a5877",
         12847 => x"80f31834",
         12848 => x"76335b7a",
         12849 => x"832e0981",
         12850 => x"06933875",
         12851 => x"902a5e7d",
         12852 => x"80ec1834",
         12853 => x"7d882a56",
         12854 => x"7580ed18",
         12855 => x"347f5781",
         12856 => x"0b831834",
         12857 => x"7808aa3d",
         12858 => x"08b23d08",
         12859 => x"575c5674",
         12860 => x"ff2e9538",
         12861 => x"74527851",
         12862 => x"fefbdb3f",
         12863 => x"84bb8408",
         12864 => x"5584bb84",
         12865 => x"0880f538",
         12866 => x"b8165c98",
         12867 => x"19085780",
         12868 => x"5ab41608",
         12869 => x"772eb438",
         12870 => x"8316337a",
         12871 => x"595f7e7a",
         12872 => x"2e098106",
         12873 => x"81a83881",
         12874 => x"547653b8",
         12875 => x"16528116",
         12876 => x"3351fee2",
         12877 => x"f63f84bb",
         12878 => x"8408802e",
         12879 => x"8538ff57",
         12880 => x"815876b4",
         12881 => x"170c7755",
         12882 => x"77aa389c",
         12883 => x"19085ae5",
         12884 => x"7a34810b",
         12885 => x"83173490",
         12886 => x"19087b27",
         12887 => x"a5388052",
         12888 => x"7851fefc",
         12889 => x"e73f84bb",
         12890 => x"84085584",
         12891 => x"bb840880",
         12892 => x"2eff9838",
         12893 => x"82567484",
         12894 => x"2ef9e138",
         12895 => x"745674f9",
         12896 => x"db387f51",
         12897 => x"fee5d63f",
         12898 => x"84bb8408",
         12899 => x"84bb840c",
         12900 => x"b13d0d04",
         12901 => x"820b84bb",
         12902 => x"840cb13d",
         12903 => x"0d049518",
         12904 => x"33941933",
         12905 => x"71982b71",
         12906 => x"902b0778",
         12907 => x"0758565c",
         12908 => x"fd8d3984",
         12909 => x"bb840884",
         12910 => x"2efbfe38",
         12911 => x"84bb8408",
         12912 => x"802efea0",
         12913 => x"387584bb",
         12914 => x"840cb13d",
         12915 => x"0d048154",
         12916 => x"b4160853",
         12917 => x"7b528116",
         12918 => x"3351fee2",
         12919 => x"cd3f8158",
         12920 => x"84bb8408",
         12921 => x"7a2e0981",
         12922 => x"06fedb38",
         12923 => x"84bb8408",
         12924 => x"831734b4",
         12925 => x"1608a817",
         12926 => x"083184bb",
         12927 => x"84085955",
         12928 => x"74a01708",
         12929 => x"27fea038",
         12930 => x"8216335d",
         12931 => x"7c822e09",
         12932 => x"8106fe93",
         12933 => x"388154b4",
         12934 => x"1608a017",
         12935 => x"0805537b",
         12936 => x"52811633",
         12937 => x"51fee282",
         12938 => x"3f7958fd",
         12939 => x"fa398154",
         12940 => x"b4170853",
         12941 => x"b8177053",
         12942 => x"81183352",
         12943 => x"5bfee1ea",
         12944 => x"3f815c84",
         12945 => x"bb8408fc",
         12946 => x"c93884bb",
         12947 => x"84088318",
         12948 => x"34b41708",
         12949 => x"a8180831",
         12950 => x"84bb8408",
         12951 => x"5d5574a0",
         12952 => x"180827fc",
         12953 => x"8e388217",
         12954 => x"335d7c82",
         12955 => x"2e098106",
         12956 => x"fc813881",
         12957 => x"54b41708",
         12958 => x"a0180805",
         12959 => x"537a5281",
         12960 => x"173351fe",
         12961 => x"e1a43f79",
         12962 => x"5cfbe839",
         12963 => x"ec3d0d02",
         12964 => x"80df0533",
         12965 => x"02840580",
         12966 => x"e3053356",
         12967 => x"57825396",
         12968 => x"3dcc0552",
         12969 => x"973d51ff",
         12970 => x"a3913f84",
         12971 => x"bb840856",
         12972 => x"84bb8408",
         12973 => x"802e8a38",
         12974 => x"7584bb84",
         12975 => x"0c963d0d",
         12976 => x"04785a66",
         12977 => x"52963dd0",
         12978 => x"0551ff97",
         12979 => x"903f84bb",
         12980 => x"84085684",
         12981 => x"bb8408e0",
         12982 => x"380280cf",
         12983 => x"053381a0",
         12984 => x"06548656",
         12985 => x"73d23874",
         12986 => x"a7066171",
         12987 => x"098b1233",
         12988 => x"71067a74",
         12989 => x"06075156",
         12990 => x"5755738b",
         12991 => x"17347855",
         12992 => x"810b8316",
         12993 => x"347851fe",
         12994 => x"e2d33f84",
         12995 => x"bb840884",
         12996 => x"bb840c96",
         12997 => x"3d0d04ec",
         12998 => x"3d0d6757",
         12999 => x"8253963d",
         13000 => x"cc055297",
         13001 => x"3d51ffa2",
         13002 => x"923f84bb",
         13003 => x"84085584",
         13004 => x"bb840880",
         13005 => x"2e8a3874",
         13006 => x"84bb840c",
         13007 => x"963d0d04",
         13008 => x"785a6652",
         13009 => x"963dd005",
         13010 => x"51ff9691",
         13011 => x"3f84bb84",
         13012 => x"085584bb",
         13013 => x"8408e038",
         13014 => x"0280cf05",
         13015 => x"3381a006",
         13016 => x"56865575",
         13017 => x"d2386084",
         13018 => x"18228619",
         13019 => x"2271902b",
         13020 => x"07595956",
         13021 => x"76961734",
         13022 => x"76882a55",
         13023 => x"74971734",
         13024 => x"76902a58",
         13025 => x"77981734",
         13026 => x"76982a54",
         13027 => x"73991734",
         13028 => x"7857810b",
         13029 => x"83183478",
         13030 => x"51fee1c1",
         13031 => x"3f84bb84",
         13032 => x"0884bb84",
         13033 => x"0c963d0d",
         13034 => x"04e83d0d",
         13035 => x"6b6d5d5b",
         13036 => x"80539a3d",
         13037 => x"cc05529b",
         13038 => x"3d51ffa0",
         13039 => x"fe3f84bb",
         13040 => x"840884bb",
         13041 => x"84083070",
         13042 => x"84bb8408",
         13043 => x"07802551",
         13044 => x"56577a80",
         13045 => x"2e8b3881",
         13046 => x"7076065a",
         13047 => x"567881a4",
         13048 => x"38763070",
         13049 => x"78078025",
         13050 => x"565b7b80",
         13051 => x"2e818c38",
         13052 => x"81707606",
         13053 => x"5a587880",
         13054 => x"2e818038",
         13055 => x"7ca41108",
         13056 => x"5856805a",
         13057 => x"b4160877",
         13058 => x"2e82f638",
         13059 => x"8316337a",
         13060 => x"5a55747a",
         13061 => x"2e098106",
         13062 => x"81983881",
         13063 => x"547653b8",
         13064 => x"16528116",
         13065 => x"3351fedd",
         13066 => x"823f84bb",
         13067 => x"8408802e",
         13068 => x"8538ff57",
         13069 => x"815976b4",
         13070 => x"170c7857",
         13071 => x"78bd387c",
         13072 => x"70335658",
         13073 => x"80c35674",
         13074 => x"832e8b38",
         13075 => x"80e45674",
         13076 => x"842e8338",
         13077 => x"a7567518",
         13078 => x"b8058311",
         13079 => x"33821233",
         13080 => x"71902b71",
         13081 => x"882b0781",
         13082 => x"14337072",
         13083 => x"07882b75",
         13084 => x"33710762",
         13085 => x"0c5f5d5e",
         13086 => x"57595676",
         13087 => x"84bb840c",
         13088 => x"9a3d0d04",
         13089 => x"7c5e8040",
         13090 => x"80528e3d",
         13091 => x"705255fe",
         13092 => x"f4c43f84",
         13093 => x"bb840857",
         13094 => x"84bb8408",
         13095 => x"802e818d",
         13096 => x"3876842e",
         13097 => x"098106fe",
         13098 => x"b838807b",
         13099 => x"348057fe",
         13100 => x"b0397754",
         13101 => x"b4160853",
         13102 => x"b8167053",
         13103 => x"81173352",
         13104 => x"5bfedce6",
         13105 => x"3f775984",
         13106 => x"bb84087a",
         13107 => x"2e098106",
         13108 => x"fee83884",
         13109 => x"bb840883",
         13110 => x"1734b416",
         13111 => x"08a81708",
         13112 => x"3184bb84",
         13113 => x"085a5574",
         13114 => x"a0170827",
         13115 => x"fead3882",
         13116 => x"16335574",
         13117 => x"822e0981",
         13118 => x"06fea038",
         13119 => x"7754b416",
         13120 => x"08a01708",
         13121 => x"05537a52",
         13122 => x"81163351",
         13123 => x"fedc9b3f",
         13124 => x"79598154",
         13125 => x"7653b816",
         13126 => x"52811633",
         13127 => x"51fedb8b",
         13128 => x"3f84bb84",
         13129 => x"08802efe",
         13130 => x"8d38fe86",
         13131 => x"39755274",
         13132 => x"51fef8f4",
         13133 => x"3f84bb84",
         13134 => x"085784bb",
         13135 => x"8408fee1",
         13136 => x"3884bb84",
         13137 => x"0884bb84",
         13138 => x"08665c59",
         13139 => x"59791881",
         13140 => x"197c1b57",
         13141 => x"59567533",
         13142 => x"75348119",
         13143 => x"598a7827",
         13144 => x"ec388b70",
         13145 => x"1c575880",
         13146 => x"76347780",
         13147 => x"2efcf238",
         13148 => x"ff187b11",
         13149 => x"70335c57",
         13150 => x"5879a02e",
         13151 => x"ea38fce1",
         13152 => x"397957fd",
         13153 => x"ba39e13d",
         13154 => x"0d8253a1",
         13155 => x"3dffb405",
         13156 => x"52a23d51",
         13157 => x"ff9da43f",
         13158 => x"84bb8408",
         13159 => x"5684bb84",
         13160 => x"0882a638",
         13161 => x"8f3d5d8b",
         13162 => x"7d5755a0",
         13163 => x"76708105",
         13164 => x"5834ff15",
         13165 => x"5574f438",
         13166 => x"74a33d08",
         13167 => x"70337081",
         13168 => x"ff065b58",
         13169 => x"585a9f78",
         13170 => x"2781b738",
         13171 => x"a23d903d",
         13172 => x"5c5c7581",
         13173 => x"ff068118",
         13174 => x"57557481",
         13175 => x"f538757c",
         13176 => x"0c7483ff",
         13177 => x"ff2681ff",
         13178 => x"387451a1",
         13179 => x"953f83b5",
         13180 => x"5284bb84",
         13181 => x"08519fdc",
         13182 => x"3f84bb84",
         13183 => x"0883ffff",
         13184 => x"06577680",
         13185 => x"2e81e038",
         13186 => x"83e8940b",
         13187 => x"83e89433",
         13188 => x"7081ff06",
         13189 => x"5b565878",
         13190 => x"802e81d6",
         13191 => x"38745678",
         13192 => x"772e9938",
         13193 => x"81187033",
         13194 => x"7081ff06",
         13195 => x"57575874",
         13196 => x"802e8938",
         13197 => x"74772e09",
         13198 => x"8106e938",
         13199 => x"7581ff06",
         13200 => x"597881a3",
         13201 => x"3881ff77",
         13202 => x"2781f838",
         13203 => x"79892681",
         13204 => x"963881ff",
         13205 => x"77278f38",
         13206 => x"76882a55",
         13207 => x"747b7081",
         13208 => x"055d3481",
         13209 => x"1a5a767b",
         13210 => x"7081055d",
         13211 => x"34811aa3",
         13212 => x"3d087033",
         13213 => x"7081ff06",
         13214 => x"5b58585a",
         13215 => x"779f26fe",
         13216 => x"d1388f3d",
         13217 => x"33578656",
         13218 => x"7681e52e",
         13219 => x"bc387980",
         13220 => x"2e993802",
         13221 => x"b7055679",
         13222 => x"1670335c",
         13223 => x"5c7aa02e",
         13224 => x"09810687",
         13225 => x"38ff1a5a",
         13226 => x"79ed387d",
         13227 => x"45804780",
         13228 => x"52953d70",
         13229 => x"5256fef0",
         13230 => x"9d3f84bb",
         13231 => x"84085584",
         13232 => x"bb840880",
         13233 => x"2eb43874",
         13234 => x"567584bb",
         13235 => x"840ca13d",
         13236 => x"0d0483b5",
         13237 => x"5274519e",
         13238 => x"e73f84bb",
         13239 => x"840883ff",
         13240 => x"ff065574",
         13241 => x"fdf83886",
         13242 => x"567584bb",
         13243 => x"840ca13d",
         13244 => x"0d0483e8",
         13245 => x"943356fe",
         13246 => x"c3398152",
         13247 => x"7551fef5",
         13248 => x"a73f84bb",
         13249 => x"84085584",
         13250 => x"bb840880",
         13251 => x"c1387980",
         13252 => x"2e82c438",
         13253 => x"8b6c7e59",
         13254 => x"57557670",
         13255 => x"81055833",
         13256 => x"76708105",
         13257 => x"5834ff15",
         13258 => x"5574ef38",
         13259 => x"7d5d810b",
         13260 => x"831e347d",
         13261 => x"51fedaa5",
         13262 => x"3f84bb84",
         13263 => x"08557456",
         13264 => x"ff87398a",
         13265 => x"7a27fe8a",
         13266 => x"388656ff",
         13267 => x"9c3984bb",
         13268 => x"8408842e",
         13269 => x"098106fe",
         13270 => x"ee388055",
         13271 => x"79752efe",
         13272 => x"e6387508",
         13273 => x"75537652",
         13274 => x"58feeeea",
         13275 => x"3f84bb84",
         13276 => x"085784bb",
         13277 => x"8408752e",
         13278 => x"09810681",
         13279 => x"843884bb",
         13280 => x"8408b819",
         13281 => x"5c5a9816",
         13282 => x"08578059",
         13283 => x"b4180877",
         13284 => x"2eb23883",
         13285 => x"18335574",
         13286 => x"792e0981",
         13287 => x"0681d738",
         13288 => x"81547653",
         13289 => x"b8185281",
         13290 => x"183351fe",
         13291 => x"d5fd3f84",
         13292 => x"bb840880",
         13293 => x"2e8538ff",
         13294 => x"57815976",
         13295 => x"b4190c78",
         13296 => x"5778be38",
         13297 => x"789c1708",
         13298 => x"7033575a",
         13299 => x"577481e5",
         13300 => x"2e819e38",
         13301 => x"74307080",
         13302 => x"25780756",
         13303 => x"5c74802e",
         13304 => x"81d73881",
         13305 => x"1a5a7981",
         13306 => x"2ea53881",
         13307 => x"527551fe",
         13308 => x"efda3f84",
         13309 => x"bb840857",
         13310 => x"84bb8408",
         13311 => x"802eff86",
         13312 => x"38875576",
         13313 => x"842efdbf",
         13314 => x"38765576",
         13315 => x"fdb938a0",
         13316 => x"6c575580",
         13317 => x"76708105",
         13318 => x"5834ff15",
         13319 => x"5574f438",
         13320 => x"6b56880b",
         13321 => x"8b17348b",
         13322 => x"6c7e5957",
         13323 => x"55767081",
         13324 => x"05583376",
         13325 => x"70810558",
         13326 => x"34ff1555",
         13327 => x"74802efd",
         13328 => x"eb387670",
         13329 => x"81055833",
         13330 => x"76708105",
         13331 => x"5834ff15",
         13332 => x"5574da38",
         13333 => x"fdd6396b",
         13334 => x"5ae57a34",
         13335 => x"7d5d810b",
         13336 => x"831e347d",
         13337 => x"51fed7f5",
         13338 => x"3f84bb84",
         13339 => x"0855fdce",
         13340 => x"398157fe",
         13341 => x"df398154",
         13342 => x"b4180853",
         13343 => x"7a528118",
         13344 => x"3351fed5",
         13345 => x"a53f84bb",
         13346 => x"8408792e",
         13347 => x"09810680",
         13348 => x"c33884bb",
         13349 => x"84088319",
         13350 => x"34b41808",
         13351 => x"a8190831",
         13352 => x"5c7ba019",
         13353 => x"08278a38",
         13354 => x"82183355",
         13355 => x"74822eb1",
         13356 => x"3884bb84",
         13357 => x"0859fde8",
         13358 => x"39745a81",
         13359 => x"527551fe",
         13360 => x"ee8a3f84",
         13361 => x"bb840857",
         13362 => x"84bb8408",
         13363 => x"802efdb6",
         13364 => x"38feae39",
         13365 => x"81705859",
         13366 => x"78802efd",
         13367 => x"e738fea1",
         13368 => x"398154b4",
         13369 => x"1808a019",
         13370 => x"0805537a",
         13371 => x"52811833",
         13372 => x"51fed4b6",
         13373 => x"3ffda939",
         13374 => x"f23d0d60",
         13375 => x"62028805",
         13376 => x"80cb0533",
         13377 => x"5e5b5789",
         13378 => x"5676802e",
         13379 => x"9f387608",
         13380 => x"5574802e",
         13381 => x"97387433",
         13382 => x"5473802e",
         13383 => x"8f388615",
         13384 => x"22841822",
         13385 => x"59597878",
         13386 => x"2e81c238",
         13387 => x"8054735f",
         13388 => x"7581a538",
         13389 => x"91173356",
         13390 => x"75819d38",
         13391 => x"79802e81",
         13392 => x"a2388c17",
         13393 => x"08819c38",
         13394 => x"90173370",
         13395 => x"812a8106",
         13396 => x"565d7480",
         13397 => x"2e818c38",
         13398 => x"7e8a1122",
         13399 => x"70892b70",
         13400 => x"557c5457",
         13401 => x"5c59fd86",
         13402 => x"bc3fff15",
         13403 => x"7a067030",
         13404 => x"7072079f",
         13405 => x"2a84bb84",
         13406 => x"0805901c",
         13407 => x"08794253",
         13408 => x"5f555881",
         13409 => x"78278838",
         13410 => x"9c190878",
         13411 => x"26833882",
         13412 => x"58777856",
         13413 => x"5b805974",
         13414 => x"527651fe",
         13415 => x"d8c03f81",
         13416 => x"157f5555",
         13417 => x"9c140875",
         13418 => x"26833882",
         13419 => x"5584bb84",
         13420 => x"08812e81",
         13421 => x"dc3884bb",
         13422 => x"8408ff2e",
         13423 => x"81d83884",
         13424 => x"bb840881",
         13425 => x"c5388119",
         13426 => x"59787d2e",
         13427 => x"bb387478",
         13428 => x"2e098106",
         13429 => x"c2388756",
         13430 => x"75547384",
         13431 => x"bb840c90",
         13432 => x"3d0d0487",
         13433 => x"0b84bb84",
         13434 => x"0c903d0d",
         13435 => x"04811533",
         13436 => x"51fed0e5",
         13437 => x"3f84bb84",
         13438 => x"08810654",
         13439 => x"73fead38",
         13440 => x"73770855",
         13441 => x"56fea739",
         13442 => x"7b802e81",
         13443 => x"8e387a7d",
         13444 => x"56587c80",
         13445 => x"2eab3881",
         13446 => x"18547481",
         13447 => x"2e80e638",
         13448 => x"73537752",
         13449 => x"7e51fede",
         13450 => x"963f84bb",
         13451 => x"84085684",
         13452 => x"bb8408ff",
         13453 => x"a3387781",
         13454 => x"19ff1757",
         13455 => x"595e74d7",
         13456 => x"387e7e90",
         13457 => x"120c557b",
         13458 => x"802eff8c",
         13459 => x"387a8818",
         13460 => x"0c798c18",
         13461 => x"0c901733",
         13462 => x"80c0075c",
         13463 => x"7b901834",
         13464 => x"9c1508fe",
         13465 => x"05941608",
         13466 => x"585a767a",
         13467 => x"26fee938",
         13468 => x"767d3194",
         13469 => x"160c8415",
         13470 => x"3381075d",
         13471 => x"7c841634",
         13472 => x"7554fed6",
         13473 => x"39ff54ff",
         13474 => x"9739745b",
         13475 => x"8059febe",
         13476 => x"398254fe",
         13477 => x"c5398154",
         13478 => x"fec039ff",
         13479 => x"1b5effa1",
         13480 => x"3984bb90",
         13481 => x"08e33d0d",
         13482 => x"a33d08a5",
         13483 => x"3d080288",
         13484 => x"05818705",
         13485 => x"3344425f",
         13486 => x"ff0ba23d",
         13487 => x"08705f5b",
         13488 => x"4079802e",
         13489 => x"858a3879",
         13490 => x"7081055b",
         13491 => x"33709f26",
         13492 => x"565675ba",
         13493 => x"2e859b38",
         13494 => x"74ed3875",
         13495 => x"ba2e8592",
         13496 => x"3884e2e0",
         13497 => x"33568076",
         13498 => x"2484e538",
         13499 => x"75101084",
         13500 => x"e2cc0570",
         13501 => x"08565a74",
         13502 => x"802e8438",
         13503 => x"80753475",
         13504 => x"1684baf8",
         13505 => x"113384ba",
         13506 => x"f9123340",
         13507 => x"5b5d8152",
         13508 => x"7951fece",
         13509 => x"e23f84bb",
         13510 => x"840881ff",
         13511 => x"06708106",
         13512 => x"5d568357",
         13513 => x"7b84ab38",
         13514 => x"75822a81",
         13515 => x"06408a57",
         13516 => x"7f849f38",
         13517 => x"9f3dfc05",
         13518 => x"53835279",
         13519 => x"51fed0e9",
         13520 => x"3f84bb84",
         13521 => x"08849838",
         13522 => x"6d557480",
         13523 => x"2e849038",
         13524 => x"74828080",
         13525 => x"26848838",
         13526 => x"ff157506",
         13527 => x"557483ff",
         13528 => x"387e802e",
         13529 => x"88388480",
         13530 => x"7f2683f8",
         13531 => x"387e8180",
         13532 => x"0a2683f0",
         13533 => x"38ff1f7f",
         13534 => x"06557483",
         13535 => x"e7387e89",
         13536 => x"2aa63d08",
         13537 => x"892a7089",
         13538 => x"2b77594c",
         13539 => x"475b6080",
         13540 => x"2e85ab38",
         13541 => x"65307080",
         13542 => x"25770756",
         13543 => x"5f915774",
         13544 => x"83b0387d",
         13545 => x"802e84df",
         13546 => x"38815474",
         13547 => x"53605279",
         13548 => x"51fecdf7",
         13549 => x"3f815784",
         13550 => x"bb840883",
         13551 => x"95386083",
         13552 => x"ff053361",
         13553 => x"83fe0533",
         13554 => x"71882b07",
         13555 => x"59568e57",
         13556 => x"7782d4d5",
         13557 => x"2e098106",
         13558 => x"82f8387d",
         13559 => x"90296105",
         13560 => x"83b21133",
         13561 => x"44586280",
         13562 => x"2e82e738",
         13563 => x"83b61883",
         13564 => x"11338212",
         13565 => x"3371902b",
         13566 => x"71882b07",
         13567 => x"81143370",
         13568 => x"7207882b",
         13569 => x"75337107",
         13570 => x"83ba1f83",
         13571 => x"11338212",
         13572 => x"3371902b",
         13573 => x"71882b07",
         13574 => x"81143370",
         13575 => x"7207882b",
         13576 => x"75337107",
         13577 => x"5ca23d0c",
         13578 => x"42a33d0c",
         13579 => x"a33d0c44",
         13580 => x"4e544559",
         13581 => x"4f415a4b",
         13582 => x"784d8e57",
         13583 => x"80ff7927",
         13584 => x"82903893",
         13585 => x"577a8180",
         13586 => x"26828738",
         13587 => x"61812a70",
         13588 => x"81064549",
         13589 => x"63802e83",
         13590 => x"f9386187",
         13591 => x"06456482",
         13592 => x"2e893861",
         13593 => x"81064766",
         13594 => x"83f43883",
         13595 => x"6e70304a",
         13596 => x"46437a58",
         13597 => x"62832e8a",
         13598 => x"c2387aae",
         13599 => x"38788c2a",
         13600 => x"57810b83",
         13601 => x"e8a82256",
         13602 => x"5874802e",
         13603 => x"9d387477",
         13604 => x"26983883",
         13605 => x"e8a85677",
         13606 => x"10821770",
         13607 => x"22575758",
         13608 => x"74802e86",
         13609 => x"38767527",
         13610 => x"ee387752",
         13611 => x"7851fcff",
         13612 => x"f43f84bb",
         13613 => x"84081084",
         13614 => x"055584bb",
         13615 => x"84089ff5",
         13616 => x"26963881",
         13617 => x"0b84bb84",
         13618 => x"081084bb",
         13619 => x"84080571",
         13620 => x"11722a83",
         13621 => x"05574c43",
         13622 => x"83ff1589",
         13623 => x"2a5d815c",
         13624 => x"a0477b1f",
         13625 => x"7d116805",
         13626 => x"6611ff05",
         13627 => x"706b0672",
         13628 => x"31584e57",
         13629 => x"4462832e",
         13630 => x"89b83874",
         13631 => x"1d5d7790",
         13632 => x"29167060",
         13633 => x"31565774",
         13634 => x"792682f2",
         13635 => x"38787c31",
         13636 => x"7d317853",
         13637 => x"70683152",
         13638 => x"56fcff89",
         13639 => x"3f84bb84",
         13640 => x"08406283",
         13641 => x"2e89f638",
         13642 => x"62822e09",
         13643 => x"810682dd",
         13644 => x"3883fff5",
         13645 => x"0b84bb84",
         13646 => x"082782ac",
         13647 => x"387a89f9",
         13648 => x"38771855",
         13649 => x"7480c026",
         13650 => x"89ef3874",
         13651 => x"5bfea339",
         13652 => x"8b577684",
         13653 => x"bb840c9f",
         13654 => x"3d0d84bb",
         13655 => x"900c0481",
         13656 => x"4efbfe39",
         13657 => x"930b84bb",
         13658 => x"840c9f3d",
         13659 => x"0d84bb90",
         13660 => x"0c047c33",
         13661 => x"d0117081",
         13662 => x"ff065757",
         13663 => x"57748926",
         13664 => x"9138821d",
         13665 => x"7781ff06",
         13666 => x"d0055d58",
         13667 => x"777a2e81",
         13668 => x"b238800b",
         13669 => x"83e6f45f",
         13670 => x"5c7d087d",
         13671 => x"575b7a70",
         13672 => x"81055c33",
         13673 => x"76708105",
         13674 => x"5833ff9f",
         13675 => x"12455957",
         13676 => x"62992689",
         13677 => x"38e01770",
         13678 => x"81ff0658",
         13679 => x"44ff9f18",
         13680 => x"45649926",
         13681 => x"8938e018",
         13682 => x"7081ff06",
         13683 => x"59467630",
         13684 => x"709f2a5a",
         13685 => x"4776782e",
         13686 => x"09810685",
         13687 => x"3878ffbe",
         13688 => x"38757a32",
         13689 => x"70307072",
         13690 => x"079f2a7b",
         13691 => x"075d4a4a",
         13692 => x"7a802e80",
         13693 => x"ce38811c",
         13694 => x"841f5f5c",
         13695 => x"837c25ff",
         13696 => x"98387f56",
         13697 => x"f9e0399f",
         13698 => x"3df80553",
         13699 => x"81527951",
         13700 => x"fecb963f",
         13701 => x"815784bb",
         13702 => x"8408feb6",
         13703 => x"3861832a",
         13704 => x"770684bb",
         13705 => x"84084056",
         13706 => x"758338bf",
         13707 => x"5f6c558e",
         13708 => x"577e7526",
         13709 => x"fe9c3874",
         13710 => x"7f3159fb",
         13711 => x"fb398156",
         13712 => x"fad2397b",
         13713 => x"8324ffba",
         13714 => x"387b7aa3",
         13715 => x"3d0c56f9",
         13716 => x"95396181",
         13717 => x"06489357",
         13718 => x"67802efd",
         13719 => x"f538826e",
         13720 => x"70304a46",
         13721 => x"43fc8b39",
         13722 => x"84bb8408",
         13723 => x"9ff5269d",
         13724 => x"387a8b38",
         13725 => x"77185b81",
         13726 => x"807b27fb",
         13727 => x"f5388e57",
         13728 => x"7684bb84",
         13729 => x"0c9f3d0d",
         13730 => x"84bb900c",
         13731 => x"04805562",
         13732 => x"812e8699",
         13733 => x"389ff560",
         13734 => x"278b3874",
         13735 => x"81065b8e",
         13736 => x"577afdae",
         13737 => x"38848061",
         13738 => x"57558076",
         13739 => x"70810558",
         13740 => x"34ff1555",
         13741 => x"74f4388b",
         13742 => x"6183e6c0",
         13743 => x"59575576",
         13744 => x"70810558",
         13745 => x"33767081",
         13746 => x"055834ff",
         13747 => x"155574ef",
         13748 => x"38608b05",
         13749 => x"45746534",
         13750 => x"82618c05",
         13751 => x"3477618d",
         13752 => x"05347b83",
         13753 => x"ffff064b",
         13754 => x"6a618e05",
         13755 => x"346a882a",
         13756 => x"5c7b618f",
         13757 => x"05348161",
         13758 => x"90053462",
         13759 => x"83327030",
         13760 => x"5a488061",
         13761 => x"91053478",
         13762 => x"9e2a8206",
         13763 => x"49686192",
         13764 => x"05346c56",
         13765 => x"7583ffff",
         13766 => x"2686ad38",
         13767 => x"7583ffff",
         13768 => x"06557461",
         13769 => x"93053474",
         13770 => x"882a4c6b",
         13771 => x"61940534",
         13772 => x"f8619505",
         13773 => x"34bf6198",
         13774 => x"05348061",
         13775 => x"990534ff",
         13776 => x"619a0534",
         13777 => x"80619b05",
         13778 => x"347e619c",
         13779 => x"05347e88",
         13780 => x"2a486761",
         13781 => x"9d05347e",
         13782 => x"902a4c6b",
         13783 => x"619e0534",
         13784 => x"7e982a84",
         13785 => x"bb900c84",
         13786 => x"bb900861",
         13787 => x"9f053462",
         13788 => x"832e85f7",
         13789 => x"388061a7",
         13790 => x"05348061",
         13791 => x"a80534a1",
         13792 => x"61a90534",
         13793 => x"80cc61aa",
         13794 => x"05347c83",
         13795 => x"ffff0655",
         13796 => x"74619605",
         13797 => x"3474882a",
         13798 => x"4b6a6197",
         13799 => x"0534ff80",
         13800 => x"61a40534",
         13801 => x"a961a605",
         13802 => x"349361ab",
         13803 => x"0583e6cc",
         13804 => x"59575576",
         13805 => x"70810558",
         13806 => x"33767081",
         13807 => x"055834ff",
         13808 => x"155574ef",
         13809 => x"386083fe",
         13810 => x"054980d5",
         13811 => x"69346083",
         13812 => x"ff054bff",
         13813 => x"aa6b3481",
         13814 => x"547e5360",
         13815 => x"527951fe",
         13816 => x"c6c83f81",
         13817 => x"5784bb84",
         13818 => x"08fae738",
         13819 => x"60175c62",
         13820 => x"832e879c",
         13821 => x"38696157",
         13822 => x"55807670",
         13823 => x"81055834",
         13824 => x"ff155574",
         13825 => x"f4386375",
         13826 => x"415b6283",
         13827 => x"2e86c038",
         13828 => x"87fffff8",
         13829 => x"5762812e",
         13830 => x"8338f857",
         13831 => x"76613476",
         13832 => x"882a7c45",
         13833 => x"55746470",
         13834 => x"81054634",
         13835 => x"76902a59",
         13836 => x"78647081",
         13837 => x"05463476",
         13838 => x"982a5675",
         13839 => x"64347c57",
         13840 => x"65597666",
         13841 => x"26833876",
         13842 => x"5978547a",
         13843 => x"53605279",
         13844 => x"51fec5d6",
         13845 => x"3f84bb84",
         13846 => x"0885e638",
         13847 => x"84806157",
         13848 => x"55807670",
         13849 => x"81055834",
         13850 => x"ff155574",
         13851 => x"f438781b",
         13852 => x"777a3158",
         13853 => x"5b76c938",
         13854 => x"7f810540",
         13855 => x"7f802eff",
         13856 => x"89387756",
         13857 => x"62832e83",
         13858 => x"38665665",
         13859 => x"55756626",
         13860 => x"83387555",
         13861 => x"74547a53",
         13862 => x"60527951",
         13863 => x"fec58b3f",
         13864 => x"84bb8408",
         13865 => x"859b3874",
         13866 => x"1b767631",
         13867 => x"575b75db",
         13868 => x"388c5862",
         13869 => x"832e9338",
         13870 => x"86586c83",
         13871 => x"ffff268a",
         13872 => x"38845862",
         13873 => x"822e8338",
         13874 => x"81587d84",
         13875 => x"c1386183",
         13876 => x"2a81065e",
         13877 => x"7d81b338",
         13878 => x"84806156",
         13879 => x"59807570",
         13880 => x"81055734",
         13881 => x"ff195978",
         13882 => x"f43880d5",
         13883 => x"6934ffaa",
         13884 => x"6b346083",
         13885 => x"be054778",
         13886 => x"67348167",
         13887 => x"81053481",
         13888 => x"67820534",
         13889 => x"78678305",
         13890 => x"34776784",
         13891 => x"05346c43",
         13892 => x"80fdc152",
         13893 => x"621f51fc",
         13894 => x"f78b3ffe",
         13895 => x"67850534",
         13896 => x"84bb8408",
         13897 => x"822abf07",
         13898 => x"57766786",
         13899 => x"053484bb",
         13900 => x"84086787",
         13901 => x"05347e61",
         13902 => x"83c60534",
         13903 => x"676183c7",
         13904 => x"05346b61",
         13905 => x"83c80534",
         13906 => x"84bb9008",
         13907 => x"6183c905",
         13908 => x"34626183",
         13909 => x"ca053462",
         13910 => x"882a4564",
         13911 => x"6183cb05",
         13912 => x"3462902a",
         13913 => x"58776183",
         13914 => x"cc053462",
         13915 => x"982a5f7e",
         13916 => x"6183cd05",
         13917 => x"34815478",
         13918 => x"53605279",
         13919 => x"51fec3aa",
         13920 => x"3f815784",
         13921 => x"bb8408f7",
         13922 => x"c9388053",
         13923 => x"80527951",
         13924 => x"fec4963f",
         13925 => x"815784bb",
         13926 => x"8408f7b6",
         13927 => x"3884bb84",
         13928 => x"0884bb84",
         13929 => x"0c9f3d0d",
         13930 => x"84bb900c",
         13931 => x"046255f9",
         13932 => x"e439741c",
         13933 => x"6416455c",
         13934 => x"f6c4397a",
         13935 => x"ae387891",
         13936 => x"2a57810b",
         13937 => x"83e8b822",
         13938 => x"56587480",
         13939 => x"2e9d3874",
         13940 => x"77269838",
         13941 => x"83e8b856",
         13942 => x"77108217",
         13943 => x"70225757",
         13944 => x"5874802e",
         13945 => x"86387675",
         13946 => x"27ee3877",
         13947 => x"527851fc",
         13948 => x"f5b33f84",
         13949 => x"bb840810",
         13950 => x"10848705",
         13951 => x"70892a5e",
         13952 => x"5ca05c80",
         13953 => x"0b84bb84",
         13954 => x"08fc808a",
         13955 => x"055847fd",
         13956 => x"fff00a77",
         13957 => x"27f5cb38",
         13958 => x"8e57f8e4",
         13959 => x"3984bb84",
         13960 => x"0883fff5",
         13961 => x"26f8e638",
         13962 => x"7af8d338",
         13963 => x"77812a5b",
         13964 => x"7af4bf38",
         13965 => x"8e57f8c8",
         13966 => x"39688106",
         13967 => x"4463802e",
         13968 => x"f8af3883",
         13969 => x"43f4ab39",
         13970 => x"7561a005",
         13971 => x"3475882a",
         13972 => x"496861a1",
         13973 => x"05347590",
         13974 => x"2a5b7a61",
         13975 => x"a2053475",
         13976 => x"982a5776",
         13977 => x"61a30534",
         13978 => x"f9c63980",
         13979 => x"6180c305",
         13980 => x"34806180",
         13981 => x"c40534a1",
         13982 => x"6180c505",
         13983 => x"3480cc61",
         13984 => x"80c60534",
         13985 => x"7c61a405",
         13986 => x"347c882a",
         13987 => x"5c7b61a5",
         13988 => x"05347c90",
         13989 => x"2a597861",
         13990 => x"a605347c",
         13991 => x"982a5675",
         13992 => x"61a70534",
         13993 => x"8261ac05",
         13994 => x"348061ad",
         13995 => x"05348061",
         13996 => x"ae053480",
         13997 => x"61af0534",
         13998 => x"8161b005",
         13999 => x"348061b1",
         14000 => x"05348661",
         14001 => x"b2053480",
         14002 => x"61b30534",
         14003 => x"ff806180",
         14004 => x"c00534a9",
         14005 => x"6180c205",
         14006 => x"34936180",
         14007 => x"c70583e6",
         14008 => x"e0595755",
         14009 => x"76708105",
         14010 => x"58337670",
         14011 => x"81055834",
         14012 => x"ff155574",
         14013 => x"802ef9cd",
         14014 => x"38767081",
         14015 => x"05583376",
         14016 => x"70810558",
         14017 => x"34ff1555",
         14018 => x"74da38f9",
         14019 => x"b8398154",
         14020 => x"80536052",
         14021 => x"7951febf",
         14022 => x"923f8157",
         14023 => x"84bb8408",
         14024 => x"f4b0387d",
         14025 => x"90296105",
         14026 => x"42776283",
         14027 => x"b2053476",
         14028 => x"5484bb84",
         14029 => x"08536052",
         14030 => x"7951febf",
         14031 => x"ed3ffcc3",
         14032 => x"39810b84",
         14033 => x"bb840c9f",
         14034 => x"3d0d84bb",
         14035 => x"900c04f8",
         14036 => x"61347b4a",
         14037 => x"ff6a7081",
         14038 => x"054c34ff",
         14039 => x"6a708105",
         14040 => x"4c34ff6a",
         14041 => x"34ff6184",
         14042 => x"0534ff61",
         14043 => x"850534ff",
         14044 => x"61860534",
         14045 => x"ff618705",
         14046 => x"34ff6188",
         14047 => x"0534ff61",
         14048 => x"890534ff",
         14049 => x"618a0534",
         14050 => x"8f65347c",
         14051 => x"57f9b139",
         14052 => x"7654861f",
         14053 => x"53605279",
         14054 => x"51febf8e",
         14055 => x"3f848061",
         14056 => x"56578075",
         14057 => x"70810557",
         14058 => x"34ff1757",
         14059 => x"76f43860",
         14060 => x"5c80d27c",
         14061 => x"7081055e",
         14062 => x"347b5580",
         14063 => x"d2757081",
         14064 => x"05573480",
         14065 => x"e1757081",
         14066 => x"05573480",
         14067 => x"c1753480",
         14068 => x"f26183e4",
         14069 => x"053480f2",
         14070 => x"6183e505",
         14071 => x"3480c161",
         14072 => x"83e60534",
         14073 => x"80e16183",
         14074 => x"e705347f",
         14075 => x"ff055b7a",
         14076 => x"6183e805",
         14077 => x"347a882a",
         14078 => x"59786183",
         14079 => x"e905347a",
         14080 => x"902a5675",
         14081 => x"6183ea05",
         14082 => x"347a982a",
         14083 => x"407f6183",
         14084 => x"eb053482",
         14085 => x"6183ec05",
         14086 => x"34766183",
         14087 => x"ed053476",
         14088 => x"6183ee05",
         14089 => x"34766183",
         14090 => x"ef053480",
         14091 => x"d56934ff",
         14092 => x"aa6b3481",
         14093 => x"54871f53",
         14094 => x"60527951",
         14095 => x"febdeb3f",
         14096 => x"8154811f",
         14097 => x"53605279",
         14098 => x"51febdde",
         14099 => x"3f696157",
         14100 => x"55f7a639",
         14101 => x"f43d0d7e",
         14102 => x"615b5b80",
         14103 => x"7b61ff05",
         14104 => x"5a575776",
         14105 => x"7825b838",
         14106 => x"8d3d598e",
         14107 => x"3df80554",
         14108 => x"81537852",
         14109 => x"7951ff9b",
         14110 => x"cc3f7b81",
         14111 => x"2e098106",
         14112 => x"9e388d3d",
         14113 => x"3355748d",
         14114 => x"2e903874",
         14115 => x"76708105",
         14116 => x"58348117",
         14117 => x"57748a2e",
         14118 => x"86387777",
         14119 => x"24cd3880",
         14120 => x"76347a55",
         14121 => x"76833876",
         14122 => x"557484bb",
         14123 => x"840c8e3d",
         14124 => x"0d04f73d",
         14125 => x"0d7b0284",
         14126 => x"05b30533",
         14127 => x"5957778a",
         14128 => x"2e80d538",
         14129 => x"84170856",
         14130 => x"8076249e",
         14131 => x"38881708",
         14132 => x"77178c05",
         14133 => x"56597775",
         14134 => x"34811655",
         14135 => x"74bb248e",
         14136 => x"38748418",
         14137 => x"0c811988",
         14138 => x"180c8b3d",
         14139 => x"0d048b3d",
         14140 => x"fc055474",
         14141 => x"538c1752",
         14142 => x"760851ff",
         14143 => x"9fa73f74",
         14144 => x"7a327030",
         14145 => x"7072079f",
         14146 => x"2a703084",
         14147 => x"1b0c811c",
         14148 => x"881b0c5a",
         14149 => x"5656d339",
         14150 => x"8d527651",
         14151 => x"ff943fff",
         14152 => x"a339e33d",
         14153 => x"0d0280ff",
         14154 => x"05338d3d",
         14155 => x"585880cc",
         14156 => x"77575580",
         14157 => x"76708105",
         14158 => x"5834ff15",
         14159 => x"5574f438",
         14160 => x"a13d0877",
         14161 => x"0c778a2e",
         14162 => x"80f7387c",
         14163 => x"56807624",
         14164 => x"80c0387d",
         14165 => x"77178c05",
         14166 => x"56597775",
         14167 => x"34811655",
         14168 => x"74bb24b8",
         14169 => x"38748418",
         14170 => x"0c811988",
         14171 => x"180c7c55",
         14172 => x"8075249e",
         14173 => x"389f3dff",
         14174 => x"ac115575",
         14175 => x"54c00552",
         14176 => x"760851ff",
         14177 => x"9e9f3f84",
         14178 => x"bb840886",
         14179 => x"387c7a2e",
         14180 => x"ba38ff0b",
         14181 => x"84bb840c",
         14182 => x"9f3d0d04",
         14183 => x"9f3dffb0",
         14184 => x"11557554",
         14185 => x"c0055276",
         14186 => x"0851ff9d",
         14187 => x"f83f747b",
         14188 => x"32703070",
         14189 => x"72079f2a",
         14190 => x"7030525a",
         14191 => x"5656ffa5",
         14192 => x"398d5276",
         14193 => x"51fdeb3f",
         14194 => x"ff81397d",
         14195 => x"84bb840c",
         14196 => x"9f3d0d04",
         14197 => x"fd3d0d75",
         14198 => x"0284059a",
         14199 => x"05225253",
         14200 => x"80527280",
         14201 => x"ff269038",
         14202 => x"7283ffff",
         14203 => x"06527184",
         14204 => x"bb840c85",
         14205 => x"3d0d0483",
         14206 => x"ffff7327",
         14207 => x"547083b5",
         14208 => x"2e098106",
         14209 => x"e9387380",
         14210 => x"2ee43883",
         14211 => x"e8c82251",
         14212 => x"72712e9c",
         14213 => x"38811270",
         14214 => x"83ffff06",
         14215 => x"53547180",
         14216 => x"ff268d38",
         14217 => x"711083e8",
         14218 => x"c8057022",
         14219 => x"5151e139",
         14220 => x"81801270",
         14221 => x"81ff0684",
         14222 => x"bb840c53",
         14223 => x"853d0d04",
         14224 => x"fe3d0d02",
         14225 => x"92052202",
         14226 => x"84059605",
         14227 => x"22535180",
         14228 => x"537080ff",
         14229 => x"268c3870",
         14230 => x"537284bb",
         14231 => x"840c843d",
         14232 => x"0d047183",
         14233 => x"b52e0981",
         14234 => x"06ef3870",
         14235 => x"81ff26e9",
         14236 => x"38701083",
         14237 => x"e6c80570",
         14238 => x"2284bb84",
         14239 => x"0c51843d",
         14240 => x"0d04fb3d",
         14241 => x"0d775170",
         14242 => x"83ffff26",
         14243 => x"80e13870",
         14244 => x"83ffff06",
         14245 => x"83eac856",
         14246 => x"56759fff",
         14247 => x"2680d938",
         14248 => x"74708205",
         14249 => x"56227571",
         14250 => x"30708025",
         14251 => x"737a2607",
         14252 => x"54565353",
         14253 => x"70b73871",
         14254 => x"70820553",
         14255 => x"22727188",
         14256 => x"2a545681",
         14257 => x"ff067014",
         14258 => x"52547076",
         14259 => x"24b13871",
         14260 => x"cf387310",
         14261 => x"15707082",
         14262 => x"05522254",
         14263 => x"73307080",
         14264 => x"25757926",
         14265 => x"07535552",
         14266 => x"70802ecb",
         14267 => x"38755170",
         14268 => x"84bb840c",
         14269 => x"873d0d04",
         14270 => x"83eebc55",
         14271 => x"ffa23971",
         14272 => x"8826ea38",
         14273 => x"71101083",
         14274 => x"caf00554",
         14275 => x"730804c7",
         14276 => x"a0167083",
         14277 => x"ffff0657",
         14278 => x"517551d3",
         14279 => x"39ffb016",
         14280 => x"7083ffff",
         14281 => x"065751f1",
         14282 => x"39881670",
         14283 => x"83ffff06",
         14284 => x"5751e639",
         14285 => x"e6167083",
         14286 => x"ffff0657",
         14287 => x"51db39d0",
         14288 => x"167083ff",
         14289 => x"ff065751",
         14290 => x"d039e016",
         14291 => x"7083ffff",
         14292 => x"065751c5",
         14293 => x"39f01670",
         14294 => x"83ffff06",
         14295 => x"5751ffb9",
         14296 => x"39757331",
         14297 => x"81067671",
         14298 => x"317083ff",
         14299 => x"ff065852",
         14300 => x"55ffa639",
         14301 => x"75733110",
         14302 => x"75057022",
         14303 => x"5252feef",
         14304 => x"39000000",
         14305 => x"00ffffff",
         14306 => x"ff00ffff",
         14307 => x"ffff00ff",
         14308 => x"ffffff00",
         14309 => x"0000198b",
         14310 => x"00001980",
         14311 => x"00001975",
         14312 => x"0000196a",
         14313 => x"0000195f",
         14314 => x"00001954",
         14315 => x"00001949",
         14316 => x"0000193e",
         14317 => x"00001933",
         14318 => x"00001928",
         14319 => x"0000191d",
         14320 => x"00001912",
         14321 => x"00001907",
         14322 => x"000018fc",
         14323 => x"000018f1",
         14324 => x"000018e6",
         14325 => x"000018db",
         14326 => x"000018d0",
         14327 => x"000018c5",
         14328 => x"000018ba",
         14329 => x"00001eca",
         14330 => x"00001f64",
         14331 => x"00001f64",
         14332 => x"00001f64",
         14333 => x"00001f64",
         14334 => x"00001f64",
         14335 => x"00001f64",
         14336 => x"00001f64",
         14337 => x"00001f64",
         14338 => x"00001f64",
         14339 => x"00001f64",
         14340 => x"00001f64",
         14341 => x"00001f64",
         14342 => x"00001f64",
         14343 => x"00001f64",
         14344 => x"00001f64",
         14345 => x"00001f64",
         14346 => x"00001f64",
         14347 => x"00001f64",
         14348 => x"00001f64",
         14349 => x"00001f64",
         14350 => x"00001f64",
         14351 => x"00001f64",
         14352 => x"00001f64",
         14353 => x"00001f64",
         14354 => x"00001f64",
         14355 => x"00001f64",
         14356 => x"00001f64",
         14357 => x"00001f64",
         14358 => x"00001f64",
         14359 => x"00001f64",
         14360 => x"00001f64",
         14361 => x"00001f64",
         14362 => x"00001f64",
         14363 => x"00001f64",
         14364 => x"00001f64",
         14365 => x"00001f64",
         14366 => x"00001f64",
         14367 => x"00001f64",
         14368 => x"00001f64",
         14369 => x"00001f64",
         14370 => x"00001f64",
         14371 => x"00001f64",
         14372 => x"00002481",
         14373 => x"00001f64",
         14374 => x"00001f64",
         14375 => x"00001f64",
         14376 => x"00001f64",
         14377 => x"00001f64",
         14378 => x"00001f64",
         14379 => x"00001f64",
         14380 => x"00001f64",
         14381 => x"00001f64",
         14382 => x"00001f64",
         14383 => x"00001f64",
         14384 => x"00001f64",
         14385 => x"00001f64",
         14386 => x"00001f64",
         14387 => x"00001f64",
         14388 => x"00001f64",
         14389 => x"00002417",
         14390 => x"00002316",
         14391 => x"00001f64",
         14392 => x"0000229a",
         14393 => x"000024b8",
         14394 => x"00002377",
         14395 => x"0000223c",
         14396 => x"000021de",
         14397 => x"00001f64",
         14398 => x"00001f64",
         14399 => x"00001f64",
         14400 => x"00001f64",
         14401 => x"00001f64",
         14402 => x"00001f64",
         14403 => x"00001f64",
         14404 => x"00001f64",
         14405 => x"00001f64",
         14406 => x"00001f64",
         14407 => x"00001f64",
         14408 => x"00001f64",
         14409 => x"00001f64",
         14410 => x"00001f64",
         14411 => x"00001f64",
         14412 => x"00001f64",
         14413 => x"00001f64",
         14414 => x"00001f64",
         14415 => x"00001f64",
         14416 => x"00001f64",
         14417 => x"00001f64",
         14418 => x"00001f64",
         14419 => x"00001f64",
         14420 => x"00001f64",
         14421 => x"00001f64",
         14422 => x"00001f64",
         14423 => x"00001f64",
         14424 => x"00001f64",
         14425 => x"00001f64",
         14426 => x"00001f64",
         14427 => x"00001f64",
         14428 => x"00001f64",
         14429 => x"00001f64",
         14430 => x"00001f64",
         14431 => x"00001f64",
         14432 => x"00001f64",
         14433 => x"00001f64",
         14434 => x"00001f64",
         14435 => x"00001f64",
         14436 => x"00001f64",
         14437 => x"00001f64",
         14438 => x"00001f64",
         14439 => x"00001f64",
         14440 => x"00001f64",
         14441 => x"00001f64",
         14442 => x"00001f64",
         14443 => x"00001f64",
         14444 => x"00001f64",
         14445 => x"00001f64",
         14446 => x"00001f64",
         14447 => x"00001f64",
         14448 => x"00001f64",
         14449 => x"000021bb",
         14450 => x"00002180",
         14451 => x"00001f64",
         14452 => x"00001f64",
         14453 => x"00001f64",
         14454 => x"00001f64",
         14455 => x"00001f64",
         14456 => x"00001f64",
         14457 => x"00001f64",
         14458 => x"00001f64",
         14459 => x"00002173",
         14460 => x"00002168",
         14461 => x"00001f64",
         14462 => x"00002150",
         14463 => x"00001f64",
         14464 => x"00002161",
         14465 => x"00002156",
         14466 => x"00002149",
         14467 => x"00003233",
         14468 => x"0000324b",
         14469 => x"00003257",
         14470 => x"00003263",
         14471 => x"0000326f",
         14472 => x"0000323f",
         14473 => x"00003c10",
         14474 => x"00003a9a",
         14475 => x"00003962",
         14476 => x"00003690",
         14477 => x"00003bac",
         14478 => x"000034fd",
         14479 => x"000037fc",
         14480 => x"000036b5",
         14481 => x"00003a44",
         14482 => x"000036e4",
         14483 => x"00003759",
         14484 => x"0000398b",
         14485 => x"000034fd",
         14486 => x"00003962",
         14487 => x"0000386c",
         14488 => x"000037fc",
         14489 => x"000034fd",
         14490 => x"000034fd",
         14491 => x"00003759",
         14492 => x"000036e4",
         14493 => x"000036b5",
         14494 => x"00003690",
         14495 => x"00004744",
         14496 => x"0000475d",
         14497 => x"00004782",
         14498 => x"000047a3",
         14499 => x"00004704",
         14500 => x"000047c8",
         14501 => x"0000471d",
         14502 => x"0000486d",
         14503 => x"0000482a",
         14504 => x"0000482a",
         14505 => x"0000482a",
         14506 => x"0000482a",
         14507 => x"0000482a",
         14508 => x"0000482a",
         14509 => x"00004803",
         14510 => x"0000482a",
         14511 => x"0000482a",
         14512 => x"0000482a",
         14513 => x"0000482a",
         14514 => x"0000482a",
         14515 => x"0000482a",
         14516 => x"0000482a",
         14517 => x"0000482a",
         14518 => x"0000482a",
         14519 => x"0000482a",
         14520 => x"0000482a",
         14521 => x"0000482a",
         14522 => x"0000482a",
         14523 => x"0000482a",
         14524 => x"0000482a",
         14525 => x"0000482a",
         14526 => x"0000482a",
         14527 => x"0000482a",
         14528 => x"0000482a",
         14529 => x"0000482a",
         14530 => x"0000482a",
         14531 => x"0000482a",
         14532 => x"00004942",
         14533 => x"00004930",
         14534 => x"0000491d",
         14535 => x"0000490a",
         14536 => x"00004834",
         14537 => x"000048f8",
         14538 => x"000048e5",
         14539 => x"0000484d",
         14540 => x"0000482a",
         14541 => x"0000484d",
         14542 => x"000048d5",
         14543 => x"00004952",
         14544 => x"0000487e",
         14545 => x"0000485c",
         14546 => x"000048c3",
         14547 => x"000048b1",
         14548 => x"0000489f",
         14549 => x"00004890",
         14550 => x"0000482a",
         14551 => x"00004834",
         14552 => x"000054d0",
         14553 => x"0000563f",
         14554 => x"00005611",
         14555 => x"00005568",
         14556 => x"00005545",
         14557 => x"00005524",
         14558 => x"000054fa",
         14559 => x"000056ca",
         14560 => x"00005351",
         14561 => x"000056a4",
         14562 => x"00005893",
         14563 => x"00005351",
         14564 => x"00005351",
         14565 => x"00005351",
         14566 => x"00005351",
         14567 => x"00005351",
         14568 => x"00005351",
         14569 => x"0000566d",
         14570 => x"0000587b",
         14571 => x"00005732",
         14572 => x"00005351",
         14573 => x"00005351",
         14574 => x"00005351",
         14575 => x"00005351",
         14576 => x"00005351",
         14577 => x"00005351",
         14578 => x"00005351",
         14579 => x"00005351",
         14580 => x"00005351",
         14581 => x"00005351",
         14582 => x"00005351",
         14583 => x"00005351",
         14584 => x"00005351",
         14585 => x"00005351",
         14586 => x"00005351",
         14587 => x"00005351",
         14588 => x"00005351",
         14589 => x"00005351",
         14590 => x"00005351",
         14591 => x"000055ef",
         14592 => x"00005351",
         14593 => x"00005351",
         14594 => x"00005351",
         14595 => x"00005592",
         14596 => x"000054a1",
         14597 => x"00005443",
         14598 => x"00005351",
         14599 => x"00005351",
         14600 => x"00005351",
         14601 => x"00005351",
         14602 => x"00005428",
         14603 => x"00005351",
         14604 => x"0000540b",
         14605 => x"00005a74",
         14606 => x"000059e9",
         14607 => x"000059e9",
         14608 => x"000059e9",
         14609 => x"000059e9",
         14610 => x"000059e9",
         14611 => x"000059e9",
         14612 => x"000059c4",
         14613 => x"000059e9",
         14614 => x"000059e9",
         14615 => x"000059e9",
         14616 => x"000059e9",
         14617 => x"000059e9",
         14618 => x"000059e9",
         14619 => x"000059e9",
         14620 => x"000059e9",
         14621 => x"000059e9",
         14622 => x"000059e9",
         14623 => x"000059e9",
         14624 => x"000059e9",
         14625 => x"000059e9",
         14626 => x"000059e9",
         14627 => x"000059e9",
         14628 => x"000059e9",
         14629 => x"000059e9",
         14630 => x"000059e9",
         14631 => x"000059e9",
         14632 => x"000059e9",
         14633 => x"000059e9",
         14634 => x"000059e9",
         14635 => x"00005a86",
         14636 => x"00005ace",
         14637 => x"00005abb",
         14638 => x"00005aa8",
         14639 => x"00005a96",
         14640 => x"00005b59",
         14641 => x"00005b46",
         14642 => x"00005b36",
         14643 => x"000059e9",
         14644 => x"00005b26",
         14645 => x"00005b16",
         14646 => x"00005b04",
         14647 => x"00005af2",
         14648 => x"00005ae0",
         14649 => x"00005a51",
         14650 => x"00005a40",
         14651 => x"00005a2f",
         14652 => x"00005a18",
         14653 => x"000059e9",
         14654 => x"00005a62",
         14655 => x"00006443",
         14656 => x"0000629f",
         14657 => x"0000629f",
         14658 => x"0000629f",
         14659 => x"0000629f",
         14660 => x"0000629f",
         14661 => x"0000629f",
         14662 => x"0000629f",
         14663 => x"0000629f",
         14664 => x"0000629f",
         14665 => x"0000629f",
         14666 => x"0000629f",
         14667 => x"0000629f",
         14668 => x"0000629f",
         14669 => x"00005fc1",
         14670 => x"0000629f",
         14671 => x"0000629f",
         14672 => x"0000629f",
         14673 => x"0000629f",
         14674 => x"0000629f",
         14675 => x"0000629f",
         14676 => x"0000648d",
         14677 => x"0000629f",
         14678 => x"0000629f",
         14679 => x"00006418",
         14680 => x"0000629f",
         14681 => x"0000642f",
         14682 => x"00005fa0",
         14683 => x"00006401",
         14684 => x"0000df74",
         14685 => x"0000df61",
         14686 => x"0000df55",
         14687 => x"0000df4a",
         14688 => x"0000df3f",
         14689 => x"0000df34",
         14690 => x"0000df29",
         14691 => x"0000df1d",
         14692 => x"0000df0f",
         14693 => x"00000e01",
         14694 => x"00000bfd",
         14695 => x"00000bfd",
         14696 => x"00000f49",
         14697 => x"00000bfd",
         14698 => x"00000bfd",
         14699 => x"00000bfd",
         14700 => x"00000bfd",
         14701 => x"00000bfd",
         14702 => x"00000bfd",
         14703 => x"00000bfd",
         14704 => x"00000dfd",
         14705 => x"00000bfd",
         14706 => x"00000f7f",
         14707 => x"00000f0d",
         14708 => x"00000bfd",
         14709 => x"00000bfd",
         14710 => x"00000bfd",
         14711 => x"00000bfd",
         14712 => x"00000bfd",
         14713 => x"00000bfd",
         14714 => x"00000bfd",
         14715 => x"00000bfd",
         14716 => x"00000bfd",
         14717 => x"00000bfd",
         14718 => x"00000bfd",
         14719 => x"00000bfd",
         14720 => x"00000bfd",
         14721 => x"00000bfd",
         14722 => x"00000bfd",
         14723 => x"00000bfd",
         14724 => x"00000bfd",
         14725 => x"00000bfd",
         14726 => x"00000bfd",
         14727 => x"00000bfd",
         14728 => x"00000bfd",
         14729 => x"00000bfd",
         14730 => x"00000bfd",
         14731 => x"00000bfd",
         14732 => x"00000bfd",
         14733 => x"00000bfd",
         14734 => x"00000bfd",
         14735 => x"00000bfd",
         14736 => x"00000bfd",
         14737 => x"00000bfd",
         14738 => x"00000bfd",
         14739 => x"00000bfd",
         14740 => x"00000bfd",
         14741 => x"00000bfd",
         14742 => x"00000bfd",
         14743 => x"00000bfd",
         14744 => x"00000f1d",
         14745 => x"00000bfd",
         14746 => x"00000bfd",
         14747 => x"00000bfd",
         14748 => x"00000bfd",
         14749 => x"00000e17",
         14750 => x"00000bfd",
         14751 => x"00000bfd",
         14752 => x"00000bfd",
         14753 => x"00000bfd",
         14754 => x"00000bfd",
         14755 => x"00000bfd",
         14756 => x"00000bfd",
         14757 => x"00000bfd",
         14758 => x"00000bfd",
         14759 => x"00000bfd",
         14760 => x"00000e2b",
         14761 => x"00000ee1",
         14762 => x"00000eb8",
         14763 => x"00000eb8",
         14764 => x"00000eb8",
         14765 => x"00000bfd",
         14766 => x"00000ee1",
         14767 => x"00000bfd",
         14768 => x"00000bfd",
         14769 => x"00000eff",
         14770 => x"00000bfd",
         14771 => x"00000bfd",
         14772 => x"00000c16",
         14773 => x"00000e0f",
         14774 => x"00000bfd",
         14775 => x"00000bfd",
         14776 => x"00000f58",
         14777 => x"00000bfd",
         14778 => x"00000c18",
         14779 => x"00000bfd",
         14780 => x"00000bfd",
         14781 => x"00000e17",
         14782 => x"64696e69",
         14783 => x"74000000",
         14784 => x"64696f63",
         14785 => x"746c0000",
         14786 => x"66696e69",
         14787 => x"74000000",
         14788 => x"666c6f61",
         14789 => x"64000000",
         14790 => x"66657865",
         14791 => x"63000000",
         14792 => x"6d636c65",
         14793 => x"61720000",
         14794 => x"6d636f70",
         14795 => x"79000000",
         14796 => x"6d646966",
         14797 => x"66000000",
         14798 => x"6d64756d",
         14799 => x"70000000",
         14800 => x"6d656200",
         14801 => x"6d656800",
         14802 => x"6d657700",
         14803 => x"68696400",
         14804 => x"68696500",
         14805 => x"68666400",
         14806 => x"68666500",
         14807 => x"63616c6c",
         14808 => x"00000000",
         14809 => x"6a6d7000",
         14810 => x"72657374",
         14811 => x"61727400",
         14812 => x"72657365",
         14813 => x"74000000",
         14814 => x"696e666f",
         14815 => x"00000000",
         14816 => x"74657374",
         14817 => x"00000000",
         14818 => x"636c7300",
         14819 => x"7a383000",
         14820 => x"74626173",
         14821 => x"69630000",
         14822 => x"6d626173",
         14823 => x"69630000",
         14824 => x"6b696c6f",
         14825 => x"00000000",
         14826 => x"65640000",
         14827 => x"556e6b6e",
         14828 => x"6f776e20",
         14829 => x"6572726f",
         14830 => x"722e0000",
         14831 => x"50617261",
         14832 => x"6d657465",
         14833 => x"72732069",
         14834 => x"6e636f72",
         14835 => x"72656374",
         14836 => x"2e000000",
         14837 => x"546f6f20",
         14838 => x"6d616e79",
         14839 => x"206f7065",
         14840 => x"6e206669",
         14841 => x"6c65732e",
         14842 => x"00000000",
         14843 => x"496e7375",
         14844 => x"66666963",
         14845 => x"69656e74",
         14846 => x"206d656d",
         14847 => x"6f72792e",
         14848 => x"00000000",
         14849 => x"46696c65",
         14850 => x"20697320",
         14851 => x"6c6f636b",
         14852 => x"65642e00",
         14853 => x"54696d65",
         14854 => x"6f75742c",
         14855 => x"206f7065",
         14856 => x"72617469",
         14857 => x"6f6e2063",
         14858 => x"616e6365",
         14859 => x"6c6c6564",
         14860 => x"2e000000",
         14861 => x"466f726d",
         14862 => x"61742061",
         14863 => x"626f7274",
         14864 => x"65642e00",
         14865 => x"4e6f2063",
         14866 => x"6f6d7061",
         14867 => x"7469626c",
         14868 => x"65206669",
         14869 => x"6c657379",
         14870 => x"7374656d",
         14871 => x"20666f75",
         14872 => x"6e64206f",
         14873 => x"6e206469",
         14874 => x"736b2e00",
         14875 => x"4469736b",
         14876 => x"206e6f74",
         14877 => x"20656e61",
         14878 => x"626c6564",
         14879 => x"2e000000",
         14880 => x"44726976",
         14881 => x"65206e75",
         14882 => x"6d626572",
         14883 => x"20697320",
         14884 => x"696e7661",
         14885 => x"6c69642e",
         14886 => x"00000000",
         14887 => x"53442069",
         14888 => x"73207772",
         14889 => x"69746520",
         14890 => x"70726f74",
         14891 => x"65637465",
         14892 => x"642e0000",
         14893 => x"46696c65",
         14894 => x"2068616e",
         14895 => x"646c6520",
         14896 => x"696e7661",
         14897 => x"6c69642e",
         14898 => x"00000000",
         14899 => x"46696c65",
         14900 => x"20616c72",
         14901 => x"65616479",
         14902 => x"20657869",
         14903 => x"7374732e",
         14904 => x"00000000",
         14905 => x"41636365",
         14906 => x"73732064",
         14907 => x"656e6965",
         14908 => x"642e0000",
         14909 => x"496e7661",
         14910 => x"6c696420",
         14911 => x"66696c65",
         14912 => x"6e616d65",
         14913 => x"2e000000",
         14914 => x"4e6f2070",
         14915 => x"61746820",
         14916 => x"666f756e",
         14917 => x"642e0000",
         14918 => x"4e6f2066",
         14919 => x"696c6520",
         14920 => x"666f756e",
         14921 => x"642e0000",
         14922 => x"4469736b",
         14923 => x"206e6f74",
         14924 => x"20726561",
         14925 => x"64792e00",
         14926 => x"496e7465",
         14927 => x"726e616c",
         14928 => x"20657272",
         14929 => x"6f722e00",
         14930 => x"4469736b",
         14931 => x"20457272",
         14932 => x"6f720000",
         14933 => x"53756363",
         14934 => x"6573732e",
         14935 => x"00000000",
         14936 => x"0a256c75",
         14937 => x"20627974",
         14938 => x"65732025",
         14939 => x"73206174",
         14940 => x"20256c75",
         14941 => x"20627974",
         14942 => x"65732f73",
         14943 => x"65632e0a",
         14944 => x"00000000",
         14945 => x"72656164",
         14946 => x"00000000",
         14947 => x"2530386c",
         14948 => x"58000000",
         14949 => x"3a202000",
         14950 => x"25303258",
         14951 => x"00000000",
         14952 => x"207c0000",
         14953 => x"7c000000",
         14954 => x"20200000",
         14955 => x"25303458",
         14956 => x"00000000",
         14957 => x"20202020",
         14958 => x"20202020",
         14959 => x"00000000",
         14960 => x"7a4f5300",
         14961 => x"2a2a2025",
         14962 => x"73202800",
         14963 => x"32352f30",
         14964 => x"372f3230",
         14965 => x"32310000",
         14966 => x"76312e33",
         14967 => x"32000000",
         14968 => x"205a5055",
         14969 => x"2c207265",
         14970 => x"76202530",
         14971 => x"32782920",
         14972 => x"25732025",
         14973 => x"73202a2a",
         14974 => x"0a0a0000",
         14975 => x"4f533a00",
         14976 => x"20202020",
         14977 => x"42617365",
         14978 => x"20416464",
         14979 => x"72657373",
         14980 => x"20202020",
         14981 => x"20202020",
         14982 => x"20202020",
         14983 => x"203d2025",
         14984 => x"30386c78",
         14985 => x"0a000000",
         14986 => x"20202020",
         14987 => x"41707020",
         14988 => x"41646472",
         14989 => x"65737320",
         14990 => x"20202020",
         14991 => x"20202020",
         14992 => x"20202020",
         14993 => x"203d2025",
         14994 => x"30386c78",
         14995 => x"0a000000",
         14996 => x"5a505520",
         14997 => x"496e7465",
         14998 => x"72727570",
         14999 => x"74204861",
         15000 => x"6e646c65",
         15001 => x"72000000",
         15002 => x"55415254",
         15003 => x"31205458",
         15004 => x"20696e74",
         15005 => x"65727275",
         15006 => x"70740000",
         15007 => x"55415254",
         15008 => x"31205258",
         15009 => x"20696e74",
         15010 => x"65727275",
         15011 => x"70740000",
         15012 => x"55415254",
         15013 => x"30205458",
         15014 => x"20696e74",
         15015 => x"65727275",
         15016 => x"70740000",
         15017 => x"55415254",
         15018 => x"30205258",
         15019 => x"20696e74",
         15020 => x"65727275",
         15021 => x"70740000",
         15022 => x"494f4354",
         15023 => x"4c205752",
         15024 => x"20696e74",
         15025 => x"65727275",
         15026 => x"70740000",
         15027 => x"494f4354",
         15028 => x"4c205244",
         15029 => x"20696e74",
         15030 => x"65727275",
         15031 => x"70740000",
         15032 => x"50533220",
         15033 => x"696e7465",
         15034 => x"72727570",
         15035 => x"74000000",
         15036 => x"54696d65",
         15037 => x"7220696e",
         15038 => x"74657272",
         15039 => x"75707400",
         15040 => x"53657474",
         15041 => x"696e6720",
         15042 => x"75702074",
         15043 => x"696d6572",
         15044 => x"2e2e2e00",
         15045 => x"456e6162",
         15046 => x"6c696e67",
         15047 => x"2074696d",
         15048 => x"65722e2e",
         15049 => x"2e000000",
         15050 => x"6175746f",
         15051 => x"65786563",
         15052 => x"2e626174",
         15053 => x"00000000",
         15054 => x"7a4f535f",
         15055 => x"7a70752e",
         15056 => x"68737400",
         15057 => x"4661696c",
         15058 => x"65642074",
         15059 => x"6f20696e",
         15060 => x"69746961",
         15061 => x"6c697365",
         15062 => x"20736420",
         15063 => x"63617264",
         15064 => x"20302c20",
         15065 => x"706c6561",
         15066 => x"73652069",
         15067 => x"6e697420",
         15068 => x"6d616e75",
         15069 => x"616c6c79",
         15070 => x"2e000000",
         15071 => x"2a200000",
         15072 => x"25643a5c",
         15073 => x"25730000",
         15074 => x"303a0000",
         15075 => x"42616420",
         15076 => x"636f6d6d",
         15077 => x"616e642e",
         15078 => x"00000000",
         15079 => x"5a505500",
         15080 => x"62696e00",
         15081 => x"25643a5c",
         15082 => x"25735c25",
         15083 => x"732e2573",
         15084 => x"00000000",
         15085 => x"436f6c64",
         15086 => x"20726562",
         15087 => x"6f6f7469",
         15088 => x"6e672e2e",
         15089 => x"2e000000",
         15090 => x"52657374",
         15091 => x"61727469",
         15092 => x"6e672061",
         15093 => x"70706c69",
         15094 => x"63617469",
         15095 => x"6f6e2e2e",
         15096 => x"2e000000",
         15097 => x"43616c6c",
         15098 => x"696e6720",
         15099 => x"636f6465",
         15100 => x"20402025",
         15101 => x"30386c78",
         15102 => x"202e2e2e",
         15103 => x"0a000000",
         15104 => x"43616c6c",
         15105 => x"20726574",
         15106 => x"75726e65",
         15107 => x"6420636f",
         15108 => x"64652028",
         15109 => x"2564292e",
         15110 => x"0a000000",
         15111 => x"45786563",
         15112 => x"7574696e",
         15113 => x"6720636f",
         15114 => x"64652040",
         15115 => x"20253038",
         15116 => x"6c78202e",
         15117 => x"2e2e0a00",
         15118 => x"2530386c",
         15119 => x"58202530",
         15120 => x"386c582d",
         15121 => x"00000000",
         15122 => x"2530386c",
         15123 => x"58202530",
         15124 => x"34582d00",
         15125 => x"436f6d70",
         15126 => x"6172696e",
         15127 => x"672e2e2e",
         15128 => x"00000000",
         15129 => x"2530386c",
         15130 => x"78282530",
         15131 => x"3878292d",
         15132 => x"3e253038",
         15133 => x"6c782825",
         15134 => x"30387829",
         15135 => x"0a000000",
         15136 => x"436f7079",
         15137 => x"696e672e",
         15138 => x"2e2e0000",
         15139 => x"2530386c",
         15140 => x"58202530",
         15141 => x"32582d00",
         15142 => x"436c6561",
         15143 => x"72696e67",
         15144 => x"2e2e2e2e",
         15145 => x"00000000",
         15146 => x"44756d70",
         15147 => x"204d656d",
         15148 => x"6f727900",
         15149 => x"0a436f6d",
         15150 => x"706c6574",
         15151 => x"652e0000",
         15152 => x"25643a5c",
         15153 => x"25735c25",
         15154 => x"73000000",
         15155 => x"4d656d6f",
         15156 => x"72792065",
         15157 => x"78686175",
         15158 => x"73746564",
         15159 => x"2c206361",
         15160 => x"6e6e6f74",
         15161 => x"2070726f",
         15162 => x"63657373",
         15163 => x"20636f6d",
         15164 => x"6d616e64",
         15165 => x"2e000000",
         15166 => x"3f3f3f00",
         15167 => x"25642f25",
         15168 => x"642f2564",
         15169 => x"2025643a",
         15170 => x"25643a25",
         15171 => x"642e2564",
         15172 => x"25640a00",
         15173 => x"536f4320",
         15174 => x"436f6e66",
         15175 => x"69677572",
         15176 => x"6174696f",
         15177 => x"6e000000",
         15178 => x"3a0a4465",
         15179 => x"76696365",
         15180 => x"7320696d",
         15181 => x"706c656d",
         15182 => x"656e7465",
         15183 => x"643a0000",
         15184 => x"41646472",
         15185 => x"65737365",
         15186 => x"733a0000",
         15187 => x"20202020",
         15188 => x"43505520",
         15189 => x"52657365",
         15190 => x"74205665",
         15191 => x"63746f72",
         15192 => x"20416464",
         15193 => x"72657373",
         15194 => x"203d2025",
         15195 => x"3038580a",
         15196 => x"00000000",
         15197 => x"20202020",
         15198 => x"43505520",
         15199 => x"4d656d6f",
         15200 => x"72792053",
         15201 => x"74617274",
         15202 => x"20416464",
         15203 => x"72657373",
         15204 => x"203d2025",
         15205 => x"3038580a",
         15206 => x"00000000",
         15207 => x"20202020",
         15208 => x"53746163",
         15209 => x"6b205374",
         15210 => x"61727420",
         15211 => x"41646472",
         15212 => x"65737320",
         15213 => x"20202020",
         15214 => x"203d2025",
         15215 => x"3038580a",
         15216 => x"00000000",
         15217 => x"4d697363",
         15218 => x"3a000000",
         15219 => x"20202020",
         15220 => x"5a505520",
         15221 => x"49642020",
         15222 => x"20202020",
         15223 => x"20202020",
         15224 => x"20202020",
         15225 => x"20202020",
         15226 => x"203d2025",
         15227 => x"3034580a",
         15228 => x"00000000",
         15229 => x"20202020",
         15230 => x"53797374",
         15231 => x"656d2043",
         15232 => x"6c6f636b",
         15233 => x"20467265",
         15234 => x"71202020",
         15235 => x"20202020",
         15236 => x"203d2025",
         15237 => x"642e2530",
         15238 => x"34644d48",
         15239 => x"7a0a0000",
         15240 => x"20202020",
         15241 => x"57697368",
         15242 => x"626f6e65",
         15243 => x"20534452",
         15244 => x"414d2043",
         15245 => x"6c6f636b",
         15246 => x"20467265",
         15247 => x"713d2025",
         15248 => x"642e2530",
         15249 => x"34644d48",
         15250 => x"7a0a0000",
         15251 => x"20202020",
         15252 => x"53445241",
         15253 => x"4d20436c",
         15254 => x"6f636b20",
         15255 => x"46726571",
         15256 => x"20202020",
         15257 => x"20202020",
         15258 => x"203d2025",
         15259 => x"642e2530",
         15260 => x"34644d48",
         15261 => x"7a0a0000",
         15262 => x"20202020",
         15263 => x"53504900",
         15264 => x"20202020",
         15265 => x"50533200",
         15266 => x"20202020",
         15267 => x"494f4354",
         15268 => x"4c000000",
         15269 => x"20202020",
         15270 => x"57422049",
         15271 => x"32430000",
         15272 => x"20202020",
         15273 => x"57495348",
         15274 => x"424f4e45",
         15275 => x"20425553",
         15276 => x"00000000",
         15277 => x"20202020",
         15278 => x"494e5452",
         15279 => x"20435452",
         15280 => x"4c202843",
         15281 => x"68616e6e",
         15282 => x"656c733d",
         15283 => x"25303264",
         15284 => x"292e0a00",
         15285 => x"20202020",
         15286 => x"54494d45",
         15287 => x"52312020",
         15288 => x"20202854",
         15289 => x"696d6572",
         15290 => x"7320203d",
         15291 => x"25303264",
         15292 => x"292e0a00",
         15293 => x"20202020",
         15294 => x"53442043",
         15295 => x"41524420",
         15296 => x"20202844",
         15297 => x"65766963",
         15298 => x"6573203d",
         15299 => x"25303264",
         15300 => x"292e0a00",
         15301 => x"20202020",
         15302 => x"52414d20",
         15303 => x"20202020",
         15304 => x"20202825",
         15305 => x"3038583a",
         15306 => x"25303858",
         15307 => x"292e0a00",
         15308 => x"20202020",
         15309 => x"4252414d",
         15310 => x"20202020",
         15311 => x"20202825",
         15312 => x"3038583a",
         15313 => x"25303858",
         15314 => x"292e0a00",
         15315 => x"20202020",
         15316 => x"494e534e",
         15317 => x"20425241",
         15318 => x"4d202825",
         15319 => x"3038583a",
         15320 => x"25303858",
         15321 => x"292e0a00",
         15322 => x"20202020",
         15323 => x"53445241",
         15324 => x"4d202020",
         15325 => x"20202825",
         15326 => x"3038583a",
         15327 => x"25303858",
         15328 => x"292e0a00",
         15329 => x"20202020",
         15330 => x"57422053",
         15331 => x"4452414d",
         15332 => x"20202825",
         15333 => x"3038583a",
         15334 => x"25303858",
         15335 => x"292e0a00",
         15336 => x"20286672",
         15337 => x"6f6d2053",
         15338 => x"6f432063",
         15339 => x"6f6e6669",
         15340 => x"67290000",
         15341 => x"556e6b6e",
         15342 => x"6f776e00",
         15343 => x"45564f6d",
         15344 => x"00000000",
         15345 => x"536d616c",
         15346 => x"6c000000",
         15347 => x"4d656469",
         15348 => x"756d0000",
         15349 => x"466c6578",
         15350 => x"00000000",
         15351 => x"45564f00",
         15352 => x"0000f13c",
         15353 => x"01000000",
         15354 => x"00000002",
         15355 => x"0000f138",
         15356 => x"01000000",
         15357 => x"00000003",
         15358 => x"0000f134",
         15359 => x"01000000",
         15360 => x"00000004",
         15361 => x"0000f130",
         15362 => x"01000000",
         15363 => x"00000005",
         15364 => x"0000f12c",
         15365 => x"01000000",
         15366 => x"00000006",
         15367 => x"0000f128",
         15368 => x"01000000",
         15369 => x"00000007",
         15370 => x"0000f124",
         15371 => x"01000000",
         15372 => x"00000001",
         15373 => x"0000f120",
         15374 => x"01000000",
         15375 => x"00000008",
         15376 => x"0000f11c",
         15377 => x"01000000",
         15378 => x"0000000b",
         15379 => x"0000f118",
         15380 => x"01000000",
         15381 => x"00000009",
         15382 => x"0000f114",
         15383 => x"01000000",
         15384 => x"0000000a",
         15385 => x"0000f110",
         15386 => x"04000000",
         15387 => x"0000000d",
         15388 => x"0000f10c",
         15389 => x"04000000",
         15390 => x"0000000c",
         15391 => x"0000f108",
         15392 => x"04000000",
         15393 => x"0000000e",
         15394 => x"0000f104",
         15395 => x"03000000",
         15396 => x"0000000f",
         15397 => x"0000f100",
         15398 => x"04000000",
         15399 => x"0000000f",
         15400 => x"0000f0fc",
         15401 => x"04000000",
         15402 => x"00000010",
         15403 => x"0000f0f8",
         15404 => x"04000000",
         15405 => x"00000011",
         15406 => x"0000f0f4",
         15407 => x"03000000",
         15408 => x"00000012",
         15409 => x"0000f0f0",
         15410 => x"03000000",
         15411 => x"00000013",
         15412 => x"0000f0ec",
         15413 => x"03000000",
         15414 => x"00000014",
         15415 => x"0000f0e8",
         15416 => x"03000000",
         15417 => x"00000015",
         15418 => x"1b5b4400",
         15419 => x"1b5b4300",
         15420 => x"1b5b4200",
         15421 => x"1b5b4100",
         15422 => x"1b5b367e",
         15423 => x"1b5b357e",
         15424 => x"1b5b347e",
         15425 => x"1b304600",
         15426 => x"1b5b337e",
         15427 => x"1b5b327e",
         15428 => x"1b5b317e",
         15429 => x"10000000",
         15430 => x"0e000000",
         15431 => x"0d000000",
         15432 => x"0b000000",
         15433 => x"08000000",
         15434 => x"06000000",
         15435 => x"05000000",
         15436 => x"04000000",
         15437 => x"03000000",
         15438 => x"02000000",
         15439 => x"01000000",
         15440 => x"48697374",
         15441 => x"6f727920",
         15442 => x"68656170",
         15443 => x"3a253038",
         15444 => x"6c780a00",
         15445 => x"43616e6e",
         15446 => x"6f74206f",
         15447 => x"70656e2f",
         15448 => x"63726561",
         15449 => x"74652068",
         15450 => x"6973746f",
         15451 => x"72792066",
         15452 => x"696c652c",
         15453 => x"20646973",
         15454 => x"61626c69",
         15455 => x"6e672e00",
         15456 => x"68697374",
         15457 => x"6f727900",
         15458 => x"68697374",
         15459 => x"00000000",
         15460 => x"21000000",
         15461 => x"48697374",
         15462 => x"6f727920",
         15463 => x"62756666",
         15464 => x"65724025",
         15465 => x"30386c78",
         15466 => x"0a000000",
         15467 => x"2530366c",
         15468 => x"75202025",
         15469 => x"730a0000",
         15470 => x"4661696c",
         15471 => x"65642074",
         15472 => x"6f207265",
         15473 => x"73657420",
         15474 => x"74686520",
         15475 => x"68697374",
         15476 => x"6f727920",
         15477 => x"66696c65",
         15478 => x"20746f20",
         15479 => x"454f462e",
         15480 => x"00000000",
         15481 => x"3e25730a",
         15482 => x"00000000",
         15483 => x"1b5b317e",
         15484 => x"00000000",
         15485 => x"1b5b4100",
         15486 => x"1b5b4200",
         15487 => x"1b5b4300",
         15488 => x"1b5b4400",
         15489 => x"1b5b3130",
         15490 => x"7e000000",
         15491 => x"1b5b3131",
         15492 => x"7e000000",
         15493 => x"1b5b3132",
         15494 => x"7e000000",
         15495 => x"1b5b3133",
         15496 => x"7e000000",
         15497 => x"1b5b3134",
         15498 => x"7e000000",
         15499 => x"1b5b3135",
         15500 => x"7e000000",
         15501 => x"1b5b3137",
         15502 => x"7e000000",
         15503 => x"1b5b3138",
         15504 => x"7e000000",
         15505 => x"1b5b3139",
         15506 => x"7e000000",
         15507 => x"1b5b3230",
         15508 => x"7e000000",
         15509 => x"1b5b327e",
         15510 => x"00000000",
         15511 => x"1b5b337e",
         15512 => x"00000000",
         15513 => x"1b5b4600",
         15514 => x"1b5b357e",
         15515 => x"00000000",
         15516 => x"1b5b367e",
         15517 => x"00000000",
         15518 => x"583a2564",
         15519 => x"2c25642c",
         15520 => x"25642c25",
         15521 => x"642c2564",
         15522 => x"2c25643a",
         15523 => x"25303278",
         15524 => x"00000000",
         15525 => x"443a2564",
         15526 => x"2d25642d",
         15527 => x"25643a25",
         15528 => x"633a2564",
         15529 => x"2c25642c",
         15530 => x"25643a00",
         15531 => x"25642c00",
         15532 => x"4b3a2564",
         15533 => x"3a000000",
         15534 => x"25303278",
         15535 => x"2c000000",
         15536 => x"25635b25",
         15537 => x"643b2564",
         15538 => x"52000000",
         15539 => x"5265706f",
         15540 => x"72742043",
         15541 => x"7572736f",
         15542 => x"723a0000",
         15543 => x"55703a25",
         15544 => x"30327820",
         15545 => x"25303278",
         15546 => x"00000000",
         15547 => x"44773a25",
         15548 => x"30327820",
         15549 => x"25303278",
         15550 => x"00000000",
         15551 => x"48643a25",
         15552 => x"30327820",
         15553 => x"00000000",
         15554 => x"4e6f2074",
         15555 => x"65737420",
         15556 => x"64656669",
         15557 => x"6e65642e",
         15558 => x"00000000",
         15559 => x"53440000",
         15560 => x"222a3a3c",
         15561 => x"3e3f7c7f",
         15562 => x"00000000",
         15563 => x"2b2c3b3d",
         15564 => x"5b5d0000",
         15565 => x"46415400",
         15566 => x"46415433",
         15567 => x"32000000",
         15568 => x"ebfe904d",
         15569 => x"53444f53",
         15570 => x"352e3000",
         15571 => x"4e4f204e",
         15572 => x"414d4520",
         15573 => x"20202046",
         15574 => x"41542020",
         15575 => x"20202000",
         15576 => x"4e4f204e",
         15577 => x"414d4520",
         15578 => x"20202046",
         15579 => x"41543332",
         15580 => x"20202000",
         15581 => x"0000f31c",
         15582 => x"00000000",
         15583 => x"00000000",
         15584 => x"00000000",
         15585 => x"01030507",
         15586 => x"090e1012",
         15587 => x"1416181c",
         15588 => x"1e000000",
         15589 => x"809a4541",
         15590 => x"8e418f80",
         15591 => x"45454549",
         15592 => x"49498e8f",
         15593 => x"9092924f",
         15594 => x"994f5555",
         15595 => x"59999a9b",
         15596 => x"9c9d9e9f",
         15597 => x"41494f55",
         15598 => x"a5a5a6a7",
         15599 => x"a8a9aaab",
         15600 => x"acadaeaf",
         15601 => x"b0b1b2b3",
         15602 => x"b4b5b6b7",
         15603 => x"b8b9babb",
         15604 => x"bcbdbebf",
         15605 => x"c0c1c2c3",
         15606 => x"c4c5c6c7",
         15607 => x"c8c9cacb",
         15608 => x"cccdcecf",
         15609 => x"d0d1d2d3",
         15610 => x"d4d5d6d7",
         15611 => x"d8d9dadb",
         15612 => x"dcdddedf",
         15613 => x"e0e1e2e3",
         15614 => x"e4e5e6e7",
         15615 => x"e8e9eaeb",
         15616 => x"ecedeeef",
         15617 => x"f0f1f2f3",
         15618 => x"f4f5f6f7",
         15619 => x"f8f9fafb",
         15620 => x"fcfdfeff",
         15621 => x"2b2e2c3b",
         15622 => x"3d5b5d2f",
         15623 => x"5c222a3a",
         15624 => x"3c3e3f7c",
         15625 => x"7f000000",
         15626 => x"00010004",
         15627 => x"00100040",
         15628 => x"01000200",
         15629 => x"00000000",
         15630 => x"00010002",
         15631 => x"00040008",
         15632 => x"00100020",
         15633 => x"00000000",
         15634 => x"00c700fc",
         15635 => x"00e900e2",
         15636 => x"00e400e0",
         15637 => x"00e500e7",
         15638 => x"00ea00eb",
         15639 => x"00e800ef",
         15640 => x"00ee00ec",
         15641 => x"00c400c5",
         15642 => x"00c900e6",
         15643 => x"00c600f4",
         15644 => x"00f600f2",
         15645 => x"00fb00f9",
         15646 => x"00ff00d6",
         15647 => x"00dc00a2",
         15648 => x"00a300a5",
         15649 => x"20a70192",
         15650 => x"00e100ed",
         15651 => x"00f300fa",
         15652 => x"00f100d1",
         15653 => x"00aa00ba",
         15654 => x"00bf2310",
         15655 => x"00ac00bd",
         15656 => x"00bc00a1",
         15657 => x"00ab00bb",
         15658 => x"25912592",
         15659 => x"25932502",
         15660 => x"25242561",
         15661 => x"25622556",
         15662 => x"25552563",
         15663 => x"25512557",
         15664 => x"255d255c",
         15665 => x"255b2510",
         15666 => x"25142534",
         15667 => x"252c251c",
         15668 => x"2500253c",
         15669 => x"255e255f",
         15670 => x"255a2554",
         15671 => x"25692566",
         15672 => x"25602550",
         15673 => x"256c2567",
         15674 => x"25682564",
         15675 => x"25652559",
         15676 => x"25582552",
         15677 => x"2553256b",
         15678 => x"256a2518",
         15679 => x"250c2588",
         15680 => x"2584258c",
         15681 => x"25902580",
         15682 => x"03b100df",
         15683 => x"039303c0",
         15684 => x"03a303c3",
         15685 => x"00b503c4",
         15686 => x"03a60398",
         15687 => x"03a903b4",
         15688 => x"221e03c6",
         15689 => x"03b52229",
         15690 => x"226100b1",
         15691 => x"22652264",
         15692 => x"23202321",
         15693 => x"00f72248",
         15694 => x"00b02219",
         15695 => x"00b7221a",
         15696 => x"207f00b2",
         15697 => x"25a000a0",
         15698 => x"0061031a",
         15699 => x"00e00317",
         15700 => x"00f80307",
         15701 => x"00ff0001",
         15702 => x"01780100",
         15703 => x"01300132",
         15704 => x"01060139",
         15705 => x"0110014a",
         15706 => x"012e0179",
         15707 => x"01060180",
         15708 => x"004d0243",
         15709 => x"01810182",
         15710 => x"01820184",
         15711 => x"01840186",
         15712 => x"01870187",
         15713 => x"0189018a",
         15714 => x"018b018b",
         15715 => x"018d018e",
         15716 => x"018f0190",
         15717 => x"01910191",
         15718 => x"01930194",
         15719 => x"01f60196",
         15720 => x"01970198",
         15721 => x"0198023d",
         15722 => x"019b019c",
         15723 => x"019d0220",
         15724 => x"019f01a0",
         15725 => x"01a001a2",
         15726 => x"01a201a4",
         15727 => x"01a401a6",
         15728 => x"01a701a7",
         15729 => x"01a901aa",
         15730 => x"01ab01ac",
         15731 => x"01ac01ae",
         15732 => x"01af01af",
         15733 => x"01b101b2",
         15734 => x"01b301b3",
         15735 => x"01b501b5",
         15736 => x"01b701b8",
         15737 => x"01b801ba",
         15738 => x"01bb01bc",
         15739 => x"01bc01be",
         15740 => x"01f701c0",
         15741 => x"01c101c2",
         15742 => x"01c301c4",
         15743 => x"01c501c4",
         15744 => x"01c701c8",
         15745 => x"01c701ca",
         15746 => x"01cb01ca",
         15747 => x"01cd0110",
         15748 => x"01dd0001",
         15749 => x"018e01de",
         15750 => x"011201f3",
         15751 => x"000301f1",
         15752 => x"01f401f4",
         15753 => x"01f80128",
         15754 => x"02220112",
         15755 => x"023a0009",
         15756 => x"2c65023b",
         15757 => x"023b023d",
         15758 => x"2c66023f",
         15759 => x"02400241",
         15760 => x"02410246",
         15761 => x"010a0253",
         15762 => x"00400181",
         15763 => x"01860255",
         15764 => x"0189018a",
         15765 => x"0258018f",
         15766 => x"025a0190",
         15767 => x"025c025d",
         15768 => x"025e025f",
         15769 => x"01930261",
         15770 => x"02620194",
         15771 => x"02640265",
         15772 => x"02660267",
         15773 => x"01970196",
         15774 => x"026a2c62",
         15775 => x"026c026d",
         15776 => x"026e019c",
         15777 => x"02700271",
         15778 => x"019d0273",
         15779 => x"0274019f",
         15780 => x"02760277",
         15781 => x"02780279",
         15782 => x"027a027b",
         15783 => x"027c2c64",
         15784 => x"027e027f",
         15785 => x"01a60281",
         15786 => x"028201a9",
         15787 => x"02840285",
         15788 => x"02860287",
         15789 => x"01ae0244",
         15790 => x"01b101b2",
         15791 => x"0245028d",
         15792 => x"028e028f",
         15793 => x"02900291",
         15794 => x"01b7037b",
         15795 => x"000303fd",
         15796 => x"03fe03ff",
         15797 => x"03ac0004",
         15798 => x"03860388",
         15799 => x"0389038a",
         15800 => x"03b10311",
         15801 => x"03c20002",
         15802 => x"03a303a3",
         15803 => x"03c40308",
         15804 => x"03cc0003",
         15805 => x"038c038e",
         15806 => x"038f03d8",
         15807 => x"011803f2",
         15808 => x"000a03f9",
         15809 => x"03f303f4",
         15810 => x"03f503f6",
         15811 => x"03f703f7",
         15812 => x"03f903fa",
         15813 => x"03fa0430",
         15814 => x"03200450",
         15815 => x"07100460",
         15816 => x"0122048a",
         15817 => x"013604c1",
         15818 => x"010e04cf",
         15819 => x"000104c0",
         15820 => x"04d00144",
         15821 => x"05610426",
         15822 => x"00000000",
         15823 => x"1d7d0001",
         15824 => x"2c631e00",
         15825 => x"01961ea0",
         15826 => x"015a1f00",
         15827 => x"06081f10",
         15828 => x"06061f20",
         15829 => x"06081f30",
         15830 => x"06081f40",
         15831 => x"06061f51",
         15832 => x"00071f59",
         15833 => x"1f521f5b",
         15834 => x"1f541f5d",
         15835 => x"1f561f5f",
         15836 => x"1f600608",
         15837 => x"1f70000e",
         15838 => x"1fba1fbb",
         15839 => x"1fc81fc9",
         15840 => x"1fca1fcb",
         15841 => x"1fda1fdb",
         15842 => x"1ff81ff9",
         15843 => x"1fea1feb",
         15844 => x"1ffa1ffb",
         15845 => x"1f800608",
         15846 => x"1f900608",
         15847 => x"1fa00608",
         15848 => x"1fb00004",
         15849 => x"1fb81fb9",
         15850 => x"1fb21fbc",
         15851 => x"1fcc0001",
         15852 => x"1fc31fd0",
         15853 => x"06021fe0",
         15854 => x"06021fe5",
         15855 => x"00011fec",
         15856 => x"1ff30001",
         15857 => x"1ffc214e",
         15858 => x"00012132",
         15859 => x"21700210",
         15860 => x"21840001",
         15861 => x"218324d0",
         15862 => x"051a2c30",
         15863 => x"042f2c60",
         15864 => x"01022c67",
         15865 => x"01062c75",
         15866 => x"01022c80",
         15867 => x"01642d00",
         15868 => x"0826ff41",
         15869 => x"031a0000",
         15870 => x"00000000",
         15871 => x"0000e6f8",
         15872 => x"01020100",
         15873 => x"00000000",
         15874 => x"00000000",
         15875 => x"0000e700",
         15876 => x"01040100",
         15877 => x"00000000",
         15878 => x"00000000",
         15879 => x"0000e708",
         15880 => x"01140300",
         15881 => x"00000000",
         15882 => x"00000000",
         15883 => x"0000e710",
         15884 => x"012b0300",
         15885 => x"00000000",
         15886 => x"00000000",
         15887 => x"0000e718",
         15888 => x"01300300",
         15889 => x"00000000",
         15890 => x"00000000",
         15891 => x"0000e720",
         15892 => x"013c0400",
         15893 => x"00000000",
         15894 => x"00000000",
         15895 => x"0000e728",
         15896 => x"013d0400",
         15897 => x"00000000",
         15898 => x"00000000",
         15899 => x"0000e730",
         15900 => x"013f0400",
         15901 => x"00000000",
         15902 => x"00000000",
         15903 => x"0000e738",
         15904 => x"01400400",
         15905 => x"00000000",
         15906 => x"00000000",
         15907 => x"0000e740",
         15908 => x"01410400",
         15909 => x"00000000",
         15910 => x"00000000",
         15911 => x"0000e744",
         15912 => x"01420400",
         15913 => x"00000000",
         15914 => x"00000000",
         15915 => x"0000e748",
         15916 => x"01430400",
         15917 => x"00000000",
         15918 => x"00000000",
         15919 => x"0000e74c",
         15920 => x"01500500",
         15921 => x"00000000",
         15922 => x"00000000",
         15923 => x"0000e750",
         15924 => x"01510500",
         15925 => x"00000000",
         15926 => x"00000000",
         15927 => x"0000e754",
         15928 => x"01540500",
         15929 => x"00000000",
         15930 => x"00000000",
         15931 => x"0000e758",
         15932 => x"01550500",
         15933 => x"00000000",
         15934 => x"00000000",
         15935 => x"0000e75c",
         15936 => x"01790700",
         15937 => x"00000000",
         15938 => x"00000000",
         15939 => x"0000e764",
         15940 => x"01780700",
         15941 => x"00000000",
         15942 => x"00000000",
         15943 => x"0000e768",
         15944 => x"01820800",
         15945 => x"00000000",
         15946 => x"00000000",
         15947 => x"0000e770",
         15948 => x"01830800",
         15949 => x"00000000",
         15950 => x"00000000",
         15951 => x"0000e778",
         15952 => x"01850800",
         15953 => x"00000000",
         15954 => x"00000000",
         15955 => x"0000e780",
         15956 => x"01870800",
         15957 => x"00000000",
         15958 => x"00000000",
         15959 => x"0000e788",
         15960 => x"01880800",
         15961 => x"00000000",
         15962 => x"00000000",
         15963 => x"0000e78c",
         15964 => x"01890800",
         15965 => x"00000000",
         15966 => x"00000000",
         15967 => x"0000e790",
         15968 => x"018c0900",
         15969 => x"00000000",
         15970 => x"00000000",
         15971 => x"0000e798",
         15972 => x"018d0900",
         15973 => x"00000000",
         15974 => x"00000000",
         15975 => x"0000e7a0",
         15976 => x"018e0900",
         15977 => x"00000000",
         15978 => x"00000000",
         15979 => x"0000e7a8",
         15980 => x"018f0900",
         15981 => x"00000000",
         15982 => x"00000000",
         15983 => x"00000000",
         15984 => x"00000000",
         15985 => x"00007fff",
         15986 => x"00000000",
         15987 => x"00007fff",
         15988 => x"00010000",
         15989 => x"00007fff",
         15990 => x"00010000",
         15991 => x"00810000",
         15992 => x"01000000",
         15993 => x"017fffff",
         15994 => x"00000000",
         15995 => x"00000000",
         15996 => x"00007800",
         15997 => x"00000000",
         15998 => x"05f5e100",
         15999 => x"05f5e100",
         16000 => x"05f5e100",
         16001 => x"00000000",
         16002 => x"01010101",
         16003 => x"01010101",
         16004 => x"01011001",
         16005 => x"01000000",
         16006 => x"00000000",
         16007 => x"00000000",
         16008 => x"00000000",
         16009 => x"00000000",
         16010 => x"00000000",
         16011 => x"00000000",
         16012 => x"00000000",
         16013 => x"00000000",
         16014 => x"00000000",
         16015 => x"00000000",
         16016 => x"00000000",
         16017 => x"00000000",
         16018 => x"00000000",
         16019 => x"00000000",
         16020 => x"00000000",
         16021 => x"00000000",
         16022 => x"00000000",
         16023 => x"00000000",
         16024 => x"00000000",
         16025 => x"00000000",
         16026 => x"00000000",
         16027 => x"00000000",
         16028 => x"00000000",
         16029 => x"00000000",
         16030 => x"0000f180",
         16031 => x"01000000",
         16032 => x"0000f188",
         16033 => x"01000000",
         16034 => x"0000f190",
         16035 => x"02000000",
         16036 => x"0001fd80",
         16037 => x"1bfc5ffd",
         16038 => x"f03b3a0d",
         16039 => x"797a405b",
         16040 => x"5df0f0f0",
         16041 => x"71727374",
         16042 => x"75767778",
         16043 => x"696a6b6c",
         16044 => x"6d6e6f70",
         16045 => x"61626364",
         16046 => x"65666768",
         16047 => x"31323334",
         16048 => x"35363738",
         16049 => x"5cf32d20",
         16050 => x"30392c2e",
         16051 => x"f67ff3f4",
         16052 => x"f1f23f2f",
         16053 => x"08f0f0f0",
         16054 => x"f0f0f0f0",
         16055 => x"80818283",
         16056 => x"84f0f0f0",
         16057 => x"1bfc58fd",
         16058 => x"f03a3b0d",
         16059 => x"595a405b",
         16060 => x"5df0f0f0",
         16061 => x"51525354",
         16062 => x"55565758",
         16063 => x"494a4b4c",
         16064 => x"4d4e4f50",
         16065 => x"41424344",
         16066 => x"45464748",
         16067 => x"31323334",
         16068 => x"35363738",
         16069 => x"5cf32d20",
         16070 => x"30392c2e",
         16071 => x"f67ff3f4",
         16072 => x"f1f23f2f",
         16073 => x"08f0f0f0",
         16074 => x"f0f0f0f0",
         16075 => x"80818283",
         16076 => x"84f0f0f0",
         16077 => x"1bfc58fd",
         16078 => x"f02b2a0d",
         16079 => x"595a607b",
         16080 => x"7df0f0f0",
         16081 => x"51525354",
         16082 => x"55565758",
         16083 => x"494a4b4c",
         16084 => x"4d4e4f50",
         16085 => x"41424344",
         16086 => x"45464748",
         16087 => x"21222324",
         16088 => x"25262728",
         16089 => x"7c7e3d20",
         16090 => x"20293c3e",
         16091 => x"f7e2e0e1",
         16092 => x"f9f83f2f",
         16093 => x"fbf0f0f0",
         16094 => x"f0f0f0f0",
         16095 => x"85868788",
         16096 => x"89f0f0f0",
         16097 => x"1bfe1efa",
         16098 => x"f0f0f0f0",
         16099 => x"191a001b",
         16100 => x"1df0f0f0",
         16101 => x"11121314",
         16102 => x"15161718",
         16103 => x"090a0b0c",
         16104 => x"0d0e0f10",
         16105 => x"01020304",
         16106 => x"05060708",
         16107 => x"f0f0f0f0",
         16108 => x"f0f0f0f0",
         16109 => x"f01ef0f0",
         16110 => x"f01ff0f0",
         16111 => x"f0f0f0f0",
         16112 => x"f0f0f01c",
         16113 => x"f0f0f0f0",
         16114 => x"f0f0f0f0",
         16115 => x"80818283",
         16116 => x"84f0f0f0",
         16117 => x"bff0cfc9",
         16118 => x"f0b54dcd",
         16119 => x"3577d7b3",
         16120 => x"b7f0f0f0",
         16121 => x"7c704131",
         16122 => x"39a678dd",
         16123 => x"3d5d6c56",
         16124 => x"1d33d5b1",
         16125 => x"466ed948",
         16126 => x"74434c73",
         16127 => x"3f367e3b",
         16128 => x"7a1e5fa2",
         16129 => x"d39fd100",
         16130 => x"9da3d0b9",
         16131 => x"c6c5c2c1",
         16132 => x"c3c4bbbe",
         16133 => x"f0f0f0f0",
         16134 => x"f0f0f0f0",
         16135 => x"80818283",
         16136 => x"84f0f0f0",
         16137 => x"00000000",
         16138 => x"00000000",
         16139 => x"00000000",
         16140 => x"00000000",
         16141 => x"00000000",
         16142 => x"00000000",
         16143 => x"00000000",
         16144 => x"00000000",
         16145 => x"00000000",
         16146 => x"00000000",
         16147 => x"00000000",
         16148 => x"00000000",
         16149 => x"00000000",
         16150 => x"00000000",
         16151 => x"00000000",
         16152 => x"00000000",
         16153 => x"00000000",
         16154 => x"00000000",
         16155 => x"00000000",
         16156 => x"00000000",
         16157 => x"00000000",
         16158 => x"00000000",
         16159 => x"00000000",
         16160 => x"00000000",
         16161 => x"00000000",
         16162 => x"00010000",
         16163 => x"00000000",
         16164 => x"f8000000",
         16165 => x"0000f1ec",
         16166 => x"f3000000",
         16167 => x"0000f1f4",
         16168 => x"f4000000",
         16169 => x"0000f1f8",
         16170 => x"f1000000",
         16171 => x"0000f1fc",
         16172 => x"f2000000",
         16173 => x"0000f200",
         16174 => x"80000000",
         16175 => x"0000f204",
         16176 => x"81000000",
         16177 => x"0000f20c",
         16178 => x"82000000",
         16179 => x"0000f214",
         16180 => x"83000000",
         16181 => x"0000f21c",
         16182 => x"84000000",
         16183 => x"0000f224",
         16184 => x"85000000",
         16185 => x"0000f22c",
         16186 => x"86000000",
         16187 => x"0000f234",
         16188 => x"87000000",
         16189 => x"0000f23c",
         16190 => x"88000000",
         16191 => x"0000f244",
         16192 => x"89000000",
         16193 => x"0000f24c",
         16194 => x"f6000000",
         16195 => x"0000f254",
         16196 => x"7f000000",
         16197 => x"0000f25c",
         16198 => x"f9000000",
         16199 => x"0000f264",
         16200 => x"e0000000",
         16201 => x"0000f268",
         16202 => x"e1000000",
         16203 => x"0000f270",
         16204 => x"71000000",
         16205 => x"00000000",
         16206 => x"00000000",
         16207 => x"00000000",
         16208 => x"00000000",
         16209 => x"00000000",
         16210 => x"00000000",
         16211 => x"00000000",
         16212 => x"00000000",
         16213 => x"00000000",
         16214 => x"00000000",
         16215 => x"00000000",
         16216 => x"00000000",
         16217 => x"00000000",
         16218 => x"00000000",
         16219 => x"00000000",
         16220 => x"00000000",
         16221 => x"00000000",
         16222 => x"00000000",
         16223 => x"00000000",
         16224 => x"00000000",
         16225 => x"00000000",
         16226 => x"00000000",
         16227 => x"00000000",
         16228 => x"00000000",
         16229 => x"00000000",
         16230 => x"00000000",
         16231 => x"00000000",
         16232 => x"00000000",
         16233 => x"00000000",
         16234 => x"00000000",
         16235 => x"00000000",
         16236 => x"00000000",
         16237 => x"00000000",
         16238 => x"00000000",
         16239 => x"00000000",
         16240 => x"00000000",
         16241 => x"00000000",
         16242 => x"00000000",
         16243 => x"00000000",
         16244 => x"00000000",
         16245 => x"00000000",
         16246 => x"00000000",
         16247 => x"00000000",
         16248 => x"00000000",
         16249 => x"00000000",
         16250 => x"00000000",
         16251 => x"00000000",
         16252 => x"00000000",
         16253 => x"00000000",
         16254 => x"00000000",
         16255 => x"00000000",
         16256 => x"00000000",
         16257 => x"00000000",
         16258 => x"00000000",
         16259 => x"00000000",
         16260 => x"00000000",
         16261 => x"00000000",
         16262 => x"00000000",
         16263 => x"00000000",
         16264 => x"00000000",
         16265 => x"00000000",
         16266 => x"00000000",
         16267 => x"00000000",
         16268 => x"00000000",
         16269 => x"00000000",
         16270 => x"00000000",
         16271 => x"00000000",
         16272 => x"00000000",
         16273 => x"00000000",
         16274 => x"00000000",
         16275 => x"00000000",
         16276 => x"00000000",
         16277 => x"00000000",
         16278 => x"00000000",
         16279 => x"00000000",
         16280 => x"00000000",
         16281 => x"00000000",
         16282 => x"00000000",
         16283 => x"00000000",
         16284 => x"00000000",
         16285 => x"00000000",
         16286 => x"00000000",
         16287 => x"00000000",
         16288 => x"00000000",
         16289 => x"00000000",
         16290 => x"00000000",
         16291 => x"00000000",
         16292 => x"00000000",
         16293 => x"00000000",
         16294 => x"00000000",
         16295 => x"00000000",
         16296 => x"00000000",
         16297 => x"00000000",
         16298 => x"00000000",
         16299 => x"00000000",
         16300 => x"00000000",
         16301 => x"00000000",
         16302 => x"00000000",
         16303 => x"00000000",
         16304 => x"00000000",
         16305 => x"00000000",
         16306 => x"00000000",
         16307 => x"00000000",
         16308 => x"00000000",
         16309 => x"00000000",
         16310 => x"00000000",
         16311 => x"00000000",
         16312 => x"00000000",
         16313 => x"00000000",
         16314 => x"00000000",
         16315 => x"00000000",
         16316 => x"00000000",
         16317 => x"00000000",
         16318 => x"00000000",
         16319 => x"00000000",
         16320 => x"00000000",
         16321 => x"00000000",
         16322 => x"00000000",
         16323 => x"00000000",
         16324 => x"00000000",
         16325 => x"00000000",
         16326 => x"00000000",
         16327 => x"00000000",
         16328 => x"00000000",
         16329 => x"00000000",
         16330 => x"00000000",
         16331 => x"00000000",
         16332 => x"00000000",
         16333 => x"00000000",
         16334 => x"00000000",
         16335 => x"00000000",
         16336 => x"00000000",
         16337 => x"00000000",
         16338 => x"00000000",
         16339 => x"00000000",
         16340 => x"00000000",
         16341 => x"00000000",
         16342 => x"00000000",
         16343 => x"00000000",
         16344 => x"00000000",
         16345 => x"00000000",
         16346 => x"00000000",
         16347 => x"00000000",
         16348 => x"00000000",
         16349 => x"00000000",
         16350 => x"00000000",
         16351 => x"00000000",
         16352 => x"00000000",
         16353 => x"00000000",
         16354 => x"00000000",
         16355 => x"00000000",
         16356 => x"00000000",
         16357 => x"00000000",
         16358 => x"00000000",
         16359 => x"00000000",
         16360 => x"00000000",
         16361 => x"00000000",
         16362 => x"00000000",
         16363 => x"00000000",
         16364 => x"00000000",
         16365 => x"00000000",
         16366 => x"00000000",
         16367 => x"00000000",
         16368 => x"00000000",
         16369 => x"00000000",
         16370 => x"00000000",
         16371 => x"00000000",
         16372 => x"00000000",
         16373 => x"00000000",
         16374 => x"00000000",
         16375 => x"00000000",
         16376 => x"00000000",
         16377 => x"00000000",
         16378 => x"00000000",
         16379 => x"00000000",
         16380 => x"00000000",
         16381 => x"00000000",
         16382 => x"00000000",
         16383 => x"00000000",
         16384 => x"00000000",
         16385 => x"00000000",
         16386 => x"00000000",
         16387 => x"00000000",
         16388 => x"00000000",
         16389 => x"00000000",
         16390 => x"00000000",
         16391 => x"00000000",
         16392 => x"00000000",
         16393 => x"00000000",
         16394 => x"00000000",
         16395 => x"00000000",
         16396 => x"00000000",
         16397 => x"00000000",
         16398 => x"00000000",
         16399 => x"00000000",
         16400 => x"00000000",
         16401 => x"00000000",
         16402 => x"00000000",
         16403 => x"00000000",
         16404 => x"00000000",
         16405 => x"00000000",
         16406 => x"00000000",
         16407 => x"00000000",
         16408 => x"00000000",
         16409 => x"00000000",
         16410 => x"00000000",
         16411 => x"00000000",
         16412 => x"00000000",
         16413 => x"00000000",
         16414 => x"00000000",
         16415 => x"00000000",
         16416 => x"00000000",
         16417 => x"00000000",
         16418 => x"00000000",
         16419 => x"00000000",
         16420 => x"00000000",
         16421 => x"00000000",
         16422 => x"00000000",
         16423 => x"00000000",
         16424 => x"00000000",
         16425 => x"00000000",
         16426 => x"00000000",
         16427 => x"00000000",
         16428 => x"00000000",
         16429 => x"00000000",
         16430 => x"00000000",
         16431 => x"00000000",
         16432 => x"00000000",
         16433 => x"00000000",
         16434 => x"00000000",
         16435 => x"00000000",
         16436 => x"00000000",
         16437 => x"00000000",
         16438 => x"00000000",
         16439 => x"00000000",
         16440 => x"00000000",
         16441 => x"00000000",
         16442 => x"00000000",
         16443 => x"00000000",
         16444 => x"00000000",
         16445 => x"00000000",
         16446 => x"00000000",
         16447 => x"00000000",
         16448 => x"00000000",
         16449 => x"00000000",
         16450 => x"00000000",
         16451 => x"00000000",
         16452 => x"00000000",
         16453 => x"00000000",
         16454 => x"00000000",
         16455 => x"00000000",
         16456 => x"00000000",
         16457 => x"00000000",
         16458 => x"00000000",
         16459 => x"00000000",
         16460 => x"00000000",
         16461 => x"00000000",
         16462 => x"00000000",
         16463 => x"00000000",
         16464 => x"00000000",
         16465 => x"00000000",
         16466 => x"00000000",
         16467 => x"00000000",
         16468 => x"00000000",
         16469 => x"00000000",
         16470 => x"00000000",
         16471 => x"00000000",
         16472 => x"00000000",
         16473 => x"00000000",
         16474 => x"00000000",
         16475 => x"00000000",
         16476 => x"00000000",
         16477 => x"00000000",
         16478 => x"00000000",
         16479 => x"00000000",
         16480 => x"00000000",
         16481 => x"00000000",
         16482 => x"00000000",
         16483 => x"00000000",
         16484 => x"00000000",
         16485 => x"00000000",
         16486 => x"00000000",
         16487 => x"00000000",
         16488 => x"00000000",
         16489 => x"00000000",
         16490 => x"00000000",
         16491 => x"00000000",
         16492 => x"00000000",
         16493 => x"00000000",
         16494 => x"00000000",
         16495 => x"00000000",
         16496 => x"00000000",
         16497 => x"00000000",
         16498 => x"00000000",
         16499 => x"00000000",
         16500 => x"00000000",
         16501 => x"00000000",
         16502 => x"00000000",
         16503 => x"00000000",
         16504 => x"00000000",
         16505 => x"00000000",
         16506 => x"00000000",
         16507 => x"00000000",
         16508 => x"00000000",
         16509 => x"00000000",
         16510 => x"00000000",
         16511 => x"00000000",
         16512 => x"00000000",
         16513 => x"00000000",
         16514 => x"00000000",
         16515 => x"00000000",
         16516 => x"00000000",
         16517 => x"00000000",
         16518 => x"00000000",
         16519 => x"00000000",
         16520 => x"00000000",
         16521 => x"00000000",
         16522 => x"00000000",
         16523 => x"00000000",
         16524 => x"00000000",
         16525 => x"00000000",
         16526 => x"00000000",
         16527 => x"00000000",
         16528 => x"00000000",
         16529 => x"00000000",
         16530 => x"00000000",
         16531 => x"00000000",
         16532 => x"00000000",
         16533 => x"00000000",
         16534 => x"00000000",
         16535 => x"00000000",
         16536 => x"00000000",
         16537 => x"00000000",
         16538 => x"00000000",
         16539 => x"00000000",
         16540 => x"00000000",
         16541 => x"00000000",
         16542 => x"00000000",
         16543 => x"00000000",
         16544 => x"00000000",
         16545 => x"00000000",
         16546 => x"00000000",
         16547 => x"00000000",
         16548 => x"00000000",
         16549 => x"00000000",
         16550 => x"00000000",
         16551 => x"00000000",
         16552 => x"00000000",
         16553 => x"00000000",
         16554 => x"00000000",
         16555 => x"00000000",
         16556 => x"00000000",
         16557 => x"00000000",
         16558 => x"00000000",
         16559 => x"00000000",
         16560 => x"00000000",
         16561 => x"00000000",
         16562 => x"00000000",
         16563 => x"00000000",
         16564 => x"00000000",
         16565 => x"00000000",
         16566 => x"00000000",
         16567 => x"00000000",
         16568 => x"00000000",
         16569 => x"00000000",
         16570 => x"00000000",
         16571 => x"00000000",
         16572 => x"00000000",
         16573 => x"00000000",
         16574 => x"00000000",
         16575 => x"00000000",
         16576 => x"00000000",
         16577 => x"00000000",
         16578 => x"00000000",
         16579 => x"00000000",
         16580 => x"00000000",
         16581 => x"00000000",
         16582 => x"00000000",
         16583 => x"00000000",
         16584 => x"00000000",
         16585 => x"00000000",
         16586 => x"00000000",
         16587 => x"00000000",
         16588 => x"00000000",
         16589 => x"00000000",
         16590 => x"00000000",
         16591 => x"00000000",
         16592 => x"00000000",
         16593 => x"00000000",
         16594 => x"00000000",
         16595 => x"00000000",
         16596 => x"00000000",
         16597 => x"00000000",
         16598 => x"00000000",
         16599 => x"00000000",
         16600 => x"00000000",
         16601 => x"00000000",
         16602 => x"00000000",
         16603 => x"00000000",
         16604 => x"00000000",
         16605 => x"00000000",
         16606 => x"00000000",
         16607 => x"00000000",
         16608 => x"00000000",
         16609 => x"00000000",
         16610 => x"00000000",
         16611 => x"00000000",
         16612 => x"00000000",
         16613 => x"00000000",
         16614 => x"00000000",
         16615 => x"00000000",
         16616 => x"00000000",
         16617 => x"00000000",
         16618 => x"00000000",
         16619 => x"00000000",
         16620 => x"00000000",
         16621 => x"00000000",
         16622 => x"00000000",
         16623 => x"00000000",
         16624 => x"00000000",
         16625 => x"00000000",
         16626 => x"00000000",
         16627 => x"00000000",
         16628 => x"00000000",
         16629 => x"00000000",
         16630 => x"00000000",
         16631 => x"00000000",
         16632 => x"00000000",
         16633 => x"00000000",
         16634 => x"00000000",
         16635 => x"00000000",
         16636 => x"00000000",
         16637 => x"00000000",
         16638 => x"00000000",
         16639 => x"00000000",
         16640 => x"00000000",
         16641 => x"00000000",
         16642 => x"00000000",
         16643 => x"00000000",
         16644 => x"00000000",
         16645 => x"00000000",
         16646 => x"00000000",
         16647 => x"00000000",
         16648 => x"00000000",
         16649 => x"00000000",
         16650 => x"00000000",
         16651 => x"00000000",
         16652 => x"00000000",
         16653 => x"00000000",
         16654 => x"00000000",
         16655 => x"00000000",
         16656 => x"00000000",
         16657 => x"00000000",
         16658 => x"00000000",
         16659 => x"00000000",
         16660 => x"00000000",
         16661 => x"00000000",
         16662 => x"00000000",
         16663 => x"00000000",
         16664 => x"00000000",
         16665 => x"00000000",
         16666 => x"00000000",
         16667 => x"00000000",
         16668 => x"00000000",
         16669 => x"00000000",
         16670 => x"00000000",
         16671 => x"00000000",
         16672 => x"00000000",
         16673 => x"00000000",
         16674 => x"00000000",
         16675 => x"00000000",
         16676 => x"00000000",
         16677 => x"00000000",
         16678 => x"00000000",
         16679 => x"00000000",
         16680 => x"00000000",
         16681 => x"00000000",
         16682 => x"00000000",
         16683 => x"00000000",
         16684 => x"00000000",
         16685 => x"00000000",
         16686 => x"00000000",
         16687 => x"00000000",
         16688 => x"00000000",
         16689 => x"00000000",
         16690 => x"00000000",
         16691 => x"00000000",
         16692 => x"00000000",
         16693 => x"00000000",
         16694 => x"00000000",
         16695 => x"00000000",
         16696 => x"00000000",
         16697 => x"00000000",
         16698 => x"00000000",
         16699 => x"00000000",
         16700 => x"00000000",
         16701 => x"00000000",
         16702 => x"00000000",
         16703 => x"00000000",
         16704 => x"00000000",
         16705 => x"00000000",
         16706 => x"00000000",
         16707 => x"00000000",
         16708 => x"00000000",
         16709 => x"00000000",
         16710 => x"00000000",
         16711 => x"00000000",
         16712 => x"00000000",
         16713 => x"00000000",
         16714 => x"00000000",
         16715 => x"00000000",
         16716 => x"00000000",
         16717 => x"00000000",
         16718 => x"00000000",
         16719 => x"00000000",
         16720 => x"00000000",
         16721 => x"00000000",
         16722 => x"00000000",
         16723 => x"00000000",
         16724 => x"00000000",
         16725 => x"00000000",
         16726 => x"00000000",
         16727 => x"00000000",
         16728 => x"00000000",
         16729 => x"00000000",
         16730 => x"00000000",
         16731 => x"00000000",
         16732 => x"00000000",
         16733 => x"00000000",
         16734 => x"00000000",
         16735 => x"00000000",
         16736 => x"00000000",
         16737 => x"00000000",
         16738 => x"00000000",
         16739 => x"00000000",
         16740 => x"00000000",
         16741 => x"00000000",
         16742 => x"00000000",
         16743 => x"00000000",
         16744 => x"00000000",
         16745 => x"00000000",
         16746 => x"00000000",
         16747 => x"00000000",
         16748 => x"00000000",
         16749 => x"00000000",
         16750 => x"00000000",
         16751 => x"00000000",
         16752 => x"00000000",
         16753 => x"00000000",
         16754 => x"00000000",
         16755 => x"00000000",
         16756 => x"00000000",
         16757 => x"00000000",
         16758 => x"00000000",
         16759 => x"00000000",
         16760 => x"00000000",
         16761 => x"00000000",
         16762 => x"00000000",
         16763 => x"00000000",
         16764 => x"00000000",
         16765 => x"00000000",
         16766 => x"00000000",
         16767 => x"00000000",
         16768 => x"00000000",
         16769 => x"00000000",
         16770 => x"00000000",
         16771 => x"00000000",
         16772 => x"00000000",
         16773 => x"00000000",
         16774 => x"00000000",
         16775 => x"00000000",
         16776 => x"00000000",
         16777 => x"00000000",
         16778 => x"00000000",
         16779 => x"00000000",
         16780 => x"00000000",
         16781 => x"00000000",
         16782 => x"00000000",
         16783 => x"00000000",
         16784 => x"00000000",
         16785 => x"00000000",
         16786 => x"00000000",
         16787 => x"00000000",
         16788 => x"00000000",
         16789 => x"00000000",
         16790 => x"00000000",
         16791 => x"00000000",
         16792 => x"00000000",
         16793 => x"00000000",
         16794 => x"00000000",
         16795 => x"00000000",
         16796 => x"00000000",
         16797 => x"00000000",
         16798 => x"00000000",
         16799 => x"00000000",
         16800 => x"00000000",
         16801 => x"00000000",
         16802 => x"00000000",
         16803 => x"00000000",
         16804 => x"00000000",
         16805 => x"00000000",
         16806 => x"00000000",
         16807 => x"00000000",
         16808 => x"00000000",
         16809 => x"00000000",
         16810 => x"00000000",
         16811 => x"00000000",
         16812 => x"00000000",
         16813 => x"00000000",
         16814 => x"00000000",
         16815 => x"00000000",
         16816 => x"00000000",
         16817 => x"00000000",
         16818 => x"00000000",
         16819 => x"00000000",
         16820 => x"00000000",
         16821 => x"00000000",
         16822 => x"00000000",
         16823 => x"00000000",
         16824 => x"00000000",
         16825 => x"00000000",
         16826 => x"00000000",
         16827 => x"00000000",
         16828 => x"00000000",
         16829 => x"00000000",
         16830 => x"00000000",
         16831 => x"00000000",
         16832 => x"00000000",
         16833 => x"00000000",
         16834 => x"00000000",
         16835 => x"00000000",
         16836 => x"00000000",
         16837 => x"00000000",
         16838 => x"00000000",
         16839 => x"00000000",
         16840 => x"00000000",
         16841 => x"00000000",
         16842 => x"00000000",
         16843 => x"00000000",
         16844 => x"00000000",
         16845 => x"00000000",
         16846 => x"00000000",
         16847 => x"00000000",
         16848 => x"00000000",
         16849 => x"00000000",
         16850 => x"00000000",
         16851 => x"00000000",
         16852 => x"00000000",
         16853 => x"00000000",
         16854 => x"00000000",
         16855 => x"00000000",
         16856 => x"00000000",
         16857 => x"00000000",
         16858 => x"00000000",
         16859 => x"00000000",
         16860 => x"00000000",
         16861 => x"00000000",
         16862 => x"00000000",
         16863 => x"00000000",
         16864 => x"00000000",
         16865 => x"00000000",
         16866 => x"00000000",
         16867 => x"00000000",
         16868 => x"00000000",
         16869 => x"00000000",
         16870 => x"00000000",
         16871 => x"00000000",
         16872 => x"00000000",
         16873 => x"00000000",
         16874 => x"00000000",
         16875 => x"00000000",
         16876 => x"00000000",
         16877 => x"00000000",
         16878 => x"00000000",
         16879 => x"00000000",
         16880 => x"00000000",
         16881 => x"00000000",
         16882 => x"00000000",
         16883 => x"00000000",
         16884 => x"00000000",
         16885 => x"00000000",
         16886 => x"00000000",
         16887 => x"00000000",
         16888 => x"00000000",
         16889 => x"00000000",
         16890 => x"00000000",
         16891 => x"00000000",
         16892 => x"00000000",
         16893 => x"00000000",
         16894 => x"00000000",
         16895 => x"00000000",
         16896 => x"00000000",
         16897 => x"00000000",
         16898 => x"00000000",
         16899 => x"00000000",
         16900 => x"00000000",
         16901 => x"00000000",
         16902 => x"00000000",
         16903 => x"00000000",
         16904 => x"00000000",
         16905 => x"00000000",
         16906 => x"00000000",
         16907 => x"00000000",
         16908 => x"00000000",
         16909 => x"00000000",
         16910 => x"00000000",
         16911 => x"00000000",
         16912 => x"00000000",
         16913 => x"00000000",
         16914 => x"00000000",
         16915 => x"00000000",
         16916 => x"00000000",
         16917 => x"00000000",
         16918 => x"00000000",
         16919 => x"00000000",
         16920 => x"00000000",
         16921 => x"00000000",
         16922 => x"00000000",
         16923 => x"00000000",
         16924 => x"00000000",
         16925 => x"00000000",
         16926 => x"00000000",
         16927 => x"00000000",
         16928 => x"00000000",
         16929 => x"00000000",
         16930 => x"00000000",
         16931 => x"00000000",
         16932 => x"00000000",
         16933 => x"00000000",
         16934 => x"00000000",
         16935 => x"00000000",
         16936 => x"00000000",
         16937 => x"00000000",
         16938 => x"00000000",
         16939 => x"00000000",
         16940 => x"00000000",
         16941 => x"00000000",
         16942 => x"00000000",
         16943 => x"00000000",
         16944 => x"00000000",
         16945 => x"00000000",
         16946 => x"00000000",
         16947 => x"00000000",
         16948 => x"00000000",
         16949 => x"00000000",
         16950 => x"00000000",
         16951 => x"00000000",
         16952 => x"00000000",
         16953 => x"00000000",
         16954 => x"00000000",
         16955 => x"00000000",
         16956 => x"00000000",
         16957 => x"00000000",
         16958 => x"00000000",
         16959 => x"00000000",
         16960 => x"00000000",
         16961 => x"00000000",
         16962 => x"00000000",
         16963 => x"00000000",
         16964 => x"00000000",
         16965 => x"00000000",
         16966 => x"00000000",
         16967 => x"00000000",
         16968 => x"00000000",
         16969 => x"00000000",
         16970 => x"00000000",
         16971 => x"00000000",
         16972 => x"00000000",
         16973 => x"00000000",
         16974 => x"00000000",
         16975 => x"00000000",
         16976 => x"00000000",
         16977 => x"00000000",
         16978 => x"00000000",
         16979 => x"00000000",
         16980 => x"00000000",
         16981 => x"00000000",
         16982 => x"00000000",
         16983 => x"00000000",
         16984 => x"00000000",
         16985 => x"00000000",
         16986 => x"00000000",
         16987 => x"00000000",
         16988 => x"00000000",
         16989 => x"00000000",
         16990 => x"00000000",
         16991 => x"00000000",
         16992 => x"00000000",
         16993 => x"00000000",
         16994 => x"00000000",
         16995 => x"00000000",
         16996 => x"00000000",
         16997 => x"00000000",
         16998 => x"00000000",
         16999 => x"00000000",
         17000 => x"00000000",
         17001 => x"00000000",
         17002 => x"00000000",
         17003 => x"00000000",
         17004 => x"00000000",
         17005 => x"00000000",
         17006 => x"00000000",
         17007 => x"00000000",
         17008 => x"00000000",
         17009 => x"00000000",
         17010 => x"00000000",
         17011 => x"00000000",
         17012 => x"00000000",
         17013 => x"00000000",
         17014 => x"00000000",
         17015 => x"00000000",
         17016 => x"00000000",
         17017 => x"00000000",
         17018 => x"00000000",
         17019 => x"00000000",
         17020 => x"00000000",
         17021 => x"00000000",
         17022 => x"00000000",
         17023 => x"00000000",
         17024 => x"00000000",
         17025 => x"00000000",
         17026 => x"00000000",
         17027 => x"00000000",
         17028 => x"00000000",
         17029 => x"00000000",
         17030 => x"00000000",
         17031 => x"00000000",
         17032 => x"00000000",
         17033 => x"00000000",
         17034 => x"00000000",
         17035 => x"00000000",
         17036 => x"00000000",
         17037 => x"00000000",
         17038 => x"00000000",
         17039 => x"00000000",
         17040 => x"00000000",
         17041 => x"00000000",
         17042 => x"00000000",
         17043 => x"00000000",
         17044 => x"00000000",
         17045 => x"00000000",
         17046 => x"00000000",
         17047 => x"00000000",
         17048 => x"00000000",
         17049 => x"00000000",
         17050 => x"00000000",
         17051 => x"00000000",
         17052 => x"00000000",
         17053 => x"00000000",
         17054 => x"00000000",
         17055 => x"00000000",
         17056 => x"00000000",
         17057 => x"00000000",
         17058 => x"00000000",
         17059 => x"00000000",
         17060 => x"00000000",
         17061 => x"00000000",
         17062 => x"00000000",
         17063 => x"00000000",
         17064 => x"00000000",
         17065 => x"00000000",
         17066 => x"00000000",
         17067 => x"00000000",
         17068 => x"00000000",
         17069 => x"00000000",
         17070 => x"00000000",
         17071 => x"00000000",
         17072 => x"00000000",
         17073 => x"00000000",
         17074 => x"00000000",
         17075 => x"00000000",
         17076 => x"00000000",
         17077 => x"00000000",
         17078 => x"00000000",
         17079 => x"00000000",
         17080 => x"00000000",
         17081 => x"00000000",
         17082 => x"00000000",
         17083 => x"00000000",
         17084 => x"00000000",
         17085 => x"00000000",
         17086 => x"00000000",
         17087 => x"00000000",
         17088 => x"00000000",
         17089 => x"00000000",
         17090 => x"00000000",
         17091 => x"00000000",
         17092 => x"00000000",
         17093 => x"00000000",
         17094 => x"00000000",
         17095 => x"00000000",
         17096 => x"00000000",
         17097 => x"00000000",
         17098 => x"00000000",
         17099 => x"00000000",
         17100 => x"00000000",
         17101 => x"00000000",
         17102 => x"00000000",
         17103 => x"00000000",
         17104 => x"00000000",
         17105 => x"00000000",
         17106 => x"00000000",
         17107 => x"00000000",
         17108 => x"00000000",
         17109 => x"00000000",
         17110 => x"00000000",
         17111 => x"00000000",
         17112 => x"00000000",
         17113 => x"00000000",
         17114 => x"00000000",
         17115 => x"00000000",
         17116 => x"00000000",
         17117 => x"00000000",
         17118 => x"00000000",
         17119 => x"00000000",
         17120 => x"00000000",
         17121 => x"00000000",
         17122 => x"00000000",
         17123 => x"00000000",
         17124 => x"00000000",
         17125 => x"00000000",
         17126 => x"00000000",
         17127 => x"00000000",
         17128 => x"00000000",
         17129 => x"00000000",
         17130 => x"00000000",
         17131 => x"00000000",
         17132 => x"00000000",
         17133 => x"00000000",
         17134 => x"00000000",
         17135 => x"00000000",
         17136 => x"00000000",
         17137 => x"00000000",
         17138 => x"00000000",
         17139 => x"00000000",
         17140 => x"00000000",
         17141 => x"00000000",
         17142 => x"00000000",
         17143 => x"00000000",
         17144 => x"00000000",
         17145 => x"00000000",
         17146 => x"00000000",
         17147 => x"00000000",
         17148 => x"00000000",
         17149 => x"00000000",
         17150 => x"00000000",
         17151 => x"00000000",
         17152 => x"00000000",
         17153 => x"00000000",
         17154 => x"00000000",
         17155 => x"00000000",
         17156 => x"00000000",
         17157 => x"00000000",
         17158 => x"00000000",
         17159 => x"00000000",
         17160 => x"00000000",
         17161 => x"00000000",
         17162 => x"00000000",
         17163 => x"00000000",
         17164 => x"00000000",
         17165 => x"00000000",
         17166 => x"00000000",
         17167 => x"00000000",
         17168 => x"00000000",
         17169 => x"00000000",
         17170 => x"00000000",
         17171 => x"00000000",
         17172 => x"00000000",
         17173 => x"00000000",
         17174 => x"00000000",
         17175 => x"00000000",
         17176 => x"00000000",
         17177 => x"00000000",
         17178 => x"00000000",
         17179 => x"00000000",
         17180 => x"00000000",
         17181 => x"00000000",
         17182 => x"00000000",
         17183 => x"00000000",
         17184 => x"00000000",
         17185 => x"00000000",
         17186 => x"00000000",
         17187 => x"00000000",
         17188 => x"00000000",
         17189 => x"00000000",
         17190 => x"00000000",
         17191 => x"00000000",
         17192 => x"00000000",
         17193 => x"00000000",
         17194 => x"00000000",
         17195 => x"00000000",
         17196 => x"00000000",
         17197 => x"00000000",
         17198 => x"00000000",
         17199 => x"00000000",
         17200 => x"00000000",
         17201 => x"00000000",
         17202 => x"00000000",
         17203 => x"00000000",
         17204 => x"00000000",
         17205 => x"00000000",
         17206 => x"00000000",
         17207 => x"00000000",
         17208 => x"00000000",
         17209 => x"00000000",
         17210 => x"00000000",
         17211 => x"00000000",
         17212 => x"00000000",
         17213 => x"00000000",
         17214 => x"00000000",
         17215 => x"00000000",
         17216 => x"00000000",
         17217 => x"00000000",
         17218 => x"00000000",
         17219 => x"00000000",
         17220 => x"00000000",
         17221 => x"00000000",
         17222 => x"00000000",
         17223 => x"00000000",
         17224 => x"00000000",
         17225 => x"00000000",
         17226 => x"00000000",
         17227 => x"00000000",
         17228 => x"00000000",
         17229 => x"00000000",
         17230 => x"00000000",
         17231 => x"00000000",
         17232 => x"00000000",
         17233 => x"00000000",
         17234 => x"00000000",
         17235 => x"00000000",
         17236 => x"00000000",
         17237 => x"00000000",
         17238 => x"00000000",
         17239 => x"00000000",
         17240 => x"00000000",
         17241 => x"00000000",
         17242 => x"00000000",
         17243 => x"00000000",
         17244 => x"00000000",
         17245 => x"00000000",
         17246 => x"00000000",
         17247 => x"00000000",
         17248 => x"00000000",
         17249 => x"00000000",
         17250 => x"00000000",
         17251 => x"00000000",
         17252 => x"00000000",
         17253 => x"00000000",
         17254 => x"00000000",
         17255 => x"00000000",
         17256 => x"00000000",
         17257 => x"00000000",
         17258 => x"00000000",
         17259 => x"00000000",
         17260 => x"00000000",
         17261 => x"00000000",
         17262 => x"00000000",
         17263 => x"00000000",
         17264 => x"00000000",
         17265 => x"00000000",
         17266 => x"00000000",
         17267 => x"00000000",
         17268 => x"00000000",
         17269 => x"00000000",
         17270 => x"00000000",
         17271 => x"00000000",
         17272 => x"00000000",
         17273 => x"00000000",
         17274 => x"00000000",
         17275 => x"00000000",
         17276 => x"00000000",
         17277 => x"00000000",
         17278 => x"00000000",
         17279 => x"00000000",
         17280 => x"00000000",
         17281 => x"00000000",
         17282 => x"00000000",
         17283 => x"00000000",
         17284 => x"00000000",
         17285 => x"00000000",
         17286 => x"00000000",
         17287 => x"00000000",
         17288 => x"00000000",
         17289 => x"00000000",
         17290 => x"00000000",
         17291 => x"00000000",
         17292 => x"00000000",
         17293 => x"00000000",
         17294 => x"00000000",
         17295 => x"00000000",
         17296 => x"00000000",
         17297 => x"00000000",
         17298 => x"00000000",
         17299 => x"00000000",
         17300 => x"00000000",
         17301 => x"00000000",
         17302 => x"00000000",
         17303 => x"00000000",
         17304 => x"00000000",
         17305 => x"00000000",
         17306 => x"00000000",
         17307 => x"00000000",
         17308 => x"00000000",
         17309 => x"00000000",
         17310 => x"00000000",
         17311 => x"00000000",
         17312 => x"00000000",
         17313 => x"00000000",
         17314 => x"00000000",
         17315 => x"00000000",
         17316 => x"00000000",
         17317 => x"00000000",
         17318 => x"00000000",
         17319 => x"00000000",
         17320 => x"00000000",
         17321 => x"00000000",
         17322 => x"00000000",
         17323 => x"00000000",
         17324 => x"00000000",
         17325 => x"00000000",
         17326 => x"00000000",
         17327 => x"00000000",
         17328 => x"00000000",
         17329 => x"00000000",
         17330 => x"00000000",
         17331 => x"00000000",
         17332 => x"00000000",
         17333 => x"00000000",
         17334 => x"00000000",
         17335 => x"00000000",
         17336 => x"00000000",
         17337 => x"00000000",
         17338 => x"00000000",
         17339 => x"00000000",
         17340 => x"00000000",
         17341 => x"00000000",
         17342 => x"00000000",
         17343 => x"00000000",
         17344 => x"00000000",
         17345 => x"00000000",
         17346 => x"00000000",
         17347 => x"00000000",
         17348 => x"00000000",
         17349 => x"00000000",
         17350 => x"00000000",
         17351 => x"00000000",
         17352 => x"00000000",
         17353 => x"00000000",
         17354 => x"00000000",
         17355 => x"00000000",
         17356 => x"00000000",
         17357 => x"00000000",
         17358 => x"00000000",
         17359 => x"00000000",
         17360 => x"00000000",
         17361 => x"00000000",
         17362 => x"00000000",
         17363 => x"00000000",
         17364 => x"00000000",
         17365 => x"00000000",
         17366 => x"00000000",
         17367 => x"00000000",
         17368 => x"00000000",
         17369 => x"00000000",
         17370 => x"00000000",
         17371 => x"00000000",
         17372 => x"00000000",
         17373 => x"00000000",
         17374 => x"00000000",
         17375 => x"00000000",
         17376 => x"00000000",
         17377 => x"00000000",
         17378 => x"00000000",
         17379 => x"00000000",
         17380 => x"00000000",
         17381 => x"00000000",
         17382 => x"00000000",
         17383 => x"00000000",
         17384 => x"00000000",
         17385 => x"00000000",
         17386 => x"00000000",
         17387 => x"00000000",
         17388 => x"00000000",
         17389 => x"00000000",
         17390 => x"00000000",
         17391 => x"00000000",
         17392 => x"00000000",
         17393 => x"00000000",
         17394 => x"00000000",
         17395 => x"00000000",
         17396 => x"00000000",
         17397 => x"00000000",
         17398 => x"00000000",
         17399 => x"00000000",
         17400 => x"00000000",
         17401 => x"00000000",
         17402 => x"00000000",
         17403 => x"00000000",
         17404 => x"00000000",
         17405 => x"00000000",
         17406 => x"00000000",
         17407 => x"00000000",
         17408 => x"00000000",
         17409 => x"00000000",
         17410 => x"00000000",
         17411 => x"00000000",
         17412 => x"00000000",
         17413 => x"00000000",
         17414 => x"00000000",
         17415 => x"00000000",
         17416 => x"00000000",
         17417 => x"00000000",
         17418 => x"00000000",
         17419 => x"00000000",
         17420 => x"00000000",
         17421 => x"00000000",
         17422 => x"00000000",
         17423 => x"00000000",
         17424 => x"00000000",
         17425 => x"00000000",
         17426 => x"00000000",
         17427 => x"00000000",
         17428 => x"00000000",
         17429 => x"00000000",
         17430 => x"00000000",
         17431 => x"00000000",
         17432 => x"00000000",
         17433 => x"00000000",
         17434 => x"00000000",
         17435 => x"00000000",
         17436 => x"00000000",
         17437 => x"00000000",
         17438 => x"00000000",
         17439 => x"00000000",
         17440 => x"00000000",
         17441 => x"00000000",
         17442 => x"00000000",
         17443 => x"00000000",
         17444 => x"00000000",
         17445 => x"00000000",
         17446 => x"00000000",
         17447 => x"00000000",
         17448 => x"00000000",
         17449 => x"00000000",
         17450 => x"00000000",
         17451 => x"00000000",
         17452 => x"00000000",
         17453 => x"00000000",
         17454 => x"00000000",
         17455 => x"00000000",
         17456 => x"00000000",
         17457 => x"00000000",
         17458 => x"00000000",
         17459 => x"00000000",
         17460 => x"00000000",
         17461 => x"00000000",
         17462 => x"00000000",
         17463 => x"00000000",
         17464 => x"00000000",
         17465 => x"00000000",
         17466 => x"00000000",
         17467 => x"00000000",
         17468 => x"00000000",
         17469 => x"00000000",
         17470 => x"00000000",
         17471 => x"00000000",
         17472 => x"00000000",
         17473 => x"00000000",
         17474 => x"00000000",
         17475 => x"00000000",
         17476 => x"00000000",
         17477 => x"00000000",
         17478 => x"00000000",
         17479 => x"00000000",
         17480 => x"00000000",
         17481 => x"00000000",
         17482 => x"00000000",
         17483 => x"00000000",
         17484 => x"00000000",
         17485 => x"00000000",
         17486 => x"00000000",
         17487 => x"00000000",
         17488 => x"00000000",
         17489 => x"00000000",
         17490 => x"00000000",
         17491 => x"00000000",
         17492 => x"00000000",
         17493 => x"00000000",
         17494 => x"00000000",
         17495 => x"00000000",
         17496 => x"00000000",
         17497 => x"00000000",
         17498 => x"00000000",
         17499 => x"00000000",
         17500 => x"00000000",
         17501 => x"00000000",
         17502 => x"00000000",
         17503 => x"00000000",
         17504 => x"00000000",
         17505 => x"00000000",
         17506 => x"00000000",
         17507 => x"00000000",
         17508 => x"00000000",
         17509 => x"00000000",
         17510 => x"00000000",
         17511 => x"00000000",
         17512 => x"00000000",
         17513 => x"00000000",
         17514 => x"00000000",
         17515 => x"00000000",
         17516 => x"00000000",
         17517 => x"00000000",
         17518 => x"00000000",
         17519 => x"00000000",
         17520 => x"00000000",
         17521 => x"00000000",
         17522 => x"00000000",
         17523 => x"00000000",
         17524 => x"00000000",
         17525 => x"00000000",
         17526 => x"00000000",
         17527 => x"00000000",
         17528 => x"00000000",
         17529 => x"00000000",
         17530 => x"00000000",
         17531 => x"00000000",
         17532 => x"00000000",
         17533 => x"00000000",
         17534 => x"00000000",
         17535 => x"00000000",
         17536 => x"00000000",
         17537 => x"00000000",
         17538 => x"00000000",
         17539 => x"00000000",
         17540 => x"00000000",
         17541 => x"00000000",
         17542 => x"00000000",
         17543 => x"00000000",
         17544 => x"00000000",
         17545 => x"00000000",
         17546 => x"00000000",
         17547 => x"00000000",
         17548 => x"00000000",
         17549 => x"00000000",
         17550 => x"00000000",
         17551 => x"00000000",
         17552 => x"00000000",
         17553 => x"00000000",
         17554 => x"00000000",
         17555 => x"00000000",
         17556 => x"00000000",
         17557 => x"00000000",
         17558 => x"00000000",
         17559 => x"00000000",
         17560 => x"00000000",
         17561 => x"00000000",
         17562 => x"00000000",
         17563 => x"00000000",
         17564 => x"00000000",
         17565 => x"00000000",
         17566 => x"00000000",
         17567 => x"00000000",
         17568 => x"00000000",
         17569 => x"00000000",
         17570 => x"00000000",
         17571 => x"00000000",
         17572 => x"00000000",
         17573 => x"00000000",
         17574 => x"00000000",
         17575 => x"00000000",
         17576 => x"00000000",
         17577 => x"00000000",
         17578 => x"00000000",
         17579 => x"00000000",
         17580 => x"00000000",
         17581 => x"00000000",
         17582 => x"00000000",
         17583 => x"00000000",
         17584 => x"00000000",
         17585 => x"00000000",
         17586 => x"00000000",
         17587 => x"00000000",
         17588 => x"00000000",
         17589 => x"00000000",
         17590 => x"00000000",
         17591 => x"00000000",
         17592 => x"00000000",
         17593 => x"00000000",
         17594 => x"00000000",
         17595 => x"00000000",
         17596 => x"00000000",
         17597 => x"00000000",
         17598 => x"00000000",
         17599 => x"00000000",
         17600 => x"00000000",
         17601 => x"00000000",
         17602 => x"00000000",
         17603 => x"00000000",
         17604 => x"00000000",
         17605 => x"00000000",
         17606 => x"00000000",
         17607 => x"00000000",
         17608 => x"00000000",
         17609 => x"00000000",
         17610 => x"00000000",
         17611 => x"00000000",
         17612 => x"00000000",
         17613 => x"00000000",
         17614 => x"00000000",
         17615 => x"00000000",
         17616 => x"00000000",
         17617 => x"00000000",
         17618 => x"00000000",
         17619 => x"00000000",
         17620 => x"00000000",
         17621 => x"00000000",
         17622 => x"00000000",
         17623 => x"00000000",
         17624 => x"00000000",
         17625 => x"00000000",
         17626 => x"00000000",
         17627 => x"00000000",
         17628 => x"00000000",
         17629 => x"00000000",
         17630 => x"00000000",
         17631 => x"00000000",
         17632 => x"00000000",
         17633 => x"00000000",
         17634 => x"00000000",
         17635 => x"00000000",
         17636 => x"00000000",
         17637 => x"00000000",
         17638 => x"00000000",
         17639 => x"00000000",
         17640 => x"00000000",
         17641 => x"00000000",
         17642 => x"00000000",
         17643 => x"00000000",
         17644 => x"00000000",
         17645 => x"00000000",
         17646 => x"00000000",
         17647 => x"00000000",
         17648 => x"00000000",
         17649 => x"00000000",
         17650 => x"00000000",
         17651 => x"00000000",
         17652 => x"00000000",
         17653 => x"00000000",
         17654 => x"00000000",
         17655 => x"00000000",
         17656 => x"00000000",
         17657 => x"00000000",
         17658 => x"00000000",
         17659 => x"00000000",
         17660 => x"00000000",
         17661 => x"00000000",
         17662 => x"00000000",
         17663 => x"00000000",
         17664 => x"00000000",
         17665 => x"00000000",
         17666 => x"00000000",
         17667 => x"00000000",
         17668 => x"00000000",
         17669 => x"00000000",
         17670 => x"00000000",
         17671 => x"00000000",
         17672 => x"00000000",
         17673 => x"00000000",
         17674 => x"00000000",
         17675 => x"00000000",
         17676 => x"00000000",
         17677 => x"00000000",
         17678 => x"00000000",
         17679 => x"00000000",
         17680 => x"00000000",
         17681 => x"00000000",
         17682 => x"00000000",
         17683 => x"00000000",
         17684 => x"00000000",
         17685 => x"00000000",
         17686 => x"00000000",
         17687 => x"00000000",
         17688 => x"00000000",
         17689 => x"00000000",
         17690 => x"00000000",
         17691 => x"00000000",
         17692 => x"00000000",
         17693 => x"00000000",
         17694 => x"00000000",
         17695 => x"00000000",
         17696 => x"00000000",
         17697 => x"00000000",
         17698 => x"00000000",
         17699 => x"00000000",
         17700 => x"00000000",
         17701 => x"00000000",
         17702 => x"00000000",
         17703 => x"00000000",
         17704 => x"00000000",
         17705 => x"00000000",
         17706 => x"00000000",
         17707 => x"00000000",
         17708 => x"00000000",
         17709 => x"00000000",
         17710 => x"00000000",
         17711 => x"00000000",
         17712 => x"00000000",
         17713 => x"00000000",
         17714 => x"00000000",
         17715 => x"00000000",
         17716 => x"00000000",
         17717 => x"00000000",
         17718 => x"00000000",
         17719 => x"00000000",
         17720 => x"00000000",
         17721 => x"00000000",
         17722 => x"00000000",
         17723 => x"00000000",
         17724 => x"00000000",
         17725 => x"00000000",
         17726 => x"00000000",
         17727 => x"00000000",
         17728 => x"00000000",
         17729 => x"00000000",
         17730 => x"00000000",
         17731 => x"00000000",
         17732 => x"00000000",
         17733 => x"00000000",
         17734 => x"00000000",
         17735 => x"00000000",
         17736 => x"00000000",
         17737 => x"00000000",
         17738 => x"00000000",
         17739 => x"00000000",
         17740 => x"00000000",
         17741 => x"00000000",
         17742 => x"00000000",
         17743 => x"00000000",
         17744 => x"00000000",
         17745 => x"00000000",
         17746 => x"00000000",
         17747 => x"00000000",
         17748 => x"00000000",
         17749 => x"00000000",
         17750 => x"00000000",
         17751 => x"00000000",
         17752 => x"00000000",
         17753 => x"00000000",
         17754 => x"00000000",
         17755 => x"00000000",
         17756 => x"00000000",
         17757 => x"00000000",
         17758 => x"00000000",
         17759 => x"00000000",
         17760 => x"00000000",
         17761 => x"00000000",
         17762 => x"00000000",
         17763 => x"00000000",
         17764 => x"00000000",
         17765 => x"00000000",
         17766 => x"00000000",
         17767 => x"00000000",
         17768 => x"00000000",
         17769 => x"00000000",
         17770 => x"00000000",
         17771 => x"00000000",
         17772 => x"00000000",
         17773 => x"00000000",
         17774 => x"00000000",
         17775 => x"00000000",
         17776 => x"00000000",
         17777 => x"00000000",
         17778 => x"00000000",
         17779 => x"00000000",
         17780 => x"00000000",
         17781 => x"00000000",
         17782 => x"00000000",
         17783 => x"00000000",
         17784 => x"00000000",
         17785 => x"00000000",
         17786 => x"00000000",
         17787 => x"00000000",
         17788 => x"00000000",
         17789 => x"00000000",
         17790 => x"00000000",
         17791 => x"00000000",
         17792 => x"00000000",
         17793 => x"00000000",
         17794 => x"00000000",
         17795 => x"00000000",
         17796 => x"00000000",
         17797 => x"00000000",
         17798 => x"00000000",
         17799 => x"00000000",
         17800 => x"00000000",
         17801 => x"00000000",
         17802 => x"00000000",
         17803 => x"00000000",
         17804 => x"00000000",
         17805 => x"00000000",
         17806 => x"00000000",
         17807 => x"00000000",
         17808 => x"00000000",
         17809 => x"00000000",
         17810 => x"00000000",
         17811 => x"00000000",
         17812 => x"00000000",
         17813 => x"00000000",
         17814 => x"00000000",
         17815 => x"00000000",
         17816 => x"00000000",
         17817 => x"00000000",
         17818 => x"00000000",
         17819 => x"00000000",
         17820 => x"00000000",
         17821 => x"00000000",
         17822 => x"00000000",
         17823 => x"00000000",
         17824 => x"00000000",
         17825 => x"00000000",
         17826 => x"00000000",
         17827 => x"00000000",
         17828 => x"00000000",
         17829 => x"00000000",
         17830 => x"00000000",
         17831 => x"00000000",
         17832 => x"00000000",
         17833 => x"00000000",
         17834 => x"00000000",
         17835 => x"00000000",
         17836 => x"00000000",
         17837 => x"00000000",
         17838 => x"00000000",
         17839 => x"00000000",
         17840 => x"00000000",
         17841 => x"00000000",
         17842 => x"00000000",
         17843 => x"00000000",
         17844 => x"00000000",
         17845 => x"00000000",
         17846 => x"00000000",
         17847 => x"00000000",
         17848 => x"00000000",
         17849 => x"00000000",
         17850 => x"00000000",
         17851 => x"00000000",
         17852 => x"00000000",
         17853 => x"00000000",
         17854 => x"00000000",
         17855 => x"00000000",
         17856 => x"00000000",
         17857 => x"00000000",
         17858 => x"00000000",
         17859 => x"00000000",
         17860 => x"00000000",
         17861 => x"00000000",
         17862 => x"00000000",
         17863 => x"00000000",
         17864 => x"00000000",
         17865 => x"00000000",
         17866 => x"00000000",
         17867 => x"00000000",
         17868 => x"00000000",
         17869 => x"00000000",
         17870 => x"00000000",
         17871 => x"00000000",
         17872 => x"00000000",
         17873 => x"00000000",
         17874 => x"00000000",
         17875 => x"00000000",
         17876 => x"00000000",
         17877 => x"00000000",
         17878 => x"00000000",
         17879 => x"00000000",
         17880 => x"00000000",
         17881 => x"00000000",
         17882 => x"00000000",
         17883 => x"00000000",
         17884 => x"00000000",
         17885 => x"00000000",
         17886 => x"00000000",
         17887 => x"00000000",
         17888 => x"00000000",
         17889 => x"00000000",
         17890 => x"00000000",
         17891 => x"00000000",
         17892 => x"00000000",
         17893 => x"00000000",
         17894 => x"00000000",
         17895 => x"00000000",
         17896 => x"00000000",
         17897 => x"00000000",
         17898 => x"00000000",
         17899 => x"00000000",
         17900 => x"00000000",
         17901 => x"00000000",
         17902 => x"00000000",
         17903 => x"00000000",
         17904 => x"00000000",
         17905 => x"00000000",
         17906 => x"00000000",
         17907 => x"00000000",
         17908 => x"00000000",
         17909 => x"00000000",
         17910 => x"00000000",
         17911 => x"00000000",
         17912 => x"00000000",
         17913 => x"00000000",
         17914 => x"00000000",
         17915 => x"00000000",
         17916 => x"00000000",
         17917 => x"00000000",
         17918 => x"00000000",
         17919 => x"00000000",
         17920 => x"00000000",
         17921 => x"00000000",
         17922 => x"00000000",
         17923 => x"00000000",
         17924 => x"00000000",
         17925 => x"00000000",
         17926 => x"00000000",
         17927 => x"00000000",
         17928 => x"00000000",
         17929 => x"00000000",
         17930 => x"00000000",
         17931 => x"00000000",
         17932 => x"00000000",
         17933 => x"00000000",
         17934 => x"00000000",
         17935 => x"00000000",
         17936 => x"00000000",
         17937 => x"00000000",
         17938 => x"00000000",
         17939 => x"00000000",
         17940 => x"00000000",
         17941 => x"00000000",
         17942 => x"00000000",
         17943 => x"00000000",
         17944 => x"00000000",
         17945 => x"00000000",
         17946 => x"00000000",
         17947 => x"00000000",
         17948 => x"00000000",
         17949 => x"00000000",
         17950 => x"00000000",
         17951 => x"00000000",
         17952 => x"00000000",
         17953 => x"00000000",
         17954 => x"00000000",
         17955 => x"00000000",
         17956 => x"00000000",
         17957 => x"00000000",
         17958 => x"00000000",
         17959 => x"00000000",
         17960 => x"00000000",
         17961 => x"00000000",
         17962 => x"00000000",
         17963 => x"00000000",
         17964 => x"00000000",
         17965 => x"00000000",
         17966 => x"00000000",
         17967 => x"00000000",
         17968 => x"00000000",
         17969 => x"00000000",
         17970 => x"00000000",
         17971 => x"00000000",
         17972 => x"00000000",
         17973 => x"00000000",
         17974 => x"00000000",
         17975 => x"00000000",
         17976 => x"00000000",
         17977 => x"00000000",
         17978 => x"00000000",
         17979 => x"00000000",
         17980 => x"00000000",
         17981 => x"00000000",
         17982 => x"00000000",
         17983 => x"00000000",
         17984 => x"00000000",
         17985 => x"00000000",
         17986 => x"00000000",
         17987 => x"00000000",
         17988 => x"00000000",
         17989 => x"00000000",
         17990 => x"00000000",
         17991 => x"00000000",
         17992 => x"00000000",
         17993 => x"00000000",
         17994 => x"00000000",
         17995 => x"00000000",
         17996 => x"00000000",
         17997 => x"00000000",
         17998 => x"00000000",
         17999 => x"00000000",
         18000 => x"00000000",
         18001 => x"00000000",
         18002 => x"00000000",
         18003 => x"00000000",
         18004 => x"00000000",
         18005 => x"00000000",
         18006 => x"00000000",
         18007 => x"00000000",
         18008 => x"00000000",
         18009 => x"00000000",
         18010 => x"00000000",
         18011 => x"00000000",
         18012 => x"00000000",
         18013 => x"00000000",
         18014 => x"00000000",
         18015 => x"00000000",
         18016 => x"00000000",
         18017 => x"00000000",
         18018 => x"00000000",
         18019 => x"00000000",
         18020 => x"00000000",
         18021 => x"00000000",
         18022 => x"00000000",
         18023 => x"00000000",
         18024 => x"00000000",
         18025 => x"00000000",
         18026 => x"00000000",
         18027 => x"00000000",
         18028 => x"00000000",
         18029 => x"00000000",
         18030 => x"00000000",
         18031 => x"00000000",
         18032 => x"00000000",
         18033 => x"00000000",
         18034 => x"00000000",
         18035 => x"00000000",
         18036 => x"00000000",
         18037 => x"00000000",
         18038 => x"00000000",
         18039 => x"00000000",
         18040 => x"00000000",
         18041 => x"00000000",
         18042 => x"00000000",
         18043 => x"00000000",
         18044 => x"00000000",
         18045 => x"00000000",
         18046 => x"00000000",
         18047 => x"00000000",
         18048 => x"00000000",
         18049 => x"00000000",
         18050 => x"00000000",
         18051 => x"00000000",
         18052 => x"00000000",
         18053 => x"00000000",
         18054 => x"00000000",
         18055 => x"00000000",
         18056 => x"00000000",
         18057 => x"00000000",
         18058 => x"00000000",
         18059 => x"00000000",
         18060 => x"00000000",
         18061 => x"00000000",
         18062 => x"00000000",
         18063 => x"00000000",
         18064 => x"00000000",
         18065 => x"00000000",
         18066 => x"00000000",
         18067 => x"00000000",
         18068 => x"00000000",
         18069 => x"00000000",
         18070 => x"00000000",
         18071 => x"00000000",
         18072 => x"00000000",
         18073 => x"00000000",
         18074 => x"00000000",
         18075 => x"00000000",
         18076 => x"00000000",
         18077 => x"00000000",
         18078 => x"00000000",
         18079 => x"00000000",
         18080 => x"00000000",
         18081 => x"00000000",
         18082 => x"00000000",
         18083 => x"00000000",
         18084 => x"00000000",
         18085 => x"00000000",
         18086 => x"00000000",
         18087 => x"00000000",
         18088 => x"00000000",
         18089 => x"00000000",
         18090 => x"00000000",
         18091 => x"00000000",
         18092 => x"00000000",
         18093 => x"00000000",
         18094 => x"00000000",
         18095 => x"00000000",
         18096 => x"00000000",
         18097 => x"00000000",
         18098 => x"00000000",
         18099 => x"00000000",
         18100 => x"00000000",
         18101 => x"00000000",
         18102 => x"00000000",
         18103 => x"00000000",
         18104 => x"00000000",
         18105 => x"00000000",
         18106 => x"00000000",
         18107 => x"00000000",
         18108 => x"00000000",
         18109 => x"00000000",
         18110 => x"00000000",
         18111 => x"00000000",
         18112 => x"00000000",
         18113 => x"00000000",
         18114 => x"00000000",
         18115 => x"00000000",
         18116 => x"00000000",
         18117 => x"00000000",
         18118 => x"00000000",
         18119 => x"00000000",
         18120 => x"00000000",
         18121 => x"00000000",
         18122 => x"00000000",
         18123 => x"00000000",
         18124 => x"00000000",
         18125 => x"00000000",
         18126 => x"00000000",
         18127 => x"00000000",
         18128 => x"00000000",
         18129 => x"00000000",
         18130 => x"00000000",
         18131 => x"00000000",
         18132 => x"00000000",
         18133 => x"00000000",
         18134 => x"00000000",
         18135 => x"00000000",
         18136 => x"00000000",
         18137 => x"00000000",
         18138 => x"00000000",
         18139 => x"00000000",
         18140 => x"00000000",
         18141 => x"00000000",
         18142 => x"00000000",
         18143 => x"00000000",
         18144 => x"00000000",
         18145 => x"00000000",
         18146 => x"00000000",
         18147 => x"00000000",
         18148 => x"00000000",
         18149 => x"00000000",
         18150 => x"00000000",
         18151 => x"00000000",
         18152 => x"00000000",
         18153 => x"00000000",
         18154 => x"00000000",
         18155 => x"00000000",
         18156 => x"00000000",
         18157 => x"00000000",
         18158 => x"00000000",
         18159 => x"00000000",
         18160 => x"00000000",
         18161 => x"00000000",
         18162 => x"00000000",
         18163 => x"00000000",
         18164 => x"00000000",
         18165 => x"00000000",
         18166 => x"00000000",
         18167 => x"00000000",
         18168 => x"00000000",
         18169 => x"00000000",
         18170 => x"00000000",
         18171 => x"00000000",
         18172 => x"00000000",
         18173 => x"00000000",
         18174 => x"00000000",
         18175 => x"00000000",
         18176 => x"00000000",
         18177 => x"00000000",
         18178 => x"00000000",
         18179 => x"00000000",
         18180 => x"00000000",
         18181 => x"00000000",
         18182 => x"00000000",
         18183 => x"00000000",
         18184 => x"00000000",
         18185 => x"00000000",
         18186 => x"00000000",
         18187 => x"00000000",
         18188 => x"00000000",
         18189 => x"00000000",
         18190 => x"00000000",
         18191 => x"00000000",
         18192 => x"00000000",
         18193 => x"00000000",
         18194 => x"00000000",
         18195 => x"00000000",
         18196 => x"00000000",
         18197 => x"00000000",
         18198 => x"00000000",
         18199 => x"00000000",
         18200 => x"00000000",
         18201 => x"00000000",
         18202 => x"00000000",
         18203 => x"00000000",
         18204 => x"00000000",
         18205 => x"00003219",
         18206 => x"50000100",
         18207 => x"00000000",
         18208 => x"cce0f2f3",
         18209 => x"cecff6f7",
         18210 => x"f8f9fafb",
         18211 => x"fcfdfeff",
         18212 => x"e1c1c2c3",
         18213 => x"c4c5c6e2",
         18214 => x"e3e4e5e6",
         18215 => x"ebeeeff4",
         18216 => x"00616263",
         18217 => x"64656667",
         18218 => x"68696b6a",
         18219 => x"2f2a2e2d",
         18220 => x"20212223",
         18221 => x"24252627",
         18222 => x"28294f2c",
         18223 => x"512b5749",
         18224 => x"55010203",
         18225 => x"04050607",
         18226 => x"08090a0b",
         18227 => x"0c0d0e0f",
         18228 => x"10111213",
         18229 => x"14151617",
         18230 => x"18191a52",
         18231 => x"5954be3c",
         18232 => x"c7818283",
         18233 => x"84858687",
         18234 => x"88898a8b",
         18235 => x"8c8d8e8f",
         18236 => x"90919293",
         18237 => x"94959697",
         18238 => x"98999abc",
         18239 => x"8040a5c0",
         18240 => x"00000000",
         18241 => x"00000000",
         18242 => x"00000000",
         18243 => x"00000000",
         18244 => x"00000000",
         18245 => x"00000000",
         18246 => x"00000000",
         18247 => x"00000000",
         18248 => x"00000000",
         18249 => x"00000000",
         18250 => x"00000000",
         18251 => x"00000000",
         18252 => x"00000000",
         18253 => x"00000000",
         18254 => x"00000000",
         18255 => x"00000000",
         18256 => x"00000000",
         18257 => x"00000000",
         18258 => x"00000000",
         18259 => x"00000000",
         18260 => x"00000000",
         18261 => x"00000000",
         18262 => x"00000000",
         18263 => x"00000000",
         18264 => x"00000000",
         18265 => x"00000000",
         18266 => x"00000000",
         18267 => x"00000000",
         18268 => x"00000000",
         18269 => x"00000000",
         18270 => x"00020003",
         18271 => x"00040101",
         18272 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

